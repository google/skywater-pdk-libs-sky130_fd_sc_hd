* File: sky130_fd_sc_hd__sdfsbp_1.pxi.spice
* Created: Thu Aug 27 14:46:25 2020
* 
x_PM_SKY130_FD_SC_HD__SDFSBP_1%SCD N_SCD_c_283_n N_SCD_c_287_n N_SCD_c_284_n
+ N_SCD_M1039_g N_SCD_c_288_n N_SCD_M1021_g N_SCD_c_289_n SCD SCD
+ PM_SKY130_FD_SC_HD__SDFSBP_1%SCD
x_PM_SKY130_FD_SC_HD__SDFSBP_1%SCE N_SCE_M1012_g N_SCE_c_319_n N_SCE_M1002_g
+ N_SCE_M1026_g N_SCE_M1013_g SCE N_SCE_c_322_n N_SCE_c_342_n N_SCE_c_357_p
+ N_SCE_c_323_n N_SCE_c_324_n PM_SKY130_FD_SC_HD__SDFSBP_1%SCE
x_PM_SKY130_FD_SC_HD__SDFSBP_1%D N_D_c_421_n N_D_M1022_g N_D_M1004_g D D
+ N_D_c_424_n PM_SKY130_FD_SC_HD__SDFSBP_1%D
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_319_21# N_A_319_21#_M1013_s N_A_319_21#_M1026_s
+ N_A_319_21#_M1031_g N_A_319_21#_M1001_g N_A_319_21#_c_464_n
+ N_A_319_21#_c_465_n N_A_319_21#_c_466_n N_A_319_21#_c_467_n
+ N_A_319_21#_c_471_n N_A_319_21#_c_472_n PM_SKY130_FD_SC_HD__SDFSBP_1%A_319_21#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%CLK N_CLK_M1034_g N_CLK_c_536_n N_CLK_M1000_g
+ N_CLK_c_537_n N_CLK_c_542_n N_CLK_c_543_n CLK CLK CLK CLK N_CLK_c_540_n
+ N_CLK_c_541_n PM_SKY130_FD_SC_HD__SDFSBP_1%CLK
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_643_369# N_A_643_369#_M1000_s
+ N_A_643_369#_M1034_s N_A_643_369#_M1030_g N_A_643_369#_c_614_n
+ N_A_643_369#_M1036_g N_A_643_369#_c_615_n N_A_643_369#_c_616_n
+ N_A_643_369#_M1023_g N_A_643_369#_M1035_g N_A_643_369#_M1017_g
+ N_A_643_369#_M1015_g N_A_643_369#_c_618_n N_A_643_369#_c_647_n
+ N_A_643_369#_c_619_n N_A_643_369#_c_634_n N_A_643_369#_c_635_n
+ N_A_643_369#_c_620_n N_A_643_369#_c_621_n N_A_643_369#_c_710_p
+ N_A_643_369#_c_622_n N_A_643_369#_c_623_n N_A_643_369#_c_624_n
+ N_A_643_369#_c_625_n N_A_643_369#_c_626_n N_A_643_369#_c_627_n
+ N_A_643_369#_c_628_n N_A_643_369#_c_629_n N_A_643_369#_c_640_n
+ N_A_643_369#_c_641_n N_A_643_369#_c_642_n N_A_643_369#_c_643_n
+ N_A_643_369#_c_644_n N_A_643_369#_c_758_p N_A_643_369#_c_630_n
+ N_A_643_369#_c_645_n N_A_643_369#_c_646_n
+ PM_SKY130_FD_SC_HD__SDFSBP_1%A_643_369#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_809_369# N_A_809_369#_M1036_d
+ N_A_809_369#_M1030_d N_A_809_369#_c_919_n N_A_809_369#_c_909_n
+ N_A_809_369#_c_920_n N_A_809_369#_M1007_g N_A_809_369#_M1024_g
+ N_A_809_369#_M1006_g N_A_809_369#_c_922_n N_A_809_369#_M1040_g
+ N_A_809_369#_c_924_n N_A_809_369#_c_925_n N_A_809_369#_c_926_n
+ N_A_809_369#_c_1049_p N_A_809_369#_c_912_n N_A_809_369#_c_913_n
+ N_A_809_369#_c_914_n N_A_809_369#_c_915_n N_A_809_369#_c_916_n
+ N_A_809_369#_c_917_n N_A_809_369#_c_918_n
+ PM_SKY130_FD_SC_HD__SDFSBP_1%A_809_369#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_1129_21# N_A_1129_21#_M1009_s
+ N_A_1129_21#_M1008_d N_A_1129_21#_M1025_g N_A_1129_21#_M1037_g
+ N_A_1129_21#_c_1098_n N_A_1129_21#_c_1099_n N_A_1129_21#_c_1092_n
+ N_A_1129_21#_c_1100_n N_A_1129_21#_c_1101_n N_A_1129_21#_c_1093_n
+ N_A_1129_21#_c_1171_p N_A_1129_21#_c_1094_n N_A_1129_21#_c_1095_n
+ N_A_1129_21#_c_1096_n PM_SKY130_FD_SC_HD__SDFSBP_1%A_1129_21#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_997_413# N_A_997_413#_M1023_d
+ N_A_997_413#_M1007_d N_A_997_413#_c_1188_n N_A_997_413#_M1008_g
+ N_A_997_413#_c_1189_n N_A_997_413#_c_1190_n N_A_997_413#_M1009_g
+ N_A_997_413#_M1014_g N_A_997_413#_M1016_g N_A_997_413#_c_1191_n
+ N_A_997_413#_c_1192_n N_A_997_413#_c_1216_n N_A_997_413#_c_1203_n
+ N_A_997_413#_c_1193_n N_A_997_413#_c_1194_n N_A_997_413#_c_1195_n
+ N_A_997_413#_c_1196_n N_A_997_413#_c_1197_n N_A_997_413#_c_1198_n
+ N_A_997_413#_c_1199_n PM_SKY130_FD_SC_HD__SDFSBP_1%A_997_413#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%SET_B N_SET_B_M1032_g N_SET_B_M1041_g
+ N_SET_B_c_1344_n N_SET_B_M1028_g N_SET_B_M1010_g N_SET_B_c_1342_n
+ N_SET_B_c_1347_n N_SET_B_c_1348_n N_SET_B_c_1349_n N_SET_B_c_1350_n SET_B
+ N_SET_B_c_1352_n N_SET_B_c_1353_n N_SET_B_c_1354_n N_SET_B_c_1355_n
+ N_SET_B_c_1356_n N_SET_B_c_1357_n PM_SKY130_FD_SC_HD__SDFSBP_1%SET_B
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_1770_295# N_A_1770_295#_M1020_d
+ N_A_1770_295#_M1038_d N_A_1770_295#_M1011_g N_A_1770_295#_c_1495_n
+ N_A_1770_295#_c_1496_n N_A_1770_295#_M1018_g N_A_1770_295#_c_1488_n
+ N_A_1770_295#_c_1489_n N_A_1770_295#_c_1490_n N_A_1770_295#_c_1491_n
+ N_A_1770_295#_c_1499_n N_A_1770_295#_c_1500_n N_A_1770_295#_c_1492_n
+ N_A_1770_295#_c_1493_n N_A_1770_295#_c_1501_n
+ PM_SKY130_FD_SC_HD__SDFSBP_1%A_1770_295#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_1587_329# N_A_1587_329#_M1006_d
+ N_A_1587_329#_M1017_d N_A_1587_329#_M1028_d N_A_1587_329#_M1038_g
+ N_A_1587_329#_M1020_g N_A_1587_329#_c_1588_n N_A_1587_329#_c_1589_n
+ N_A_1587_329#_M1005_g N_A_1587_329#_M1029_g N_A_1587_329#_c_1590_n
+ N_A_1587_329#_M1033_g N_A_1587_329#_M1027_g N_A_1587_329#_c_1604_n
+ N_A_1587_329#_c_1592_n N_A_1587_329#_c_1593_n N_A_1587_329#_c_1615_n
+ N_A_1587_329#_c_1616_n N_A_1587_329#_c_1607_n N_A_1587_329#_c_1594_n
+ N_A_1587_329#_c_1608_n N_A_1587_329#_c_1595_n N_A_1587_329#_c_1596_n
+ N_A_1587_329#_c_1597_n N_A_1587_329#_c_1610_n N_A_1587_329#_c_1643_n
+ N_A_1587_329#_c_1611_n N_A_1587_329#_c_1612_n N_A_1587_329#_c_1653_n
+ N_A_1587_329#_c_1598_n PM_SKY130_FD_SC_HD__SDFSBP_1%A_1587_329#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_2412_47# N_A_2412_47#_M1033_s
+ N_A_2412_47#_M1027_s N_A_2412_47#_M1019_g N_A_2412_47#_M1003_g
+ N_A_2412_47#_c_1756_n N_A_2412_47#_c_1761_n N_A_2412_47#_c_1757_n
+ N_A_2412_47#_c_1758_n N_A_2412_47#_c_1772_n N_A_2412_47#_c_1759_n
+ PM_SKY130_FD_SC_HD__SDFSBP_1%A_2412_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_27_369# N_A_27_369#_M1021_s N_A_27_369#_M1001_d
+ N_A_27_369#_c_1803_n N_A_27_369#_c_1804_n N_A_27_369#_c_1805_n
+ N_A_27_369#_c_1811_n N_A_27_369#_c_1818_n N_A_27_369#_c_1806_n
+ PM_SKY130_FD_SC_HD__SDFSBP_1%A_27_369#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%VPWR N_VPWR_M1021_d N_VPWR_M1026_d N_VPWR_M1034_d
+ N_VPWR_M1037_d N_VPWR_M1032_d N_VPWR_M1011_d N_VPWR_M1038_s N_VPWR_M1029_s
+ N_VPWR_M1027_d N_VPWR_c_1852_n N_VPWR_c_1853_n N_VPWR_c_1854_n N_VPWR_c_1855_n
+ N_VPWR_c_1856_n N_VPWR_c_1857_n N_VPWR_c_1858_n N_VPWR_c_1859_n
+ N_VPWR_c_1860_n N_VPWR_c_1861_n N_VPWR_c_1862_n N_VPWR_c_1863_n
+ N_VPWR_c_1864_n VPWR N_VPWR_c_1865_n N_VPWR_c_1866_n N_VPWR_c_1867_n
+ N_VPWR_c_1868_n N_VPWR_c_1869_n N_VPWR_c_1870_n N_VPWR_c_1851_n
+ N_VPWR_c_1872_n N_VPWR_c_1873_n N_VPWR_c_1874_n N_VPWR_c_1875_n
+ N_VPWR_c_1876_n N_VPWR_c_1877_n N_VPWR_c_1878_n N_VPWR_c_1879_n VPWR
+ PM_SKY130_FD_SC_HD__SDFSBP_1%VPWR
x_PM_SKY130_FD_SC_HD__SDFSBP_1%A_181_47# N_A_181_47#_M1012_d N_A_181_47#_M1023_s
+ N_A_181_47#_M1004_d N_A_181_47#_M1007_s N_A_181_47#_c_2068_n
+ N_A_181_47#_c_2056_n N_A_181_47#_c_2061_n N_A_181_47#_c_2062_n
+ N_A_181_47#_c_2057_n N_A_181_47#_c_2071_n N_A_181_47#_c_2058_n
+ N_A_181_47#_c_2059_n N_A_181_47#_c_2064_n N_A_181_47#_c_2065_n
+ N_A_181_47#_c_2060_n N_A_181_47#_c_2067_n
+ PM_SKY130_FD_SC_HD__SDFSBP_1%A_181_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_1%Q_N N_Q_N_M1005_d N_Q_N_M1029_d Q_N Q_N Q_N Q_N
+ Q_N Q_N N_Q_N_c_2204_n PM_SKY130_FD_SC_HD__SDFSBP_1%Q_N
x_PM_SKY130_FD_SC_HD__SDFSBP_1%Q N_Q_M1019_d N_Q_M1003_d Q Q Q Q Q Q
+ N_Q_c_2223_n Q Q PM_SKY130_FD_SC_HD__SDFSBP_1%Q
x_PM_SKY130_FD_SC_HD__SDFSBP_1%VGND N_VGND_M1039_s N_VGND_M1031_d N_VGND_M1013_d
+ N_VGND_M1000_d N_VGND_M1025_d N_VGND_M1041_d N_VGND_M1010_d N_VGND_M1005_s
+ N_VGND_M1033_d N_VGND_c_2244_n N_VGND_c_2245_n N_VGND_c_2246_n N_VGND_c_2247_n
+ N_VGND_c_2248_n N_VGND_c_2249_n N_VGND_c_2250_n N_VGND_c_2251_n
+ N_VGND_c_2252_n N_VGND_c_2253_n N_VGND_c_2254_n N_VGND_c_2255_n
+ N_VGND_c_2256_n N_VGND_c_2257_n VGND N_VGND_c_2258_n N_VGND_c_2259_n
+ N_VGND_c_2260_n N_VGND_c_2261_n N_VGND_c_2262_n N_VGND_c_2263_n
+ N_VGND_c_2264_n N_VGND_c_2265_n N_VGND_c_2266_n N_VGND_c_2267_n
+ N_VGND_c_2268_n VGND PM_SKY130_FD_SC_HD__SDFSBP_1%VGND
cc_1 VNB N_SCD_c_283_n 0.0597753f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.325
cc_2 VNB N_SCD_c_284_n 0.0176456f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB SCD 0.02094f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_4 VNB N_SCE_M1012_g 0.0306921f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_5 VNB N_SCE_c_319_n 0.019383f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_6 VNB N_SCE_M1013_g 0.0380618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB SCE 0.00752716f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_8 VNB N_SCE_c_322_n 0.00910746f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_9 VNB N_SCE_c_323_n 0.0289071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_324_n 0.00122333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D_c_421_n 0.0164669f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.325
cc_12 VNB N_D_M1004_g 0.00862768f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.77
cc_13 VNB D 0.00527848f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_14 VNB N_D_c_424_n 0.0252553f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_15 VNB N_A_319_21#_M1031_g 0.0301639f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_16 VNB N_A_319_21#_c_464_n 0.00437998f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_17 VNB N_A_319_21#_c_465_n 0.0389075f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_18 VNB N_A_319_21#_c_466_n 0.0143935f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=0.85
cc_19 VNB N_A_319_21#_c_467_n 0.00705881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_CLK_c_536_n 0.017089f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_21 VNB N_CLK_c_537_n 0.0143095f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_22 VNB CLK 0.010708f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_23 VNB CLK 0.0136397f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=0.85
cc_24 VNB N_CLK_c_540_n 0.0164797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_CLK_c_541_n 0.0133943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_643_369#_c_614_n 0.0171953f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_27 VNB N_A_643_369#_c_615_n 0.051233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_643_369#_c_616_n 0.0170002f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_29 VNB N_A_643_369#_M1015_g 0.0234798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_643_369#_c_618_n 0.00552567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_643_369#_c_619_n 0.00133463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_643_369#_c_620_n 0.00586703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_643_369#_c_621_n 0.00228328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_643_369#_c_622_n 0.00316033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_643_369#_c_623_n 0.0160923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_643_369#_c_624_n 0.00196678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_643_369#_c_625_n 0.0263191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_643_369#_c_626_n 0.0103075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_643_369#_c_627_n 2.44915e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_643_369#_c_628_n 0.00417414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_643_369#_c_629_n 0.0283056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_643_369#_c_630_n 0.0110155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_809_369#_c_909_n 0.0426125f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_44 VNB N_A_809_369#_M1024_g 0.0306428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_809_369#_M1006_g 0.0362967f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=0.85
cc_46 VNB N_A_809_369#_c_912_n 0.0183981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_809_369#_c_913_n 0.00270322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_809_369#_c_914_n 0.00326418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_809_369#_c_915_n 0.0040767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_809_369#_c_916_n 0.00213039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_809_369#_c_917_n 0.0170178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_809_369#_c_918_n 0.00465628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1129_21#_M1025_g 0.0184566f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_54 VNB N_A_1129_21#_c_1092_n 0.00698964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1129_21#_c_1093_n 0.00466108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1129_21#_c_1094_n 0.00277762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1129_21#_c_1095_n 0.0285343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1129_21#_c_1096_n 0.0122702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_997_413#_c_1188_n 0.0189941f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_60 VNB N_A_997_413#_c_1189_n 0.0121485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_997_413#_c_1190_n 0.0163752f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_62 VNB N_A_997_413#_c_1191_n 0.0230071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_997_413#_c_1192_n 0.00674904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_997_413#_c_1193_n 0.00491887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_997_413#_c_1194_n 0.00176087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_997_413#_c_1195_n 0.00237739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_997_413#_c_1196_n 0.00479464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_997_413#_c_1197_n 0.0186258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_997_413#_c_1198_n 0.0109983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_997_413#_c_1199_n 0.0190763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_SET_B_M1041_g 0.0363083f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_72 VNB N_SET_B_M1010_g 0.0460164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_SET_B_c_1342_n 0.00804866f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=0.85
cc_74 VNB N_A_1770_295#_M1018_g 0.0227627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1770_295#_c_1488_n 0.00709852f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_76 VNB N_A_1770_295#_c_1489_n 8.65854e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1770_295#_c_1490_n 0.0290239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1770_295#_c_1491_n 0.00955884f $X=-0.19 $Y=-0.24 $X2=0.215
+ $Y2=1.53
cc_79 VNB N_A_1770_295#_c_1492_n 0.0078261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1770_295#_c_1493_n 0.00312069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1587_329#_c_1588_n 0.0476297f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_82 VNB N_A_1587_329#_c_1589_n 0.0238274f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_83 VNB N_A_1587_329#_c_1590_n 0.0485498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1587_329#_M1033_g 0.0331715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1587_329#_c_1592_n 0.004935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1587_329#_c_1593_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1587_329#_c_1594_n 0.00402188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1587_329#_c_1595_n 0.00287883f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1587_329#_c_1596_n 0.00685423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1587_329#_c_1597_n 0.0381676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1587_329#_c_1598_n 0.0206125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2412_47#_c_1756_n 0.00667692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_2412_47#_c_1757_n 0.00393517f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_94 VNB N_A_2412_47#_c_1758_n 0.0234543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2412_47#_c_1759_n 0.019962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VPWR_c_1851_n 0.554392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_181_47#_c_2056_n 0.00555327f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_98 VNB N_A_181_47#_c_2057_n 0.00327209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_181_47#_c_2058_n 9.84301e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_181_47#_c_2059_n 0.00128389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_181_47#_c_2060_n 0.00342661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_Q_N_c_2204_n 0.00698648f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=0.85
cc_103 VNB Q 0.00666696f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_104 VNB N_Q_c_2223_n 0.0152331f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.16
cc_105 VNB Q 0.022394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_2244_n 0.010916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2245_n 0.0174985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2246_n 0.0047534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2247_n 0.00603716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2248_n 4.108e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2249_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2250_n 0.00706343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2251_n 0.00606125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2252_n 0.0345333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2253_n 0.00343497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2254_n 0.0173287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2255_n 0.00529866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2256_n 0.0666076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2257_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2258_n 0.0153362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2259_n 0.055057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2260_n 0.0199057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2261_n 0.0332726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2262_n 0.0180194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2263_n 0.636166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2264_n 0.00409993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2265_n 0.0170817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2266_n 0.0166279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2267_n 0.00403597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2268_n 0.00394313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VPB N_SCD_c_283_n 0.00536633f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.325
cc_132 VPB N_SCD_c_287_n 0.0192739f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.62
cc_133 VPB N_SCD_c_288_n 0.0190089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.77
cc_134 VPB N_SCD_c_289_n 0.0260603f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_135 VPB SCD 0.0148824f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_136 VPB N_SCE_c_319_n 0.0131457f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_137 VPB N_SCE_M1002_g 0.0316859f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_138 VPB N_SCE_M1026_g 0.0507489f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_139 VPB SCE 0.00508528f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_140 VPB N_SCE_c_323_n 0.00635923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_SCE_c_324_n 0.0041855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_D_M1004_g 0.0334021f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.77
cc_143 VPB D 0.00612245f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_144 VPB N_A_319_21#_M1001_g 0.0422977f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_145 VPB N_A_319_21#_c_464_n 0.0098512f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_146 VPB N_A_319_21#_c_465_n 0.0139989f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_147 VPB N_A_319_21#_c_471_n 0.0040706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_319_21#_c_472_n 0.0119991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_CLK_c_542_n 0.0119079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_CLK_c_543_n 0.0309801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB CLK 0.00940396f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_152 VPB CLK 0.0079789f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_153 VPB N_CLK_c_540_n 0.0104614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_643_369#_M1030_g 0.0354172f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.695
cc_155 VPB N_A_643_369#_M1035_g 0.019201f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.16
cc_156 VPB N_A_643_369#_M1017_g 0.0242872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_643_369#_c_634_n 0.00144932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_643_369#_c_635_n 0.00165593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_643_369#_c_622_n 0.00314891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_643_369#_c_623_n 0.0105554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_643_369#_c_624_n 0.00131691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_643_369#_c_625_n 0.00502458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_643_369#_c_640_n 0.00472415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_643_369#_c_641_n 0.00584226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_643_369#_c_642_n 3.73476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_643_369#_c_643_n 0.00736633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_643_369#_c_644_n 0.00213153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_643_369#_c_645_n 0.0321882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_643_369#_c_646_n 0.00192244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_809_369#_c_919_n 0.0244169f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_171 VPB N_A_809_369#_c_920_n 0.0174418f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_172 VPB N_A_809_369#_M1006_g 0.0158967f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_173 VPB N_A_809_369#_c_922_n 0.0358849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_809_369#_M1040_g 0.0213215f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_175 VPB N_A_809_369#_c_924_n 0.0283114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_809_369#_c_925_n 0.00485301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_809_369#_c_926_n 0.00934509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_809_369#_c_914_n 0.00121793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_809_369#_c_915_n 3.90977e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_809_369#_c_916_n 0.00497366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_809_369#_c_917_n 0.0169522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1129_21#_M1037_g 0.0212875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1129_21#_c_1098_n 0.00176545f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_184 VPB N_A_1129_21#_c_1099_n 0.0370307f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_185 VPB N_A_1129_21#_c_1100_n 0.00551022f $X=-0.19 $Y=1.305 $X2=0.215
+ $Y2=1.53
cc_186 VPB N_A_1129_21#_c_1101_n 7.28078e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1129_21#_c_1096_n 0.0163815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_997_413#_c_1188_n 0.0093243f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_189 VPB N_A_997_413#_M1008_g 0.0472573f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.695
cc_190 VPB N_A_997_413#_M1016_g 0.0258061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_997_413#_c_1203_n 0.0126708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_997_413#_c_1193_n 0.00574591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_997_413#_c_1194_n 0.00282717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_997_413#_c_1195_n 0.00137632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_997_413#_c_1196_n 9.88491e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_997_413#_c_1197_n 0.00385999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_SET_B_M1032_g 0.0241123f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_198 VPB N_SET_B_c_1344_n 0.0190225f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_199 VPB N_SET_B_M1010_g 0.00750549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_SET_B_c_1342_n 0.00780115f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_201 VPB N_SET_B_c_1347_n 0.0322945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_SET_B_c_1348_n 0.0114467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_SET_B_c_1349_n 0.0103946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_SET_B_c_1350_n 0.0195847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB SET_B 0.00709599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_SET_B_c_1352_n 0.0153414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_SET_B_c_1353_n 0.00440092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_1354_n 0.00615367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_SET_B_c_1355_n 0.00370111f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_SET_B_c_1356_n 0.027252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_SET_B_c_1357_n 0.00813525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1770_295#_M1011_g 0.0382432f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.695
cc_213 VPB N_A_1770_295#_c_1495_n 0.0290745f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.695
cc_214 VPB N_A_1770_295#_c_1496_n 0.00653126f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_A_1770_295#_c_1488_n 0.0114128f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_216 VPB N_A_1770_295#_c_1491_n 0.00758554f $X=-0.19 $Y=1.305 $X2=0.215
+ $Y2=1.53
cc_217 VPB N_A_1770_295#_c_1499_n 6.44545e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1770_295#_c_1500_n 0.0200503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_1770_295#_c_1501_n 3.55501e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1587_329#_M1038_g 0.0262794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1587_329#_c_1588_n 0.0235554f $X=-0.19 $Y=1.305 $X2=0.327
+ $Y2=1.16
cc_222 VPB N_A_1587_329#_M1029_g 0.0274517f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_223 VPB N_A_1587_329#_c_1590_n 0.0242972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1587_329#_M1027_g 0.0439943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1587_329#_c_1604_n 0.0183001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1587_329#_c_1592_n 3.18387e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1587_329#_c_1593_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1587_329#_c_1607_n 0.00981719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_1587_329#_c_1608_n 0.00404031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_1587_329#_c_1597_n 9.35315e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_1587_329#_c_1610_n 0.00677623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_1587_329#_c_1611_n 0.0286225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_1587_329#_c_1612_n 0.0023123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_2412_47#_M1003_g 0.0238987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_2412_47#_c_1761_n 0.0120731f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_236 VPB N_A_2412_47#_c_1757_n 0.00506288f $X=-0.19 $Y=1.305 $X2=0.215
+ $Y2=1.53
cc_237 VPB N_A_2412_47#_c_1758_n 0.00557918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_27_369#_c_1803_n 0.0170416f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_239 VPB N_A_27_369#_c_1804_n 0.00111532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_27_369#_c_1805_n 0.00941534f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_241 VPB N_A_27_369#_c_1806_n 0.00262476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1852_n 0.00231024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1853_n 0.00982031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1854_n 4.05231e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1855_n 0.00562973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1856_n 0.00274169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1857_n 0.00492674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1858_n 0.00655454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1859_n 0.0343864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1860_n 0.00468577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1861_n 0.0463443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1862_n 0.00651315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1863_n 0.0508433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1864_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1865_n 0.0143786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1866_n 0.0154837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1867_n 0.0296156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1868_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1869_n 0.0173058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1870_n 0.0179894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1851_n 0.0864307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1872_n 0.00353358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1873_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1874_n 0.0199409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1875_n 0.0192332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1876_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1877_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1878_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1879_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_A_181_47#_c_2061_n 0.00388704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_A_181_47#_c_2062_n 0.00300602f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.16
cc_272 VPB N_A_181_47#_c_2057_n 0.00201708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_A_181_47#_c_2064_n 0.0319385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_A_181_47#_c_2065_n 0.0031324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_A_181_47#_c_2060_n 0.00329791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_A_181_47#_c_2067_n 0.00436874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_Q_N_c_2204_n 0.0107498f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_278 VPB Q 0.0311129f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_279 VPB Q 0.00899783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB Q 0.00666696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 N_SCD_c_283_n N_SCE_M1012_g 0.00595043f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_282 N_SCD_c_284_n N_SCE_M1012_g 0.0478814f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_283 SCD N_SCE_M1012_g 2.58702e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_284 N_SCD_c_283_n N_SCE_c_319_n 0.0200825f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_285 SCD N_SCE_c_319_n 3.42084e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_286 N_SCD_c_287_n N_SCE_M1002_g 0.00461989f $X=0.32 $Y=1.62 $X2=0 $Y2=0
cc_287 N_SCD_c_289_n N_SCE_M1002_g 0.0325519f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_288 SCD N_SCE_M1002_g 2.05572e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_289 N_SCD_c_283_n SCE 0.00609912f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_290 N_SCD_c_289_n SCE 5.18368e-19 $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_291 SCD SCE 0.0601261f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_292 SCD N_SCE_c_342_n 0.00158449f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_293 N_SCD_c_288_n N_A_27_369#_c_1804_n 0.0143471f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_294 N_SCD_c_283_n N_A_27_369#_c_1805_n 5.05332e-19 $X=0.32 $Y=1.325 $X2=0
+ $Y2=0
cc_295 N_SCD_c_289_n N_A_27_369#_c_1805_n 0.00301379f $X=0.47 $Y=1.695 $X2=0
+ $Y2=0
cc_296 SCD N_A_27_369#_c_1805_n 0.0229297f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_297 N_SCD_c_288_n N_A_27_369#_c_1811_n 4.53479e-19 $X=0.47 $Y=1.77 $X2=0
+ $Y2=0
cc_298 N_SCD_c_288_n N_VPWR_c_1852_n 0.00861999f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_299 N_SCD_c_288_n N_VPWR_c_1865_n 0.00346207f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_300 N_SCD_c_288_n N_VPWR_c_1851_n 0.00509645f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_301 N_SCD_c_284_n N_A_181_47#_c_2068_n 7.32861e-19 $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_302 N_SCD_c_283_n N_VGND_c_2245_n 0.00470012f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_303 N_SCD_c_284_n N_VGND_c_2245_n 0.018456f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_304 SCD N_VGND_c_2245_n 0.022355f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_305 N_SCD_c_284_n N_VGND_c_2252_n 0.00251889f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_306 N_SCD_c_284_n N_VGND_c_2263_n 0.00453995f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_307 SCD N_VGND_c_2263_n 0.00100835f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_308 N_SCE_M1012_g N_D_c_421_n 0.0148575f $X=0.83 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_309 N_SCE_c_319_n N_D_M1004_g 0.091197f $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_310 SCE N_D_M1004_g 6.20161e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_311 N_SCE_M1012_g D 0.00298976f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_312 N_SCE_c_319_n D 0.00289923f $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_313 SCE D 0.0530853f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_314 N_SCE_c_322_n D 0.0236806f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_315 N_SCE_c_342_n D 0.00219399f $X=0.84 $Y=1.19 $X2=0 $Y2=0
cc_316 N_SCE_M1012_g N_D_c_424_n 0.0194421f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_317 SCE N_D_c_424_n 3.44852e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_318 N_SCE_c_322_n N_D_c_424_n 0.00134139f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_319 N_SCE_M1026_g N_A_319_21#_c_464_n 0.00659955f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_320 N_SCE_M1013_g N_A_319_21#_c_464_n 0.00270542f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_321 N_SCE_c_322_n N_A_319_21#_c_464_n 0.0170338f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_322 N_SCE_c_357_p N_A_319_21#_c_464_n 6.89964e-19 $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_323 N_SCE_c_323_n N_A_319_21#_c_464_n 0.00254863f $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_SCE_c_324_n N_A_319_21#_c_464_n 0.0398188f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_325 N_SCE_c_322_n N_A_319_21#_c_465_n 0.00655791f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_326 N_SCE_c_323_n N_A_319_21#_c_465_n 0.0167027f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_327 N_SCE_c_324_n N_A_319_21#_c_465_n 6.5476e-19 $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_328 N_SCE_M1013_g N_A_319_21#_c_466_n 0.0052874f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_329 N_SCE_c_322_n N_A_319_21#_c_466_n 0.00905152f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_330 N_SCE_c_357_p N_A_319_21#_c_466_n 0.00100397f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_331 N_SCE_c_323_n N_A_319_21#_c_466_n 0.0028405f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_332 N_SCE_c_324_n N_A_319_21#_c_466_n 0.00947756f $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_SCE_M1013_g N_A_319_21#_c_467_n 0.00282117f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_334 N_SCE_M1026_g N_A_319_21#_c_472_n 0.00209962f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_335 N_SCE_c_323_n N_A_319_21#_c_472_n 4.82439e-19 $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_SCE_c_324_n N_A_319_21#_c_472_n 0.0105043f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_337 N_SCE_M1013_g N_CLK_c_537_n 0.00166043f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_338 N_SCE_M1013_g CLK 0.00585565f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_339 N_SCE_M1026_g CLK 0.00946284f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_340 N_SCE_c_324_n CLK 5.93234e-19 $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_341 N_SCE_M1026_g CLK 0.00157541f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_342 N_SCE_c_357_p CLK 0.0017785f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_343 N_SCE_c_323_n CLK 0.00323603f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_344 N_SCE_c_324_n CLK 0.034472f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_345 N_SCE_M1026_g N_CLK_c_540_n 0.00124122f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_346 N_SCE_c_323_n N_CLK_c_540_n 0.00327928f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_347 N_SCE_c_324_n N_CLK_c_540_n 3.62704e-19 $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_348 N_SCE_c_323_n N_CLK_c_541_n 0.00166043f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_349 N_SCE_M1026_g N_A_643_369#_c_647_n 0.00432238f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_350 N_SCE_M1013_g N_A_643_369#_c_619_n 0.00346504f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_SCE_M1013_g N_A_643_369#_c_621_n 5.16475e-19 $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_352 N_SCE_c_319_n N_A_27_369#_c_1804_n 7.48208e-19 $X=0.89 $Y=1.415 $X2=0
+ $Y2=0
cc_353 N_SCE_M1002_g N_A_27_369#_c_1804_n 0.0119179f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_354 SCE N_A_27_369#_c_1804_n 0.0186134f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_355 N_SCE_c_322_n N_A_27_369#_c_1804_n 0.00670567f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_356 N_SCE_c_342_n N_A_27_369#_c_1804_n 0.00141303f $X=0.84 $Y=1.19 $X2=0
+ $Y2=0
cc_357 N_SCE_M1002_g N_A_27_369#_c_1811_n 0.00502132f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_358 N_SCE_M1002_g N_A_27_369#_c_1818_n 0.00435752f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_359 N_SCE_M1002_g N_VPWR_c_1852_n 0.00279634f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_360 N_SCE_M1026_g N_VPWR_c_1853_n 0.00506557f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_361 N_SCE_M1002_g N_VPWR_c_1861_n 0.00418507f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_362 N_SCE_M1026_g N_VPWR_c_1861_n 0.00585385f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_363 N_SCE_M1002_g N_VPWR_c_1851_n 0.0055978f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_364 N_SCE_M1026_g N_VPWR_c_1851_n 0.0132032f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_365 N_SCE_M1012_g N_A_181_47#_c_2068_n 0.00520504f $X=0.83 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_SCE_c_322_n N_A_181_47#_c_2068_n 0.00829441f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_SCE_c_322_n N_A_181_47#_c_2071_n 0.0041843f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_SCE_c_322_n N_A_181_47#_c_2058_n 0.00449403f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_369 N_SCE_M1026_g N_A_181_47#_c_2064_n 0.00616318f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_370 N_SCE_c_322_n N_A_181_47#_c_2064_n 0.0490896f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_371 N_SCE_c_357_p N_A_181_47#_c_2064_n 0.0249445f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_372 N_SCE_c_323_n N_A_181_47#_c_2064_n 4.55029e-19 $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_SCE_c_324_n N_A_181_47#_c_2064_n 0.017162f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_374 N_SCE_c_322_n N_A_181_47#_c_2065_n 0.0258818f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_375 N_SCE_c_322_n N_A_181_47#_c_2060_n 0.0180487f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_376 N_SCE_M1012_g N_VGND_c_2245_n 0.00256902f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_377 N_SCE_M1013_g N_VGND_c_2246_n 0.00254064f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_378 N_SCE_c_322_n N_VGND_c_2246_n 0.00127321f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_379 N_SCE_M1013_g N_VGND_c_2247_n 0.0108433f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_380 N_SCE_c_324_n N_VGND_c_2247_n 2.63385e-19 $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_381 N_SCE_M1012_g N_VGND_c_2252_n 0.00540919f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_382 N_SCE_M1013_g N_VGND_c_2254_n 0.00486043f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_383 N_SCE_M1012_g N_VGND_c_2263_n 0.00743398f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_384 N_SCE_M1013_g N_VGND_c_2263_n 0.00965187f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_385 SCE N_VGND_c_2263_n 0.0111022f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_386 N_D_c_421_n N_A_319_21#_M1031_g 0.030873f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_387 D N_A_319_21#_M1031_g 3.19952e-19 $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_388 N_D_c_424_n N_A_319_21#_M1031_g 0.0201233f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_389 N_D_M1004_g N_A_319_21#_c_465_n 0.05672f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_390 D N_A_319_21#_c_465_n 0.00149798f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_391 N_D_M1004_g N_A_27_369#_c_1804_n 0.00142933f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_392 D N_A_27_369#_c_1804_n 0.00436538f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_393 N_D_M1004_g N_A_27_369#_c_1811_n 0.00434757f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_394 N_D_M1004_g N_A_27_369#_c_1806_n 0.0121184f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_395 D N_A_27_369#_c_1806_n 0.00493017f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_396 N_D_M1004_g N_VPWR_c_1861_n 0.00357877f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_397 N_D_M1004_g N_VPWR_c_1851_n 0.00515774f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_398 N_D_c_421_n N_A_181_47#_c_2068_n 0.010779f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_399 D N_A_181_47#_c_2068_n 0.0155023f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_400 N_D_c_424_n N_A_181_47#_c_2068_n 2.6926e-19 $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_401 N_D_M1004_g N_A_181_47#_c_2071_n 0.00302647f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_402 D N_A_181_47#_c_2071_n 0.00236045f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_403 N_D_c_421_n N_A_181_47#_c_2058_n 0.00235822f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_404 D N_A_181_47#_c_2065_n 0.00763197f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_405 N_D_c_421_n N_A_181_47#_c_2060_n 0.0012254f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_406 N_D_M1004_g N_A_181_47#_c_2060_n 0.00526995f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_407 D N_A_181_47#_c_2060_n 0.0668229f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_408 N_D_c_424_n N_A_181_47#_c_2060_n 0.00189474f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_409 N_D_c_421_n N_VGND_c_2252_n 0.00363059f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_410 N_D_c_421_n N_VGND_c_2263_n 0.00528803f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_411 N_A_319_21#_c_466_n CLK 0.00850801f $X=2.387 $Y=0.715 $X2=0 $Y2=0
cc_412 N_A_319_21#_c_472_n CLK 0.00581744f $X=2.4 $Y=1.99 $X2=0 $Y2=0
cc_413 N_A_319_21#_c_472_n N_A_27_369#_M1001_d 0.00524371f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_414 N_A_319_21#_M1001_g N_A_27_369#_c_1806_n 0.0091819f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_415 N_A_319_21#_c_471_n N_A_27_369#_c_1806_n 0.0148151f $X=2.395 $Y=1.927
+ $X2=0 $Y2=0
cc_416 N_A_319_21#_c_472_n N_A_27_369#_c_1806_n 0.0132953f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_417 N_A_319_21#_M1001_g N_VPWR_c_1861_n 0.00357877f $X=1.67 $Y=2.165 $X2=0
+ $Y2=0
cc_418 N_A_319_21#_c_471_n N_VPWR_c_1861_n 0.0154197f $X=2.395 $Y=1.927 $X2=0
+ $Y2=0
cc_419 N_A_319_21#_c_472_n N_VPWR_c_1861_n 0.00432835f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_420 N_A_319_21#_M1026_s N_VPWR_c_1851_n 0.00261392f $X=2.275 $Y=1.845 $X2=0
+ $Y2=0
cc_421 N_A_319_21#_M1001_g N_VPWR_c_1851_n 0.00657041f $X=1.67 $Y=2.165 $X2=0
+ $Y2=0
cc_422 N_A_319_21#_c_471_n N_VPWR_c_1851_n 0.00941222f $X=2.395 $Y=1.927 $X2=0
+ $Y2=0
cc_423 N_A_319_21#_c_472_n N_VPWR_c_1851_n 0.00699224f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_424 N_A_319_21#_M1001_g N_A_181_47#_c_2071_n 0.0048545f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_425 N_A_319_21#_c_472_n N_A_181_47#_c_2071_n 0.0170257f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_426 N_A_319_21#_M1031_g N_A_181_47#_c_2058_n 0.0130996f $X=1.67 $Y=0.445
+ $X2=0 $Y2=0
cc_427 N_A_319_21#_c_467_n N_A_181_47#_c_2058_n 0.00478561f $X=2.43 $Y=0.44
+ $X2=0 $Y2=0
cc_428 N_A_319_21#_c_464_n N_A_181_47#_c_2064_n 0.0169458f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_429 N_A_319_21#_c_465_n N_A_181_47#_c_2064_n 0.00172463f $X=1.95 $Y=1.16
+ $X2=0 $Y2=0
cc_430 N_A_319_21#_c_472_n N_A_181_47#_c_2064_n 0.0111897f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_431 N_A_319_21#_M1001_g N_A_181_47#_c_2065_n 0.00423017f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_432 N_A_319_21#_c_464_n N_A_181_47#_c_2065_n 0.0027962f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_433 N_A_319_21#_M1031_g N_A_181_47#_c_2060_n 0.00584437f $X=1.67 $Y=0.445
+ $X2=0 $Y2=0
cc_434 N_A_319_21#_M1001_g N_A_181_47#_c_2060_n 0.0107523f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_435 N_A_319_21#_c_464_n N_A_181_47#_c_2060_n 0.0614598f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_436 N_A_319_21#_c_465_n N_A_181_47#_c_2060_n 0.0084262f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_437 N_A_319_21#_c_466_n N_A_181_47#_c_2060_n 0.0152187f $X=2.387 $Y=0.715
+ $X2=0 $Y2=0
cc_438 N_A_319_21#_c_467_n N_A_181_47#_c_2060_n 2.89284e-19 $X=2.43 $Y=0.44
+ $X2=0 $Y2=0
cc_439 N_A_319_21#_c_472_n N_A_181_47#_c_2060_n 0.00797602f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_440 N_A_319_21#_M1031_g N_VGND_c_2246_n 0.00570299f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_A_319_21#_c_465_n N_VGND_c_2246_n 0.00128608f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_442 N_A_319_21#_c_466_n N_VGND_c_2246_n 0.010779f $X=2.387 $Y=0.715 $X2=0
+ $Y2=0
cc_443 N_A_319_21#_c_467_n N_VGND_c_2246_n 0.0166348f $X=2.43 $Y=0.44 $X2=0
+ $Y2=0
cc_444 N_A_319_21#_M1031_g N_VGND_c_2252_n 0.00453652f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_445 N_A_319_21#_c_466_n N_VGND_c_2254_n 0.00401857f $X=2.387 $Y=0.715 $X2=0
+ $Y2=0
cc_446 N_A_319_21#_c_467_n N_VGND_c_2254_n 0.0171533f $X=2.43 $Y=0.44 $X2=0
+ $Y2=0
cc_447 N_A_319_21#_M1013_s N_VGND_c_2263_n 0.00382897f $X=2.305 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_A_319_21#_M1031_g N_VGND_c_2263_n 0.00851114f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_319_21#_c_466_n N_VGND_c_2263_n 0.00745898f $X=2.387 $Y=0.715 $X2=0
+ $Y2=0
cc_450 N_A_319_21#_c_467_n N_VGND_c_2263_n 0.00964668f $X=2.43 $Y=0.44 $X2=0
+ $Y2=0
cc_451 N_CLK_c_542_n N_A_643_369#_M1030_g 0.00717124f $X=3.52 $Y=1.62 $X2=0
+ $Y2=0
cc_452 N_CLK_c_543_n N_A_643_369#_M1030_g 0.0306795f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_453 CLK N_A_643_369#_M1030_g 2.31516e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_454 N_CLK_c_536_n N_A_643_369#_c_614_n 0.0138064f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_455 N_CLK_c_537_n N_A_643_369#_c_618_n 0.00767217f $X=3.58 $Y=0.805 $X2=0
+ $Y2=0
cc_456 CLK N_A_643_369#_c_647_n 3.35151e-19 $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_457 N_CLK_c_536_n N_A_643_369#_c_619_n 0.00270983f $X=3.58 $Y=0.73 $X2=0
+ $Y2=0
cc_458 N_CLK_c_543_n N_A_643_369#_c_634_n 0.0147667f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_459 CLK N_A_643_369#_c_634_n 0.00781016f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_460 N_CLK_c_543_n N_A_643_369#_c_635_n 3.33785e-19 $X=3.52 $Y=1.77 $X2=0
+ $Y2=0
cc_461 CLK N_A_643_369#_c_635_n 0.0150671f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_462 CLK N_A_643_369#_c_635_n 0.0114033f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_463 N_CLK_c_540_n N_A_643_369#_c_635_n 6.22831e-19 $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_464 N_CLK_c_536_n N_A_643_369#_c_620_n 0.00396355f $X=3.58 $Y=0.73 $X2=0
+ $Y2=0
cc_465 N_CLK_c_537_n N_A_643_369#_c_620_n 0.00637134f $X=3.58 $Y=0.805 $X2=0
+ $Y2=0
cc_466 CLK N_A_643_369#_c_620_n 0.00793982f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_467 N_CLK_c_541_n N_A_643_369#_c_620_n 0.00151794f $X=3.43 $Y=1.09 $X2=0
+ $Y2=0
cc_468 N_CLK_c_537_n N_A_643_369#_c_621_n 0.00352145f $X=3.58 $Y=0.805 $X2=0
+ $Y2=0
cc_469 CLK N_A_643_369#_c_621_n 0.0136403f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_470 CLK N_A_643_369#_c_621_n 0.016055f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_471 N_CLK_c_540_n N_A_643_369#_c_621_n 8.54762e-19 $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_472 N_CLK_c_541_n N_A_643_369#_c_621_n 5.61645e-19 $X=3.43 $Y=1.09 $X2=0
+ $Y2=0
cc_473 N_CLK_c_542_n N_A_643_369#_c_622_n 3.32736e-19 $X=3.52 $Y=1.62 $X2=0
+ $Y2=0
cc_474 N_CLK_c_543_n N_A_643_369#_c_622_n 0.00192453f $X=3.52 $Y=1.77 $X2=0
+ $Y2=0
cc_475 CLK N_A_643_369#_c_622_n 0.0052596f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_476 CLK N_A_643_369#_c_622_n 0.00543392f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_477 CLK N_A_643_369#_c_622_n 0.042042f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_478 N_CLK_c_541_n N_A_643_369#_c_622_n 0.00366024f $X=3.43 $Y=1.09 $X2=0
+ $Y2=0
cc_479 CLK N_A_643_369#_c_623_n 3.7897e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_480 N_CLK_c_540_n N_A_643_369#_c_623_n 0.0213743f $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_481 N_CLK_c_543_n N_A_643_369#_c_642_n 4.69296e-19 $X=3.52 $Y=1.77 $X2=0
+ $Y2=0
cc_482 N_CLK_c_541_n N_A_643_369#_c_630_n 0.0064798f $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_483 CLK N_VPWR_M1026_d 0.00205233f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_484 N_CLK_c_543_n N_VPWR_c_1853_n 0.00413466f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_485 CLK N_VPWR_c_1853_n 0.00968055f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_486 N_CLK_c_543_n N_VPWR_c_1854_n 0.00818001f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_487 N_CLK_c_543_n N_VPWR_c_1866_n 0.0046653f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_488 CLK N_VPWR_c_1866_n 8.13541e-19 $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_489 N_CLK_c_543_n N_VPWR_c_1851_n 0.00562323f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_490 CLK N_VPWR_c_1851_n 0.0019648f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_491 N_CLK_c_542_n N_A_181_47#_c_2064_n 0.00245154f $X=3.52 $Y=1.62 $X2=0
+ $Y2=0
cc_492 N_CLK_c_543_n N_A_181_47#_c_2064_n 0.00182678f $X=3.52 $Y=1.77 $X2=0
+ $Y2=0
cc_493 CLK N_A_181_47#_c_2064_n 5.20642e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_494 CLK N_A_181_47#_c_2064_n 0.00542825f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_495 CLK N_A_181_47#_c_2064_n 0.0328531f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_496 N_CLK_c_536_n N_VGND_c_2247_n 0.00215264f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_497 CLK N_VGND_c_2247_n 0.0103825f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_498 N_CLK_c_536_n N_VGND_c_2248_n 0.00757678f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_499 N_CLK_c_536_n N_VGND_c_2258_n 0.00362954f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_500 N_CLK_c_537_n N_VGND_c_2258_n 2.82692e-19 $X=3.58 $Y=0.805 $X2=0 $Y2=0
cc_501 CLK N_VGND_c_2258_n 0.00110113f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_502 N_CLK_c_536_n N_VGND_c_2263_n 0.00567184f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_503 CLK N_VGND_c_2263_n 0.0024143f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_504 N_A_643_369#_c_641_n N_A_809_369#_M1030_d 0.00106464f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_505 N_A_643_369#_c_642_n N_A_809_369#_M1030_d 4.96569e-19 $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_506 N_A_643_369#_M1030_g N_A_809_369#_c_919_n 0.0121191f $X=3.97 $Y=2.165
+ $X2=0 $Y2=0
cc_507 N_A_643_369#_c_641_n N_A_809_369#_c_919_n 0.00109505f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_508 N_A_643_369#_c_645_n N_A_809_369#_c_919_n 0.0032436f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_509 N_A_643_369#_c_645_n N_A_809_369#_c_909_n 0.0085606f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_510 N_A_643_369#_c_646_n N_A_809_369#_c_909_n 2.0638e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_511 N_A_643_369#_c_616_n N_A_809_369#_M1024_g 0.0193318f $X=4.94 $Y=0.73
+ $X2=0 $Y2=0
cc_512 N_A_643_369#_M1017_g N_A_809_369#_M1006_g 0.0143377f $X=7.86 $Y=2.065
+ $X2=0 $Y2=0
cc_513 N_A_643_369#_M1015_g N_A_809_369#_M1006_g 0.0168783f $X=8.96 $Y=0.445
+ $X2=0 $Y2=0
cc_514 N_A_643_369#_c_624_n N_A_809_369#_M1006_g 0.00455669f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_515 N_A_643_369#_c_625_n N_A_809_369#_M1006_g 0.021266f $X=7.92 $Y=1.16 $X2=0
+ $Y2=0
cc_516 N_A_643_369#_c_626_n N_A_809_369#_M1006_g 0.0158174f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_517 N_A_643_369#_c_628_n N_A_809_369#_M1006_g 0.00137775f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_518 N_A_643_369#_c_629_n N_A_809_369#_M1006_g 0.0115051f $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_519 N_A_643_369#_c_640_n N_A_809_369#_M1006_g 0.00173186f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_520 N_A_643_369#_M1017_g N_A_809_369#_c_922_n 0.00438518f $X=7.86 $Y=2.065
+ $X2=0 $Y2=0
cc_521 N_A_643_369#_c_626_n N_A_809_369#_c_922_n 0.00124012f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_522 N_A_643_369#_c_640_n N_A_809_369#_c_922_n 8.84937e-19 $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_523 N_A_643_369#_M1017_g N_A_809_369#_M1040_g 0.0127652f $X=7.86 $Y=2.065
+ $X2=0 $Y2=0
cc_524 N_A_643_369#_c_640_n N_A_809_369#_M1040_g 0.00111273f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_525 N_A_643_369#_M1035_g N_A_809_369#_c_924_n 0.0161622f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_526 N_A_643_369#_c_641_n N_A_809_369#_c_924_n 0.00560081f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_527 N_A_643_369#_c_644_n N_A_809_369#_c_924_n 7.24988e-19 $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_528 N_A_643_369#_c_645_n N_A_809_369#_c_924_n 0.00461659f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_529 N_A_643_369#_c_646_n N_A_809_369#_c_924_n 5.74415e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_530 N_A_643_369#_c_641_n N_A_809_369#_c_925_n 0.00228522f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_531 N_A_643_369#_M1030_g N_A_809_369#_c_926_n 0.0100044f $X=3.97 $Y=2.165
+ $X2=0 $Y2=0
cc_532 N_A_643_369#_c_710_p N_A_809_369#_c_926_n 0.0121614f $X=3.865 $Y=1.775
+ $X2=0 $Y2=0
cc_533 N_A_643_369#_c_641_n N_A_809_369#_c_926_n 0.0190932f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_534 N_A_643_369#_c_642_n N_A_809_369#_c_926_n 0.00348404f $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_535 N_A_643_369#_c_615_n N_A_809_369#_c_912_n 0.00100605f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_536 N_A_643_369#_c_624_n N_A_809_369#_c_912_n 0.0170797f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_537 N_A_643_369#_c_625_n N_A_809_369#_c_912_n 0.00419944f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_538 N_A_643_369#_c_626_n N_A_809_369#_c_912_n 0.0147683f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_539 N_A_643_369#_c_640_n N_A_809_369#_c_912_n 0.00221057f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_540 N_A_643_369#_c_641_n N_A_809_369#_c_912_n 0.0075219f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_541 N_A_643_369#_c_643_n N_A_809_369#_c_912_n 0.0472312f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_542 N_A_643_369#_c_644_n N_A_809_369#_c_912_n 0.0126603f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_543 N_A_643_369#_c_646_n N_A_809_369#_c_912_n 6.70475e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_544 N_A_643_369#_c_615_n N_A_809_369#_c_913_n 0.00234075f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_545 N_A_643_369#_c_622_n N_A_809_369#_c_913_n 0.00138833f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_546 N_A_643_369#_c_615_n N_A_809_369#_c_914_n 0.00183262f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_547 N_A_643_369#_c_623_n N_A_809_369#_c_914_n 0.0031868f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_548 N_A_643_369#_c_624_n N_A_809_369#_c_915_n 0.00187989f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_549 N_A_643_369#_c_625_n N_A_809_369#_c_915_n 4.43515e-19 $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_550 N_A_643_369#_c_626_n N_A_809_369#_c_915_n 0.00465135f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_551 N_A_643_369#_c_628_n N_A_809_369#_c_915_n 0.00559275f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_552 N_A_643_369#_c_629_n N_A_809_369#_c_915_n 0.00344514f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_553 N_A_643_369#_M1017_g N_A_809_369#_c_916_n 0.00113007f $X=7.86 $Y=2.065
+ $X2=0 $Y2=0
cc_554 N_A_643_369#_c_624_n N_A_809_369#_c_916_n 0.0133976f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_555 N_A_643_369#_c_625_n N_A_809_369#_c_916_n 8.43582e-19 $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_556 N_A_643_369#_c_626_n N_A_809_369#_c_916_n 0.0144046f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_557 N_A_643_369#_c_628_n N_A_809_369#_c_916_n 0.00843986f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_558 N_A_643_369#_c_629_n N_A_809_369#_c_916_n 0.00117437f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_559 N_A_643_369#_c_640_n N_A_809_369#_c_916_n 0.0178429f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_560 N_A_643_369#_c_615_n N_A_809_369#_c_917_n 0.0487935f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_561 N_A_643_369#_c_622_n N_A_809_369#_c_917_n 3.00848e-19 $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_562 N_A_643_369#_c_623_n N_A_809_369#_c_917_n 0.0203131f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_563 N_A_643_369#_c_614_n N_A_809_369#_c_918_n 0.00458005f $X=4 $Y=0.73 $X2=0
+ $Y2=0
cc_564 N_A_643_369#_c_615_n N_A_809_369#_c_918_n 0.0132045f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_565 N_A_643_369#_c_620_n N_A_809_369#_c_918_n 0.0129402f $X=3.735 $Y=0.8
+ $X2=0 $Y2=0
cc_566 N_A_643_369#_c_622_n N_A_809_369#_c_918_n 0.0649873f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_567 N_A_643_369#_c_630_n N_A_809_369#_c_918_n 0.0031868f $X=3.917 $Y=1.09
+ $X2=0 $Y2=0
cc_568 N_A_643_369#_M1035_g N_A_1129_21#_M1037_g 0.0211742f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_569 N_A_643_369#_c_643_n N_A_1129_21#_M1037_g 0.00304183f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_570 N_A_643_369#_c_643_n N_A_1129_21#_c_1098_n 0.0108654f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_571 N_A_643_369#_c_643_n N_A_1129_21#_c_1099_n 0.0039051f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_572 N_A_643_369#_c_645_n N_A_1129_21#_c_1099_n 0.0130435f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_573 N_A_643_369#_c_640_n N_A_1129_21#_c_1100_n 7.99648e-19 $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_574 N_A_643_369#_c_643_n N_A_1129_21#_c_1100_n 0.0238856f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_575 N_A_643_369#_c_643_n N_A_1129_21#_c_1101_n 0.00322176f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_576 N_A_643_369#_c_643_n N_A_997_413#_M1008_g 0.00365451f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_577 N_A_643_369#_M1017_g N_A_997_413#_M1016_g 0.080634f $X=7.86 $Y=2.065
+ $X2=0 $Y2=0
cc_578 N_A_643_369#_c_624_n N_A_997_413#_M1016_g 0.00111359f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_579 N_A_643_369#_c_640_n N_A_997_413#_M1016_g 0.0186626f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_580 N_A_643_369#_c_758_p N_A_997_413#_M1016_g 0.00166818f $X=7.59 $Y=1.87
+ $X2=0 $Y2=0
cc_581 N_A_643_369#_c_615_n N_A_997_413#_c_1192_n 0.0042049f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_582 N_A_643_369#_c_616_n N_A_997_413#_c_1192_n 0.00613402f $X=4.94 $Y=0.73
+ $X2=0 $Y2=0
cc_583 N_A_643_369#_M1035_g N_A_997_413#_c_1216_n 0.0121756f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_584 N_A_643_369#_c_641_n N_A_997_413#_c_1216_n 0.00379337f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_585 N_A_643_369#_c_643_n N_A_997_413#_c_1216_n 0.00492445f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_586 N_A_643_369#_c_644_n N_A_997_413#_c_1216_n 0.00506476f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_587 N_A_643_369#_c_645_n N_A_997_413#_c_1216_n 9.46198e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_588 N_A_643_369#_c_646_n N_A_997_413#_c_1216_n 0.0108411f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_589 N_A_643_369#_M1035_g N_A_997_413#_c_1203_n 0.00392912f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_590 N_A_643_369#_c_643_n N_A_997_413#_c_1203_n 0.0149262f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_591 N_A_643_369#_c_644_n N_A_997_413#_c_1203_n 0.00307458f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_592 N_A_643_369#_c_645_n N_A_997_413#_c_1203_n 0.00212617f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_593 N_A_643_369#_c_646_n N_A_997_413#_c_1203_n 0.0263544f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_594 N_A_643_369#_c_641_n N_A_997_413#_c_1193_n 0.00396196f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_595 N_A_643_369#_c_643_n N_A_997_413#_c_1193_n 0.00354029f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_596 N_A_643_369#_c_644_n N_A_997_413#_c_1193_n 0.0032583f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_597 N_A_643_369#_c_645_n N_A_997_413#_c_1193_n 0.00293864f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_598 N_A_643_369#_c_646_n N_A_997_413#_c_1193_n 0.014754f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_599 N_A_643_369#_c_643_n N_A_997_413#_c_1194_n 0.00736646f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_600 N_A_643_369#_c_624_n N_A_997_413#_c_1196_n 0.0257532f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_601 N_A_643_369#_c_625_n N_A_997_413#_c_1196_n 0.00191578f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_602 N_A_643_369#_c_640_n N_A_997_413#_c_1196_n 0.0237306f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_603 N_A_643_369#_c_624_n N_A_997_413#_c_1197_n 3.8924e-19 $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_604 N_A_643_369#_c_625_n N_A_997_413#_c_1197_n 0.0210994f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_605 N_A_643_369#_c_640_n N_A_997_413#_c_1197_n 0.00266154f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_606 N_A_643_369#_c_640_n N_A_997_413#_c_1198_n 0.00583817f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_607 N_A_643_369#_c_643_n N_A_997_413#_c_1198_n 0.00170959f $X=7.445 $Y=1.87
+ $X2=0 $Y2=0
cc_608 N_A_643_369#_c_624_n N_A_997_413#_c_1199_n 0.00180149f $X=7.92 $Y=1.16
+ $X2=0 $Y2=0
cc_609 N_A_643_369#_c_627_n N_A_997_413#_c_1199_n 0.00302498f $X=8.005 $Y=0.795
+ $X2=0 $Y2=0
cc_610 N_A_643_369#_c_643_n N_SET_B_M1032_g 0.00451304f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_611 N_A_643_369#_c_640_n SET_B 0.0213138f $X=7.835 $Y=1.725 $X2=0 $Y2=0
cc_612 N_A_643_369#_c_643_n SET_B 0.00815691f $X=7.445 $Y=1.87 $X2=0 $Y2=0
cc_613 N_A_643_369#_M1017_g N_SET_B_c_1352_n 6.92361e-19 $X=7.86 $Y=2.065 $X2=0
+ $Y2=0
cc_614 N_A_643_369#_c_624_n N_SET_B_c_1352_n 0.00478454f $X=7.92 $Y=1.16 $X2=0
+ $Y2=0
cc_615 N_A_643_369#_c_625_n N_SET_B_c_1352_n 7.93137e-19 $X=7.92 $Y=1.16 $X2=0
+ $Y2=0
cc_616 N_A_643_369#_c_626_n N_SET_B_c_1352_n 0.00555644f $X=8.81 $Y=0.795 $X2=0
+ $Y2=0
cc_617 N_A_643_369#_c_628_n N_SET_B_c_1352_n 4.06665e-19 $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_618 N_A_643_369#_c_629_n N_SET_B_c_1352_n 0.00119869f $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_619 N_A_643_369#_c_640_n N_SET_B_c_1352_n 0.0309316f $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_620 N_A_643_369#_c_643_n N_SET_B_c_1352_n 0.0446385f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_621 N_A_643_369#_c_758_p N_SET_B_c_1352_n 0.0249445f $X=7.59 $Y=1.87 $X2=0
+ $Y2=0
cc_622 N_A_643_369#_c_640_n N_SET_B_c_1353_n 2.70806e-19 $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_623 N_A_643_369#_c_643_n N_SET_B_c_1353_n 0.0264998f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_624 N_A_643_369#_c_628_n N_SET_B_c_1354_n 0.00332589f $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_625 N_A_643_369#_c_628_n N_SET_B_c_1355_n 0.0106848f $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_626 N_A_643_369#_c_629_n N_SET_B_c_1355_n 3.93267e-19 $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_627 N_A_643_369#_c_640_n N_SET_B_c_1356_n 0.00378468f $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_628 N_A_643_369#_c_643_n N_SET_B_c_1356_n 0.00379442f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_629 N_A_643_369#_c_640_n N_SET_B_c_1357_n 0.00102452f $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_630 N_A_643_369#_c_628_n N_A_1770_295#_c_1496_n 3.03e-19 $X=8.9 $Y=1.08 $X2=0
+ $Y2=0
cc_631 N_A_643_369#_c_629_n N_A_1770_295#_c_1496_n 0.0108867f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_632 N_A_643_369#_M1015_g N_A_1770_295#_M1018_g 0.0359432f $X=8.96 $Y=0.445
+ $X2=0 $Y2=0
cc_633 N_A_643_369#_c_626_n N_A_1770_295#_M1018_g 0.00204989f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_634 N_A_643_369#_M1015_g N_A_1770_295#_c_1489_n 3.90915e-19 $X=8.96 $Y=0.445
+ $X2=0 $Y2=0
cc_635 N_A_643_369#_c_626_n N_A_1770_295#_c_1489_n 0.00242692f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_636 N_A_643_369#_c_628_n N_A_1770_295#_c_1489_n 0.0159294f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_637 N_A_643_369#_c_628_n N_A_1770_295#_c_1490_n 0.00202708f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_638 N_A_643_369#_c_629_n N_A_1770_295#_c_1490_n 0.0359432f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_639 N_A_643_369#_c_628_n N_A_1770_295#_c_1499_n 0.00363474f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_640 N_A_643_369#_c_626_n N_A_1587_329#_M1006_d 0.00279878f $X=8.81 $Y=0.795
+ $X2=-0.19 $Y2=-0.24
cc_641 N_A_643_369#_c_640_n N_A_1587_329#_M1017_d 0.00444765f $X=7.835 $Y=1.725
+ $X2=0 $Y2=0
cc_642 N_A_643_369#_M1017_g N_A_1587_329#_c_1615_n 0.00140068f $X=7.86 $Y=2.065
+ $X2=0 $Y2=0
cc_643 N_A_643_369#_M1015_g N_A_1587_329#_c_1616_n 0.0106703f $X=8.96 $Y=0.445
+ $X2=0 $Y2=0
cc_644 N_A_643_369#_c_626_n N_A_1587_329#_c_1616_n 0.0274979f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_645 N_A_643_369#_c_629_n N_A_1587_329#_c_1616_n 3.14717e-19 $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_646 N_A_643_369#_c_626_n N_A_1587_329#_c_1594_n 0.00509298f $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_647 N_A_643_369#_c_626_n N_A_1587_329#_c_1595_n 3.76722e-19 $X=8.81 $Y=0.795
+ $X2=0 $Y2=0
cc_648 N_A_643_369#_c_628_n N_A_1587_329#_c_1612_n 8.16162e-19 $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_649 N_A_643_369#_c_629_n N_A_1587_329#_c_1612_n 0.00144538f $X=8.9 $Y=1.08
+ $X2=0 $Y2=0
cc_650 N_A_643_369#_c_634_n N_VPWR_M1034_d 7.20981e-19 $X=3.735 $Y=1.865 $X2=0
+ $Y2=0
cc_651 N_A_643_369#_c_710_p N_VPWR_M1034_d 0.00104088f $X=3.865 $Y=1.775 $X2=0
+ $Y2=0
cc_652 N_A_643_369#_c_642_n N_VPWR_M1034_d 0.00130251f $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_653 N_A_643_369#_c_640_n N_VPWR_M1032_d 0.00676884f $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_654 N_A_643_369#_c_643_n N_VPWR_M1032_d 2.72657e-19 $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_655 N_A_643_369#_c_647_n N_VPWR_c_1853_n 0.0118221f $X=3.34 $Y=2.16 $X2=0
+ $Y2=0
cc_656 N_A_643_369#_M1030_g N_VPWR_c_1854_n 0.00823695f $X=3.97 $Y=2.165 $X2=0
+ $Y2=0
cc_657 N_A_643_369#_c_634_n N_VPWR_c_1854_n 0.00350403f $X=3.735 $Y=1.865 $X2=0
+ $Y2=0
cc_658 N_A_643_369#_c_710_p N_VPWR_c_1854_n 0.005559f $X=3.865 $Y=1.775 $X2=0
+ $Y2=0
cc_659 N_A_643_369#_c_642_n N_VPWR_c_1854_n 0.00178155f $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_660 N_A_643_369#_c_643_n N_VPWR_c_1855_n 0.00119067f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_661 N_A_643_369#_M1030_g N_VPWR_c_1863_n 0.0046653f $X=3.97 $Y=2.165 $X2=0
+ $Y2=0
cc_662 N_A_643_369#_M1035_g N_VPWR_c_1863_n 0.00357877f $X=5.33 $Y=2.275 $X2=0
+ $Y2=0
cc_663 N_A_643_369#_c_647_n N_VPWR_c_1866_n 0.00597665f $X=3.34 $Y=2.16 $X2=0
+ $Y2=0
cc_664 N_A_643_369#_M1034_s N_VPWR_c_1851_n 0.00391264f $X=3.215 $Y=1.845 $X2=0
+ $Y2=0
cc_665 N_A_643_369#_M1030_g N_VPWR_c_1851_n 0.0053279f $X=3.97 $Y=2.165 $X2=0
+ $Y2=0
cc_666 N_A_643_369#_M1035_g N_VPWR_c_1851_n 0.00539327f $X=5.33 $Y=2.275 $X2=0
+ $Y2=0
cc_667 N_A_643_369#_c_647_n N_VPWR_c_1851_n 0.00593257f $X=3.34 $Y=2.16 $X2=0
+ $Y2=0
cc_668 N_A_643_369#_c_634_n N_VPWR_c_1851_n 0.00605909f $X=3.735 $Y=1.865 $X2=0
+ $Y2=0
cc_669 N_A_643_369#_c_710_p N_VPWR_c_1851_n 0.00132255f $X=3.865 $Y=1.775 $X2=0
+ $Y2=0
cc_670 N_A_643_369#_c_640_n N_VPWR_c_1851_n 0.0036075f $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_671 N_A_643_369#_c_641_n N_VPWR_c_1851_n 0.0529551f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_672 N_A_643_369#_c_642_n N_VPWR_c_1851_n 0.0150349f $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_673 N_A_643_369#_c_643_n N_VPWR_c_1851_n 0.091386f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_674 N_A_643_369#_c_644_n N_VPWR_c_1851_n 0.0156394f $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_675 N_A_643_369#_c_758_p N_VPWR_c_1851_n 0.0143849f $X=7.59 $Y=1.87 $X2=0
+ $Y2=0
cc_676 N_A_643_369#_M1017_g N_VPWR_c_1875_n 0.0199371f $X=7.86 $Y=2.065 $X2=0
+ $Y2=0
cc_677 N_A_643_369#_c_640_n N_VPWR_c_1875_n 0.0431194f $X=7.835 $Y=1.725 $X2=0
+ $Y2=0
cc_678 N_A_643_369#_c_643_n N_VPWR_c_1875_n 0.00805283f $X=7.445 $Y=1.87 $X2=0
+ $Y2=0
cc_679 N_A_643_369#_c_758_p N_VPWR_c_1875_n 0.00338024f $X=7.59 $Y=1.87 $X2=0
+ $Y2=0
cc_680 N_A_643_369#_c_615_n N_A_181_47#_c_2056_n 0.00755734f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_681 N_A_643_369#_c_616_n N_A_181_47#_c_2056_n 0.00248143f $X=4.94 $Y=0.73
+ $X2=0 $Y2=0
cc_682 N_A_643_369#_c_641_n N_A_181_47#_c_2061_n 6.0342e-19 $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_683 N_A_643_369#_c_645_n N_A_181_47#_c_2061_n 2.97233e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_684 N_A_643_369#_c_646_n N_A_181_47#_c_2061_n 0.00145132f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_685 N_A_643_369#_M1035_g N_A_181_47#_c_2062_n 2.14528e-19 $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_686 N_A_643_369#_c_641_n N_A_181_47#_c_2062_n 0.0164833f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_687 N_A_643_369#_c_644_n N_A_181_47#_c_2062_n 0.00280193f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_688 N_A_643_369#_c_645_n N_A_181_47#_c_2062_n 0.00239438f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_689 N_A_643_369#_c_646_n N_A_181_47#_c_2062_n 0.0106469f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_690 N_A_643_369#_c_615_n N_A_181_47#_c_2059_n 0.00896128f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_691 N_A_643_369#_M1030_g N_A_181_47#_c_2064_n 0.00390687f $X=3.97 $Y=2.165
+ $X2=0 $Y2=0
cc_692 N_A_643_369#_c_618_n N_A_181_47#_c_2064_n 0.00230404f $X=3.992 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_A_643_369#_c_634_n N_A_181_47#_c_2064_n 0.0104627f $X=3.735 $Y=1.865
+ $X2=0 $Y2=0
cc_694 N_A_643_369#_c_635_n N_A_181_47#_c_2064_n 0.00440811f $X=3.425 $Y=1.865
+ $X2=0 $Y2=0
cc_695 N_A_643_369#_c_620_n N_A_181_47#_c_2064_n 0.00559677f $X=3.735 $Y=0.8
+ $X2=0 $Y2=0
cc_696 N_A_643_369#_c_621_n N_A_181_47#_c_2064_n 7.07979e-19 $X=3.455 $Y=0.8
+ $X2=0 $Y2=0
cc_697 N_A_643_369#_c_622_n N_A_181_47#_c_2064_n 0.021893f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_698 N_A_643_369#_c_623_n N_A_181_47#_c_2064_n 4.51301e-19 $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_699 N_A_643_369#_c_641_n N_A_181_47#_c_2064_n 0.0490514f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_700 N_A_643_369#_c_642_n N_A_181_47#_c_2064_n 0.0254571f $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_701 N_A_643_369#_c_641_n N_A_181_47#_c_2067_n 0.0264737f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_702 N_A_643_369#_c_645_n N_A_181_47#_c_2067_n 0.00127036f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_703 N_A_643_369#_c_646_n N_A_181_47#_c_2067_n 0.00208921f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_704 N_A_643_369#_c_640_n A_1514_329# 4.80034e-19 $X=7.835 $Y=1.725 $X2=-0.19
+ $Y2=-0.24
cc_705 N_A_643_369#_c_758_p A_1514_329# 0.00159144f $X=7.59 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_706 N_A_643_369#_c_619_n N_VGND_c_2247_n 0.0184198f $X=3.37 $Y=0.44 $X2=0
+ $Y2=0
cc_707 N_A_643_369#_c_614_n N_VGND_c_2248_n 0.00822761f $X=4 $Y=0.73 $X2=0 $Y2=0
cc_708 N_A_643_369#_c_620_n N_VGND_c_2248_n 0.0207423f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_709 N_A_643_369#_c_623_n N_VGND_c_2248_n 4.22312e-19 $X=3.91 $Y=1.255 $X2=0
+ $Y2=0
cc_710 N_A_643_369#_M1015_g N_VGND_c_2256_n 0.00362032f $X=8.96 $Y=0.445 $X2=0
+ $Y2=0
cc_711 N_A_643_369#_c_626_n N_VGND_c_2256_n 0.00572424f $X=8.81 $Y=0.795 $X2=0
+ $Y2=0
cc_712 N_A_643_369#_c_627_n N_VGND_c_2256_n 0.00289816f $X=8.005 $Y=0.795 $X2=0
+ $Y2=0
cc_713 N_A_643_369#_c_619_n N_VGND_c_2258_n 0.0125902f $X=3.37 $Y=0.44 $X2=0
+ $Y2=0
cc_714 N_A_643_369#_c_620_n N_VGND_c_2258_n 0.00247138f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_715 N_A_643_369#_c_614_n N_VGND_c_2259_n 0.00471416f $X=4 $Y=0.73 $X2=0 $Y2=0
cc_716 N_A_643_369#_c_615_n N_VGND_c_2259_n 0.00382237f $X=4.865 $Y=0.805 $X2=0
+ $Y2=0
cc_717 N_A_643_369#_c_616_n N_VGND_c_2259_n 0.00564131f $X=4.94 $Y=0.73 $X2=0
+ $Y2=0
cc_718 N_A_643_369#_c_620_n N_VGND_c_2259_n 8.20832e-19 $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_719 N_A_643_369#_M1000_s N_VGND_c_2263_n 0.00323692f $X=3.245 $Y=0.235 $X2=0
+ $Y2=0
cc_720 N_A_643_369#_c_614_n N_VGND_c_2263_n 0.00836944f $X=4 $Y=0.73 $X2=0 $Y2=0
cc_721 N_A_643_369#_c_615_n N_VGND_c_2263_n 0.00372099f $X=4.865 $Y=0.805 $X2=0
+ $Y2=0
cc_722 N_A_643_369#_c_616_n N_VGND_c_2263_n 0.0115324f $X=4.94 $Y=0.73 $X2=0
+ $Y2=0
cc_723 N_A_643_369#_M1015_g N_VGND_c_2263_n 0.00559388f $X=8.96 $Y=0.445 $X2=0
+ $Y2=0
cc_724 N_A_643_369#_c_619_n N_VGND_c_2263_n 0.00703355f $X=3.37 $Y=0.44 $X2=0
+ $Y2=0
cc_725 N_A_643_369#_c_620_n N_VGND_c_2263_n 0.00665853f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_726 N_A_643_369#_c_626_n N_VGND_c_2263_n 0.01133f $X=8.81 $Y=0.795 $X2=0
+ $Y2=0
cc_727 N_A_643_369#_c_627_n N_VGND_c_2263_n 0.00489372f $X=8.005 $Y=0.795 $X2=0
+ $Y2=0
cc_728 N_A_643_369#_c_627_n N_VGND_c_2266_n 0.00854165f $X=8.005 $Y=0.795 $X2=0
+ $Y2=0
cc_729 N_A_643_369#_c_626_n A_1514_47# 0.00430463f $X=8.81 $Y=0.795 $X2=-0.19
+ $Y2=-0.24
cc_730 N_A_643_369#_c_627_n A_1514_47# 0.00655491f $X=8.005 $Y=0.795 $X2=-0.19
+ $Y2=-0.24
cc_731 N_A_809_369#_M1024_g N_A_1129_21#_M1025_g 0.0610902f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_732 N_A_809_369#_c_912_n N_A_1129_21#_c_1098_n 5.84337e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_733 N_A_809_369#_c_912_n N_A_1129_21#_c_1092_n 0.00810105f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_734 N_A_809_369#_M1024_g N_A_1129_21#_c_1094_n 0.00121075f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_735 N_A_809_369#_c_912_n N_A_1129_21#_c_1094_n 0.00959352f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_736 N_A_809_369#_c_912_n N_A_1129_21#_c_1095_n 0.00455149f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_737 N_A_809_369#_M1024_g N_A_1129_21#_c_1096_n 0.00652836f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_738 N_A_809_369#_c_912_n N_A_1129_21#_c_1096_n 0.0025903f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_739 N_A_809_369#_c_912_n N_A_997_413#_c_1188_n 0.0012497f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_740 N_A_809_369#_c_909_n N_A_997_413#_c_1192_n 0.0138219f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_741 N_A_809_369#_M1024_g N_A_997_413#_c_1192_n 0.0212478f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_742 N_A_809_369#_c_912_n N_A_997_413#_c_1192_n 0.0327595f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_743 N_A_809_369#_c_909_n N_A_997_413#_c_1193_n 0.00618953f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_744 N_A_809_369#_c_912_n N_A_997_413#_c_1193_n 0.0236092f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_745 N_A_809_369#_c_917_n N_A_997_413#_c_1193_n 3.67923e-19 $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_746 N_A_809_369#_c_912_n N_A_997_413#_c_1194_n 0.0155265f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_747 N_A_809_369#_c_912_n N_A_997_413#_c_1195_n 0.0118734f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_748 N_A_809_369#_c_912_n N_A_997_413#_c_1196_n 0.0155535f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_749 N_A_809_369#_c_912_n N_A_997_413#_c_1198_n 0.0332506f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_750 N_A_809_369#_M1006_g N_A_997_413#_c_1199_n 0.00957282f $X=8.34 $Y=0.555
+ $X2=0 $Y2=0
cc_751 N_A_809_369#_c_912_n SET_B 7.79765e-19 $X=8.365 $Y=1.19 $X2=0 $Y2=0
cc_752 N_A_809_369#_M1006_g N_SET_B_c_1352_n 0.00162265f $X=8.34 $Y=0.555 $X2=0
+ $Y2=0
cc_753 N_A_809_369#_c_922_n N_SET_B_c_1352_n 0.00252692f $X=8.485 $Y=1.905 $X2=0
+ $Y2=0
cc_754 N_A_809_369#_c_912_n N_SET_B_c_1352_n 0.117877f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_755 N_A_809_369#_c_915_n N_SET_B_c_1352_n 0.0255536f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_756 N_A_809_369#_c_916_n N_SET_B_c_1352_n 0.0151558f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_757 N_A_809_369#_c_912_n N_SET_B_c_1353_n 0.0264108f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_758 N_A_809_369#_c_922_n N_SET_B_c_1354_n 6.80577e-19 $X=8.485 $Y=1.905 $X2=0
+ $Y2=0
cc_759 N_A_809_369#_c_916_n N_SET_B_c_1354_n 0.00255044f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_760 N_A_809_369#_M1006_g N_SET_B_c_1355_n 3.72311e-19 $X=8.34 $Y=0.555 $X2=0
+ $Y2=0
cc_761 N_A_809_369#_c_922_n N_SET_B_c_1355_n 5.60869e-19 $X=8.485 $Y=1.905 $X2=0
+ $Y2=0
cc_762 N_A_809_369#_c_916_n N_SET_B_c_1355_n 0.0123114f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_763 N_A_809_369#_M1040_g N_A_1770_295#_M1011_g 0.0304309f $X=8.485 $Y=2.275
+ $X2=0 $Y2=0
cc_764 N_A_809_369#_M1006_g N_A_1770_295#_c_1496_n 0.00277264f $X=8.34 $Y=0.555
+ $X2=0 $Y2=0
cc_765 N_A_809_369#_c_922_n N_A_1770_295#_c_1496_n 0.0208879f $X=8.485 $Y=1.905
+ $X2=0 $Y2=0
cc_766 N_A_809_369#_c_916_n N_A_1770_295#_c_1496_n 0.00205278f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_767 N_A_809_369#_c_915_n N_A_1770_295#_c_1488_n 0.00116813f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_768 N_A_809_369#_c_916_n N_A_1770_295#_c_1488_n 0.00344735f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_769 N_A_809_369#_c_922_n N_A_1587_329#_c_1615_n 0.00463493f $X=8.485 $Y=1.905
+ $X2=0 $Y2=0
cc_770 N_A_809_369#_M1040_g N_A_1587_329#_c_1615_n 0.0113397f $X=8.485 $Y=2.275
+ $X2=0 $Y2=0
cc_771 N_A_809_369#_c_916_n N_A_1587_329#_c_1615_n 0.0110537f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_772 N_A_809_369#_M1006_g N_A_1587_329#_c_1616_n 0.00763795f $X=8.34 $Y=0.555
+ $X2=0 $Y2=0
cc_773 N_A_809_369#_M1040_g N_A_1587_329#_c_1612_n 0.00469548f $X=8.485 $Y=2.275
+ $X2=0 $Y2=0
cc_774 N_A_809_369#_c_916_n N_A_1587_329#_c_1612_n 7.3132e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_775 N_A_809_369#_c_920_n N_VPWR_c_1863_n 0.00585385f $X=4.91 $Y=1.99 $X2=0
+ $Y2=0
cc_776 N_A_809_369#_c_924_n N_VPWR_c_1863_n 0.00207412f $X=4.91 $Y=1.915 $X2=0
+ $Y2=0
cc_777 N_A_809_369#_c_925_n N_VPWR_c_1863_n 0.023872f $X=4.18 $Y=2.3 $X2=0 $Y2=0
cc_778 N_A_809_369#_M1040_g N_VPWR_c_1867_n 0.00358923f $X=8.485 $Y=2.275 $X2=0
+ $Y2=0
cc_779 N_A_809_369#_M1030_d N_VPWR_c_1851_n 0.00210742f $X=4.045 $Y=1.845 $X2=0
+ $Y2=0
cc_780 N_A_809_369#_c_920_n N_VPWR_c_1851_n 0.00769758f $X=4.91 $Y=1.99 $X2=0
+ $Y2=0
cc_781 N_A_809_369#_M1040_g N_VPWR_c_1851_n 0.00575532f $X=8.485 $Y=2.275 $X2=0
+ $Y2=0
cc_782 N_A_809_369#_c_924_n N_VPWR_c_1851_n 0.00134305f $X=4.91 $Y=1.915 $X2=0
+ $Y2=0
cc_783 N_A_809_369#_c_925_n N_VPWR_c_1851_n 0.00624504f $X=4.18 $Y=2.3 $X2=0
+ $Y2=0
cc_784 N_A_809_369#_M1040_g N_VPWR_c_1875_n 0.0015896f $X=8.485 $Y=2.275 $X2=0
+ $Y2=0
cc_785 N_A_809_369#_c_1049_p N_A_181_47#_c_2056_n 0.0256936f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_786 N_A_809_369#_c_919_n N_A_181_47#_c_2061_n 0.00548737f $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_787 N_A_809_369#_c_909_n N_A_181_47#_c_2061_n 0.0014889f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_788 N_A_809_369#_c_924_n N_A_181_47#_c_2061_n 0.00150693f $X=4.91 $Y=1.915
+ $X2=0 $Y2=0
cc_789 N_A_809_369#_c_926_n N_A_181_47#_c_2061_n 0.00941409f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_790 N_A_809_369#_c_912_n N_A_181_47#_c_2061_n 9.28094e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_791 N_A_809_369#_c_919_n N_A_181_47#_c_2062_n 0.00452993f $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_792 N_A_809_369#_c_920_n N_A_181_47#_c_2062_n 0.00393901f $X=4.91 $Y=1.99
+ $X2=0 $Y2=0
cc_793 N_A_809_369#_c_924_n N_A_181_47#_c_2062_n 0.0126899f $X=4.91 $Y=1.915
+ $X2=0 $Y2=0
cc_794 N_A_809_369#_c_926_n N_A_181_47#_c_2062_n 0.0646535f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_795 N_A_809_369#_c_919_n N_A_181_47#_c_2057_n 6.71081e-19 $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_796 N_A_809_369#_c_909_n N_A_181_47#_c_2057_n 0.00723713f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_797 N_A_809_369#_c_926_n N_A_181_47#_c_2057_n 0.00124944f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_798 N_A_809_369#_c_912_n N_A_181_47#_c_2057_n 0.0120122f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_799 N_A_809_369#_c_913_n N_A_181_47#_c_2057_n 0.00235599f $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_800 N_A_809_369#_c_914_n N_A_181_47#_c_2057_n 0.0217629f $X=4.37 $Y=1.19
+ $X2=0 $Y2=0
cc_801 N_A_809_369#_c_917_n N_A_181_47#_c_2057_n 0.00624074f $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_802 N_A_809_369#_c_918_n N_A_181_47#_c_2057_n 0.00789495f $X=4.327 $Y=1.09
+ $X2=0 $Y2=0
cc_803 N_A_809_369#_M1024_g N_A_181_47#_c_2059_n 8.04362e-19 $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_804 N_A_809_369#_c_912_n N_A_181_47#_c_2059_n 0.00596662f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_805 N_A_809_369#_c_913_n N_A_181_47#_c_2059_n 5.00901e-19 $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_806 N_A_809_369#_c_917_n N_A_181_47#_c_2059_n 0.00349764f $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_807 N_A_809_369#_c_918_n N_A_181_47#_c_2059_n 0.0256936f $X=4.327 $Y=1.09
+ $X2=0 $Y2=0
cc_808 N_A_809_369#_c_919_n N_A_181_47#_c_2064_n 0.0030262f $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_809 N_A_809_369#_c_926_n N_A_181_47#_c_2064_n 0.0163657f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_810 N_A_809_369#_c_912_n N_A_181_47#_c_2064_n 0.013591f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_811 N_A_809_369#_c_913_n N_A_181_47#_c_2064_n 0.0254082f $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_812 N_A_809_369#_c_914_n N_A_181_47#_c_2064_n 0.0014472f $X=4.37 $Y=1.19
+ $X2=0 $Y2=0
cc_813 N_A_809_369#_c_917_n N_A_181_47#_c_2064_n 8.3882e-19 $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_814 N_A_809_369#_c_909_n N_A_181_47#_c_2067_n 4.09059e-19 $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_815 N_A_809_369#_c_924_n N_A_181_47#_c_2067_n 4.12766e-19 $X=4.91 $Y=1.915
+ $X2=0 $Y2=0
cc_816 N_A_809_369#_c_926_n N_A_181_47#_c_2067_n 5.66756e-19 $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_817 N_A_809_369#_c_912_n N_A_181_47#_c_2067_n 0.0264737f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_818 N_A_809_369#_M1006_g N_VGND_c_2256_n 0.00431327f $X=8.34 $Y=0.555 $X2=0
+ $Y2=0
cc_819 N_A_809_369#_M1024_g N_VGND_c_2259_n 0.00592053f $X=5.36 $Y=0.445 $X2=0
+ $Y2=0
cc_820 N_A_809_369#_c_1049_p N_VGND_c_2259_n 0.014833f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_821 N_A_809_369#_M1036_d N_VGND_c_2263_n 0.00330021f $X=4.075 $Y=0.235 $X2=0
+ $Y2=0
cc_822 N_A_809_369#_M1024_g N_VGND_c_2263_n 0.00511765f $X=5.36 $Y=0.445 $X2=0
+ $Y2=0
cc_823 N_A_809_369#_M1006_g N_VGND_c_2263_n 0.00715368f $X=8.34 $Y=0.555 $X2=0
+ $Y2=0
cc_824 N_A_809_369#_c_1049_p N_VGND_c_2263_n 0.0085511f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_825 N_A_809_369#_M1006_g N_VGND_c_2266_n 0.00975709f $X=8.34 $Y=0.555 $X2=0
+ $Y2=0
cc_826 N_A_809_369#_c_912_n N_VGND_c_2266_n 0.0053776f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_827 N_A_1129_21#_c_1092_n N_A_997_413#_c_1188_n 0.00200711f $X=6.275 $Y=0.72
+ $X2=0 $Y2=0
cc_828 N_A_1129_21#_c_1100_n N_A_997_413#_c_1188_n 8.3118e-19 $X=6.55 $Y=2.02
+ $X2=0 $Y2=0
cc_829 N_A_1129_21#_c_1096_n N_A_997_413#_c_1188_n 0.0134492f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_830 N_A_1129_21#_M1037_g N_A_997_413#_M1008_g 0.0129854f $X=5.84 $Y=2.275
+ $X2=0 $Y2=0
cc_831 N_A_1129_21#_c_1098_n N_A_997_413#_M1008_g 0.00226771f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_832 N_A_1129_21#_c_1099_n N_A_997_413#_M1008_g 0.0214214f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_833 N_A_1129_21#_c_1100_n N_A_997_413#_M1008_g 0.01283f $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_834 N_A_1129_21#_c_1096_n N_A_997_413#_M1008_g 0.00590653f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_835 N_A_1129_21#_c_1096_n N_A_997_413#_c_1189_n 6.19699e-19 $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_836 N_A_1129_21#_c_1092_n N_A_997_413#_c_1190_n 0.00174171f $X=6.275 $Y=0.72
+ $X2=0 $Y2=0
cc_837 N_A_1129_21#_M1025_g N_A_997_413#_c_1191_n 9.74282e-19 $X=5.72 $Y=0.445
+ $X2=0 $Y2=0
cc_838 N_A_1129_21#_c_1092_n N_A_997_413#_c_1191_n 0.00951634f $X=6.275 $Y=0.72
+ $X2=0 $Y2=0
cc_839 N_A_1129_21#_c_1094_n N_A_997_413#_c_1191_n 0.00110159f $X=5.792 $Y=0.72
+ $X2=0 $Y2=0
cc_840 N_A_1129_21#_c_1095_n N_A_997_413#_c_1191_n 0.0086776f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_841 N_A_1129_21#_M1025_g N_A_997_413#_c_1192_n 0.00116003f $X=5.72 $Y=0.445
+ $X2=0 $Y2=0
cc_842 N_A_1129_21#_c_1094_n N_A_997_413#_c_1192_n 0.0307762f $X=5.792 $Y=0.72
+ $X2=0 $Y2=0
cc_843 N_A_1129_21#_c_1095_n N_A_997_413#_c_1192_n 0.00118264f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_844 N_A_1129_21#_c_1096_n N_A_997_413#_c_1192_n 0.00259391f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_845 N_A_1129_21#_c_1098_n N_A_997_413#_c_1203_n 0.0251699f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_846 N_A_1129_21#_c_1101_n N_A_997_413#_c_1203_n 0.010676f $X=6.095 $Y=2.02
+ $X2=0 $Y2=0
cc_847 N_A_1129_21#_c_1096_n N_A_997_413#_c_1203_n 0.0119128f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_848 N_A_1129_21#_c_1094_n N_A_997_413#_c_1193_n 0.00784248f $X=5.792 $Y=0.72
+ $X2=0 $Y2=0
cc_849 N_A_1129_21#_c_1095_n N_A_997_413#_c_1193_n 0.00297153f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_850 N_A_1129_21#_c_1098_n N_A_997_413#_c_1194_n 0.0109804f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_851 N_A_1129_21#_c_1099_n N_A_997_413#_c_1194_n 0.00260846f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_852 N_A_1129_21#_c_1092_n N_A_997_413#_c_1194_n 0.00671458f $X=6.275 $Y=0.72
+ $X2=0 $Y2=0
cc_853 N_A_1129_21#_c_1100_n N_A_997_413#_c_1194_n 0.00617396f $X=6.55 $Y=2.02
+ $X2=0 $Y2=0
cc_854 N_A_1129_21#_c_1094_n N_A_997_413#_c_1194_n 0.0109475f $X=5.792 $Y=0.72
+ $X2=0 $Y2=0
cc_855 N_A_1129_21#_c_1095_n N_A_997_413#_c_1194_n 7.94205e-19 $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_856 N_A_1129_21#_c_1096_n N_A_997_413#_c_1194_n 0.0126776f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_857 N_A_1129_21#_c_1092_n N_A_997_413#_c_1195_n 0.0218346f $X=6.275 $Y=0.72
+ $X2=0 $Y2=0
cc_858 N_A_1129_21#_c_1094_n N_A_997_413#_c_1195_n 0.00231435f $X=5.792 $Y=0.72
+ $X2=0 $Y2=0
cc_859 N_A_1129_21#_c_1095_n N_A_997_413#_c_1195_n 0.00162316f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_860 N_A_1129_21#_c_1096_n N_A_997_413#_c_1195_n 0.00183382f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_861 N_A_1129_21#_c_1100_n N_A_997_413#_c_1198_n 0.00266207f $X=6.55 $Y=2.02
+ $X2=0 $Y2=0
cc_862 N_A_1129_21#_c_1100_n N_SET_B_M1032_g 0.00492702f $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_863 N_A_1129_21#_c_1098_n SET_B 0.0050279f $X=6.01 $Y=1.74 $X2=0 $Y2=0
cc_864 N_A_1129_21#_c_1100_n SET_B 0.00846821f $X=6.55 $Y=2.02 $X2=0 $Y2=0
cc_865 N_A_1129_21#_c_1098_n N_SET_B_c_1353_n 0.00168225f $X=6.01 $Y=1.74 $X2=0
+ $Y2=0
cc_866 N_A_1129_21#_c_1100_n N_SET_B_c_1353_n 2.95185e-19 $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_867 N_A_1129_21#_c_1100_n N_SET_B_c_1356_n 9.77119e-19 $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_868 N_A_1129_21#_c_1100_n N_VPWR_M1037_d 0.00228817f $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_869 N_A_1129_21#_c_1101_n N_VPWR_M1037_d 0.00142005f $X=6.095 $Y=2.02 $X2=0
+ $Y2=0
cc_870 N_A_1129_21#_M1037_g N_VPWR_c_1855_n 0.00324191f $X=5.84 $Y=2.275 $X2=0
+ $Y2=0
cc_871 N_A_1129_21#_c_1099_n N_VPWR_c_1855_n 7.77116e-19 $X=6.01 $Y=1.74 $X2=0
+ $Y2=0
cc_872 N_A_1129_21#_c_1100_n N_VPWR_c_1855_n 0.0125888f $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_873 N_A_1129_21#_c_1101_n N_VPWR_c_1855_n 0.00947355f $X=6.095 $Y=2.02 $X2=0
+ $Y2=0
cc_874 N_A_1129_21#_M1037_g N_VPWR_c_1863_n 0.00585385f $X=5.84 $Y=2.275 $X2=0
+ $Y2=0
cc_875 N_A_1129_21#_M1008_d N_VPWR_c_1851_n 0.00271411f $X=6.505 $Y=2.065 $X2=0
+ $Y2=0
cc_876 N_A_1129_21#_M1037_g N_VPWR_c_1851_n 0.0068485f $X=5.84 $Y=2.275 $X2=0
+ $Y2=0
cc_877 N_A_1129_21#_c_1100_n N_VPWR_c_1851_n 0.0035918f $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_878 N_A_1129_21#_c_1101_n N_VPWR_c_1851_n 7.82982e-19 $X=6.095 $Y=2.02 $X2=0
+ $Y2=0
cc_879 N_A_1129_21#_c_1171_p N_VPWR_c_1851_n 0.00381852f $X=6.66 $Y=2.285 $X2=0
+ $Y2=0
cc_880 N_A_1129_21#_c_1100_n N_VPWR_c_1874_n 0.00402862f $X=6.55 $Y=2.02 $X2=0
+ $Y2=0
cc_881 N_A_1129_21#_c_1171_p N_VPWR_c_1874_n 0.0130575f $X=6.66 $Y=2.285 $X2=0
+ $Y2=0
cc_882 N_A_1129_21#_c_1092_n N_VGND_M1025_d 8.64202e-19 $X=6.275 $Y=0.72 $X2=0
+ $Y2=0
cc_883 N_A_1129_21#_c_1094_n N_VGND_M1025_d 0.00132848f $X=5.792 $Y=0.72 $X2=0
+ $Y2=0
cc_884 N_A_1129_21#_M1025_g N_VGND_c_2259_n 0.0133423f $X=5.72 $Y=0.445 $X2=0
+ $Y2=0
cc_885 N_A_1129_21#_c_1092_n N_VGND_c_2259_n 0.00919218f $X=6.275 $Y=0.72 $X2=0
+ $Y2=0
cc_886 N_A_1129_21#_c_1093_n N_VGND_c_2259_n 0.0170013f $X=6.45 $Y=0.51 $X2=0
+ $Y2=0
cc_887 N_A_1129_21#_c_1094_n N_VGND_c_2259_n 0.0212099f $X=5.792 $Y=0.72 $X2=0
+ $Y2=0
cc_888 N_A_1129_21#_c_1095_n N_VGND_c_2259_n 8.18098e-19 $X=5.81 $Y=0.93 $X2=0
+ $Y2=0
cc_889 N_A_1129_21#_M1009_s N_VGND_c_2263_n 0.00268769f $X=6.325 $Y=0.235 $X2=0
+ $Y2=0
cc_890 N_A_1129_21#_c_1092_n N_VGND_c_2263_n 0.00566344f $X=6.275 $Y=0.72 $X2=0
+ $Y2=0
cc_891 N_A_1129_21#_c_1093_n N_VGND_c_2263_n 0.00988152f $X=6.45 $Y=0.51 $X2=0
+ $Y2=0
cc_892 N_A_1129_21#_c_1094_n N_VGND_c_2263_n 0.00167167f $X=5.792 $Y=0.72 $X2=0
+ $Y2=0
cc_893 N_A_1129_21#_c_1092_n N_VGND_c_2265_n 0.00328118f $X=6.275 $Y=0.72 $X2=0
+ $Y2=0
cc_894 N_A_1129_21#_c_1093_n N_VGND_c_2265_n 0.0177262f $X=6.45 $Y=0.51 $X2=0
+ $Y2=0
cc_895 N_A_1129_21#_c_1092_n N_VGND_c_2266_n 0.0118971f $X=6.275 $Y=0.72 $X2=0
+ $Y2=0
cc_896 N_A_997_413#_M1008_g N_SET_B_M1032_g 0.0141406f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_897 N_A_997_413#_c_1189_n N_SET_B_M1041_g 0.00918774f $X=6.44 $Y=1.095 $X2=0
+ $Y2=0
cc_898 N_A_997_413#_c_1190_n N_SET_B_M1041_g 0.0503585f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_899 N_A_997_413#_c_1197_n N_SET_B_M1041_g 0.0211491f $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_900 N_A_997_413#_c_1198_n N_SET_B_M1041_g 0.0114968f $X=7.3 $Y=1.15 $X2=0
+ $Y2=0
cc_901 N_A_997_413#_c_1199_n N_SET_B_M1041_g 0.0223839f $X=7.44 $Y=0.995 $X2=0
+ $Y2=0
cc_902 N_A_997_413#_c_1188_n N_SET_B_c_1342_n 0.00844505f $X=6.43 $Y=1.365 $X2=0
+ $Y2=0
cc_903 N_A_997_413#_M1016_g N_SET_B_c_1342_n 0.00182806f $X=7.495 $Y=2.065 $X2=0
+ $Y2=0
cc_904 N_A_997_413#_c_1195_n N_SET_B_c_1342_n 6.38923e-19 $X=6.435 $Y=1.185
+ $X2=0 $Y2=0
cc_905 N_A_997_413#_c_1196_n N_SET_B_c_1342_n 0.0011077f $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_906 N_A_997_413#_c_1198_n N_SET_B_c_1342_n 0.00810141f $X=7.3 $Y=1.15 $X2=0
+ $Y2=0
cc_907 N_A_997_413#_M1008_g SET_B 0.0043986f $X=6.43 $Y=2.275 $X2=0 $Y2=0
cc_908 N_A_997_413#_M1016_g SET_B 0.00130013f $X=7.495 $Y=2.065 $X2=0 $Y2=0
cc_909 N_A_997_413#_c_1198_n SET_B 0.0245396f $X=7.3 $Y=1.15 $X2=0 $Y2=0
cc_910 N_A_997_413#_M1016_g N_SET_B_c_1352_n 0.00137751f $X=7.495 $Y=2.065 $X2=0
+ $Y2=0
cc_911 N_A_997_413#_c_1196_n N_SET_B_c_1352_n 0.00232559f $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_912 N_A_997_413#_c_1197_n N_SET_B_c_1352_n 0.00186621f $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_913 N_A_997_413#_c_1198_n N_SET_B_c_1352_n 0.00598577f $X=7.3 $Y=1.15 $X2=0
+ $Y2=0
cc_914 N_A_997_413#_M1008_g N_SET_B_c_1353_n 0.00435388f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_915 N_A_997_413#_c_1198_n N_SET_B_c_1353_n 0.00230051f $X=7.3 $Y=1.15 $X2=0
+ $Y2=0
cc_916 N_A_997_413#_M1008_g N_SET_B_c_1356_n 0.0201157f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_917 N_A_997_413#_c_1191_n N_SET_B_c_1356_n 2.44193e-19 $X=6.66 $Y=0.805 $X2=0
+ $Y2=0
cc_918 N_A_997_413#_c_1198_n N_SET_B_c_1356_n 7.14223e-19 $X=7.3 $Y=1.15 $X2=0
+ $Y2=0
cc_919 N_A_997_413#_M1008_g N_SET_B_c_1357_n 0.00297195f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_920 N_A_997_413#_M1016_g N_SET_B_c_1357_n 0.0291182f $X=7.495 $Y=2.065 $X2=0
+ $Y2=0
cc_921 N_A_997_413#_M1008_g N_VPWR_c_1855_n 0.00571865f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_922 N_A_997_413#_c_1216_n N_VPWR_c_1863_n 0.0428204f $X=5.585 $Y=2.3 $X2=0
+ $Y2=0
cc_923 N_A_997_413#_M1007_d N_VPWR_c_1851_n 0.00208736f $X=4.985 $Y=2.065 $X2=0
+ $Y2=0
cc_924 N_A_997_413#_M1008_g N_VPWR_c_1851_n 0.00610863f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_925 N_A_997_413#_c_1216_n N_VPWR_c_1851_n 0.0123083f $X=5.585 $Y=2.3 $X2=0
+ $Y2=0
cc_926 N_A_997_413#_M1008_g N_VPWR_c_1874_n 0.00422112f $X=6.43 $Y=2.275 $X2=0
+ $Y2=0
cc_927 N_A_997_413#_M1016_g N_VPWR_c_1875_n 0.0235413f $X=7.495 $Y=2.065 $X2=0
+ $Y2=0
cc_928 N_A_997_413#_c_1192_n N_A_181_47#_c_2056_n 0.0591375f $X=5.15 $Y=0.42
+ $X2=0 $Y2=0
cc_929 N_A_997_413#_c_1203_n N_A_181_47#_c_2061_n 0.00197049f $X=5.67 $Y=2.135
+ $X2=0 $Y2=0
cc_930 N_A_997_413#_c_1193_n N_A_181_47#_c_2057_n 0.0111326f $X=5.755 $Y=1.31
+ $X2=0 $Y2=0
cc_931 N_A_997_413#_c_1203_n N_A_181_47#_c_2067_n 0.00424021f $X=5.67 $Y=2.135
+ $X2=0 $Y2=0
cc_932 N_A_997_413#_c_1216_n A_1081_413# 0.0063224f $X=5.585 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_933 N_A_997_413#_c_1203_n A_1081_413# 0.0012628f $X=5.67 $Y=2.135 $X2=-0.19
+ $Y2=-0.24
cc_934 N_A_997_413#_c_1190_n N_VGND_c_2259_n 0.00201292f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_935 N_A_997_413#_c_1192_n N_VGND_c_2259_n 0.0262729f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_936 N_A_997_413#_M1023_d N_VGND_c_2263_n 0.00215201f $X=5.015 $Y=0.235 $X2=0
+ $Y2=0
cc_937 N_A_997_413#_c_1190_n N_VGND_c_2263_n 0.011139f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_938 N_A_997_413#_c_1191_n N_VGND_c_2263_n 0.00109181f $X=6.66 $Y=0.805 $X2=0
+ $Y2=0
cc_939 N_A_997_413#_c_1192_n N_VGND_c_2263_n 0.0159733f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_940 N_A_997_413#_c_1190_n N_VGND_c_2265_n 0.00583607f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_941 N_A_997_413#_c_1191_n N_VGND_c_2265_n 0.001207f $X=6.66 $Y=0.805 $X2=0
+ $Y2=0
cc_942 N_A_997_413#_c_1190_n N_VGND_c_2266_n 0.00692823f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_943 N_A_997_413#_c_1197_n N_VGND_c_2266_n 6.94553e-19 $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_944 N_A_997_413#_c_1198_n N_VGND_c_2266_n 0.0658132f $X=7.3 $Y=1.15 $X2=0
+ $Y2=0
cc_945 N_A_997_413#_c_1199_n N_VGND_c_2266_n 0.0277551f $X=7.44 $Y=0.995 $X2=0
+ $Y2=0
cc_946 N_SET_B_c_1347_n N_A_1770_295#_M1011_g 0.013067f $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_947 N_SET_B_c_1349_n N_A_1770_295#_M1011_g 6.24257e-19 $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_948 N_SET_B_c_1354_n N_A_1770_295#_M1011_g 3.69011e-19 $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_949 N_SET_B_c_1355_n N_A_1770_295#_M1011_g 0.00496572f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_950 N_SET_B_c_1349_n N_A_1770_295#_c_1495_n 0.0171616f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_951 N_SET_B_c_1350_n N_A_1770_295#_c_1495_n 0.00313671f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_952 N_SET_B_c_1354_n N_A_1770_295#_c_1495_n 0.00212943f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_953 N_SET_B_c_1355_n N_A_1770_295#_c_1495_n 0.00562733f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_954 N_SET_B_c_1354_n N_A_1770_295#_c_1496_n 0.00102336f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_955 N_SET_B_c_1355_n N_A_1770_295#_c_1496_n 0.00260561f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_956 N_SET_B_M1010_g N_A_1770_295#_M1018_g 0.0139533f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_957 N_SET_B_M1010_g N_A_1770_295#_c_1488_n 0.00611735f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_958 N_SET_B_c_1348_n N_A_1770_295#_c_1488_n 0.00313671f $X=9.9 $Y=1.58 $X2=0
+ $Y2=0
cc_959 N_SET_B_c_1354_n N_A_1770_295#_c_1488_n 0.00151827f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_960 N_SET_B_c_1355_n N_A_1770_295#_c_1488_n 0.00193706f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_961 N_SET_B_M1010_g N_A_1770_295#_c_1489_n 0.00105364f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_962 N_SET_B_M1010_g N_A_1770_295#_c_1490_n 0.0105912f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_963 N_SET_B_c_1347_n N_A_1770_295#_c_1490_n 2.21899e-19 $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_964 N_SET_B_c_1349_n N_A_1770_295#_c_1490_n 3.26955e-19 $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_965 N_SET_B_M1010_g N_A_1770_295#_c_1491_n 0.0109021f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_966 N_SET_B_c_1348_n N_A_1770_295#_c_1491_n 0.00327249f $X=9.9 $Y=1.58 $X2=0
+ $Y2=0
cc_967 N_SET_B_c_1349_n N_A_1770_295#_c_1491_n 0.0448652f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1349_n N_A_1770_295#_c_1499_n 0.0137214f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_969 N_SET_B_M1010_g N_A_1770_295#_c_1492_n 4.78445e-19 $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_970 N_SET_B_c_1347_n N_A_1587_329#_M1038_g 0.00304082f $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_971 N_SET_B_c_1350_n N_A_1587_329#_c_1604_n 0.0246322f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_972 N_SET_B_c_1352_n N_A_1587_329#_c_1615_n 0.0145826f $X=8.825 $Y=1.53 $X2=0
+ $Y2=0
cc_973 N_SET_B_M1010_g N_A_1587_329#_c_1616_n 0.002505f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_974 N_SET_B_c_1344_n N_A_1587_329#_c_1607_n 0.00755042f $X=9.57 $Y=1.985
+ $X2=0 $Y2=0
cc_975 N_SET_B_c_1347_n N_A_1587_329#_c_1607_n 0.00535795f $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1349_n N_A_1587_329#_c_1607_n 0.0437797f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_977 N_SET_B_c_1354_n N_A_1587_329#_c_1607_n 0.00107633f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_978 N_SET_B_c_1355_n N_A_1587_329#_c_1607_n 0.012295f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_979 N_SET_B_M1010_g N_A_1587_329#_c_1594_n 0.0090884f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_980 N_SET_B_M1010_g N_A_1587_329#_c_1596_n 0.0114527f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_981 N_SET_B_M1010_g N_A_1587_329#_c_1597_n 0.0246322f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_982 N_SET_B_c_1347_n N_A_1587_329#_c_1610_n 0.00607875f $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1349_n N_A_1587_329#_c_1610_n 0.0115956f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_984 N_SET_B_c_1347_n N_A_1587_329#_c_1643_n 4.48138e-19 $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_985 N_SET_B_c_1348_n N_A_1587_329#_c_1643_n 2.28373e-19 $X=9.9 $Y=1.58 $X2=0
+ $Y2=0
cc_986 N_SET_B_c_1349_n N_A_1587_329#_c_1643_n 0.0162126f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_987 N_SET_B_c_1350_n N_A_1587_329#_c_1643_n 0.0010808f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_988 N_SET_B_c_1348_n N_A_1587_329#_c_1611_n 0.0246322f $X=9.9 $Y=1.58 $X2=0
+ $Y2=0
cc_989 N_SET_B_c_1349_n N_A_1587_329#_c_1611_n 0.00121532f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_990 N_SET_B_c_1344_n N_A_1587_329#_c_1612_n 6.37057e-19 $X=9.57 $Y=1.985
+ $X2=0 $Y2=0
cc_991 N_SET_B_c_1352_n N_A_1587_329#_c_1612_n 0.00244169f $X=8.825 $Y=1.53
+ $X2=0 $Y2=0
cc_992 N_SET_B_c_1354_n N_A_1587_329#_c_1612_n 0.00212299f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_993 N_SET_B_c_1355_n N_A_1587_329#_c_1612_n 0.00347269f $X=8.97 $Y=1.53 $X2=0
+ $Y2=0
cc_994 N_SET_B_c_1347_n N_A_1587_329#_c_1653_n 0.00907673f $X=9.9 $Y=1.835 $X2=0
+ $Y2=0
cc_995 N_SET_B_c_1349_n N_A_1587_329#_c_1653_n 0.0165572f $X=9.9 $Y=1.61 $X2=0
+ $Y2=0
cc_996 N_SET_B_M1010_g N_A_1587_329#_c_1598_n 0.0135558f $X=9.96 $Y=0.445 $X2=0
+ $Y2=0
cc_997 N_SET_B_c_1344_n N_VPWR_c_1856_n 0.00777846f $X=9.57 $Y=1.985 $X2=0 $Y2=0
cc_998 N_SET_B_c_1344_n N_VPWR_c_1857_n 0.0019106f $X=9.57 $Y=1.985 $X2=0 $Y2=0
cc_999 N_SET_B_c_1344_n N_VPWR_c_1868_n 0.00341689f $X=9.57 $Y=1.985 $X2=0 $Y2=0
cc_1000 N_SET_B_c_1347_n N_VPWR_c_1868_n 0.00111314f $X=9.9 $Y=1.835 $X2=0 $Y2=0
cc_1001 N_SET_B_M1032_g N_VPWR_c_1851_n 0.00671739f $X=6.915 $Y=2.275 $X2=0
+ $Y2=0
cc_1002 N_SET_B_c_1344_n N_VPWR_c_1851_n 0.00538978f $X=9.57 $Y=1.985 $X2=0
+ $Y2=0
cc_1003 N_SET_B_c_1356_n N_VPWR_c_1851_n 4.0446e-19 $X=6.85 $Y=1.68 $X2=0 $Y2=0
cc_1004 N_SET_B_M1032_g N_VPWR_c_1874_n 0.00585385f $X=6.915 $Y=2.275 $X2=0
+ $Y2=0
cc_1005 N_SET_B_M1032_g N_VPWR_c_1875_n 0.00385005f $X=6.915 $Y=2.275 $X2=0
+ $Y2=0
cc_1006 N_SET_B_c_1352_n N_VPWR_c_1875_n 0.00101216f $X=8.825 $Y=1.53 $X2=0
+ $Y2=0
cc_1007 N_SET_B_M1010_g N_VGND_c_2249_n 0.00545251f $X=9.96 $Y=0.445 $X2=0 $Y2=0
cc_1008 N_SET_B_M1010_g N_VGND_c_2256_n 0.00585385f $X=9.96 $Y=0.445 $X2=0 $Y2=0
cc_1009 N_SET_B_M1010_g N_VGND_c_2263_n 0.0072274f $X=9.96 $Y=0.445 $X2=0 $Y2=0
cc_1010 N_SET_B_M1041_g N_VGND_c_2266_n 0.0259455f $X=7.02 $Y=0.445 $X2=0 $Y2=0
cc_1011 N_SET_B_c_1342_n N_VGND_c_2266_n 4.81194e-19 $X=7.02 $Y=1.29 $X2=0 $Y2=0
cc_1012 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1588_n 0.0017596f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1013 N_A_1770_295#_c_1492_n N_A_1587_329#_c_1588_n 0.0160404f $X=10.805
+ $Y=1.185 $X2=0 $Y2=0
cc_1014 N_A_1770_295#_c_1493_n N_A_1587_329#_c_1588_n 0.00116113f $X=10.805
+ $Y=0.397 $X2=0 $Y2=0
cc_1015 N_A_1770_295#_c_1501_n N_A_1587_329#_c_1588_n 0.0149226f $X=10.765
+ $Y=1.27 $X2=0 $Y2=0
cc_1016 N_A_1770_295#_c_1492_n N_A_1587_329#_c_1589_n 0.00230329f $X=10.805
+ $Y=1.185 $X2=0 $Y2=0
cc_1017 N_A_1770_295#_c_1500_n N_A_1587_329#_M1029_g 0.00383768f $X=10.72
+ $Y=2.285 $X2=0 $Y2=0
cc_1018 N_A_1770_295#_c_1501_n N_A_1587_329#_M1029_g 5.11687e-19 $X=10.765
+ $Y=1.27 $X2=0 $Y2=0
cc_1019 N_A_1770_295#_M1011_g N_A_1587_329#_c_1615_n 5.40489e-19 $X=8.925
+ $Y=2.275 $X2=0 $Y2=0
cc_1020 N_A_1770_295#_M1018_g N_A_1587_329#_c_1616_n 0.0123541f $X=9.32 $Y=0.445
+ $X2=0 $Y2=0
cc_1021 N_A_1770_295#_c_1489_n N_A_1587_329#_c_1616_n 0.00443217f $X=9.38
+ $Y=1.02 $X2=0 $Y2=0
cc_1022 N_A_1770_295#_c_1490_n N_A_1587_329#_c_1616_n 0.00170909f $X=9.38
+ $Y=1.02 $X2=0 $Y2=0
cc_1023 N_A_1770_295#_M1011_g N_A_1587_329#_c_1607_n 0.00683237f $X=8.925
+ $Y=2.275 $X2=0 $Y2=0
cc_1024 N_A_1770_295#_c_1495_n N_A_1587_329#_c_1607_n 0.00214711f $X=9.245
+ $Y=1.55 $X2=0 $Y2=0
cc_1025 N_A_1770_295#_M1018_g N_A_1587_329#_c_1594_n 0.00659402f $X=9.32
+ $Y=0.445 $X2=0 $Y2=0
cc_1026 N_A_1770_295#_c_1489_n N_A_1587_329#_c_1595_n 0.0118984f $X=9.38 $Y=1.02
+ $X2=0 $Y2=0
cc_1027 N_A_1770_295#_c_1490_n N_A_1587_329#_c_1595_n 0.00140267f $X=9.38
+ $Y=1.02 $X2=0 $Y2=0
cc_1028 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1595_n 0.0143582f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1029 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1596_n 0.0507947f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1030 N_A_1770_295#_c_1492_n N_A_1587_329#_c_1596_n 0.013409f $X=10.805
+ $Y=1.185 $X2=0 $Y2=0
cc_1031 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1597_n 0.0113963f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1032 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1610_n 0.00572977f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1033 N_A_1770_295#_c_1500_n N_A_1587_329#_c_1610_n 0.0139716f $X=10.72
+ $Y=2.285 $X2=0 $Y2=0
cc_1034 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1643_n 0.0162897f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1035 N_A_1770_295#_c_1500_n N_A_1587_329#_c_1643_n 0.027789f $X=10.72
+ $Y=2.285 $X2=0 $Y2=0
cc_1036 N_A_1770_295#_c_1491_n N_A_1587_329#_c_1611_n 0.0100451f $X=10.635
+ $Y=1.27 $X2=0 $Y2=0
cc_1037 N_A_1770_295#_c_1500_n N_A_1587_329#_c_1611_n 0.0215199f $X=10.72
+ $Y=2.285 $X2=0 $Y2=0
cc_1038 N_A_1770_295#_M1011_g N_A_1587_329#_c_1612_n 0.0152398f $X=8.925
+ $Y=2.275 $X2=0 $Y2=0
cc_1039 N_A_1770_295#_c_1492_n N_A_1587_329#_c_1598_n 0.0135137f $X=10.805
+ $Y=1.185 $X2=0 $Y2=0
cc_1040 N_A_1770_295#_c_1493_n N_A_1587_329#_c_1598_n 0.00407946f $X=10.805
+ $Y=0.397 $X2=0 $Y2=0
cc_1041 N_A_1770_295#_M1011_g N_VPWR_c_1856_n 0.00493655f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_1042 N_A_1770_295#_c_1500_n N_VPWR_c_1858_n 0.0622166f $X=10.72 $Y=2.285
+ $X2=0 $Y2=0
cc_1043 N_A_1770_295#_M1011_g N_VPWR_c_1867_n 0.00390259f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_1044 N_A_1770_295#_c_1500_n N_VPWR_c_1869_n 0.018001f $X=10.72 $Y=2.285 $X2=0
+ $Y2=0
cc_1045 N_A_1770_295#_M1038_d N_VPWR_c_1851_n 0.00382897f $X=10.585 $Y=2.065
+ $X2=0 $Y2=0
cc_1046 N_A_1770_295#_M1011_g N_VPWR_c_1851_n 0.00612329f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_1047 N_A_1770_295#_c_1500_n N_VPWR_c_1851_n 0.00993603f $X=10.72 $Y=2.285
+ $X2=0 $Y2=0
cc_1048 N_A_1770_295#_c_1500_n N_Q_N_c_2204_n 0.00384388f $X=10.72 $Y=2.285
+ $X2=0 $Y2=0
cc_1049 N_A_1770_295#_c_1492_n N_Q_N_c_2204_n 0.00790731f $X=10.805 $Y=1.185
+ $X2=0 $Y2=0
cc_1050 N_A_1770_295#_c_1501_n N_Q_N_c_2204_n 0.00485259f $X=10.765 $Y=1.27
+ $X2=0 $Y2=0
cc_1051 N_A_1770_295#_c_1492_n N_VGND_c_2250_n 0.0212846f $X=10.805 $Y=1.185
+ $X2=0 $Y2=0
cc_1052 N_A_1770_295#_c_1493_n N_VGND_c_2250_n 0.0183991f $X=10.805 $Y=0.397
+ $X2=0 $Y2=0
cc_1053 N_A_1770_295#_M1018_g N_VGND_c_2256_n 0.00362032f $X=9.32 $Y=0.445 $X2=0
+ $Y2=0
cc_1054 N_A_1770_295#_c_1493_n N_VGND_c_2260_n 0.0202265f $X=10.805 $Y=0.397
+ $X2=0 $Y2=0
cc_1055 N_A_1770_295#_M1020_d N_VGND_c_2263_n 0.00209344f $X=10.59 $Y=0.235
+ $X2=0 $Y2=0
cc_1056 N_A_1770_295#_M1018_g N_VGND_c_2263_n 0.00562894f $X=9.32 $Y=0.445 $X2=0
+ $Y2=0
cc_1057 N_A_1770_295#_c_1493_n N_VGND_c_2263_n 0.0124125f $X=10.805 $Y=0.397
+ $X2=0 $Y2=0
cc_1058 N_A_1587_329#_M1027_g N_A_2412_47#_M1003_g 0.0209953f $X=12.395 $Y=2.095
+ $X2=0 $Y2=0
cc_1059 N_A_1587_329#_c_1589_n N_A_2412_47#_c_1756_n 0.00140651f $X=11.455
+ $Y=0.995 $X2=0 $Y2=0
cc_1060 N_A_1587_329#_M1033_g N_A_2412_47#_c_1756_n 0.0111765f $X=12.395
+ $Y=0.445 $X2=0 $Y2=0
cc_1061 N_A_1587_329#_M1029_g N_A_2412_47#_c_1761_n 0.00214796f $X=11.455
+ $Y=1.985 $X2=0 $Y2=0
cc_1062 N_A_1587_329#_M1027_g N_A_2412_47#_c_1761_n 0.0150771f $X=12.395
+ $Y=2.095 $X2=0 $Y2=0
cc_1063 N_A_1587_329#_c_1590_n N_A_2412_47#_c_1757_n 0.00606691f $X=12.32
+ $Y=1.16 $X2=0 $Y2=0
cc_1064 N_A_1587_329#_c_1593_n N_A_2412_47#_c_1757_n 0.0219697f $X=12.395
+ $Y=1.16 $X2=0 $Y2=0
cc_1065 N_A_1587_329#_c_1593_n N_A_2412_47#_c_1758_n 0.0214963f $X=12.395
+ $Y=1.16 $X2=0 $Y2=0
cc_1066 N_A_1587_329#_c_1590_n N_A_2412_47#_c_1772_n 0.0205144f $X=12.32 $Y=1.16
+ $X2=0 $Y2=0
cc_1067 N_A_1587_329#_M1033_g N_A_2412_47#_c_1759_n 0.0174217f $X=12.395
+ $Y=0.445 $X2=0 $Y2=0
cc_1068 N_A_1587_329#_c_1610_n N_VPWR_M1038_s 0.00200513f $X=10.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1069 N_A_1587_329#_c_1607_n N_VPWR_c_1856_n 0.0228646f $X=9.695 $Y=1.98 $X2=0
+ $Y2=0
cc_1070 N_A_1587_329#_c_1612_n N_VPWR_c_1856_n 0.0120282f $X=8.85 $Y=1.98 $X2=0
+ $Y2=0
cc_1071 N_A_1587_329#_M1038_g N_VPWR_c_1857_n 0.00845001f $X=10.51 $Y=2.275
+ $X2=0 $Y2=0
cc_1072 N_A_1587_329#_c_1604_n N_VPWR_c_1857_n 8.1628e-19 $X=10.415 $Y=1.875
+ $X2=0 $Y2=0
cc_1073 N_A_1587_329#_c_1608_n N_VPWR_c_1857_n 0.0142545f $X=9.78 $Y=2.285 $X2=0
+ $Y2=0
cc_1074 N_A_1587_329#_c_1610_n N_VPWR_c_1857_n 0.024109f $X=10.245 $Y=1.98 $X2=0
+ $Y2=0
cc_1075 N_A_1587_329#_M1038_g N_VPWR_c_1858_n 0.00283108f $X=10.51 $Y=2.275
+ $X2=0 $Y2=0
cc_1076 N_A_1587_329#_c_1588_n N_VPWR_c_1858_n 0.00502715f $X=11.38 $Y=1.16
+ $X2=0 $Y2=0
cc_1077 N_A_1587_329#_M1029_g N_VPWR_c_1858_n 0.00444548f $X=11.455 $Y=1.985
+ $X2=0 $Y2=0
cc_1078 N_A_1587_329#_M1029_g N_VPWR_c_1859_n 0.00541359f $X=11.455 $Y=1.985
+ $X2=0 $Y2=0
cc_1079 N_A_1587_329#_M1027_g N_VPWR_c_1859_n 0.00585385f $X=12.395 $Y=2.095
+ $X2=0 $Y2=0
cc_1080 N_A_1587_329#_M1027_g N_VPWR_c_1860_n 0.00774293f $X=12.395 $Y=2.095
+ $X2=0 $Y2=0
cc_1081 N_A_1587_329#_c_1615_n N_VPWR_c_1867_n 0.0371085f $X=8.765 $Y=2.292
+ $X2=0 $Y2=0
cc_1082 N_A_1587_329#_c_1607_n N_VPWR_c_1867_n 0.00442379f $X=9.695 $Y=1.98
+ $X2=0 $Y2=0
cc_1083 N_A_1587_329#_c_1612_n N_VPWR_c_1867_n 0.00925064f $X=8.85 $Y=1.98 $X2=0
+ $Y2=0
cc_1084 N_A_1587_329#_c_1607_n N_VPWR_c_1868_n 0.00273399f $X=9.695 $Y=1.98
+ $X2=0 $Y2=0
cc_1085 N_A_1587_329#_c_1608_n N_VPWR_c_1868_n 0.0132839f $X=9.78 $Y=2.285 $X2=0
+ $Y2=0
cc_1086 N_A_1587_329#_c_1610_n N_VPWR_c_1868_n 0.00392551f $X=10.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1087 N_A_1587_329#_M1038_g N_VPWR_c_1869_n 0.0046653f $X=10.51 $Y=2.275 $X2=0
+ $Y2=0
cc_1088 N_A_1587_329#_M1017_d N_VPWR_c_1851_n 0.00817954f $X=7.935 $Y=1.645
+ $X2=0 $Y2=0
cc_1089 N_A_1587_329#_M1028_d N_VPWR_c_1851_n 0.00228252f $X=9.645 $Y=2.065
+ $X2=0 $Y2=0
cc_1090 N_A_1587_329#_M1038_g N_VPWR_c_1851_n 0.00929867f $X=10.51 $Y=2.275
+ $X2=0 $Y2=0
cc_1091 N_A_1587_329#_M1029_g N_VPWR_c_1851_n 0.0121537f $X=11.455 $Y=1.985
+ $X2=0 $Y2=0
cc_1092 N_A_1587_329#_M1027_g N_VPWR_c_1851_n 0.0123514f $X=12.395 $Y=2.095
+ $X2=0 $Y2=0
cc_1093 N_A_1587_329#_c_1615_n N_VPWR_c_1851_n 0.0231897f $X=8.765 $Y=2.292
+ $X2=0 $Y2=0
cc_1094 N_A_1587_329#_c_1607_n N_VPWR_c_1851_n 0.0124932f $X=9.695 $Y=1.98 $X2=0
+ $Y2=0
cc_1095 N_A_1587_329#_c_1608_n N_VPWR_c_1851_n 0.00809922f $X=9.78 $Y=2.285
+ $X2=0 $Y2=0
cc_1096 N_A_1587_329#_c_1610_n N_VPWR_c_1851_n 0.00780649f $X=10.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1097 N_A_1587_329#_c_1612_n N_VPWR_c_1851_n 0.00603799f $X=8.85 $Y=1.98 $X2=0
+ $Y2=0
cc_1098 N_A_1587_329#_c_1615_n A_1712_413# 0.00493444f $X=8.765 $Y=2.292
+ $X2=-0.19 $Y2=-0.24
cc_1099 N_A_1587_329#_c_1612_n A_1712_413# 0.00180472f $X=8.85 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_1100 N_A_1587_329#_c_1589_n N_Q_N_c_2204_n 0.0116659f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1101 N_A_1587_329#_M1029_g N_Q_N_c_2204_n 0.017611f $X=11.455 $Y=1.985 $X2=0
+ $Y2=0
cc_1102 N_A_1587_329#_c_1590_n N_Q_N_c_2204_n 0.0249928f $X=12.32 $Y=1.16 $X2=0
+ $Y2=0
cc_1103 N_A_1587_329#_c_1592_n N_Q_N_c_2204_n 0.0102263f $X=11.455 $Y=1.16 $X2=0
+ $Y2=0
cc_1104 N_A_1587_329#_M1027_g Q 4.73325e-19 $X=12.395 $Y=2.095 $X2=0 $Y2=0
cc_1105 N_A_1587_329#_c_1616_n N_VGND_c_2249_n 0.00740647f $X=9.655 $Y=0.36
+ $X2=0 $Y2=0
cc_1106 N_A_1587_329#_c_1594_n N_VGND_c_2249_n 0.00387989f $X=9.74 $Y=0.845
+ $X2=0 $Y2=0
cc_1107 N_A_1587_329#_c_1596_n N_VGND_c_2249_n 0.00778757f $X=10.38 $Y=0.93
+ $X2=0 $Y2=0
cc_1108 N_A_1587_329#_c_1597_n N_VGND_c_2249_n 0.0039218f $X=10.38 $Y=0.93 $X2=0
+ $Y2=0
cc_1109 N_A_1587_329#_c_1598_n N_VGND_c_2249_n 0.00287978f $X=10.417 $Y=0.765
+ $X2=0 $Y2=0
cc_1110 N_A_1587_329#_c_1588_n N_VGND_c_2250_n 0.00537422f $X=11.38 $Y=1.16
+ $X2=0 $Y2=0
cc_1111 N_A_1587_329#_c_1589_n N_VGND_c_2250_n 0.00444548f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1112 N_A_1587_329#_c_1598_n N_VGND_c_2250_n 0.00213038f $X=10.417 $Y=0.765
+ $X2=0 $Y2=0
cc_1113 N_A_1587_329#_M1033_g N_VGND_c_2251_n 0.00642475f $X=12.395 $Y=0.445
+ $X2=0 $Y2=0
cc_1114 N_A_1587_329#_c_1616_n N_VGND_c_2256_n 0.0730142f $X=9.655 $Y=0.36 $X2=0
+ $Y2=0
cc_1115 N_A_1587_329#_c_1597_n N_VGND_c_2260_n 9.87024e-19 $X=10.38 $Y=0.93
+ $X2=0 $Y2=0
cc_1116 N_A_1587_329#_c_1598_n N_VGND_c_2260_n 0.00539883f $X=10.417 $Y=0.765
+ $X2=0 $Y2=0
cc_1117 N_A_1587_329#_c_1589_n N_VGND_c_2261_n 0.00541359f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1118 N_A_1587_329#_M1033_g N_VGND_c_2261_n 0.00585385f $X=12.395 $Y=0.445
+ $X2=0 $Y2=0
cc_1119 N_A_1587_329#_M1006_d N_VGND_c_2263_n 0.00380013f $X=8.415 $Y=0.235
+ $X2=0 $Y2=0
cc_1120 N_A_1587_329#_c_1589_n N_VGND_c_2263_n 0.0121537f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1121 N_A_1587_329#_M1033_g N_VGND_c_2263_n 0.0121969f $X=12.395 $Y=0.445
+ $X2=0 $Y2=0
cc_1122 N_A_1587_329#_c_1616_n N_VGND_c_2263_n 0.0508216f $X=9.655 $Y=0.36 $X2=0
+ $Y2=0
cc_1123 N_A_1587_329#_c_1596_n N_VGND_c_2263_n 0.0174077f $X=10.38 $Y=0.93 $X2=0
+ $Y2=0
cc_1124 N_A_1587_329#_c_1597_n N_VGND_c_2263_n 0.00131752f $X=10.38 $Y=0.93
+ $X2=0 $Y2=0
cc_1125 N_A_1587_329#_c_1598_n N_VGND_c_2263_n 0.00805362f $X=10.417 $Y=0.765
+ $X2=0 $Y2=0
cc_1126 N_A_1587_329#_c_1616_n A_1807_47# 0.00460484f $X=9.655 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1127 N_A_1587_329#_c_1616_n A_1879_47# 0.0142908f $X=9.655 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1128 N_A_1587_329#_c_1594_n A_1879_47# 0.00689044f $X=9.74 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_1129 N_A_2412_47#_c_1761_n N_VPWR_c_1859_n 0.0149126f $X=12.185 $Y=1.93 $X2=0
+ $Y2=0
cc_1130 N_A_2412_47#_M1003_g N_VPWR_c_1860_n 0.00363679f $X=12.87 $Y=1.985 $X2=0
+ $Y2=0
cc_1131 N_A_2412_47#_c_1761_n N_VPWR_c_1860_n 0.0274302f $X=12.185 $Y=1.93 $X2=0
+ $Y2=0
cc_1132 N_A_2412_47#_c_1757_n N_VPWR_c_1860_n 0.0105531f $X=12.815 $Y=1.16 $X2=0
+ $Y2=0
cc_1133 N_A_2412_47#_c_1758_n N_VPWR_c_1860_n 0.0014049f $X=12.815 $Y=1.16 $X2=0
+ $Y2=0
cc_1134 N_A_2412_47#_M1003_g N_VPWR_c_1870_n 0.00541964f $X=12.87 $Y=1.985 $X2=0
+ $Y2=0
cc_1135 N_A_2412_47#_M1003_g N_VPWR_c_1851_n 0.0106947f $X=12.87 $Y=1.985 $X2=0
+ $Y2=0
cc_1136 N_A_2412_47#_c_1761_n N_VPWR_c_1851_n 0.00801045f $X=12.185 $Y=1.93
+ $X2=0 $Y2=0
cc_1137 N_A_2412_47#_c_1756_n N_Q_N_c_2204_n 0.0476102f $X=12.185 $Y=0.44 $X2=0
+ $Y2=0
cc_1138 N_A_2412_47#_c_1761_n N_Q_N_c_2204_n 0.073327f $X=12.185 $Y=1.93 $X2=0
+ $Y2=0
cc_1139 N_A_2412_47#_c_1772_n N_Q_N_c_2204_n 0.0206626f $X=12.165 $Y=1.16 $X2=0
+ $Y2=0
cc_1140 N_A_2412_47#_c_1759_n Q 0.00258335f $X=12.815 $Y=0.995 $X2=0 $Y2=0
cc_1141 N_A_2412_47#_M1003_g Q 0.00850773f $X=12.87 $Y=1.985 $X2=0 $Y2=0
cc_1142 N_A_2412_47#_c_1759_n N_Q_c_2223_n 0.00425287f $X=12.815 $Y=0.995 $X2=0
+ $Y2=0
cc_1143 N_A_2412_47#_M1003_g Q 0.00433918f $X=12.87 $Y=1.985 $X2=0 $Y2=0
cc_1144 N_A_2412_47#_c_1757_n Q 0.0263712f $X=12.815 $Y=1.16 $X2=0 $Y2=0
cc_1145 N_A_2412_47#_c_1758_n Q 0.00757624f $X=12.815 $Y=1.16 $X2=0 $Y2=0
cc_1146 N_A_2412_47#_c_1759_n Q 0.00416176f $X=12.815 $Y=0.995 $X2=0 $Y2=0
cc_1147 N_A_2412_47#_M1003_g Q 0.00332631f $X=12.87 $Y=1.985 $X2=0 $Y2=0
cc_1148 N_A_2412_47#_c_1761_n Q 0.00219581f $X=12.185 $Y=1.93 $X2=0 $Y2=0
cc_1149 N_A_2412_47#_c_1756_n N_VGND_c_2251_n 0.0201419f $X=12.185 $Y=0.44 $X2=0
+ $Y2=0
cc_1150 N_A_2412_47#_c_1757_n N_VGND_c_2251_n 0.017073f $X=12.815 $Y=1.16 $X2=0
+ $Y2=0
cc_1151 N_A_2412_47#_c_1758_n N_VGND_c_2251_n 0.00147264f $X=12.815 $Y=1.16
+ $X2=0 $Y2=0
cc_1152 N_A_2412_47#_c_1759_n N_VGND_c_2251_n 0.00378931f $X=12.815 $Y=0.995
+ $X2=0 $Y2=0
cc_1153 N_A_2412_47#_c_1756_n N_VGND_c_2261_n 0.0144177f $X=12.185 $Y=0.44 $X2=0
+ $Y2=0
cc_1154 N_A_2412_47#_c_1759_n N_VGND_c_2262_n 0.00542163f $X=12.815 $Y=0.995
+ $X2=0 $Y2=0
cc_1155 N_A_2412_47#_M1033_s N_VGND_c_2263_n 0.00386369f $X=12.06 $Y=0.235 $X2=0
+ $Y2=0
cc_1156 N_A_2412_47#_c_1756_n N_VGND_c_2263_n 0.00801045f $X=12.185 $Y=0.44
+ $X2=0 $Y2=0
cc_1157 N_A_2412_47#_c_1759_n N_VGND_c_2263_n 0.0106134f $X=12.815 $Y=0.995
+ $X2=0 $Y2=0
cc_1158 N_A_27_369#_c_1804_n N_VPWR_M1021_d 0.00300292f $X=0.935 $Y=1.935
+ $X2=-0.19 $Y2=1.305
cc_1159 N_A_27_369#_c_1804_n N_VPWR_c_1852_n 0.0142338f $X=0.935 $Y=1.935 $X2=0
+ $Y2=0
cc_1160 N_A_27_369#_c_1804_n N_VPWR_c_1861_n 0.00212534f $X=0.935 $Y=1.935 $X2=0
+ $Y2=0
cc_1161 N_A_27_369#_c_1818_n N_VPWR_c_1861_n 0.0098514f $X=1.105 $Y=2.36 $X2=0
+ $Y2=0
cc_1162 N_A_27_369#_c_1806_n N_VPWR_c_1861_n 0.0532339f $X=1.88 $Y=2.34 $X2=0
+ $Y2=0
cc_1163 N_A_27_369#_c_1803_n N_VPWR_c_1865_n 0.0178803f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1164 N_A_27_369#_c_1804_n N_VPWR_c_1865_n 0.00212534f $X=0.935 $Y=1.935 $X2=0
+ $Y2=0
cc_1165 N_A_27_369#_M1021_s N_VPWR_c_1851_n 0.00231948f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_1166 N_A_27_369#_M1001_d N_VPWR_c_1851_n 0.00209344f $X=1.745 $Y=1.845 $X2=0
+ $Y2=0
cc_1167 N_A_27_369#_c_1803_n N_VPWR_c_1851_n 0.00991202f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1168 N_A_27_369#_c_1804_n N_VPWR_c_1851_n 0.00897281f $X=0.935 $Y=1.935 $X2=0
+ $Y2=0
cc_1169 N_A_27_369#_c_1818_n N_VPWR_c_1851_n 0.00639401f $X=1.105 $Y=2.36 $X2=0
+ $Y2=0
cc_1170 N_A_27_369#_c_1806_n N_VPWR_c_1851_n 0.0337295f $X=1.88 $Y=2.34 $X2=0
+ $Y2=0
cc_1171 N_A_27_369#_c_1804_n A_193_369# 0.00298964f $X=0.935 $Y=1.935 $X2=-0.19
+ $Y2=1.305
cc_1172 N_A_27_369#_c_1811_n A_193_369# 0.00239321f $X=1.02 $Y=2.255 $X2=-0.19
+ $Y2=1.305
cc_1173 N_A_27_369#_c_1818_n A_193_369# 8.09413e-19 $X=1.105 $Y=2.36 $X2=-0.19
+ $Y2=1.305
cc_1174 N_A_27_369#_c_1806_n A_193_369# 3.49598e-19 $X=1.88 $Y=2.34 $X2=-0.19
+ $Y2=1.305
cc_1175 N_A_27_369#_c_1806_n N_A_181_47#_M1004_d 0.00317809f $X=1.88 $Y=2.34
+ $X2=0 $Y2=0
cc_1176 N_A_27_369#_c_1804_n N_A_181_47#_c_2071_n 0.0118796f $X=0.935 $Y=1.935
+ $X2=0 $Y2=0
cc_1177 N_A_27_369#_c_1811_n N_A_181_47#_c_2071_n 0.00335193f $X=1.02 $Y=2.255
+ $X2=0 $Y2=0
cc_1178 N_A_27_369#_c_1806_n N_A_181_47#_c_2071_n 0.0183361f $X=1.88 $Y=2.34
+ $X2=0 $Y2=0
cc_1179 N_A_27_369#_c_1806_n N_A_181_47#_c_2065_n 0.00157f $X=1.88 $Y=2.34 $X2=0
+ $Y2=0
cc_1180 N_A_27_369#_c_1804_n N_A_181_47#_c_2060_n 0.00108706f $X=0.935 $Y=1.935
+ $X2=0 $Y2=0
cc_1181 N_VPWR_c_1851_n A_193_369# 0.00168634f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1182 N_VPWR_c_1851_n N_A_181_47#_M1004_d 0.00216833f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1851_n N_A_181_47#_M1007_s 0.00194602f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1863_n N_A_181_47#_c_2062_n 0.0135531f $X=5.945 $Y=2.72 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1851_n N_A_181_47#_c_2062_n 0.00399922f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1853_n N_A_181_47#_c_2064_n 0.00822115f $X=2.82 $Y=2.34 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1851_n A_1081_413# 0.00244888f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1188 N_VPWR_c_1875_n A_1514_329# 0.00101109f $X=7.96 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1189 N_VPWR_c_1851_n A_1712_413# 0.00232248f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1190 N_VPWR_c_1851_n N_Q_N_M1029_d 0.00209319f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1191 N_VPWR_c_1859_n N_Q_N_c_2204_n 0.0210382f $X=12.575 $Y=2.72 $X2=0 $Y2=0
cc_1192 N_VPWR_c_1851_n N_Q_N_c_2204_n 0.0124268f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1193 N_VPWR_c_1851_n N_Q_M1003_d 0.00209863f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1194 N_VPWR_c_1870_n Q 0.0198578f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1195 N_VPWR_c_1851_n Q 0.0127182f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1196 N_VPWR_c_1858_n N_VGND_c_2250_n 0.00700912f $X=11.245 $Y=1.66 $X2=0
+ $Y2=0
cc_1197 N_A_181_47#_c_2068_n N_VGND_c_2245_n 0.0113707f $X=1.38 $Y=0.42 $X2=0
+ $Y2=0
cc_1198 N_A_181_47#_c_2058_n N_VGND_c_2246_n 0.0209118f $X=1.6 $Y=0.705 $X2=0
+ $Y2=0
cc_1199 N_A_181_47#_c_2068_n N_VGND_c_2252_n 0.0238306f $X=1.38 $Y=0.42 $X2=0
+ $Y2=0
cc_1200 N_A_181_47#_c_2058_n N_VGND_c_2252_n 0.0151677f $X=1.6 $Y=0.705 $X2=0
+ $Y2=0
cc_1201 N_A_181_47#_c_2056_n N_VGND_c_2259_n 0.0220997f $X=4.73 $Y=0.42 $X2=0
+ $Y2=0
cc_1202 N_A_181_47#_M1012_d N_VGND_c_2263_n 0.00216413f $X=0.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1203 N_A_181_47#_M1023_s N_VGND_c_2263_n 0.00330824f $X=4.605 $Y=0.235 $X2=0
+ $Y2=0
cc_1204 N_A_181_47#_c_2068_n N_VGND_c_2263_n 0.0177716f $X=1.38 $Y=0.42 $X2=0
+ $Y2=0
cc_1205 N_A_181_47#_c_2056_n N_VGND_c_2263_n 0.0124358f $X=4.73 $Y=0.42 $X2=0
+ $Y2=0
cc_1206 N_A_181_47#_c_2058_n N_VGND_c_2263_n 0.0110868f $X=1.6 $Y=0.705 $X2=0
+ $Y2=0
cc_1207 N_A_181_47#_c_2058_n A_265_47# 0.00402976f $X=1.6 $Y=0.705 $X2=-0.19
+ $Y2=-0.24
cc_1208 N_Q_N_c_2204_n N_VGND_c_2261_n 0.0210382f $X=11.665 $Y=0.38 $X2=0 $Y2=0
cc_1209 N_Q_N_M1005_d N_VGND_c_2263_n 0.00209319f $X=11.53 $Y=0.235 $X2=0 $Y2=0
cc_1210 N_Q_N_c_2204_n N_VGND_c_2263_n 0.0124268f $X=11.665 $Y=0.38 $X2=0 $Y2=0
cc_1211 N_Q_c_2223_n N_VGND_c_2262_n 0.019206f $X=13.08 $Y=0.4 $X2=0 $Y2=0
cc_1212 N_Q_M1019_d N_VGND_c_2263_n 0.00210124f $X=12.945 $Y=0.235 $X2=0 $Y2=0
cc_1213 N_Q_c_2223_n N_VGND_c_2263_n 0.0126519f $X=13.08 $Y=0.4 $X2=0 $Y2=0
cc_1214 N_VGND_c_2263_n A_109_47# 0.00283904f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1215 N_VGND_c_2263_n A_265_47# 0.00217974f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1216 N_VGND_c_2263_n A_1087_47# 0.00726675f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1217 N_VGND_c_2263_n A_1514_47# 0.014219f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1218 N_VGND_c_2266_n A_1514_47# 0.0105439f $X=7.63 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1219 N_VGND_c_2263_n A_1807_47# 0.00169327f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1220 N_VGND_c_2263_n A_1879_47# 0.00437636f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o21ai_1.spice
* Created: Thu Aug 27 14:35:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21ai_1.spice.pex"
.subckt sky130_fd_sc_hd__o21ai_1  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.169 PD=0.98 PS=1.82 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_47#_M1002_d N_A2_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_27_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 A_109_297# N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.26 PD=1.21 PS=2.52 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75000.9
+ A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g A_109_297# VPB PHIGHVT L=0.15 W=1 AD=0.204706
+ AS=0.105 PD=1.63529 PS=1.21 NRD=16.7253 NRS=9.8303 M=1 R=6.66667 SA=75000.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=0.7 AD=0.182
+ AS=0.143294 PD=1.92 PS=1.14471 NRD=0 NRS=7.0329 M=1 R=4.66667 SA=75001.1
+ SB=75000.2 A=0.105 P=1.7 MULT=1
DX6_noxref VNB VPB NWDIODE A=3.5631 P=7.65
*
.include "sky130_fd_sc_hd__o21ai_1.spice.SKY130_FD_SC_HD__O21AI_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a2111o_2.spice.pex
* Created: Thu Aug 27 13:58:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111O_2%A_86_235# 1 2 3 12 14 16 19 21 23 24 30 33
+ 35 37 38 41 43 47 49 50 51 55
c95 49 0 1.96852e-19 $X=1.6 $Y=1.2
r96 54 55 12.2413 $w=3.15e-07 $l=8e-08 $layer=POLY_cond $X=0.935 $Y=1.16
+ $X2=1.015 $Y2=1.16
r97 53 54 53.5556 $w=3.15e-07 $l=3.5e-07 $layer=POLY_cond $X=0.585 $Y=1.16
+ $X2=0.935 $Y2=1.16
r98 45 47 9.17251 $w=2.43e-07 $l=1.95e-07 $layer=LI1_cond $X=3.212 $Y=0.615
+ $X2=3.212 $Y2=0.42
r99 44 51 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.42 $Y=0.7 $X2=2.3
+ $Y2=0.7
r100 43 45 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.09 $Y=0.7
+ $X2=3.212 $Y2=0.615
r101 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.09 $Y=0.7
+ $X2=2.42 $Y2=0.7
r102 39 51 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.615
+ $X2=2.3 $Y2=0.7
r103 39 41 9.3636 $w=2.38e-07 $l=1.95e-07 $layer=LI1_cond $X=2.3 $Y=0.615
+ $X2=2.3 $Y2=0.42
r104 37 51 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.18 $Y=0.7 $X2=2.3
+ $Y2=0.7
r105 37 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.18 $Y=0.7
+ $X2=1.705 $Y2=0.7
r106 33 50 6.65895 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.64 $Y=1.64
+ $X2=1.64 $Y2=1.495
r107 33 35 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=1.64 $Y=1.64
+ $X2=1.64 $Y2=1.66
r108 31 49 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.6 $Y=1.325
+ $X2=1.6 $Y2=1.2
r109 31 50 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.6 $Y=1.325
+ $X2=1.6 $Y2=1.495
r110 30 49 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.6 $Y=1.075
+ $X2=1.6 $Y2=1.2
r111 29 38 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.6 $Y=0.785
+ $X2=1.705 $Y2=0.7
r112 29 30 15.316 $w=2.08e-07 $l=2.9e-07 $layer=LI1_cond $X=1.6 $Y=0.785 $X2=1.6
+ $Y2=1.075
r113 27 55 35.9587 $w=3.15e-07 $l=2.35e-07 $layer=POLY_cond $X=1.25 $Y=1.16
+ $X2=1.015 $Y2=1.16
r114 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.16 $X2=1.25 $Y2=1.16
r115 24 49 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.495 $Y=1.2
+ $X2=1.6 $Y2=1.2
r116 24 26 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=1.495 $Y=1.2
+ $X2=1.25 $Y2=1.2
r117 21 55 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=1.16
r118 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=0.56
r119 17 54 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.325
+ $X2=0.935 $Y2=1.16
r120 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.935 $Y=1.325
+ $X2=0.935 $Y2=1.985
r121 14 53 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=0.995
+ $X2=0.585 $Y2=1.16
r122 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.585 $Y=0.995
+ $X2=0.585 $Y2=0.56
r123 10 53 12.2413 $w=3.15e-07 $l=2.0106e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.585 $Y2=1.16
r124 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=1.985
r125 3 35 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.485 $X2=1.7 $Y2=1.66
r126 2 47 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.235 $X2=3.23 $Y2=0.42
r127 1 41 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.275 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%D1 3 6 8 9 10 11 17 18 19
r39 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.16
+ $X2=1.97 $Y2=1.325
r40 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.16
+ $X2=1.97 $Y2=0.995
r41 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r42 10 11 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.107 $Y=1.87
+ $X2=2.107 $Y2=2.21
r43 9 10 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.107 $Y=1.53
+ $X2=2.107 $Y2=1.87
r44 9 33 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=2.107 $Y=1.53
+ $X2=2.107 $Y2=1.325
r45 8 33 4.71133 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.325
r46 8 18 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=2.07 $Y=1.19 $X2=2.07
+ $Y2=1.16
r47 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.06 $Y=1.985
+ $X2=2.06 $Y2=1.325
r48 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.06 $Y=0.56 $X2=2.06
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%C1 3 7 8 9 10 11 17 19
r35 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.16
+ $X2=2.51 $Y2=1.325
r36 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.16
+ $X2=2.51 $Y2=0.995
r37 10 11 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=2.58 $Y=1.87
+ $X2=2.58 $Y2=2.21
r38 9 10 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=2.58 $Y=1.53 $X2=2.58
+ $Y2=1.87
r39 8 9 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.58 $Y=1.16 $X2=2.58
+ $Y2=1.53
r40 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.16 $X2=2.51 $Y2=1.16
r41 7 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.49 $Y=0.56 $X2=2.49
+ $Y2=0.995
r42 3 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.42 $Y=1.985
+ $X2=2.42 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%B1 3 7 8 9 13 15
r36 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.16
+ $X2=3.05 $Y2=1.325
r37 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.16
+ $X2=3.05 $Y2=0.995
r38 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.05 $Y=1.16 $X2=3.05
+ $Y2=1.53
r39 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.05
+ $Y=1.16 $X2=3.05 $Y2=1.16
r40 7 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.015 $Y=0.56
+ $X2=3.015 $Y2=0.995
r41 3 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.96 $Y=1.985
+ $X2=2.96 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%A1 3 6 8 9 10 16 17 18 23 29
r44 29 30 17.3251 $w=4.38e-07 $l=6.22e-07 $layer=LI1_cond $X=3.68 $Y=0.51
+ $X2=3.68 $Y2=1.132
r45 17 30 0.846205 $w=4.38e-07 $l=1.23207e-07 $layer=LI1_cond $X=3.57 $Y=1.16
+ $X2=3.68 $Y2=1.132
r46 17 23 0.843251 $w=4.08e-07 $l=3e-08 $layer=LI1_cond $X=3.57 $Y=1.16 $X2=3.57
+ $Y2=1.19
r47 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.16
+ $X2=3.59 $Y2=1.325
r48 16 18 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.59 $Y=1.16
+ $X2=3.59 $Y2=0.98
r49 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.16 $X2=3.59 $Y2=1.16
r50 10 29 6.33358 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.91 $Y=0.51 $X2=3.68
+ $Y2=0.51
r51 8 30 6.33358 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.45 $Y=1.132 $X2=3.68
+ $Y2=1.132
r52 8 9 8.79792 $w=4.08e-07 $l=3.13e-07 $layer=LI1_cond $X=3.57 $Y=1.217
+ $X2=3.57 $Y2=1.53
r53 8 23 0.758926 $w=4.08e-07 $l=2.7e-08 $layer=LI1_cond $X=3.57 $Y=1.217
+ $X2=3.57 $Y2=1.19
r54 6 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.5 $Y=1.985 $X2=3.5
+ $Y2=1.325
r55 3 18 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.5 $Y=0.56 $X2=3.5
+ $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%A2 3 6 8 9 13 14 15
r28 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.16
+ $X2=4.13 $Y2=1.325
r29 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.16
+ $X2=4.13 $Y2=0.995
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.16 $X2=4.13 $Y2=1.16
r31 8 9 7.1345 $w=5.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.23 $Y=1.19 $X2=4.23
+ $Y2=1.53
r32 8 14 0.629515 $w=5.68e-07 $l=3e-08 $layer=LI1_cond $X=4.23 $Y=1.19 $X2=4.23
+ $Y2=1.16
r33 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.04 $Y=1.985
+ $X2=4.04 $Y2=1.325
r34 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.04 $Y=0.56 $X2=4.04
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%VPWR 1 2 3 10 12 16 22 25 26 27 29 42 43 49
r56 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r58 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r59 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 37 40 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 36 39 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 34 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=2.72
+ $X2=1.19 $Y2=2.72
r65 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.315 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 33 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 30 46 5.00068 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.217 $Y2=2.72
r69 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 29 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.19 $Y2=2.72
r71 29 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 27 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 27 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 25 39 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.59 $Y=2.72
+ $X2=3.45 $Y2=2.72
r75 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=2.72
+ $X2=3.755 $Y2=2.72
r76 24 42 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.92 $Y=2.72
+ $X2=4.37 $Y2=2.72
r77 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.92 $Y=2.72
+ $X2=3.755 $Y2=2.72
r78 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=2.635
+ $X2=3.755 $Y2=2.72
r79 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.755 $Y=2.635
+ $X2=3.755 $Y2=2.34
r80 16 19 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.19 $Y=1.66
+ $X2=1.19 $Y2=2.34
r81 14 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=2.635
+ $X2=1.19 $Y2=2.72
r82 14 19 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.19 $Y=2.635
+ $X2=1.19 $Y2=2.34
r83 10 46 2.93618 $w=3.5e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.217 $Y2=2.72
r84 10 12 26.8355 $w=3.48e-07 $l=8.15e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=1.82
r85 3 22 600 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=3.575
+ $Y=1.485 $X2=3.755 $Y2=2.34
r86 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.485 $X2=1.15 $Y2=2.34
r87 2 16 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.485 $X2=1.15 $Y2=1.66
r88 1 12 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.485 $X2=0.29 $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%X 1 2 7 8 9 10 11 12 20
r17 11 12 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=1.87
+ $X2=0.75 $Y2=2.21
r18 11 31 6.35831 $w=2.88e-07 $l=1.6e-07 $layer=LI1_cond $X=0.75 $Y=1.87
+ $X2=0.75 $Y2=1.71
r19 10 31 7.15309 $w=2.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.75 $Y=1.53
+ $X2=0.75 $Y2=1.71
r20 9 10 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=1.19 $X2=0.75
+ $Y2=1.53
r21 8 9 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=0.85 $X2=0.75
+ $Y2=1.19
r22 7 8 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=0.51 $X2=0.75
+ $Y2=0.85
r23 7 20 3.57655 $w=2.88e-07 $l=9e-08 $layer=LI1_cond $X=0.75 $Y=0.51 $X2=0.75
+ $Y2=0.42
r24 2 31 300 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.485 $X2=0.72 $Y2=1.71
r25 1 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.235 $X2=0.8 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%A_607_297# 1 2 7 9 11
r21 12 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=2 $X2=3.235
+ $Y2=2
r22 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.09 $Y=2 $X2=3.4
+ $Y2=2
r23 7 14 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=2.085
+ $X2=3.235 $Y2=2
r24 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.235 $Y=2.085
+ $X2=3.235 $Y2=2.34
r25 2 11 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=4.115
+ $Y=1.485 $X2=4.255 $Y2=2
r26 1 14 600 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.485 $X2=3.235 $Y2=2
r27 1 9 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.485 $X2=3.235 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_2%VGND 1 2 3 4 13 15 19 23 25 27 30 33 35 36
+ 37 39 51 62 67
r71 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r72 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r73 57 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r74 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r75 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r76 53 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r77 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r78 51 66 5.00668 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.382
+ $Y2=0
r79 51 56 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=3.91
+ $Y2=0
r80 50 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r81 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r82 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r83 47 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r84 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r85 44 62 4.00737 $w=3.5e-07 $l=1.3e-07 $layer=LI1_cond $X=1.325 $Y=0.18
+ $X2=1.195 $Y2=0.18
r86 44 46 6.43174 $w=5.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.325 $Y=0.18
+ $X2=1.61 $Y2=0.18
r87 43 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r88 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r89 40 59 5.00068 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r90 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.69
+ $Y2=0
r91 39 62 4.00737 $w=3.5e-07 $l=2.3622e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=1.195 $Y2=0.18
r92 39 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.69
+ $Y2=0
r93 37 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r94 37 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r95 35 49 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.53
+ $Y2=0
r96 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.755
+ $Y2=0
r97 34 53 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.99
+ $Y2=0
r98 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.755
+ $Y2=0
r99 33 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.53
+ $Y2=0
r100 32 33 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0.18
+ $X2=2.01 $Y2=0.18
r101 30 46 3.04661 $w=5.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=0.18
+ $X2=1.61 $Y2=0.18
r102 30 32 2.25675 $w=5.28e-07 $l=1e-07 $layer=LI1_cond $X=1.745 $Y=0.18
+ $X2=1.845 $Y2=0.18
r103 25 66 2.93018 $w=3.5e-07 $l=1.03899e-07 $layer=LI1_cond $X=4.34 $Y=0.085
+ $X2=4.382 $Y2=0
r104 25 27 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.34 $Y=0.085
+ $X2=4.34 $Y2=0.38
r105 21 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.085
+ $X2=2.755 $Y2=0
r106 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.755 $Y=0.085
+ $X2=2.755 $Y2=0.36
r107 17 62 2.43179 $w=2.6e-07 $l=2.65e-07 $layer=LI1_cond $X=1.195 $Y=0.445
+ $X2=1.195 $Y2=0.18
r108 17 19 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=1.195 $Y=0.445
+ $X2=1.195 $Y2=0.7
r109 13 59 2.93618 $w=3.5e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.217 $Y2=0
r110 13 15 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r111 4 27 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=4.115
+ $Y=0.235 $X2=4.33 $Y2=0.38
r112 3 23 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.235 $X2=2.755 $Y2=0.36
r113 2 62 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.36
r114 2 32 182 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.845 $Y2=0.36
r115 2 19 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.7
r116 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.235 $X2=0.35 $Y2=0.38
.ends


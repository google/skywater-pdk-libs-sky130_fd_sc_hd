* File: sky130_fd_sc_hd__nor2_4.spice.pex
* Created: Thu Aug 27 14:31:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR2_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 42 43
r80 41 43 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.62 $Y=1.16 $X2=1.75
+ $Y2=1.16
r81 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r82 39 41 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.62 $Y2=1.16
r83 38 39 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r84 36 38 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.6 $Y=1.16 $X2=0.91
+ $Y2=1.16
r85 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6 $Y=1.16
+ $X2=0.6 $Y2=1.16
r86 33 36 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.6
+ $Y2=1.16
r87 30 42 51.2955 $w=1.98e-07 $l=9.25e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.62 $Y2=1.175
r88 30 37 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.6 $Y2=1.175
r89 29 37 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.6 $Y2=1.175
r90 25 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r91 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r92 22 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r93 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r94 18 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r95 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r96 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r97 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r98 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r99 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r100 8 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r101 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r102 4 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r103 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r104 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
c88 13 0 7.39456e-20 $X=2.59 $Y=1.985
r89 39 41 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.315 $Y=1.16
+ $X2=3.43 $Y2=1.16
r90 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.315
+ $Y=1.16 $X2=3.315 $Y2=1.16
r91 37 39 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.315 $Y2=1.16
r92 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=3.01 $Y2=1.16
r93 34 36 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=2.295 $Y=1.16
+ $X2=2.59 $Y2=1.16
r94 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.295
+ $Y=1.16 $X2=2.295 $Y2=1.16
r95 31 34 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.17 $Y=1.16
+ $X2=2.295 $Y2=1.16
r96 29 40 17.7455 $w=1.98e-07 $l=3.2e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=3.315 $Y2=1.175
r97 29 35 38.8182 $w=1.98e-07 $l=7e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=2.295 $Y2=1.175
r98 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r99 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.985
r100 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r101 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r102 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r103 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.985
r104 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.16
r105 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r106 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.16
r107 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.985
r108 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r109 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r110 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r111 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r112 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r113 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 36 41 46 48
c77 28 0 7.39456e-20 $X=1.96 $Y=1.665
r78 37 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=2.38
+ $X2=2.8 $Y2=2.38
r79 36 48 10.5525 $w=4.13e-07 $l=3.8e-07 $layer=LI1_cond $X=3.682 $Y=2.38
+ $X2=3.682 $Y2=2
r80 36 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.475 $Y=2.38
+ $X2=2.965 $Y2=2.38
r81 32 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=2.295 $X2=2.8
+ $Y2=2.38
r82 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.8 $Y=2.295
+ $X2=2.8 $Y2=2.02
r83 31 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=2.38
+ $X2=1.96 $Y2=2.38
r84 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=2.38
+ $X2=2.8 $Y2=2.38
r85 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.635 $Y=2.38
+ $X2=2.125 $Y2=2.38
r86 29 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.295 $X2=1.96
+ $Y2=2.38
r87 28 43 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=1.56
r88 28 29 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=2.295
r89 27 41 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.56 $X2=1.12
+ $Y2=1.56
r90 26 43 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=1.56
+ $X2=1.96 $Y2=1.56
r91 26 27 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=1.795 $Y=1.56
+ $X2=1.205 $Y2=1.56
r92 22 41 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.56
r93 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=2.3
r94 21 39 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=1.56
+ $X2=0.227 $Y2=1.56
r95 20 41 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=1.56 $X2=1.12
+ $Y2=1.56
r96 20 21 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.035 $Y=1.56
+ $X2=0.365 $Y2=1.56
r97 16 39 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=1.56
r98 16 18 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=2.3
r99 5 48 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=2
r100 4 34 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=2.02
r101 3 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.34
r102 3 43 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r103 2 41 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r104 2 24 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r105 1 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r106 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_4%VPWR 1 2 9 13 15 17 22 29 30 33 36
r56 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 30 37 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.5 $Y2=2.72
r61 27 29 149.075 $w=1.68e-07 $l=2.285e-06 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.7 $Y2=2.72
r66 23 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 22 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.5 $Y2=2.72
r68 22 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.7 $Y2=2.72
r70 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 11 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=2.635
+ $X2=1.5 $Y2=2.72
r74 11 13 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.5 $Y=2.635
+ $X2=1.5 $Y2=2
r75 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r76 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2
r77 2 13 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2
r78 1 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_4%Y 1 2 3 4 5 6 21 23 24 27 29 33 35 37 39 41
+ 45 49 51 53 55 56 59 61 63
r121 62 63 12.128 $w=5.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.855 $Y=0.905
+ $X2=3.855 $Y2=1.445
r122 54 59 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.815
+ $X2=3.22 $Y2=0.815
r123 53 62 8.17735 $w=1.8e-07 $l=2.40832e-07 $layer=LI1_cond $X=3.655 $Y=0.815
+ $X2=3.855 $Y2=0.905
r124 53 54 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.655 $Y=0.815
+ $X2=3.385 $Y2=0.815
r125 52 61 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=1.595
+ $X2=3.22 $Y2=1.595
r126 51 63 3.99943 $w=3e-07 $l=2e-07 $layer=LI1_cond $X=3.655 $Y=1.595 $X2=3.855
+ $Y2=1.595
r127 51 52 13.4452 $w=2.98e-07 $l=3.5e-07 $layer=LI1_cond $X=3.655 $Y=1.595
+ $X2=3.305 $Y2=1.595
r128 47 61 3.44808 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.22 $Y=1.745
+ $X2=3.22 $Y2=1.595
r129 47 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.22 $Y=1.745
+ $X2=3.22 $Y2=1.96
r130 43 59 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.815
r131 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.39
r132 42 56 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0.815
+ $X2=2.38 $Y2=0.815
r133 41 59 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=3.22 $Y2=0.815
r134 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=2.545 $Y2=0.815
r135 40 58 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.595
+ $X2=2.38 $Y2=1.595
r136 39 61 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=1.595
+ $X2=3.22 $Y2=1.595
r137 39 40 25.7379 $w=2.98e-07 $l=6.7e-07 $layer=LI1_cond $X=3.135 $Y=1.595
+ $X2=2.465 $Y2=1.595
r138 35 58 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.38 $Y=1.745
+ $X2=2.38 $Y2=1.595
r139 35 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.38 $Y=1.745
+ $X2=2.38 $Y2=1.96
r140 31 56 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.815
r141 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.39
r142 30 55 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r143 29 56 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=2.38 $Y2=0.815
r144 29 30 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=1.705 $Y2=0.815
r145 25 55 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r146 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r147 23 55 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r148 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r149 19 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r150 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r151 6 61 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.62
r152 6 49 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.96
r153 5 58 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.62
r154 5 37 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.96
r155 4 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.39
r156 3 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.39
r157 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r158 1 21 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 64 65
r75 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r76 62 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r77 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r78 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r79 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r80 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r81 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r82 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r83 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r84 50 68 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r85 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r86 48 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r87 48 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r88 46 61 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.45
+ $Y2=0
r89 46 47 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.697
+ $Y2=0
r90 45 64 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.91
+ $Y2=0
r91 45 47 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.697
+ $Y2=0
r92 43 58 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.53
+ $Y2=0
r93 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.8
+ $Y2=0
r94 42 61 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r95 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.8
+ $Y2=0
r96 40 55 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r97 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r98 39 58 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.53
+ $Y2=0
r99 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r100 37 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r101 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r102 36 55 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r103 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r104 32 47 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.697 $Y=0.085
+ $X2=3.697 $Y2=0
r105 32 34 12.3332 $w=2.83e-07 $l=3.05e-07 $layer=LI1_cond $X=3.697 $Y=0.085
+ $X2=3.697 $Y2=0.39
r106 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r107 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.39
r108 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r109 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r110 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r111 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r112 16 68 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r113 16 18 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r114 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.39
r115 4 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.39
r116 3 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r117 2 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r118 1 18 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.495000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.075000 3.080000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.845000 1.275000 ;
    END
  END D
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 3.925000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.355000 1.665000 2.685000 2.465000 ;
        RECT 3.370000 1.055000 3.925000 1.445000 ;
        RECT 3.595000 0.635000 3.925000 1.055000 ;
        RECT 3.595000 1.665000 3.925000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 1.185000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 2.125000 0.465000 ;
      RECT 0.935000  0.465000 1.185000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.635000 3.085000 0.905000 ;
      RECT 1.855000  1.835000 2.185000 2.635000 ;
      RECT 2.315000  0.255000 4.425000 0.465000 ;
      RECT 2.995000  1.835000 3.325000 2.635000 ;
      RECT 3.255000  0.465000 3.425000 0.885000 ;
      RECT 4.095000  0.465000 4.425000 0.905000 ;
      RECT 4.095000  1.445000 4.425000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_2
END LIBRARY

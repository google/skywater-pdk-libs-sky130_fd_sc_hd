* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
M1000 X a_311_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=5.5025e+11p ps=6.15e+06u
M1001 a_561_297# B a_489_297# VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1002 X a_311_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=5.41725e+11p ps=5.32e+06u
M1003 a_311_413# a_205_93# VGND VNB nshort w=420000u l=150000u
+  ad=2.331e+11p pd=2.79e+06u as=0p ps=0u
M1004 a_489_297# a_27_410# a_393_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.43e+11p ps=2.66e+06u
M1005 a_393_413# a_205_93# a_311_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1006 VGND a_27_410# a_311_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_311_413# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1009 a_205_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1010 VGND A a_311_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C_N a_27_410# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1012 VPWR A a_561_297# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_205_93# D_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__einvn_0.pex.spice
* Created: Tue Sep  1 19:07:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVN_0%A_30_47# 1 2 9 13 17 19 20 21 22 26 30
c61 21 0 1.7629e-19 $X=0.82 $Y=1.98
c62 19 0 1.46566e-19 $X=0.82 $Y=0.74
r63 27 30 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.905 $Y=1.16 $X2=1
+ $Y2=1.16
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.16 $X2=0.905 $Y2=1.16
r65 24 26 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.905 $Y=1.895
+ $X2=0.905 $Y2=1.16
r66 23 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.905 $Y=0.825
+ $X2=0.905 $Y2=1.16
r67 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=1.98
+ $X2=0.905 $Y2=1.895
r68 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.82 $Y=1.98 $X2=0.4
+ $Y2=1.98
r69 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=0.74
+ $X2=0.905 $Y2=0.825
r70 19 20 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.82 $Y=0.74
+ $X2=0.36 $Y2=0.74
r71 15 22 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=0.242 $Y=2.065
+ $X2=0.4 $Y2=1.98
r72 15 17 7.68295 $w=3.13e-07 $l=2.1e-07 $layer=LI1_cond $X=0.242 $Y=2.065
+ $X2=0.242 $Y2=2.275
r73 11 20 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=0.222 $Y=0.655
+ $X2=0.36 $Y2=0.74
r74 11 13 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=0.222 $Y=0.655
+ $X2=0.222 $Y2=0.445
r75 7 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=1.16
r76 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=0.445
r77 2 17 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.065 $X2=0.275 $Y2=2.275
r78 1 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_0%TE_B 3 6 9 11 13 15 16 17 18 22 23
c45 22 0 2.97245e-20 $X=0.425 $Y=1.16
r46 22 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.16
+ $X2=0.425 $Y2=1.325
r47 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.16
+ $X2=0.425 $Y2=0.995
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.425
+ $Y=1.16 $X2=0.425 $Y2=1.16
r49 17 18 7.19764 $w=5.63e-07 $l=3.4e-07 $layer=LI1_cond $X=0.367 $Y=1.19
+ $X2=0.367 $Y2=1.53
r50 17 23 0.635086 $w=5.63e-07 $l=3e-08 $layer=LI1_cond $X=0.367 $Y=1.19
+ $X2=0.367 $Y2=1.16
r51 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1 $Y=1.77 $X2=1
+ $Y2=2.165
r52 12 16 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.56 $Y=1.695
+ $X2=0.485 $Y2=1.695
r53 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=1.695
+ $X2=1 $Y2=1.77
r54 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.925 $Y=1.695
+ $X2=0.56 $Y2=1.695
r55 7 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.485 $Y=1.77
+ $X2=0.485 $Y2=1.695
r56 7 9 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.485 $Y=1.77
+ $X2=0.485 $Y2=2.275
r57 6 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.485 $Y=1.62
+ $X2=0.485 $Y2=1.695
r58 6 25 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.485 $Y=1.62
+ $X2=0.485 $Y2=1.325
r59 3 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.485 $Y=0.445
+ $X2=0.485 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_0%A 3 7 9 10 11 12 20
c27 7 0 1.46566e-19 $X=1.36 $Y=2.165
c28 3 0 1.46566e-19 $X=1.36 $Y=0.445
r29 17 20 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.36 $Y=1.16
+ $X2=1.585 $Y2=1.16
r30 11 12 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=1.627 $Y=1.53
+ $X2=1.627 $Y2=1.87
r31 10 11 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.627 $Y=1.16
+ $X2=1.627 $Y2=1.53
r32 10 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.16 $X2=1.585 $Y2=1.16
r33 9 10 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=1.627 $Y=0.85
+ $X2=1.627 $Y2=1.16
r34 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.16
r35 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.36 $Y=1.325 $X2=1.36
+ $Y2=2.165
r36 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=1.16
r37 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.36 $Y=0.995 $X2=1.36
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_0%VPWR 1 4 6 13 14 17
r28 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r29 17 20 9.87808 $w=4.18e-07 $l=3.6e-07 $layer=LI1_cond $X=0.78 $Y=2.36
+ $X2=0.78 $Y2=2.72
r30 14 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r32 11 20 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=0.78
+ $Y2=2.72
r33 11 13 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.99 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 6 20 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.57 $Y=2.72 $X2=0.78
+ $Y2=2.72
r35 6 8 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=2.72 $X2=0.23
+ $Y2=2.72
r36 4 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r37 4 8 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r38 1 17 600 $w=1.7e-07 $l=3.76298e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=2.065 $X2=0.745 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_0%Z 1 2 8 9 10
r33 20 23 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=1.245 $Y=2.295
+ $X2=1.57 $Y2=2.295
r34 13 16 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=1.245 $Y=0.425
+ $X2=1.57 $Y2=0.425
r35 10 23 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=1.61 $Y=2.295 $X2=1.57
+ $Y2=2.295
r36 9 16 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=1.61 $Y=0.425 $X2=1.57
+ $Y2=0.425
r37 8 20 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.245 $Y=2.125
+ $X2=1.245 $Y2=2.295
r38 7 13 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.245 $Y=0.595
+ $X2=1.245 $Y2=0.425
r39 7 8 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=1.245 $Y=0.595
+ $X2=1.245 $Y2=2.125
r40 2 23 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.845 $X2=1.57 $Y2=2.3
r41 1 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.57 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_0%VGND 1 4 6 13 14 18
r26 18 21 9.36061 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.76
+ $Y2=0.36
r27 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r28 14 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r29 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r30 11 18 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.76
+ $Y2=0
r31 11 13 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.61
+ $Y2=0
r32 6 18 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.76
+ $Y2=0
r33 6 8 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.23 $Y2=0
r34 4 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r35 4 8 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r36 1 21 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.74 $Y2=0.36
.ends


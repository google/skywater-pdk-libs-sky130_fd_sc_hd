* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=1.635e+12p ps=1.527e+07u
M1001 a_478_47# A2 a_730_47# VNB nshort w=650000u l=150000u
+  ad=5.2e+11p pd=5.5e+06u as=4.16e+11p ps=3.88e+06u
M1002 a_27_297# B2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.035e+12p ps=1.007e+07u
M1004 a_730_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.4925e+11p ps=5.59e+06u
M1005 a_730_47# A2 a_478_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=0p ps=0u
M1007 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.51e+11p ps=3.68e+06u
M1009 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_478_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A3 a_730_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_478_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__a21boi_2.spice
* Created: Thu Aug 27 14:00:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21boi_2.spice.pex"
.subckt sky130_fd_sc_hd__a21boi_2  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B1_N_M1001_g N_A_61_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.143762 AS=0.126 PD=0.973458 PS=1.44 NRD=60.708 NRS=9.996 M=1 R=2.8
+ SA=75000.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1001_d N_A_61_47#_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.222488 AS=0.08775 PD=1.50654 PS=0.92 NRD=18.456 NRS=0 M=1 R=4.33333
+ SA=75000.8 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_61_47#_M1008_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1004 A_637_47# N_A2_M1004_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.10725 PD=0.86 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.7 SB=75001.4
+ A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g A_637_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.06825 PD=0.93 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002 SB=75001.1
+ A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1003_d N_A1_M1010_g A_479_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75002.5 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1013 A_479_47# N_A2_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.18525 PD=0.93 PS=1.87 NRD=15.684 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_61_47#_M1011_d N_B1_N_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_217_297#_M1009_d N_A_61_47#_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1012 N_A_217_297#_M1012_d N_A_61_47#_M1012_g N_Y_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1002 N_A_217_297#_M1012_d N_A2_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1002_s N_A1_M1000_g N_A_217_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.14 PD=1.27 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_217_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_A_217_297#_M1006_d N_A2_M1006_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_38 VNB 0 5.44765e-20 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__a21boi_2.spice.SKY130_FD_SC_HD__A21BOI_2.pxi"
*
.ends
*
*

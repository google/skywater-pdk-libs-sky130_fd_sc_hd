* File: sky130_fd_sc_hd__or4_2.pex.spice
* Created: Tue Sep  1 19:28:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4_2%D 3 7 9 10 17
c28 9 0 1.84467e-19 $X=0.235 $Y=0.85
r29 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r31 9 10 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.262 $Y=0.85
+ $X2=0.262 $Y2=1.16
r32 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r34 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%C 3 7 9 11 18
r38 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=1.325
r39 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r41 11 19 5.11227 $w=6.18e-07 $l=2.65e-07 $layer=LI1_cond $X=1.155 $Y=1.305
+ $X2=0.89 $Y2=1.305
r42 9 19 3.76186 $w=6.18e-07 $l=1.95e-07 $layer=LI1_cond $X=0.695 $Y=1.305
+ $X2=0.89 $Y2=1.305
r43 7 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.95 $Y=1.695
+ $X2=0.95 $Y2=1.325
r44 3 20 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.95 $Y=0.475
+ $X2=0.95 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%B 4 7 8 9 10 11 12 17 18
c39 17 0 1.73735e-19 $X=1.37 $Y=2.28
r40 17 19 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.37 $Y=2.28
+ $X2=1.37 $Y2=2.145
r41 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=2.28 $X2=1.37 $Y2=2.28
r42 12 18 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.155 $Y=2.27
+ $X2=1.37 $Y2=2.27
r43 11 12 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=2.27
+ $X2=1.155 $Y2=2.27
r44 10 11 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=2.27
+ $X2=0.695 $Y2=2.27
r45 8 9 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.34 $Y=0.76 $X2=1.34
+ $Y2=0.91
r46 7 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.37 $Y=0.475 $X2=1.37
+ $Y2=0.76
r47 4 19 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.31 $Y=1.695
+ $X2=1.31 $Y2=2.145
r48 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.31 $Y=1.695
+ $X2=1.31 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%A 3 7 9 12 13
r42 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.16
+ $X2=1.775 $Y2=1.325
r43 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.16
+ $X2=1.775 $Y2=0.995
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.775
+ $Y=1.16 $X2=1.775 $Y2=1.16
r45 9 13 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.775 $Y2=1.16
r46 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.79 $Y=1.695
+ $X2=1.79 $Y2=1.325
r47 3 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.79 $Y=0.475
+ $X2=1.79 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%A_27_297# 1 2 3 10 12 15 17 19 22 24 28 30 31
+ 34 36 38 43 45 49 50 55 57 62
c116 55 0 1.14153e-19 $X=2.255 $Y=1.16
c117 50 0 1.73735e-19 $X=1.595 $Y=1.58
c118 43 0 1.06604e-19 $X=2.15 $Y=1.495
c119 36 0 2.82207e-20 $X=2.065 $Y=0.74
r120 61 62 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.28 $Y=1.16
+ $X2=2.7 $Y2=1.16
r121 56 61 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.28 $Y2=1.16
r122 55 58 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.202 $Y=1.16
+ $X2=2.202 $Y2=1.325
r123 55 57 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.202 $Y=1.16
+ $X2=2.202 $Y2=0.995
r124 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=1.16 $X2=2.255 $Y2=1.16
r125 50 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.595 $Y=1.58
+ $X2=1.595 $Y2=1.87
r126 45 47 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=0.247 $Y=1.685
+ $X2=0.247 $Y2=1.87
r127 43 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=1.495
+ $X2=2.15 $Y2=1.325
r128 40 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=0.825
+ $X2=2.15 $Y2=0.995
r129 39 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.58
+ $X2=1.595 $Y2=1.58
r130 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=1.58
+ $X2=2.15 $Y2=1.495
r131 38 39 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=1.58
+ $X2=1.68 $Y2=1.58
r132 37 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.74
+ $X2=1.58 $Y2=0.74
r133 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=0.74
+ $X2=2.15 $Y2=0.825
r134 36 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.065 $Y=0.74
+ $X2=1.665 $Y2=0.74
r135 32 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.655
+ $X2=1.58 $Y2=0.74
r136 32 34 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.58 $Y=0.655
+ $X2=1.58 $Y2=0.47
r137 30 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=0.74
+ $X2=1.58 $Y2=0.74
r138 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.495 $Y=0.74
+ $X2=0.795 $Y2=0.74
r139 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=0.655
+ $X2=0.795 $Y2=0.74
r140 26 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.71 $Y=0.655
+ $X2=0.71 $Y2=0.47
r141 25 47 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.41 $Y=1.87
+ $X2=0.247 $Y2=1.87
r142 24 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=1.87
+ $X2=1.595 $Y2=1.87
r143 24 25 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=1.51 $Y=1.87
+ $X2=0.41 $Y2=1.87
r144 20 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.16
r145 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.985
r146 17 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=1.16
r147 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=0.56
r148 13 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.325
+ $X2=2.28 $Y2=1.16
r149 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.28 $Y=1.325
+ $X2=2.28 $Y2=1.985
r150 10 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=0.995
+ $X2=2.28 $Y2=1.16
r151 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.28 $Y=0.995
+ $X2=2.28 $Y2=0.56
r152 3 45 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.685
r153 2 34 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.265 $X2=1.58 $Y2=0.47
r154 1 28 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=0.71 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%VPWR 1 2 9 11 13 17 19 27 33 37
c33 1 0 1.06604e-19 $X=1.865 $Y=1.485
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r37 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 28 33 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.055 $Y2=2.72
r40 28 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 27 36 3.40825 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.85 $Y=2.72
+ $X2=3.035 $Y2=2.72
r42 27 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.85 $Y=2.72 $X2=2.53
+ $Y2=2.72
r43 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r45 21 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r46 19 33 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.055 $Y2=2.72
r47 19 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 17 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 17 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r50 13 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.935 $Y=1.66
+ $X2=2.935 $Y2=2.34
r51 11 36 3.40825 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.935 $Y=2.635
+ $X2=3.035 $Y2=2.72
r52 11 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=2.635
+ $X2=2.935 $Y2=2.34
r53 7 33 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.72
r54 7 9 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2
r55 2 16 400 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.485 $X2=2.935 $Y2=2.34
r56 2 13 400 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.485 $X2=2.935 $Y2=1.66
r57 1 9 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.485 $X2=2.065 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%X 1 2 12 14 15 16
r25 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=2.542 $Y=1.632
+ $X2=2.542 $Y2=1.845
r26 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.542 $Y=1.632
+ $X2=2.542 $Y2=1.495
r27 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=2.49 $Y=0.587
+ $X2=2.595 $Y2=0.587
r28 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.595 $Y=0.76
+ $X2=2.595 $Y2=0.587
r29 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.595 $Y=0.76
+ $X2=2.595 $Y2=1.495
r30 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=1.485 $X2=2.49 $Y2=1.845
r31 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.49 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_2%VGND 1 2 3 4 13 15 19 23 25 27 29 31 36 41 50
+ 53 57
c63 31 0 1.84467e-19 $X=0.995 $Y=0
c64 27 0 2.82207e-20 $X=2.935 $Y=0.4
r65 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r66 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r67 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r68 45 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r69 45 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r70 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r71 42 53 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.025
+ $Y2=0
r72 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.53
+ $Y2=0
r73 41 56 3.40825 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.035
+ $Y2=0
r74 41 44 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.53
+ $Y2=0
r75 40 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r76 40 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r77 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r78 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.16
+ $Y2=0
r79 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.61
+ $Y2=0
r80 36 53 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.025
+ $Y2=0
r81 36 39 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.61
+ $Y2=0
r82 35 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r83 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r84 32 47 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r85 32 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r86 31 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.16
+ $Y2=0
r87 31 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.69
+ $Y2=0
r88 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r89 29 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r90 25 56 3.40825 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.935 $Y=0.085
+ $X2=3.035 $Y2=0
r91 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.935 $Y=0.085
+ $X2=2.935 $Y2=0.4
r92 21 53 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r93 21 23 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.4
r94 17 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0
r95 17 19 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0.4
r96 13 47 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r97 13 15 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.5
r98 4 27 91 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.235 $X2=2.935 $Y2=0.4
r99 3 23 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.265 $X2=2.05 $Y2=0.4
r100 2 19 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.265 $X2=1.16 $Y2=0.4
r101 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__clkdlybuf4s18_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.055000 0.550000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.255000 3.590000 0.545000 ;
        RECT 3.220000 1.760000 3.590000 2.465000 ;
        RECT 3.365000 0.545000 3.590000 1.760000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.595000  0.085000 0.910000 0.545000 ;
        RECT 2.710000  0.085000 3.040000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.595000 1.835000 0.925000 2.635000 ;
        RECT 2.710000 1.760000 3.040000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.255000 0.425000 0.715000 ;
      RECT 0.095000 0.715000 1.215000 0.885000 ;
      RECT 0.095000 1.495000 1.215000 1.665000 ;
      RECT 0.095000 1.665000 0.425000 2.465000 ;
      RECT 0.720000 0.885000 1.215000 1.495000 ;
      RECT 1.385000 0.255000 1.760000 0.825000 ;
      RECT 1.385000 1.835000 1.760000 2.465000 ;
      RECT 1.590000 0.825000 1.760000 1.055000 ;
      RECT 1.590000 1.055000 2.685000 1.250000 ;
      RECT 1.590000 1.250000 1.760000 1.835000 ;
      RECT 1.930000 0.255000 2.260000 0.715000 ;
      RECT 1.930000 0.715000 3.195000 0.885000 ;
      RECT 1.930000 1.420000 3.195000 1.590000 ;
      RECT 1.930000 1.590000 2.260000 2.465000 ;
      RECT 2.855000 0.885000 3.195000 1.420000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_1

* File: sky130_fd_sc_hd__o211a_2.spice
* Created: Thu Aug 27 14:34:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o211a_2.pex.spice"
.subckt sky130_fd_sc_hd__o211a_2  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1003 A_110_47# N_C1_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.17225 PD=0.86 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1000 N_A_182_47#_M1000_d N_B1_M1000_g A_110_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.16535 AS=0.06825 PD=1.82 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_182_47#_M1002_d N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.16535 PD=0.93 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_182_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.091 PD=0.97 PS=0.93 NRD=3.684 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1005_d N_A_27_47#_M1005_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.104 PD=0.93 PS=0.97 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1005_d N_A_27_47#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.23075 PD=0.93 PS=2.01 NRD=0 NRS=12.912 M=1 R=4.33333 SA=75001.5
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_47#_M1011_d N_B1_M1011_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.3675 AS=0.14 PD=1.735 PS=1.28 NRD=13.7703 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1007 A_373_297# N_A2_M1007_g N_A_27_47#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.3675 PD=1.21 PS=1.735 NRD=9.8303 NRS=8.8453 M=1 R=6.66667
+ SA=75001.5 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_373_297# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.105 PD=1.39 PS=1.21 NRD=9.8303 NRS=9.8303 M=1 R=6.66667 SA=75001.9
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.195 PD=1.28 PS=1.39 NRD=0 NRS=11.8003 M=1 R=6.66667 SA=75002.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1001_d N_A_27_47#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_63 VPB 0 1.13771e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__o211a_2.pxi.spice"
*
.ends
*
*

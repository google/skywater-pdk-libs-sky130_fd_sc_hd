* File: sky130_fd_sc_hd__buf_2.pex.spice
* Created: Tue Sep  1 18:59:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUF_2%A 3 7 9 15
c31 9 0 3.26313e-20 $X=0.23 $Y=1.19
r32 12 15 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.27 $Y=1.16 $X2=0.47
+ $Y2=1.16
r33 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r34 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r35 5 7 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.125
r36 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r37 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_2%A_27_47# 1 2 7 9 12 14 16 19 23 27 29 30 31 32
+ 36 38 40 45
c78 38 0 1.42894e-19 $X=0.89 $Y=1.16
c79 12 0 2.53799e-20 $X=0.945 $Y=1.985
c80 7 0 7.25139e-21 $X=0.945 $Y=0.995
r81 44 45 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.945 $Y=1.16
+ $X2=1.365 $Y2=1.16
r82 39 44 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.945 $Y2=1.16
r83 38 41 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.847 $Y=1.16
+ $X2=0.847 $Y2=1.325
r84 38 40 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.847 $Y=1.16
+ $X2=0.847 $Y2=0.995
r85 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r86 36 41 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.805 $Y=1.535
+ $X2=0.805 $Y2=1.325
r87 33 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.805 $Y=0.805
+ $X2=0.805 $Y2=0.995
r88 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.62
+ $X2=0.805 $Y2=1.535
r89 31 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.72 $Y=1.62
+ $X2=0.345 $Y2=1.62
r90 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=0.72
+ $X2=0.805 $Y2=0.805
r91 29 30 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.72 $Y=0.72
+ $X2=0.345 $Y2=0.72
r92 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.705
+ $X2=0.345 $Y2=1.62
r93 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=1.705
+ $X2=0.26 $Y2=1.96
r94 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r95 21 23 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.445
r96 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.16
r97 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.985
r98 14 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=1.16
r99 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=0.56
r100 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.325
+ $X2=0.945 $Y2=1.16
r101 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.945 $Y=1.325
+ $X2=0.945 $Y2=1.985
r102 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=1.16
r103 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r104 2 27 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.805 $X2=0.26 $Y2=1.96
r105 1 23 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_2%VPWR 1 2 9 11 13 17 19 21 27 33 37
r29 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r32 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 28 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=2.72
+ $X2=0.725 $Y2=2.72
r35 28 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.89 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 27 36 4.13816 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.49 $Y=2.72
+ $X2=1.665 $Y2=2.72
r37 27 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.49 $Y=2.72
+ $X2=1.15 $Y2=2.72
r38 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=2.72
+ $X2=0.725 $Y2=2.72
r39 19 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 17 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.56 $Y2=2.72
r41 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r42 13 16 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.62 $Y=1.66
+ $X2=1.62 $Y2=2.34
r43 11 36 3.07406 $w=2.6e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.665 $Y2=2.72
r44 11 16 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.34
r45 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2.72
r46 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=1.96
r47 2 16 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.485 $X2=1.575 $Y2=2.34
r48 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.485 $X2=1.575 $Y2=1.66
r49 1 9 300 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.805 $X2=0.725 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_2%X 1 2 10 11 12 13 14 15
r24 14 15 17.8516 $w=2.53e-07 $l=3.95e-07 $layer=LI1_cond $X=1.187 $Y=1.815
+ $X2=1.187 $Y2=2.21
r25 11 14 5.78481 $w=2.53e-07 $l=1.28e-07 $layer=LI1_cond $X=1.187 $Y=1.687
+ $X2=1.187 $Y2=1.815
r26 11 12 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=1.187 $Y=1.687
+ $X2=1.187 $Y2=1.56
r27 10 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.23 $Y=0.83
+ $X2=1.23 $Y2=1.56
r28 9 13 8.72241 $w=2.53e-07 $l=1.93e-07 $layer=LI1_cond $X=1.187 $Y=0.703
+ $X2=1.187 $Y2=0.51
r29 9 10 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=1.187 $Y=0.703
+ $X2=1.187 $Y2=0.83
r30 2 14 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.485 $X2=1.155 $Y2=1.815
r31 1 13 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_2%VGND 1 2 9 11 13 15 17 19 25 31 35
r31 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r32 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r33 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r34 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r35 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r36 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.725
+ $Y2=0
r37 26 28 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.15
+ $Y2=0
r38 25 34 4.13816 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.665
+ $Y2=0
r39 25 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.15
+ $Y2=0
r40 19 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.725
+ $Y2=0
r41 17 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r42 15 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.56
+ $Y2=0
r43 15 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r44 11 34 3.07406 $w=2.6e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.665 $Y2=0
r45 11 13 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.4
r46 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r47 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.38
r48 2 13 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.44
+ $Y=0.235 $X2=1.575 $Y2=0.4
r49 1 9 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.725 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o32ai_1.pex.spice
* Created: Thu Aug 27 14:41:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O32AI_1%B1 1 3 6 8 9 16
r29 13 16 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 9 23 7.09132 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.225 $Y=1.16
+ $X2=0.225 $Y2=0.995
r31 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r32 8 23 6.55311 $w=2.53e-07 $l=1.45e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=0.995
r33 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r34 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r35 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%B2 1 3 5 7 8
c37 5 0 8.66312e-20 $X=0.945 $Y=0.995
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=1.16 $X2=0.955 $Y2=1.16
r39 8 12 3.85832 $w=6.18e-07 $l=2e-07 $layer=LI1_cond $X=1.155 $Y=1.305
+ $X2=0.955 $Y2=1.305
r40 5 11 38.8702 $w=3.57e-07 $l=1.68953e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.937 $Y2=1.16
r41 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r42 1 11 38.8702 $w=3.57e-07 $l=2.11849e-07 $layer=POLY_cond $X=0.83 $Y=1.325
+ $X2=0.937 $Y2=1.16
r43 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.83 $Y=1.325 $X2=0.83
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%A3 1 3 6 8 12
r37 12 14 13.9604 $w=3.28e-07 $l=9.5e-08 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.59 $Y2=1.16
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r39 10 12 13.2256 $w=3.28e-07 $l=9e-08 $layer=POLY_cond $X=1.405 $Y=1.16
+ $X2=1.495 $Y2=1.16
r40 8 13 2.31499 $w=6.18e-07 $l=1.2e-07 $layer=LI1_cond $X=1.615 $Y=1.305
+ $X2=1.495 $Y2=1.305
r41 4 14 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.325
+ $X2=1.59 $Y2=1.16
r42 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.59 $Y=1.325 $X2=1.59
+ $Y2=1.985
r43 1 10 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=0.995
+ $X2=1.405 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.405 $Y=0.995
+ $X2=1.405 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%A2 3 6 8 9 10 11 17 19
r36 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.16
+ $X2=2.14 $Y2=1.325
r37 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.16
+ $X2=2.14 $Y2=0.995
r38 10 11 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.077 $Y=1.87
+ $X2=2.077 $Y2=2.21
r39 9 10 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.077 $Y=1.53
+ $X2=2.077 $Y2=1.87
r40 8 9 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.077 $Y=1.16
+ $X2=2.077 $Y2=1.53
r41 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r42 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.23 $Y=1.985
+ $X2=2.23 $Y2=1.325
r43 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.23 $Y=0.56 $X2=2.23
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%A1 3 6 8 11 13
r23 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.16
+ $X2=2.74 $Y2=1.325
r24 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.16
+ $X2=2.74 $Y2=0.995
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.16 $X2=2.74 $Y2=1.16
r26 8 12 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=2.74 $Y2=1.16
r27 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.65 $Y=1.985
+ $X2=2.65 $Y2=1.325
r28 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.65 $Y=0.56 $X2=2.65
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%VPWR 1 2 7 9 13 15 19 21 34
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r36 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r37 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 25 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 24 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r40 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 22 30 4.22982 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=2.72 $X2=0.18
+ $Y2=2.72
r42 22 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.36 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 21 33 5.87207 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.957 $Y2=2.72
r44 21 27 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 19 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 19 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 15 18 17.8105 $w=4.38e-07 $l=6.8e-07 $layer=LI1_cond $X=2.915 $Y=1.66
+ $X2=2.915 $Y2=2.34
r48 13 33 2.84639 $w=4.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.915 $Y=2.635
+ $X2=2.957 $Y2=2.72
r49 13 18 7.72661 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.915 $Y=2.635
+ $X2=2.915 $Y2=2.34
r50 9 12 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.225 $Y=1.66
+ $X2=0.225 $Y2=2.34
r51 7 30 3.05487 $w=2.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.18 $Y2=2.72
r52 7 12 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.225 $Y2=2.34
r53 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=1.485 $X2=2.86 $Y2=2.34
r54 2 15 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=1.485 $X2=2.86 $Y2=1.66
r55 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r56 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%Y 1 2 10 12 14 29
r31 14 29 3.95761 $w=6.78e-07 $l=2.25e-07 $layer=LI1_cond $X=1.155 $Y=2.125
+ $X2=1.38 $Y2=2.125
r32 12 23 2.13119 $w=6.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.615 $Y=2.125
+ $X2=0.7 $Y2=2.125
r33 12 14 7.2996 $w=6.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.74 $Y=2.125
+ $X2=1.155 $Y2=2.125
r34 12 23 0.703576 $w=6.78e-07 $l=4e-08 $layer=LI1_cond $X=0.74 $Y=2.125 $X2=0.7
+ $Y2=2.125
r35 8 12 43.7938 $w=2.58e-07 $l=9.6e-07 $layer=LI1_cond $X=0.615 $Y=0.825
+ $X2=0.615 $Y2=1.785
r36 8 10 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.615 $Y=0.825
+ $X2=0.615 $Y2=0.74
r37 2 29 150 $w=1.7e-07 $l=7.14038e-07 $layer=licon1_PDIFF $count=4 $X=0.905
+ $Y=1.485 $X2=1.38 $Y2=2
r38 1 10 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%A_27_47# 1 2 3 10 14 15 16 17 20
c38 14 0 8.66312e-20 $X=1.18 $Y=0.485
r39 18 20 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.44 $Y=0.655
+ $X2=2.44 $Y2=0.54
r40 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.355 $Y=0.74
+ $X2=2.44 $Y2=0.655
r41 16 17 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.355 $Y=0.74
+ $X2=1.345 $Y2=0.74
r42 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.18 $Y=0.655
+ $X2=1.345 $Y2=0.74
r43 14 23 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.18 $Y=0.485
+ $X2=1.18 $Y2=0.37
r44 14 15 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.18 $Y=0.485
+ $X2=1.18 $Y2=0.655
r45 10 23 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0.37
+ $X2=1.18 $Y2=0.37
r46 10 12 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.015 $Y=0.37
+ $X2=0.26 $Y2=0.37
r47 3 20 182 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.44 $Y2=0.54
r48 2 23 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.02
+ $Y=0.235 $X2=1.18 $Y2=0.38
r49 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_1%VGND 1 2 7 9 11 21 29 35 38
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r39 33 35 8.91182 $w=5.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.07 $Y=0.2
+ $X2=2.185 $Y2=0.2
r40 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r41 31 33 1.04919 $w=5.68e-07 $l=5e-08 $layer=LI1_cond $X=2.02 $Y=0.2 $X2=2.07
+ $Y2=0.2
r42 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r43 27 31 8.60337 $w=5.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.61 $Y=0.2 $X2=2.02
+ $Y2=0.2
r44 27 29 8.49214 $w=5.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=0.2
+ $X2=1.515 $Y2=0.2
r45 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r46 25 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r47 25 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r48 24 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.185
+ $Y2=0
r49 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 21 37 5.87207 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.957
+ $Y2=0
r51 21 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.53
+ $Y2=0
r52 20 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r53 19 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.515
+ $Y2=0
r54 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r55 15 19 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r56 11 20 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r57 11 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 7 37 2.84639 $w=4.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.957 $Y2=0
r59 7 9 7.72661 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.38
r60 2 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=0.235 $X2=2.86 $Y2=0.38
r61 1 31 91 $w=1.7e-07 $l=6.08194e-07 $layer=licon1_NDIFF $count=2 $X=1.48
+ $Y=0.235 $X2=2.02 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a31o_2.spice.SKY130_FD_SC_HD__A31O_2.pxi
* Created: Thu Aug 27 14:04:41 2020
* 
x_PM_SKY130_FD_SC_HD__A31O_2%A_79_21# N_A_79_21#_M1000_d N_A_79_21#_M1002_d
+ N_A_79_21#_c_59_n N_A_79_21#_M1005_g N_A_79_21#_M1003_g N_A_79_21#_c_60_n
+ N_A_79_21#_M1011_g N_A_79_21#_M1009_g N_A_79_21#_c_65_n N_A_79_21#_c_70_p
+ N_A_79_21#_c_119_p N_A_79_21#_c_61_n N_A_79_21#_c_97_p N_A_79_21#_c_74_p
+ N_A_79_21#_c_81_p N_A_79_21#_c_98_p N_A_79_21#_c_62_n
+ PM_SKY130_FD_SC_HD__A31O_2%A_79_21#
x_PM_SKY130_FD_SC_HD__A31O_2%A3 N_A3_c_147_n N_A3_M1008_g N_A3_M1001_g A3 A3
+ N_A3_c_149_n PM_SKY130_FD_SC_HD__A31O_2%A3
x_PM_SKY130_FD_SC_HD__A31O_2%A2 N_A2_M1007_g N_A2_M1010_g N_A2_c_186_n
+ N_A2_c_193_n N_A2_c_187_n N_A2_c_188_n A2 N_A2_c_189_n
+ PM_SKY130_FD_SC_HD__A31O_2%A2
x_PM_SKY130_FD_SC_HD__A31O_2%A1 N_A1_M1000_g N_A1_M1006_g N_A1_c_238_n
+ N_A1_c_239_n N_A1_c_251_n A1 N_A1_c_240_n PM_SKY130_FD_SC_HD__A31O_2%A1
x_PM_SKY130_FD_SC_HD__A31O_2%B1 N_B1_M1002_g N_B1_c_290_n N_B1_M1004_g B1 B1
+ N_B1_c_292_n PM_SKY130_FD_SC_HD__A31O_2%B1
x_PM_SKY130_FD_SC_HD__A31O_2%VPWR N_VPWR_M1003_d N_VPWR_M1009_d N_VPWR_M1010_d
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n VPWR N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_322_n
+ N_VPWR_c_332_n PM_SKY130_FD_SC_HD__A31O_2%VPWR
x_PM_SKY130_FD_SC_HD__A31O_2%X N_X_M1005_s N_X_M1003_s N_X_c_381_n N_X_c_391_n
+ N_X_c_411_p N_X_c_401_n X X X X N_X_c_383_n N_X_c_385_n
+ PM_SKY130_FD_SC_HD__A31O_2%X
x_PM_SKY130_FD_SC_HD__A31O_2%A_277_297# N_A_277_297#_M1001_d
+ N_A_277_297#_M1006_d N_A_277_297#_c_419_n N_A_277_297#_c_424_n
+ N_A_277_297#_c_420_n N_A_277_297#_c_421_n N_A_277_297#_c_439_n
+ PM_SKY130_FD_SC_HD__A31O_2%A_277_297#
x_PM_SKY130_FD_SC_HD__A31O_2%VGND N_VGND_M1005_d N_VGND_M1011_d N_VGND_M1004_d
+ N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ VGND N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n
+ PM_SKY130_FD_SC_HD__A31O_2%VGND
cc_1 VNB N_A_79_21#_c_59_n 0.0191079f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_60_n 0.0160515f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_61_n 0.00256351f $X=-0.19 $Y=-0.24 $X2=2.62 $Y2=1.495
cc_4 VNB N_A_79_21#_c_62_n 0.0336216f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_A3_c_147_n 0.0154361f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.235
cc_6 VNB A3 0.0036805f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_A3_c_149_n 0.0217003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_186_n 0.00139769f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_9 VNB N_A2_c_187_n 0.00403204f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_10 VNB N_A2_c_188_n 0.022485f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_11 VNB N_A2_c_189_n 0.0163571f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.245
cc_12 VNB N_A1_c_238_n 7.27863e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_13 VNB N_A1_c_239_n 0.0230678f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_14 VNB N_A1_c_240_n 0.0173926f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.245
cc_15 VNB N_B1_c_290_n 0.0198027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB B1 0.00904727f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_17 VNB N_B1_c_292_n 0.0472781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_18 VNB N_VPWR_c_322_n 0.136896f $X=-0.19 $Y=-0.24 $X2=2.62 $Y2=1.58
cc_19 VNB N_X_c_381_n 0.00119493f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB X 0.021429f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_21 VNB N_X_c_383_n 0.00758104f $X=-0.19 $Y=-0.24 $X2=2.96 $Y2=1.96
cc_22 VNB N_VGND_c_441_n 0.00994884f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_23 VNB N_VGND_c_442_n 0.0166098f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_24 VNB N_VGND_c_443_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_25 VNB N_VGND_c_444_n 0.00988261f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_26 VNB N_VGND_c_445_n 0.0187519f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_27 VNB N_VGND_c_446_n 0.0157645f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.58
cc_28 VNB N_VGND_c_447_n 0.0426414f $X=-0.19 $Y=-0.24 $X2=2.96 $Y2=1.96
cc_29 VNB N_VGND_c_448_n 0.00438976f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_30 VNB N_VGND_c_449_n 0.179359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_A_79_21#_M1003_g 0.0218284f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_32 VPB N_A_79_21#_M1009_g 0.0185209f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_33 VPB N_A_79_21#_c_65_n 0.0024477f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.495
cc_34 VPB N_A_79_21#_c_61_n 0.00175326f $X=-0.19 $Y=1.305 $X2=2.62 $Y2=1.495
cc_35 VPB N_A_79_21#_c_62_n 0.00457736f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_36 VPB N_A3_M1001_g 0.0191621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A3 0.00183392f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_38 VPB N_A3_c_149_n 0.00431904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A2_M1010_g 0.019823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A2_c_188_n 0.00413452f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_41 VPB N_A1_M1006_g 0.0202773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A1_c_238_n 6.43507e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_43 VPB N_A1_c_239_n 0.00444023f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_B1_M1002_g 0.0260335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB B1 0.00313953f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_46 VPB N_B1_c_292_n 0.0124317f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_47 VPB N_VPWR_c_323_n 0.011108f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_48 VPB N_VPWR_c_324_n 0.00451022f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_49 VPB N_VPWR_c_325_n 0.00166889f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_50 VPB N_VPWR_c_326_n 0.00234028f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_327_n 0.0140067f $X=-0.19 $Y=1.305 $X2=2.535 $Y2=1.58
cc_52 VPB N_VPWR_c_328_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.58
cc_53 VPB N_VPWR_c_329_n 0.0170221f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.16
cc_54 VPB N_VPWR_c_330_n 0.0305977f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=0.42
cc_55 VPB N_VPWR_c_322_n 0.0452754f $X=-0.19 $Y=1.305 $X2=2.62 $Y2=1.58
cc_56 VPB N_VPWR_c_332_n 0.00519461f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_57 VPB X 0.022467f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_58 VPB N_X_c_385_n 0.00784216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_60_n N_A3_c_147_n 0.0242109f $X=0.89 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_60 N_A_79_21#_M1009_g N_A3_M1001_g 0.0300229f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_70_p N_A3_M1001_g 0.0139369f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_60_n A3 0.00765163f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_65_n A3 0.00362039f $X=0.64 $Y=1.495 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_70_p A3 0.0228278f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_74_p A3 0.0128542f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_70_p N_A3_c_149_n 0.00136195f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_62_n N_A3_c_149_n 0.0212612f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_70_p N_A2_M1010_g 0.0110022f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_70_p N_A2_c_193_n 0.00186086f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_70_p N_A2_c_187_n 0.015782f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_70_p N_A2_c_188_n 0.0026229f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_81_p A2 3.71082e-19 $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_70_p N_A1_M1006_g 0.0116745f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_61_n N_A1_M1006_g 0.00326588f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_70_p N_A1_c_238_n 0.0104659f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_61_n N_A1_c_238_n 0.031608f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_70_p N_A1_c_239_n 0.00226733f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_61_n N_A1_c_239_n 0.00187856f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_81_p N_A1_c_239_n 8.07307e-19 $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_80 N_A_79_21#_M1000_d N_A1_c_251_n 0.00183052f $X=2.285 $Y=0.235 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_70_p N_A1_c_251_n 0.0042936f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_61_n N_A1_c_251_n 0.0125242f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_61_n A1 0.00779435f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_81_p A1 0.0059919f $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_61_n N_A1_c_240_n 0.00234585f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_81_p N_A1_c_240_n 0.00464315f $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_61_n N_B1_M1002_g 0.00910921f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_97_p N_B1_M1002_g 0.00792476f $X=2.96 $Y=1.96 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_98_p N_B1_M1002_g 0.0166342f $X=2.96 $Y=1.58 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_61_n N_B1_c_290_n 0.014726f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_81_p N_B1_c_290_n 0.00300781f $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_61_n B1 0.0364324f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_98_p B1 0.011545f $X=2.96 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_61_n N_B1_c_292_n 0.0102911f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_98_p N_B1_c_292_n 0.00521959f $X=2.96 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_70_p N_VPWR_M1009_d 0.00446832f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_70_p N_VPWR_M1010_d 0.00597469f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_79_21#_M1003_g N_VPWR_c_324_n 0.00332648f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_79_21#_M1003_g N_VPWR_c_325_n 7.226e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_79_21#_M1009_g N_VPWR_c_325_n 0.0107351f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_70_p N_VPWR_c_325_n 0.0148589f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_79_21#_M1003_g N_VPWR_c_327_n 0.00436487f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_M1009_g N_VPWR_c_327_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_97_p N_VPWR_c_330_n 0.0118139f $X=2.96 $Y=1.96 $X2=0 $Y2=0
cc_105 N_A_79_21#_M1002_d N_VPWR_c_322_n 0.00782714f $X=2.765 $Y=1.485 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_M1003_g N_VPWR_c_322_n 0.006716f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_79_21#_M1009_g N_VPWR_c_322_n 0.00789179f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_79_21#_c_97_p N_VPWR_c_322_n 0.00646998f $X=2.96 $Y=1.96 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_70_p N_X_M1003_s 6.7956e-19 $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_119_p N_X_M1003_s 0.0016062f $X=0.725 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_59_n N_X_c_381_n 0.0176327f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_74_p N_X_c_381_n 0.0116632f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_62_n N_X_c_381_n 0.00227788f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_79_21#_M1003_g N_X_c_391_n 0.0176327f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_70_p N_X_c_391_n 0.00263167f $X=2.535 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_119_p N_X_c_391_n 0.010603f $X=0.725 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_62_n N_X_c_391_n 3.39427e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_59_n X 0.0261841f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_65_n X 0.0156892f $X=0.64 $Y=1.495 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_74_p X 0.0111625f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_70_p N_A_277_297#_M1001_d 0.00629077f $X=2.535 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_122 N_A_79_21#_c_70_p N_A_277_297#_M1006_d 0.00764319f $X=2.535 $Y=1.58 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_c_98_p N_A_277_297#_M1006_d 2.98916e-19 $X=2.96 $Y=1.58 $X2=0
+ $Y2=0
cc_124 N_A_79_21#_c_70_p N_A_277_297#_c_419_n 0.014764f $X=2.535 $Y=1.58 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_c_70_p N_A_277_297#_c_420_n 0.0359551f $X=2.535 $Y=1.58 $X2=0
+ $Y2=0
cc_126 N_A_79_21#_c_70_p N_A_277_297#_c_421_n 0.0193093f $X=2.535 $Y=1.58 $X2=0
+ $Y2=0
cc_127 N_A_79_21#_c_97_p N_A_277_297#_c_421_n 0.0105708f $X=2.96 $Y=1.96 $X2=0
+ $Y2=0
cc_128 N_A_79_21#_c_59_n N_VGND_c_442_n 0.00314466f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_59_n N_VGND_c_443_n 4.77885e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_60_n N_VGND_c_443_n 0.00606866f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_59_n N_VGND_c_446_n 0.00436487f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_60_n N_VGND_c_446_n 0.00544582f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_81_p N_VGND_c_447_n 0.0183725f $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_134 N_A_79_21#_M1000_d N_VGND_c_449_n 0.00416274f $X=2.285 $Y=0.235 $X2=0
+ $Y2=0
cc_135 N_A_79_21#_c_59_n N_VGND_c_449_n 0.00681636f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_60_n N_VGND_c_449_n 0.00912034f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_81_p N_VGND_c_449_n 0.0121681f $X=2.54 $Y=0.42 $X2=0 $Y2=0
cc_138 N_A3_M1001_g N_A2_M1010_g 0.028197f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A3_c_147_n N_A2_c_186_n 7.68589e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_140 A3 N_A2_c_186_n 0.00974947f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A3_c_149_n N_A2_c_186_n 4.53861e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A3_c_147_n N_A2_c_193_n 0.00222764f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_143 A3 N_A2_c_193_n 0.00557445f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_144 A3 N_A2_c_187_n 0.0117213f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A3_c_149_n N_A2_c_187_n 0.001136f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_146 A3 N_A2_c_188_n 6.99855e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A3_c_149_n N_A2_c_188_n 0.0206289f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A3_c_147_n A2 0.00422932f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A3_c_147_n N_A2_c_189_n 0.0399056f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_150 A3 N_A2_c_189_n 2.31086e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A3_M1001_g N_VPWR_c_325_n 0.0014671f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A3_M1001_g N_VPWR_c_329_n 0.00542953f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A3_M1001_g N_VPWR_c_322_n 0.0095987f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A3_M1001_g N_A_277_297#_c_419_n 0.00218411f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A3_M1001_g N_A_277_297#_c_424_n 0.00466005f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_156 A3 N_VGND_M1011_d 0.00263007f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A3_c_147_n N_VGND_c_443_n 0.010618f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_158 A3 N_VGND_c_443_n 0.00998502f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A3_c_147_n N_VGND_c_447_n 0.00388479f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A3_c_147_n N_VGND_c_449_n 0.0067649f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_161 A3 N_VGND_c_449_n 9.73992e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A2_M1010_g N_A1_M1006_g 0.0353864f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_c_186_n N_A1_c_238_n 0.00706888f $X=1.71 $Y=1.075 $X2=0 $Y2=0
cc_164 N_A2_c_187_n N_A1_c_238_n 0.0108115f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A2_c_188_n N_A1_c_238_n 9.21181e-19 $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A2_c_189_n N_A1_c_238_n 4.06098e-19 $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_c_187_n N_A1_c_239_n 0.00109547f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A2_c_188_n N_A1_c_239_n 0.0205795f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A2_c_193_n N_A1_c_251_n 0.0127437f $X=1.71 $Y=0.78 $X2=0 $Y2=0
cc_170 N_A2_c_189_n N_A1_c_251_n 0.0012074f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_171 A2 A1 0.0142232f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_172 N_A2_c_189_n A1 0.00219906f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_186_n N_A1_c_240_n 6.73963e-19 $X=1.71 $Y=1.075 $X2=0 $Y2=0
cc_174 A2 N_A1_c_240_n 2.97717e-19 $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_175 N_A2_c_189_n N_A1_c_240_n 0.0312718f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A2_M1010_g N_VPWR_c_326_n 0.00192512f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1010_g N_VPWR_c_329_n 0.00436487f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_M1010_g N_VPWR_c_322_n 0.00605263f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_M1010_g N_A_277_297#_c_420_n 0.0103728f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_180 A2 N_VGND_c_443_n 0.00363701f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_181 N_A2_c_189_n N_VGND_c_443_n 0.00198722f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_193_n N_VGND_c_447_n 0.00138719f $X=1.71 $Y=0.78 $X2=0 $Y2=0
cc_183 A2 N_VGND_c_447_n 0.00481649f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_184 N_A2_c_189_n N_VGND_c_447_n 0.00429875f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A2_c_193_n N_VGND_c_449_n 0.00214628f $X=1.71 $Y=0.78 $X2=0 $Y2=0
cc_186 A2 N_VGND_c_449_n 0.00557356f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_187 N_A2_c_189_n N_VGND_c_449_n 0.00635939f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A2_c_193_n A_277_47# 0.0033894f $X=1.71 $Y=0.78 $X2=-0.19 $Y2=-0.24
cc_189 A2 A_277_47# 0.00426869f $X=1.53 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_190 N_A1_M1006_g N_B1_M1002_g 0.020739f $X=2.21 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A1_c_238_n N_B1_c_290_n 3.12997e-19 $X=2.27 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A1_c_251_n N_B1_c_290_n 4.82639e-19 $X=2.27 $Y=0.785 $X2=0 $Y2=0
cc_193 N_A1_c_240_n N_B1_c_290_n 0.0194383f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_238_n N_B1_c_292_n 3.26767e-19 $X=2.27 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A1_c_239_n N_B1_c_292_n 0.0202685f $X=2.27 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A1_M1006_g N_VPWR_c_326_n 0.0083152f $X=2.21 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A1_M1006_g N_VPWR_c_330_n 0.00406603f $X=2.21 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A1_M1006_g N_VPWR_c_322_n 0.00491662f $X=2.21 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A1_M1006_g N_A_277_297#_c_420_n 0.0102439f $X=2.21 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A1_c_251_n N_VGND_c_447_n 0.00225336f $X=2.27 $Y=0.785 $X2=0 $Y2=0
cc_201 A1 N_VGND_c_447_n 0.00587427f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_202 N_A1_c_240_n N_VGND_c_447_n 0.00422577f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_251_n N_VGND_c_449_n 0.00435174f $X=2.27 $Y=0.785 $X2=0 $Y2=0
cc_204 A1 N_VGND_c_449_n 0.00689293f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_205 N_A1_c_240_n N_VGND_c_449_n 0.00635347f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A1_c_251_n A_361_47# 0.00407707f $X=2.27 $Y=0.785 $X2=-0.19 $Y2=-0.24
cc_207 A1 A_361_47# 0.00465222f $X=1.99 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_208 N_B1_M1002_g N_VPWR_c_326_n 0.00120088f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1002_g N_VPWR_c_330_n 0.00555578f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1002_g N_VPWR_c_322_n 0.0109689f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1002_g N_A_277_297#_c_421_n 0.00326491f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_212 B1 N_VGND_M1004_d 0.00386298f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_213 N_B1_c_290_n N_VGND_c_445_n 0.00450677f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_214 B1 N_VGND_c_445_n 0.0150828f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_215 N_B1_c_292_n N_VGND_c_445_n 0.00231635f $X=2.98 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B1_c_290_n N_VGND_c_447_n 0.00539841f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_290_n N_VGND_c_449_n 0.0107126f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_218 B1 N_VGND_c_449_n 8.24099e-19 $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_219 N_VPWR_c_322_n N_X_M1003_s 0.00411607f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_327_n N_X_c_391_n 0.00252138f $X=0.935 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_322_n N_X_c_391_n 0.00490759f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_327_n N_X_c_401_n 0.0113346f $X=0.935 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_c_322_n N_X_c_401_n 0.00645703f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_M1003_d X 0.00270956f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_225 N_VPWR_M1003_d N_X_c_385_n 0.00293089f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_226 N_VPWR_c_323_n N_X_c_385_n 7.73122e-19 $X=0.26 $Y=2.635 $X2=0 $Y2=0
cc_227 N_VPWR_c_324_n N_X_c_385_n 0.0174235f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_228 N_VPWR_c_322_n N_X_c_385_n 0.00220706f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_322_n N_A_277_297#_M1001_d 0.00242015f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_230 N_VPWR_c_322_n N_A_277_297#_M1006_d 0.00304066f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_329_n N_A_277_297#_c_424_n 0.0119683f $X=1.815 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_322_n N_A_277_297#_c_424_n 0.00917629f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_VPWR_M1010_d N_A_277_297#_c_420_n 0.00446632f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_326_n N_A_277_297#_c_420_n 0.0174795f $X=1.98 $Y=2.26 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_329_n N_A_277_297#_c_420_n 0.00251566f $X=1.815 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_330_n N_A_277_297#_c_420_n 0.0022993f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_322_n N_A_277_297#_c_420_n 0.0104683f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_330_n N_A_277_297#_c_421_n 6.45126e-19 $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_322_n N_A_277_297#_c_421_n 0.00144032f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_330_n N_A_277_297#_c_439_n 0.0128729f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_322_n N_A_277_297#_c_439_n 0.00932279f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_X_c_383_n N_VGND_M1005_d 0.00294167f $X=0.217 $Y=0.885 $X2=-0.19
+ $Y2=-0.24
cc_243 N_X_c_383_n N_VGND_c_442_n 0.0214535f $X=0.217 $Y=0.885 $X2=0 $Y2=0
cc_244 N_X_c_381_n N_VGND_c_446_n 0.00283959f $X=0.595 $Y=0.8 $X2=0 $Y2=0
cc_245 N_X_c_411_p N_VGND_c_446_n 0.0113346f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_246 N_X_M1005_s N_VGND_c_449_n 0.00411607f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_247 N_X_c_381_n N_VGND_c_449_n 0.00580092f $X=0.595 $Y=0.8 $X2=0 $Y2=0
cc_248 N_X_c_411_p N_VGND_c_449_n 0.00645703f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_249 N_X_c_383_n N_VGND_c_449_n 0.00111111f $X=0.217 $Y=0.885 $X2=0 $Y2=0
cc_250 N_VGND_c_449_n A_277_47# 0.00728607f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_251 N_VGND_c_449_n A_361_47# 0.0083453f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

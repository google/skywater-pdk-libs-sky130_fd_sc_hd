* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
M1000 X a_1028_32# VPWR VPB phighvt w=790000u l=150000u
+  ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB phighvt w=790000u l=150000u
+  ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB phighvt w=790000u l=150000u
+  ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nshort w=650000u l=150000u
+  ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nshort w=650000u l=150000u
+  ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nshort w=650000u l=150000u
+  ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nshort w=650000u l=150000u
+  ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A LOWLVPWR LOWLVPWR phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_714_58# VGND nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB phighvt w=790000u l=150000u
+  ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ends


* File: sky130_fd_sc_hd__a31oi_4.pex.spice
* Created: Tue Sep  1 18:55:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A31OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47
r69 45 47 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.73 $Y2=1.16
r70 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.395
+ $Y=1.16 $X2=1.395 $Y2=1.16
r71 43 45 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.395 $Y2=1.16
r72 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r73 41 42 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r74 38 41 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.285 $Y=1.16
+ $X2=0.47 $Y2=1.16
r75 32 46 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.395 $Y2=1.16
r76 31 46 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.395 $Y2=1.16
r77 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=1.155 $Y2=1.16
r78 29 30 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.695 $Y2=1.16
r79 29 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r80 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r81 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r82 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r83 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r84 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r85 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r86 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r87 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r88 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r89 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r90 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r91 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r92 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r93 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r94 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r95 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47
r71 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.32 $Y=1.16 $X2=3.41
+ $Y2=1.16
r72 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=1.16 $X2=3.32 $Y2=1.16
r73 43 45 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.32 $Y2=1.16
r74 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r75 40 42 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.21 $Y=1.16
+ $X2=2.57 $Y2=1.16
r76 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.21
+ $Y=1.16 $X2=2.21 $Y2=1.16
r77 37 40 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.15 $Y=1.16 $X2=2.21
+ $Y2=1.16
r78 32 46 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.32 $Y2=1.16
r79 31 46 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=3.32 $Y2=1.16
r80 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.995 $Y2=1.16
r81 30 41 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.21 $Y2=1.16
r82 29 41 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.075 $Y=1.16
+ $X2=2.21 $Y2=1.16
r83 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r85 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r87 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r89 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r91 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r93 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r95 4 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r97 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%A1 3 7 9 11 14 16 18 21 23 25 26 28 29 30 31
+ 32 49
c70 32 0 1.91216e-19 $X=5.315 $Y=1.19
r71 48 49 11.3079 $w=3.41e-07 $l=8e-08 $layer=POLY_cond $X=5.11 $Y=1.17 $X2=5.19
+ $Y2=1.17
r72 46 48 12.7214 $w=3.41e-07 $l=9e-08 $layer=POLY_cond $X=5.02 $Y=1.17 $X2=5.11
+ $Y2=1.17
r73 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.02
+ $Y=1.16 $X2=5.02 $Y2=1.16
r74 44 46 35.3372 $w=3.41e-07 $l=2.5e-07 $layer=POLY_cond $X=4.77 $Y=1.17
+ $X2=5.02 $Y2=1.17
r75 43 44 11.3079 $w=3.41e-07 $l=8e-08 $layer=POLY_cond $X=4.69 $Y=1.17 $X2=4.77
+ $Y2=1.17
r76 42 43 48.0587 $w=3.41e-07 $l=3.4e-07 $layer=POLY_cond $X=4.35 $Y=1.17
+ $X2=4.69 $Y2=1.17
r77 41 42 11.3079 $w=3.41e-07 $l=8e-08 $layer=POLY_cond $X=4.27 $Y=1.17 $X2=4.35
+ $Y2=1.17
r78 39 41 50.8856 $w=3.41e-07 $l=3.6e-07 $layer=POLY_cond $X=3.91 $Y=1.17
+ $X2=4.27 $Y2=1.17
r79 37 39 8.48094 $w=3.41e-07 $l=6e-08 $layer=POLY_cond $X=3.85 $Y=1.17 $X2=3.91
+ $Y2=1.17
r80 32 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.315 $Y=1.16
+ $X2=5.02 $Y2=1.16
r81 31 47 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=1.16
+ $X2=5.02 $Y2=1.16
r82 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.395 $Y=1.16
+ $X2=4.855 $Y2=1.16
r83 29 30 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.91 $Y=1.16
+ $X2=4.395 $Y2=1.16
r84 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.91
+ $Y=1.16 $X2=3.91 $Y2=1.16
r85 26 49 59.3666 $w=3.41e-07 $l=4.2e-07 $layer=POLY_cond $X=5.61 $Y=1.17
+ $X2=5.19 $Y2=1.17
r86 26 28 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.61 $Y=1.01 $X2=5.61
+ $Y2=0.56
r87 23 49 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.17
r88 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r89 19 48 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.11 $Y=1.345
+ $X2=5.11 $Y2=1.17
r90 19 21 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.11 $Y=1.345
+ $X2=5.11 $Y2=1.985
r91 16 44 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.17
r92 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r93 12 43 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.69 $Y=1.345
+ $X2=4.69 $Y2=1.17
r94 12 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.69 $Y=1.345
+ $X2=4.69 $Y2=1.985
r95 9 42 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.17
r96 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
r97 5 41 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.27 $Y=1.345
+ $X2=4.27 $Y2=1.17
r98 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.27 $Y=1.345 $X2=4.27
+ $Y2=1.985
r99 1 37 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.85 $Y=1.345
+ $X2=3.85 $Y2=1.17
r100 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.85 $Y=1.345 $X2=3.85
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 31 33
+ 48 50
c76 50 0 1.91216e-19 $X=7.29 $Y=1.16
r77 49 50 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.87 $Y=1.16
+ $X2=7.29 $Y2=1.16
r78 47 49 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.77 $Y=1.16 $X2=6.87
+ $Y2=1.16
r79 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.16 $X2=6.77 $Y2=1.16
r80 45 47 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.77 $Y2=1.16
r81 43 45 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.03 $Y=1.16
+ $X2=6.45 $Y2=1.16
r82 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r83 33 48 1.41269 $w=6.33e-07 $l=7.5e-08 $layer=LI1_cond $X=6.695 $Y=1.312
+ $X2=6.77 $Y2=1.312
r84 31 33 8.66451 $w=6.33e-07 $l=4.6e-07 $layer=LI1_cond $X=6.235 $Y=1.312
+ $X2=6.695 $Y2=1.312
r85 31 44 3.86136 $w=6.33e-07 $l=2.05e-07 $layer=LI1_cond $X=6.235 $Y=1.312
+ $X2=6.03 $Y2=1.312
r86 29 44 4.80315 $w=6.33e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=1.312
+ $X2=6.03 $Y2=1.312
r87 25 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.16
r88 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.985
r89 22 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=1.16
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=0.56
r91 18 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.16
r92 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.985
r93 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=1.16
r94 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=0.56
r95 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r96 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r97 8 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r98 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r99 4 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r100 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r101 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 54 56 60 62 67 68 69 72 76 77 78 79 80
r92 72 82 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.54 $Y=2.255
+ $X2=7.54 $Y2=2.34
r93 72 74 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=7.54 $Y=2.255
+ $X2=7.54 $Y2=1.66
r94 69 71 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=5.405 $Y=2.34
+ $X2=6.66 $Y2=2.34
r95 68 82 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.415 $Y=2.34
+ $X2=7.54 $Y2=2.34
r96 68 71 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.415 $Y=2.34
+ $X2=6.66 $Y2=2.34
r97 65 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.32 $Y=2.255
+ $X2=5.405 $Y2=2.34
r98 65 67 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.32 $Y=2.255
+ $X2=5.32 $Y2=1.8
r99 64 67 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.32 $Y=1.665
+ $X2=5.32 $Y2=1.8
r100 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=1.58
+ $X2=4.48 $Y2=1.58
r101 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.235 $Y=1.58
+ $X2=5.32 $Y2=1.665
r102 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.235 $Y=1.58
+ $X2=4.565 $Y2=1.58
r103 58 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=1.665
+ $X2=4.48 $Y2=1.58
r104 58 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.48 $Y=1.665
+ $X2=4.48 $Y2=1.96
r105 57 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=1.58
+ $X2=3.62 $Y2=1.58
r106 56 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=1.58
+ $X2=4.48 $Y2=1.58
r107 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.395 $Y=1.58
+ $X2=3.705 $Y2=1.58
r108 52 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.665
+ $X2=3.62 $Y2=1.58
r109 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.62 $Y=1.665
+ $X2=3.62 $Y2=1.96
r110 51 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.58
+ $X2=2.78 $Y2=1.58
r111 50 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=1.58
+ $X2=3.62 $Y2=1.58
r112 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=1.58
+ $X2=2.865 $Y2=1.58
r113 46 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=1.665
+ $X2=2.78 $Y2=1.58
r114 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.78 $Y=1.665
+ $X2=2.78 $Y2=1.96
r115 45 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.58
+ $X2=1.94 $Y2=1.58
r116 44 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=1.58
+ $X2=2.78 $Y2=1.58
r117 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=1.58
+ $X2=2.025 $Y2=1.58
r118 40 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=1.665
+ $X2=1.94 $Y2=1.58
r119 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=1.665
+ $X2=1.94 $Y2=1.96
r120 39 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.58
+ $X2=1.1 $Y2=1.58
r121 38 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=1.58
+ $X2=1.94 $Y2=1.58
r122 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=1.58
+ $X2=1.185 $Y2=1.58
r123 34 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.665 $X2=1.1
+ $Y2=1.58
r124 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=1.665
+ $X2=1.1 $Y2=1.96
r125 32 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=1.58
+ $X2=1.1 $Y2=1.58
r126 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=1.58
+ $X2=0.345 $Y2=1.58
r127 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.345 $Y2=1.58
r128 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.96
r129 9 82 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=2.34
r130 9 74 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=1.66
r131 8 71 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=2.34
r132 7 67 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=5.185
+ $Y=1.485 $X2=5.32 $Y2=1.8
r133 6 60 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.48 $Y2=1.96
r134 5 54 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.96
r135 4 48 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.96
r136 3 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r137 2 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r138 1 30 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 43 46 47
+ 49 50 51 52 53 55 70 80 81 84 87 90
r117 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r118 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 78 81 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.59 $Y2=2.72
r122 78 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 77 80 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=7.59 $Y2=2.72
r124 77 78 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r125 75 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.9 $Y2=2.72
r126 75 77 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=5.29 $Y2=2.72
r127 74 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 74 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r130 71 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.06 $Y2=2.72
r131 71 73 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 70 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=2.72
+ $X2=4.9 $Y2=2.72
r133 70 73 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.735 $Y=2.72
+ $X2=4.37 $Y2=2.72
r134 69 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r135 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r136 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r137 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r138 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r139 63 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r140 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r142 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 55 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r144 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 53 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 53 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 51 68 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.99 $Y2=2.72
r148 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.2 $Y2=2.72
r149 49 65 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r150 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.36 $Y2=2.72
r151 48 68 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.99 $Y2=2.72
r152 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.36 $Y2=2.72
r153 46 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.15 $Y2=2.72
r154 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.52 $Y2=2.72
r155 45 65 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=2.07 $Y2=2.72
r156 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.52 $Y2=2.72
r157 41 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.9 $Y=2.635 $X2=4.9
+ $Y2=2.72
r158 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.9 $Y=2.635
+ $X2=4.9 $Y2=2.34
r159 37 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=2.635
+ $X2=4.06 $Y2=2.72
r160 37 39 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.06 $Y=2.635
+ $X2=4.06 $Y2=2
r161 36 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.72
+ $X2=3.2 $Y2=2.72
r162 35 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=4.06 $Y2=2.72
r163 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=3.365 $Y2=2.72
r164 31 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635 $X2=3.2
+ $Y2=2.72
r165 31 33 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2
r166 27 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r167 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2
r168 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r169 23 25 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2
r170 19 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r171 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2
r172 6 43 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.485 $X2=4.9 $Y2=2.34
r173 5 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.485 $X2=4.06 $Y2=2
r174 4 33 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2
r175 3 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2
r176 2 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
r177 1 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%Y 1 2 3 4 5 6 7 22 30 36 38 42 44 45 46 47
+ 48 56 58 66 69
r69 56 66 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=7.145 $Y=1.915
+ $X2=7.145 $Y2=1.87
r70 55 58 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=7.145 $Y=0.805
+ $X2=7.145 $Y2=0.85
r71 48 56 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=2 $X2=7.145
+ $Y2=1.915
r72 48 66 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=7.145 $Y=1.85
+ $X2=7.145 $Y2=1.87
r73 47 48 17.7455 $w=1.98e-07 $l=3.2e-07 $layer=LI1_cond $X=7.145 $Y=1.53
+ $X2=7.145 $Y2=1.85
r74 46 47 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=7.145 $Y=1.19
+ $X2=7.145 $Y2=1.53
r75 45 69 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.155 $Y=0.72
+ $X2=7.5 $Y2=0.72
r76 45 55 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.155 $Y=0.72
+ $X2=7.145 $Y2=0.72
r77 45 46 17.7455 $w=1.98e-07 $l=3.2e-07 $layer=LI1_cond $X=7.145 $Y=0.87
+ $X2=7.145 $Y2=1.19
r78 45 58 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=7.145 $Y=0.87
+ $X2=7.145 $Y2=0.85
r79 40 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.635 $X2=7.5
+ $Y2=0.72
r80 40 42 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.5 $Y=0.635
+ $X2=7.5 $Y2=0.42
r81 39 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0.72
+ $X2=6.66 $Y2=0.72
r82 38 55 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=7.045 $Y=0.72
+ $X2=7.145 $Y2=0.72
r83 38 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.045 $Y=0.72
+ $X2=6.745 $Y2=0.72
r84 34 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.635
+ $X2=6.66 $Y2=0.72
r85 34 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.66 $Y=0.635
+ $X2=6.66 $Y2=0.42
r86 30 48 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.045 $Y=2 $X2=7.145
+ $Y2=2
r87 30 32 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=7.045 $Y=2 $X2=6.24
+ $Y2=2
r88 27 29 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.98 $Y=0.72
+ $X2=5.82 $Y2=0.72
r89 24 27 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.72
+ $X2=4.98 $Y2=0.72
r90 22 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0.72
+ $X2=6.66 $Y2=0.72
r91 22 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.575 $Y=0.72
+ $X2=5.82 $Y2=0.72
r92 7 48 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=2
r93 6 32 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=2
r94 5 42 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.42
r95 4 36 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.42
r96 3 29 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.72
r97 2 27 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.72
r98 1 24 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 30 36 38
+ 39
r50 34 36 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.72
+ $X2=3.62 $Y2=0.72
r51 32 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.72
+ $X2=1.94 $Y2=0.72
r52 32 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.72
+ $X2=2.78 $Y2=0.72
r53 28 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.635
+ $X2=1.94 $Y2=0.72
r54 28 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.94 $Y=0.635
+ $X2=1.94 $Y2=0.42
r55 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.72 $X2=1.1
+ $Y2=0.72
r56 26 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0.72
+ $X2=1.94 $Y2=0.72
r57 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=0.72
+ $X2=1.185 $Y2=0.72
r58 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.635 $X2=1.1
+ $Y2=0.72
r59 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.1 $Y=0.635
+ $X2=1.1 $Y2=0.42
r60 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.72 $X2=1.1
+ $Y2=0.72
r61 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=0.345 $Y2=0.72
r62 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r63 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r64 5 36 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.72
r65 4 34 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.72
r66 3 30 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.42
r67 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r68 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 53
+ 54 57 60 63 66
r112 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r113 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r114 60 61 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r115 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 54 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r117 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r118 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=0 $X2=7.08
+ $Y2=0
r119 51 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.245 $Y=0 $X2=7.59
+ $Y2=0
r120 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r121 50 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r122 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r123 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.24
+ $Y2=0
r124 47 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=0
+ $X2=6.67 $Y2=0
r125 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=7.08
+ $Y2=0
r126 46 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.67
+ $Y2=0
r127 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r128 45 61 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=1.61
+ $Y2=0
r129 44 45 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r130 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r131 42 44 265.203 $w=1.68e-07 $l=4.065e-06 $layer=LI1_cond $X=1.685 $Y=0
+ $X2=5.75 $Y2=0
r132 41 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0 $X2=6.24
+ $Y2=0
r133 41 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=5.75 $Y2=0
r134 40 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r135 40 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r136 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r137 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r138 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r139 36 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r140 36 39 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.15 $Y2=0
r141 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r142 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r143 29 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r144 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r145 25 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0
r146 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0.38
r147 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=0.085
+ $X2=6.24 $Y2=0
r148 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.24 $Y=0.085
+ $X2=6.24 $Y2=0.38
r149 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r150 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.38
r151 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r152 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r153 4 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.38
r154 3 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.38
r155 2 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r156 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_4%A_445_47# 1 2 3 4 21
r29 19 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.38 $X2=5.4
+ $Y2=0.38
r30 17 19 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.2 $Y=0.38
+ $X2=4.56 $Y2=0.38
r31 14 17 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.38 $X2=3.2
+ $Y2=0.38
r32 4 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.38
r33 3 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.38
r34 2 17 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.38
r35 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.38
.ends


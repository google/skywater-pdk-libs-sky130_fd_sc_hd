* File: sky130_fd_sc_hd__sdfsbp_2.spice
* Created: Thu Aug 27 14:46:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfsbp_2.spice.pex"
.subckt sky130_fd_sc_hd__sdfsbp_2  VNB VPB SCD SCE D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1041 A_109_47# N_SCD_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1016 N_A_181_47#_M1016_d N_SCE_M1016_g A_109_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1027 A_265_47# N_D_M1027_g N_A_181_47#_M1016_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.0567 PD=0.735 PS=0.69 NRD=29.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_328_21#_M1036_g A_265_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.06615 PD=1.36 PS=0.735 NRD=0 NRS=29.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SCE_M1024_g N_A_328_21#_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_CLK_M1003_g N_A_652_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1045 N_A_818_47#_M1045_d N_A_652_47#_M1045_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_A_1006_47#_M1030_d N_A_652_47#_M1030_g N_A_181_47#_M1030_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1019 A_1090_47# N_A_818_47#_M1019_g N_A_1006_47#_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1132_21#_M1022_g A_1090_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1350_47# N_A_1006_47#_M1002_g N_A_1132_21#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_SET_B_M1037_g A_1350_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0758774 AS=0.0441 PD=0.764717 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1023 A_1517_47# N_A_1006_47#_M1023_g N_VGND_M1037_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2336 AS=0.115623 PD=1.37 PS=1.16528 NRD=58.116 NRS=9.372 M=1 R=4.26667
+ SA=75000.7 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1043 N_A_1597_329#_M1043_d N_A_818_47#_M1043_g A_1517_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.147321 AS=0.2336 PD=1.31623 PS=1.37 NRD=4.68 NRS=58.116 M=1
+ R=4.26667 SA=75001.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1018 A_1813_47# N_A_652_47#_M1018_g N_A_1597_329#_M1043_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0966792 PD=0.63 PS=0.863774 NRD=14.28 NRS=41.424 M=1
+ R=2.8 SA=75002.5 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1020 A_1885_47# N_A_1781_295#_M1020_g A_1813_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8 SA=75002.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SET_B_M1014_g A_1885_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0735 PD=0.755 PS=0.77 NRD=15.708 NRS=34.284 M=1 R=2.8
+ SA=75003.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_1781_295#_M1000_d N_A_1597_329#_M1000_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.07035 PD=1.37 PS=0.755 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_1597_329#_M1035_g N_Q_N_M1035_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1038_d N_A_1597_329#_M1038_g N_Q_N_M1035_s VNB NSHORT L=0.15
+ W=0.65 AD=0.21125 AS=0.08775 PD=1.95 PS=0.92 NRD=11.076 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_1597_329#_M1011_g N_A_2501_47#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=5.712 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1040 N_VGND_M1011_d N_A_2501_47#_M1040_g N_Q_M1040_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.08775 PD=1.18458 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1042 N_VGND_M1042_d N_A_2501_47#_M1042_g N_Q_M1040_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1025 N_VPWR_M1025_d N_SCD_M1025_g N_A_27_369#_M1025_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 A_193_369# N_SCE_M1001_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1004 N_A_181_47#_M1004_d N_D_M1004_g A_193_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1056 AS=0.0672 PD=0.97 PS=0.85 NRD=16.9223 NRS=15.3857 M=1 R=4.26667
+ SA=75001 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1032 N_A_27_369#_M1032_d N_A_328_21#_M1032_g N_A_181_47#_M1004_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.162825 AS=0.1056 PD=1.8 PS=0.97 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_VPWR_M1029_d N_SCE_M1029_g N_A_328_21#_M1029_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.162825 PD=1.8 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_652_47#_M1010_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1031 N_A_818_47#_M1031_d N_A_652_47#_M1031_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_1006_47#_M1007_d N_A_818_47#_M1007_g N_A_181_47#_M1007_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06825 AS=0.1092 PD=0.745 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1034 A_1102_413# N_A_652_47#_M1034_g N_A_1006_47#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.06825 PD=0.72 PS=0.745 NRD=44.5417 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1044 N_VPWR_M1044_d N_A_1132_21#_M1044_g A_1102_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09345 AS=0.063 PD=0.865 PS=0.72 NRD=30.4759 NRS=44.5417 M=1 R=2.8
+ SA=75001.1 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_1132_21#_M1008_d N_A_1006_47#_M1008_g N_VPWR_M1044_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0714 AS=0.09345 PD=0.76 PS=0.865 NRD=9.3772 NRS=46.886 M=1
+ R=2.8 SA=75001.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1033 N_VPWR_M1033_d N_SET_B_M1033_g N_A_1132_21#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0952 AS=0.0714 PD=0.846667 PS=0.76 NRD=18.7544 NRS=18.7544 M=1
+ R=2.8 SA=75002.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1015 A_1525_329# N_A_1006_47#_M1015_g N_VPWR_M1033_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.0882 AS=0.1904 PD=1.05 PS=1.69333 NRD=11.7215 NRS=25.7873 M=1 R=5.6
+ SA=75001.5 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1021 N_A_1597_329#_M1021_d N_A_652_47#_M1021_g A_1525_329# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2044 AS=0.0882 PD=1.76 PS=1.05 NRD=34.0022 NRS=11.7215 M=1 R=5.6
+ SA=75001.8 SB=75001 A=0.126 P=1.98 MULT=1
MM1039 A_1723_413# N_A_818_47#_M1039_g N_A_1597_329#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0609 AS=0.1022 PD=0.71 PS=0.88 NRD=42.1974 NRS=25.7873 M=1 R=2.8
+ SA=75003.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1781_295#_M1009_g A_1723_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.08505 AS=0.0609 PD=0.825 PS=0.71 NRD=60.9715 NRS=42.1974 M=1 R=2.8
+ SA=75004.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_1597_329#_M1013_d N_SET_B_M1013_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.08505 PD=1.36 PS=0.825 NRD=0 NRS=0 M=1 R=2.8 SA=75004.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_A_1781_295#_M1026_d N_A_1597_329#_M1026_g N_VPWR_M1026_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_1597_329#_M1012_g N_Q_N_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1028_d N_A_1597_329#_M1028_g N_Q_N_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.325 AS=0.135 PD=2.65 PS=1.27 NRD=11.8003 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_1597_329#_M1005_g N_A_2501_47#_M1005_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=13.8491 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1005_d N_A_2501_47#_M1006_g N_Q_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.181707 AS=0.135 PD=1.61585 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A_2501_47#_M1017_g N_Q_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.31 AS=0.135 PD=2.62 PS=1.27 NRD=8.8453 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX46_noxref VNB VPB NWDIODE A=23.4972 P=32.49
c_294 VPB 0 9.29321e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__sdfsbp_2.spice.SKY130_FD_SC_HD__SDFSBP_2.pxi"
*
.ends
*
*

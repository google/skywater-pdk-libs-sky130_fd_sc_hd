* File: sky130_fd_sc_hd__nor4_2.spice.pex
* Created: Thu Aug 27 14:32:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4_2%A 1 3 6 8 10 13 15 22
r40 20 22 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.645 $Y=1.16
+ $X2=0.91 $Y2=1.16
r41 17 20 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.645 $Y2=1.16
r42 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r43 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r44 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r45 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r46 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r47 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%B 1 3 6 8 10 13 15 22
r44 20 22 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.525 $Y=1.16
+ $X2=1.75 $Y2=1.16
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.16 $X2=1.525 $Y2=1.16
r46 17 20 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.525 $Y2=1.16
r47 15 21 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=1.525 $Y2=1.18
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325 $X2=1.33
+ $Y2=1.985
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995 $X2=1.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%C 1 3 6 8 10 13 15 21 22
c41 21 0 1.72994e-19 $X=2.94 $Y=1.16
r42 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.94 $Y=1.16
+ $X2=3.15 $Y2=1.16
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.16 $X2=2.94 $Y2=1.16
r44 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=2.94 $Y2=1.16
r45 15 21 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=2.555 $Y=1.18
+ $X2=2.94 $Y2=1.18
r46 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.16
r47 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.985
r48 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=1.16
r49 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=0.56
r50 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.16
r51 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.325 $X2=2.73
+ $Y2=1.985
r52 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=0.995
+ $X2=2.73 $Y2=1.16
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.995 $X2=2.73
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%D 1 3 6 8 10 13 15 21 22
c43 22 0 1.72994e-19 $X=3.99 $Y=1.16
r44 20 22 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.76 $Y=1.16
+ $X2=3.99 $Y2=1.16
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.16 $X2=3.76 $Y2=1.16
r46 17 20 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.57 $Y=1.16
+ $X2=3.76 $Y2=1.16
r47 15 21 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=3.475 $Y=1.18
+ $X2=3.76 $Y2=1.18
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.985
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=0.995
+ $X2=3.99 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.99 $Y=0.995
+ $X2=3.99 $Y2=0.56
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.57 $Y=1.325 $X2=3.57
+ $Y2=1.985
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=0.995
+ $X2=3.57 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.57 $Y=0.995 $X2=3.57
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%A_27_297# 1 2 3 10 12 14 18 20 27 29
r36 21 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.54
+ $X2=1.12 $Y2=1.54
r37 20 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.96 $Y2=1.54
r38 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.245 $Y2=1.54
r39 16 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=1.54
r40 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=2.3
r41 15 25 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r42 14 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=1.12 $Y2=1.54
r43 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=0.405 $Y2=1.54
r44 10 25 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r45 10 12 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r46 3 29 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r47 2 27 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r48 2 18 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r49 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r50 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%VPWR 1 6 8 10 20 21 24
r47 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 20 21 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r49 18 21 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=4.37 $Y2=2.72
r50 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 17 20 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=4.37 $Y2=2.72
r52 17 18 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 15 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r54 15 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 10 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r56 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r59 4 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r60 4 6 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r61 1 6 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%A_281_297# 1 2 9 11 12 15
r19 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.94 $Y=2.295
+ $X2=2.94 $Y2=1.96
r20 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.815 $Y=2.38
+ $X2=2.94 $Y2=2.295
r21 11 12 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=2.815 $Y=2.38
+ $X2=1.665 $Y2=2.38
r22 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.665 $Y2=2.38
r23 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.54 $Y2=1.96
r24 2 15 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=1.96
r25 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%A_475_297# 1 2 3 12 14 15 16 20 23
r35 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.2 $Y=2.295
+ $X2=4.2 $Y2=1.96
r36 17 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=2.38
+ $X2=3.36 $Y2=2.38
r37 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.075 $Y=2.38
+ $X2=4.2 $Y2=2.295
r38 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.075 $Y=2.38
+ $X2=3.485 $Y2=2.38
r39 15 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=2.295
+ $X2=3.36 $Y2=2.38
r40 14 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=1.625
+ $X2=3.36 $Y2=1.54
r41 14 15 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.36 $Y=1.625
+ $X2=3.36 $Y2=2.295
r42 13 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.645 $Y=1.54
+ $X2=2.52 $Y2=1.54
r43 12 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=1.54
+ $X2=3.36 $Y2=1.54
r44 12 13 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.235 $Y=1.54
+ $X2=2.645 $Y2=1.54
r45 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.065
+ $Y=1.485 $X2=4.2 $Y2=1.96
r46 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=2.3
r47 2 25 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=1.62
r48 1 23 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.375
+ $Y=1.485 $X2=2.52 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%Y 1 2 3 4 5 18 20 21 24 26 30 32 36 40 42 44
+ 45 46 48 50 53
r109 50 53 2.6797 $w=3.35e-07 $l=9e-08 $layer=LI1_cond $X=4.347 $Y=0.815
+ $X2=4.347 $Y2=0.905
r110 50 53 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=4.347 $Y=0.92
+ $X2=4.347 $Y2=0.905
r111 49 50 18.4047 $w=3.33e-07 $l=5.35e-07 $layer=LI1_cond $X=4.347 $Y=1.455
+ $X2=4.347 $Y2=0.92
r112 43 46 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0.815
+ $X2=3.78 $Y2=0.815
r113 42 50 4.97233 $w=1.8e-07 $l=1.67e-07 $layer=LI1_cond $X=4.18 $Y=0.815
+ $X2=4.347 $Y2=0.815
r114 42 43 14.4798 $w=1.78e-07 $l=2.35e-07 $layer=LI1_cond $X=4.18 $Y=0.815
+ $X2=3.945 $Y2=0.815
r115 41 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=1.54
+ $X2=3.78 $Y2=1.54
r116 40 49 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=4.18 $Y=1.54
+ $X2=4.347 $Y2=1.455
r117 40 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.18 $Y=1.54
+ $X2=3.905 $Y2=1.54
r118 34 46 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.78 $Y=0.725
+ $X2=3.78 $Y2=0.815
r119 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.78 $Y=0.725
+ $X2=3.78 $Y2=0.39
r120 33 45 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0.815
+ $X2=2.94 $Y2=0.815
r121 32 46 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0.815
+ $X2=3.78 $Y2=0.815
r122 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.615 $Y=0.815
+ $X2=3.105 $Y2=0.815
r123 28 45 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.94 $Y=0.725
+ $X2=2.94 $Y2=0.815
r124 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.94 $Y=0.725
+ $X2=2.94 $Y2=0.39
r125 27 44 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r126 26 45 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=2.94 $Y2=0.815
r127 26 27 65.9293 $w=1.78e-07 $l=1.07e-06 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=1.705 $Y2=0.815
r128 22 44 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r129 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r130 20 44 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r131 20 21 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r132 16 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r133 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r134 5 48 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.645
+ $Y=1.485 $X2=3.78 $Y2=1.62
r135 4 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.645
+ $Y=0.235 $X2=3.78 $Y2=0.39
r136 3 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.235 $X2=2.94 $Y2=0.39
r137 2 24 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r138 1 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_2%VGND 1 2 3 4 5 6 19 21 25 29 31 33 36 37 39
+ 40 41 55 64 70 73
r77 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r78 69 70 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0.235
+ $X2=2.605 $Y2=0.235
r79 66 69 8.40993 $w=6.38e-07 $l=4.5e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.52 $Y2=0.235
r80 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r81 63 66 2.05576 $w=6.38e-07 $l=1.1e-07 $layer=LI1_cond $X=1.96 $Y=0.235
+ $X2=2.07 $Y2=0.235
r82 63 64 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.235
+ $X2=1.875 $Y2=0.235
r83 58 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r84 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r85 55 72 4.24518 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.357
+ $Y2=0
r86 55 57 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=3.91
+ $Y2=0
r87 54 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r88 54 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r89 53 70 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.605
+ $Y2=0
r90 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r91 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r92 49 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.875
+ $Y2=0
r93 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r94 46 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r95 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r96 43 60 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r97 43 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r98 41 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r99 41 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r100 39 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.275 $Y=0
+ $X2=2.99 $Y2=0
r101 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.36
+ $Y2=0
r102 38 57 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.91 $Y2=0
r103 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.36
+ $Y2=0
r104 36 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r105 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r106 35 49 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r107 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r108 31 72 3.19266 $w=2.9e-07 $l=1.32868e-07 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.357 $Y2=0
r109 31 33 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0.39
r110 27 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=0.085
+ $X2=3.36 $Y2=0
r111 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.36 $Y=0.085
+ $X2=3.36 $Y2=0.39
r112 23 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r113 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r114 19 60 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r115 19 21 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r116 6 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.235 $X2=4.2 $Y2=0.39
r117 5 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.36 $Y2=0.39
r118 4 69 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.235 $X2=2.52 $Y2=0.39
r119 3 63 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r120 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r121 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_8.pxi.spice
* Created: Tue Sep  1 19:10:56 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%A N_A_M1004_g N_A_c_74_n N_A_M1007_g
+ N_A_M1012_g N_A_c_75_n N_A_M1018_g A A N_A_c_73_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%A_110_47# N_A_110_47#_M1004_d
+ N_A_110_47#_M1007_d N_A_110_47#_M1001_g N_A_110_47#_M1000_g
+ N_A_110_47#_M1006_g N_A_110_47#_M1002_g N_A_110_47#_M1008_g
+ N_A_110_47#_M1003_g N_A_110_47#_M1010_g N_A_110_47#_M1005_g
+ N_A_110_47#_M1014_g N_A_110_47#_M1009_g N_A_110_47#_M1016_g
+ N_A_110_47#_M1011_g N_A_110_47#_M1017_g N_A_110_47#_M1013_g
+ N_A_110_47#_c_120_n N_A_110_47#_M1019_g N_A_110_47#_M1015_g
+ N_A_110_47#_c_122_n N_A_110_47#_c_133_n N_A_110_47#_c_123_n
+ N_A_110_47#_c_146_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%A_110_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%KAPWR N_KAPWR_M1007_s N_KAPWR_M1018_s
+ N_KAPWR_M1002_s N_KAPWR_M1005_s N_KAPWR_M1011_s N_KAPWR_M1015_s
+ N_KAPWR_c_283_n N_KAPWR_c_288_n N_KAPWR_c_290_n N_KAPWR_c_300_n
+ N_KAPWR_c_302_n N_KAPWR_c_304_n N_KAPWR_c_305_n N_KAPWR_c_307_n
+ N_KAPWR_c_309_n N_KAPWR_c_310_n N_KAPWR_c_312_n N_KAPWR_c_314_n
+ N_KAPWR_c_284_n N_KAPWR_c_285_n N_KAPWR_c_316_n KAPWR N_KAPWR_c_286_n
+ N_KAPWR_c_294_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%X N_X_M1001_s N_X_M1008_s N_X_M1014_s
+ N_X_M1017_s N_X_M1000_d N_X_M1003_d N_X_M1009_d N_X_M1013_d N_X_c_391_n
+ N_X_c_392_n N_X_c_393_n N_X_c_415_n N_X_c_394_n N_X_c_395_n N_X_c_425_n
+ N_X_c_396_n N_X_c_397_n N_X_c_434_n N_X_c_398_n N_X_c_439_n N_X_c_399_n
+ N_X_c_445_n N_X_c_400_n N_X_c_451_n X X X
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%X
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%VGND N_VGND_M1004_s N_VGND_M1012_s
+ N_VGND_M1006_d N_VGND_M1010_d N_VGND_M1016_d N_VGND_M1019_d N_VGND_c_544_n
+ N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n N_VGND_c_549_n
+ N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n
+ N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n VGND
+ N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n N_VGND_c_562_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%VPWR VPWR N_VPWR_c_629_n
+ N_VPWR_c_628_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%VPWR
cc_1 VNB N_A_M1004_g 0.0280927f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_M1012_g 0.0234436f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_3 VNB A 0.0260861f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_A_c_73_n 0.0669956f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.155
cc_5 VNB N_A_110_47#_M1001_g 0.0260664f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_6 VNB N_A_110_47#_M1006_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_110_47#_M1008_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_110_47#_M1010_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_110_47#_M1014_g 0.0241252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_110_47#_M1016_g 0.0241164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_110_47#_M1017_g 0.023767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_110_47#_c_120_n 0.151577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_110_47#_M1019_g 0.0320587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_110_47#_c_122_n 0.00445674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_c_123_n 0.00442652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_391_n 0.00160391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_392_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_393_n 0.00419804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_394_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_395_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_396_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_397_n 0.00400554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_398_n 0.0013724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_399_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_400_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0301966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_544_n 0.0112866f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.155
cc_28 VNB N_VGND_c_545_n 0.00454665f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_29 VNB N_VGND_c_546_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_547_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.16
cc_31 VNB N_VGND_c_548_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_549_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_550_n 0.0177301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_551_n 0.0160902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_552_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_553_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_554_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_555_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_556_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_557_n 0.0154599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_558_n 0.00574315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_559_n 0.0166984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_560_n 0.0126445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_561_n 0.266016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_562_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_628_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_47 VPB N_A_c_74_n 0.0192408f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.41
cc_48 VPB N_A_c_75_n 0.0145802f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.41
cc_49 VPB A 0.00123221f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_50 VPB N_A_c_73_n 0.0273976f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.155
cc_51 VPB N_A_110_47#_M1000_g 0.0190615f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_52 VPB N_A_110_47#_M1002_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_53 VPB N_A_110_47#_M1003_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.16
cc_54 VPB N_A_110_47#_M1005_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_110_47#_M1009_g 0.0187459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_110_47#_M1011_g 0.0187139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_110_47#_M1013_g 0.0173762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_110_47#_c_120_n 0.0250755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_110_47#_M1015_g 0.0224494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_110_47#_c_133_n 0.00140018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_110_47#_c_123_n 0.00331269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_KAPWR_c_283_n 0.00916947f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_63 VPB N_KAPWR_c_284_n 0.0196104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_KAPWR_c_285_n 0.0172609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_KAPWR_c_286_n 0.0316932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB X 0.010431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB X 0.0105833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_629_n 0.138209f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.9
cc_69 VPB N_VPWR_c_628_n 0.0446842f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.445
cc_70 N_A_M1012_g N_A_110_47#_M1001_g 0.0206811f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_c_75_n N_A_110_47#_M1000_g 0.0206811f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_c_73_n N_A_110_47#_c_120_n 0.0206811f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_A_110_47#_c_122_n 0.0030957f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1012_g N_A_110_47#_c_122_n 0.00356184f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_75 A N_A_110_47#_c_122_n 0.0277994f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_c_73_n N_A_110_47#_c_122_n 0.0116674f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_77 N_A_c_74_n N_A_110_47#_c_133_n 0.00314473f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_75_n N_A_110_47#_c_133_n 0.00318278f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_73_n N_A_110_47#_c_133_n 0.00945812f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_80 N_A_c_73_n N_A_110_47#_c_123_n 0.0213857f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_81 A N_A_110_47#_c_146_n 0.0198893f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A_c_73_n N_A_110_47#_c_146_n 0.00950927f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_83 N_A_c_74_n N_KAPWR_c_283_n 8.41569e-19 $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_74_n N_KAPWR_c_288_n 0.00707826f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_75_n N_KAPWR_c_288_n 0.00707826f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_75_n N_KAPWR_c_290_n 6.76362e-19 $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_74_n N_KAPWR_c_286_n 0.00416048f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_88 A N_KAPWR_c_286_n 0.0206626f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_c_73_n N_KAPWR_c_286_n 0.00767867f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_90 N_A_c_75_n N_KAPWR_c_294_n 0.00123279f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_91 A N_VGND_c_544_n 0.00101698f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_M1004_g N_VGND_c_545_n 0.00339198f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_93 A N_VGND_c_545_n 0.0191362f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_94 N_A_c_73_n N_VGND_c_545_n 0.00113059f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_95 N_A_M1012_g N_VGND_c_546_n 0.00168046f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_M1004_g N_VGND_c_559_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_M1012_g N_VGND_c_559_n 0.00585385f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_M1004_g N_VGND_c_561_n 0.011499f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_M1012_g N_VGND_c_561_n 0.0106694f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_100 A N_VGND_c_561_n 0.00301823f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_101 N_A_c_74_n N_VPWR_c_629_n 0.00585385f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_75_n N_VPWR_c_629_n 0.00585385f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_74_n N_VPWR_c_628_n 0.00626028f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_75_n N_VPWR_c_628_n 0.00531811f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_110_47#_c_133_n N_KAPWR_c_283_n 0.00151781f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_106 N_A_110_47#_M1007_d N_KAPWR_c_288_n 0.00115925f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_107 N_A_110_47#_c_133_n N_KAPWR_c_288_n 0.0252733f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_108 N_A_110_47#_M1000_g N_KAPWR_c_290_n 6.76362e-19 $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_110_47#_c_133_n N_KAPWR_c_290_n 0.00152672f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_110 N_A_110_47#_M1002_g N_KAPWR_c_300_n 0.00115346f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_110_47#_M1003_g N_KAPWR_c_300_n 0.00115346f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_110_47#_M1000_g N_KAPWR_c_302_n 0.00707826f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_110_47#_M1002_g N_KAPWR_c_302_n 0.00267097f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_110_47#_M1002_g N_KAPWR_c_304_n 6.44793e-19 $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_110_47#_M1005_g N_KAPWR_c_305_n 0.00114528f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_110_47#_M1009_g N_KAPWR_c_305_n 0.00114528f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_110_47#_M1003_g N_KAPWR_c_307_n 0.00285301f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_110_47#_M1005_g N_KAPWR_c_307_n 0.00248894f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_110_47#_M1005_g N_KAPWR_c_309_n 6.91139e-19 $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_110_47#_M1011_g N_KAPWR_c_310_n 0.00115346f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_110_47#_M1013_g N_KAPWR_c_310_n 0.00115346f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_110_47#_M1009_g N_KAPWR_c_312_n 0.00285301f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_110_47#_M1011_g N_KAPWR_c_312_n 0.00285301f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_110_47#_M1013_g N_KAPWR_c_314_n 6.44661e-19 $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_110_47#_M1015_g N_KAPWR_c_285_n 0.00379528f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_110_47#_M1013_g N_KAPWR_c_316_n 0.00266891f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_110_47#_M1015_g N_KAPWR_c_316_n 0.0028508f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_110_47#_c_133_n N_KAPWR_c_286_n 0.00777957f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_129 N_A_110_47#_M1000_g N_KAPWR_c_294_n 0.00123279f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_110_47#_c_133_n N_KAPWR_c_294_n 0.0082174f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_131 N_A_110_47#_c_123_n N_KAPWR_c_294_n 0.0158218f $X=3.245 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_110_47#_M1001_g N_X_c_391_n 0.00120255f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_110_47#_M1006_g N_X_c_391_n 0.00120255f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A_110_47#_c_122_n N_X_c_391_n 0.00257148f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_110_47#_M1006_g N_X_c_392_n 0.0119364f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_110_47#_M1008_g N_X_c_392_n 0.0122327f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_110_47#_c_120_n N_X_c_392_n 0.00267078f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_138 N_A_110_47#_c_123_n N_X_c_392_n 0.0429599f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_110_47#_M1001_g N_X_c_393_n 0.00289158f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_110_47#_c_120_n N_X_c_393_n 0.00277135f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_141 N_A_110_47#_c_122_n N_X_c_393_n 0.00599637f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_110_47#_c_123_n N_X_c_393_n 0.0213686f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_110_47#_M1002_g N_X_c_415_n 0.0113563f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_110_47#_M1003_g N_X_c_415_n 0.0113034f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_110_47#_c_120_n N_X_c_415_n 0.00232005f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_146 N_A_110_47#_c_123_n N_X_c_415_n 0.0385727f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_110_47#_M1008_g N_X_c_394_n 0.00120255f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_110_47#_M1010_g N_X_c_394_n 0.00120255f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_110_47#_M1010_g N_X_c_395_n 0.0122792f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_110_47#_M1014_g N_X_c_395_n 0.0122792f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A_110_47#_c_120_n N_X_c_395_n 0.00267078f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_152 N_A_110_47#_c_123_n N_X_c_395_n 0.0429599f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_110_47#_M1005_g N_X_c_425_n 0.0113432f $X=2.625 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_110_47#_M1009_g N_X_c_425_n 0.0113694f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_110_47#_c_120_n N_X_c_425_n 0.00232005f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_156 N_A_110_47#_c_123_n N_X_c_425_n 0.0385727f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_110_47#_M1014_g N_X_c_396_n 0.00120255f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_110_47#_M1016_g N_X_c_396_n 0.00120255f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_110_47#_M1016_g N_X_c_397_n 0.0122792f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_110_47#_c_120_n N_X_c_397_n 0.00320502f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_161 N_A_110_47#_c_123_n N_X_c_397_n 0.0133842f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_110_47#_M1011_g N_X_c_434_n 0.0113694f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_110_47#_c_120_n N_X_c_434_n 0.00278134f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_164 N_A_110_47#_c_123_n N_X_c_434_n 0.0121568f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_110_47#_M1017_g N_X_c_398_n 0.00120255f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_110_47#_M1019_g N_X_c_398_n 0.00221636f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A_110_47#_M1000_g N_X_c_439_n 0.00112492f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_110_47#_M1002_g N_X_c_439_n 0.00112492f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_110_47#_c_120_n N_X_c_439_n 0.00238948f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_170 N_A_110_47#_c_123_n N_X_c_439_n 0.0168441f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_110_47#_c_120_n N_X_c_399_n 0.00277135f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_172 N_A_110_47#_c_123_n N_X_c_399_n 0.0213686f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_110_47#_M1003_g N_X_c_445_n 0.00112492f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_110_47#_M1005_g N_X_c_445_n 0.00112341f $X=2.625 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_110_47#_c_120_n N_X_c_445_n 0.00238948f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_176 N_A_110_47#_c_123_n N_X_c_445_n 0.0168441f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_110_47#_c_120_n N_X_c_400_n 0.00277135f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_178 N_A_110_47#_c_123_n N_X_c_400_n 0.0213686f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_110_47#_M1009_g N_X_c_451_n 0.00112341f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_110_47#_M1011_g N_X_c_451_n 0.00112492f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_110_47#_c_120_n N_X_c_451_n 0.00238948f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_182 N_A_110_47#_c_123_n N_X_c_451_n 0.0168441f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_110_47#_M1016_g X 0.00116814f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_110_47#_M1011_g X 0.00448672f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_110_47#_M1017_g X 0.0116551f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_110_47#_M1013_g X 0.0053012f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_110_47#_c_120_n X 0.0458412f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_188 N_A_110_47#_M1019_g X 0.0136957f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_110_47#_M1015_g X 0.00773738f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_110_47#_c_123_n X 0.0208936f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_110_47#_M1013_g X 0.0108558f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_110_47#_M1015_g X 0.0128711f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_110_47#_M1001_g N_VGND_c_546_n 0.00168046f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_110_47#_c_123_n N_VGND_c_546_n 0.00869033f $X=3.245 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_110_47#_M1006_g N_VGND_c_547_n 0.00161372f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A_110_47#_M1008_g N_VGND_c_547_n 0.00161372f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_197 N_A_110_47#_M1010_g N_VGND_c_548_n 0.00161372f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_198 N_A_110_47#_M1014_g N_VGND_c_548_n 0.00161372f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_199 N_A_110_47#_M1016_g N_VGND_c_549_n 0.00161372f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_A_110_47#_M1017_g N_VGND_c_549_n 0.00161372f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_110_47#_M1019_g N_VGND_c_550_n 0.00341923f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_110_47#_M1001_g N_VGND_c_551_n 0.00585385f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_110_47#_M1006_g N_VGND_c_551_n 0.00439206f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_110_47#_M1008_g N_VGND_c_553_n 0.00439206f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_110_47#_M1010_g N_VGND_c_553_n 0.00439206f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_110_47#_M1014_g N_VGND_c_555_n 0.00439206f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_110_47#_M1016_g N_VGND_c_555_n 0.00439206f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_110_47#_M1017_g N_VGND_c_557_n 0.00439071f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_110_47#_M1019_g N_VGND_c_557_n 0.00439071f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_210 N_A_110_47#_c_122_n N_VGND_c_559_n 0.0137163f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_110_47#_M1004_d N_VGND_c_561_n 0.00336236f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_212 N_A_110_47#_M1001_g N_VGND_c_561_n 0.0106694f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_213 N_A_110_47#_M1006_g N_VGND_c_561_n 0.00590932f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_214 N_A_110_47#_M1008_g N_VGND_c_561_n 0.00590932f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_110_47#_M1010_g N_VGND_c_561_n 0.00590932f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_110_47#_M1014_g N_VGND_c_561_n 0.00590932f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_110_47#_M1016_g N_VGND_c_561_n 0.00590932f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_110_47#_M1017_g N_VGND_c_561_n 0.00590684f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_A_110_47#_M1019_g N_VGND_c_561_n 0.00700101f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_110_47#_c_122_n N_VGND_c_561_n 0.00950576f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_110_47#_M1000_g N_VPWR_c_629_n 0.00585385f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_110_47#_M1002_g N_VPWR_c_629_n 0.00585385f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_110_47#_M1003_g N_VPWR_c_629_n 0.00585385f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_110_47#_M1005_g N_VPWR_c_629_n 0.00585385f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_110_47#_M1009_g N_VPWR_c_629_n 0.00585385f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_110_47#_M1011_g N_VPWR_c_629_n 0.00585385f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_110_47#_M1013_g N_VPWR_c_629_n 0.00585385f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_110_47#_M1015_g N_VPWR_c_629_n 0.00585385f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_110_47#_c_133_n N_VPWR_c_629_n 0.0141362f $X=0.69 $Y=1.69 $X2=0 $Y2=0
cc_230 N_A_110_47#_M1007_d N_VPWR_c_628_n 0.00127217f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_231 N_A_110_47#_M1000_g N_VPWR_c_628_n 0.00531811f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_110_47#_M1002_g N_VPWR_c_628_n 0.0052918f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_110_47#_M1003_g N_VPWR_c_628_n 0.0052918f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_110_47#_M1005_g N_VPWR_c_628_n 0.0052918f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_110_47#_M1009_g N_VPWR_c_628_n 0.0052918f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_110_47#_M1011_g N_VPWR_c_628_n 0.0052918f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_110_47#_M1013_g N_VPWR_c_628_n 0.0052918f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_110_47#_M1015_g N_VPWR_c_628_n 0.00642806f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A_110_47#_c_133_n N_VPWR_c_628_n 0.00231204f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_240 N_KAPWR_c_302_n N_X_M1000_d 4.89441e-19 $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_241 N_KAPWR_c_307_n N_X_M1003_d 2.61752e-19 $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_242 N_KAPWR_c_312_n N_X_M1009_d 2.61752e-19 $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_243 N_KAPWR_c_316_n N_X_M1013_d 2.61539e-19 $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_244 N_KAPWR_M1002_s N_X_c_415_n 0.00325489f $X=1.84 $Y=1.485 $X2=0 $Y2=0
cc_245 N_KAPWR_c_300_n N_X_c_415_n 0.0128604f $X=1.975 $Y=2.21 $X2=0 $Y2=0
cc_246 N_KAPWR_c_302_n N_X_c_415_n 0.00466059f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_247 N_KAPWR_c_304_n N_X_c_415_n 0.00245411f $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_248 N_KAPWR_c_307_n N_X_c_415_n 0.00497471f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_249 N_KAPWR_M1005_s N_X_c_425_n 0.00325883f $X=2.7 $Y=1.485 $X2=0 $Y2=0
cc_250 N_KAPWR_c_305_n N_X_c_425_n 0.0127908f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_251 N_KAPWR_c_307_n N_X_c_425_n 0.00434646f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_252 N_KAPWR_c_309_n N_X_c_425_n 0.0023936f $X=2.97 $Y=2.21 $X2=0 $Y2=0
cc_253 N_KAPWR_c_312_n N_X_c_425_n 0.00532372f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_254 N_KAPWR_M1011_s N_X_c_434_n 0.0035494f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_255 N_KAPWR_c_310_n N_X_c_434_n 0.0110447f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_256 N_KAPWR_c_312_n N_X_c_434_n 0.00497471f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_257 N_KAPWR_c_314_n N_X_c_434_n 0.00136985f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_258 N_KAPWR_c_290_n N_X_c_439_n 0.00152822f $X=1.265 $Y=2.21 $X2=0 $Y2=0
cc_259 N_KAPWR_c_300_n N_X_c_439_n 0.00822181f $X=1.975 $Y=2.21 $X2=0 $Y2=0
cc_260 N_KAPWR_c_302_n N_X_c_439_n 0.0260313f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_261 N_KAPWR_c_304_n N_X_c_439_n 0.00153797f $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_262 N_KAPWR_c_294_n N_X_c_439_n 0.00822181f $X=1.12 $Y=1.69 $X2=0 $Y2=0
cc_263 N_KAPWR_c_300_n N_X_c_445_n 0.00822181f $X=1.975 $Y=2.21 $X2=0 $Y2=0
cc_264 N_KAPWR_c_304_n N_X_c_445_n 7.53589e-19 $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_265 N_KAPWR_c_305_n N_X_c_445_n 0.0082718f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_266 N_KAPWR_c_307_n N_X_c_445_n 0.0260214f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_267 N_KAPWR_c_309_n N_X_c_445_n 6.95463e-19 $X=2.97 $Y=2.21 $X2=0 $Y2=0
cc_268 N_KAPWR_c_305_n N_X_c_451_n 0.0082718f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_269 N_KAPWR_c_309_n N_X_c_451_n 4.70067e-19 $X=2.97 $Y=2.21 $X2=0 $Y2=0
cc_270 N_KAPWR_c_310_n N_X_c_451_n 0.00822181f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_271 N_KAPWR_c_312_n N_X_c_451_n 0.0260214f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_272 N_KAPWR_c_314_n N_X_c_451_n 0.00175189f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_273 N_KAPWR_M1011_s X 2.31797e-19 $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_274 N_KAPWR_M1015_s X 0.00332068f $X=4.42 $Y=1.485 $X2=0 $Y2=0
cc_275 N_KAPWR_c_310_n X 0.0101047f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_276 N_KAPWR_c_314_n X 0.00274884f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_277 N_KAPWR_c_284_n X 0.00408548f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_278 N_KAPWR_c_285_n X 0.0290295f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_279 N_KAPWR_c_316_n X 0.0369801f $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_280 N_KAPWR_c_283_n N_VPWR_c_629_n 0.0012443f $X=0.405 $Y=2.24 $X2=0 $Y2=0
cc_281 N_KAPWR_c_288_n N_VPWR_c_629_n 0.00102631f $X=0.975 $Y=2.21 $X2=0 $Y2=0
cc_282 N_KAPWR_c_290_n N_VPWR_c_629_n 0.00102914f $X=1.265 $Y=2.21 $X2=0 $Y2=0
cc_283 N_KAPWR_c_300_n N_VPWR_c_629_n 0.0147733f $X=1.975 $Y=2.21 $X2=0 $Y2=0
cc_284 N_KAPWR_c_302_n N_VPWR_c_629_n 0.00102995f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_285 N_KAPWR_c_304_n N_VPWR_c_629_n 0.00102658f $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_286 N_KAPWR_c_305_n N_VPWR_c_629_n 0.0147484f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_287 N_KAPWR_c_307_n N_VPWR_c_629_n 0.00102756f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_288 N_KAPWR_c_310_n N_VPWR_c_629_n 0.0147733f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_289 N_KAPWR_c_312_n N_VPWR_c_629_n 0.00187779f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_290 N_KAPWR_c_314_n N_VPWR_c_629_n 0.00102581f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_291 N_KAPWR_c_284_n N_VPWR_c_629_n 0.00141328f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_292 N_KAPWR_c_285_n N_VPWR_c_629_n 0.0188086f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_293 N_KAPWR_c_316_n N_VPWR_c_629_n 0.00103071f $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_294 N_KAPWR_c_286_n N_VPWR_c_629_n 0.0190549f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_295 N_KAPWR_c_294_n N_VPWR_c_629_n 0.0149375f $X=1.12 $Y=1.69 $X2=0 $Y2=0
cc_296 N_KAPWR_M1007_s N_VPWR_c_628_n 0.00114006f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_297 N_KAPWR_M1018_s N_VPWR_c_628_n 0.00123133f $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_298 N_KAPWR_M1002_s N_VPWR_c_628_n 0.00123133f $X=1.84 $Y=1.485 $X2=0 $Y2=0
cc_299 N_KAPWR_M1005_s N_VPWR_c_628_n 0.00122337f $X=2.7 $Y=1.485 $X2=0 $Y2=0
cc_300 N_KAPWR_M1011_s N_VPWR_c_628_n 0.00123133f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_301 N_KAPWR_M1015_s N_VPWR_c_628_n 0.00114006f $X=4.42 $Y=1.485 $X2=0 $Y2=0
cc_302 N_KAPWR_c_283_n N_VPWR_c_628_n 0.507437f $X=0.405 $Y=2.24 $X2=0 $Y2=0
cc_303 N_KAPWR_c_300_n N_VPWR_c_628_n 0.00234462f $X=1.975 $Y=2.21 $X2=0 $Y2=0
cc_304 N_KAPWR_c_305_n N_VPWR_c_628_n 0.00236391f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_305 N_KAPWR_c_310_n N_VPWR_c_628_n 0.00234462f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_306 N_KAPWR_c_285_n N_VPWR_c_628_n 0.00266268f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_307 N_KAPWR_c_286_n N_VPWR_c_628_n 0.00271943f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_308 N_KAPWR_c_294_n N_VPWR_c_628_n 0.00239458f $X=1.12 $Y=1.69 $X2=0 $Y2=0
cc_309 N_X_c_392_n N_VGND_c_547_n 0.0164628f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_310 N_X_c_395_n N_VGND_c_548_n 0.0164628f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_311 N_X_c_397_n N_VGND_c_549_n 0.0129787f $X=3.76 $Y=0.82 $X2=0 $Y2=0
cc_312 X N_VGND_c_549_n 0.00403581f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_313 X N_VGND_c_550_n 0.0243348f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_314 N_X_c_391_n N_VGND_c_551_n 0.0128416f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_315 N_X_c_392_n N_VGND_c_551_n 0.00224999f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_316 N_X_c_392_n N_VGND_c_553_n 0.00224999f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_317 N_X_c_394_n N_VGND_c_553_n 0.0128416f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_318 N_X_c_395_n N_VGND_c_553_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_319 N_X_c_395_n N_VGND_c_555_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_320 N_X_c_396_n N_VGND_c_555_n 0.0128416f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_321 N_X_c_397_n N_VGND_c_555_n 0.00224999f $X=3.76 $Y=0.82 $X2=0 $Y2=0
cc_322 N_X_c_398_n N_VGND_c_557_n 0.0129027f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_323 X N_VGND_c_557_n 0.00498855f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_324 N_X_M1001_s N_VGND_c_561_n 0.00268444f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_325 N_X_M1008_s N_VGND_c_561_n 0.00234574f $X=2.27 $Y=0.235 $X2=0 $Y2=0
cc_326 N_X_M1014_s N_VGND_c_561_n 0.00234574f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_M1017_s N_VGND_c_561_n 0.00234544f $X=3.99 $Y=0.235 $X2=0 $Y2=0
cc_328 N_X_c_391_n N_VGND_c_561_n 0.00979224f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_329 N_X_c_392_n N_VGND_c_561_n 0.00829353f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_330 N_X_c_394_n N_VGND_c_561_n 0.00979224f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_331 N_X_c_395_n N_VGND_c_561_n 0.00829353f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_332 N_X_c_396_n N_VGND_c_561_n 0.00979224f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_333 N_X_c_397_n N_VGND_c_561_n 0.00436967f $X=3.76 $Y=0.82 $X2=0 $Y2=0
cc_334 N_X_c_398_n N_VGND_c_561_n 0.00981584f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_335 X N_VGND_c_561_n 0.00944699f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_336 N_X_c_439_n N_VPWR_c_629_n 0.0144808f $X=1.55 $Y=1.69 $X2=0 $Y2=0
cc_337 N_X_c_445_n N_VPWR_c_629_n 0.0144808f $X=2.41 $Y=1.69 $X2=0 $Y2=0
cc_338 N_X_c_451_n N_VPWR_c_629_n 0.0144808f $X=3.27 $Y=1.69 $X2=0 $Y2=0
cc_339 X N_VPWR_c_629_n 0.0144808f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_340 N_X_M1000_d N_VPWR_c_628_n 0.00123188f $X=1.41 $Y=1.485 $X2=0 $Y2=0
cc_341 N_X_M1003_d N_VPWR_c_628_n 0.00123188f $X=2.27 $Y=1.485 $X2=0 $Y2=0
cc_342 N_X_M1009_d N_VPWR_c_628_n 0.00123188f $X=3.13 $Y=1.485 $X2=0 $Y2=0
cc_343 N_X_M1013_d N_VPWR_c_628_n 0.00123188f $X=3.99 $Y=1.485 $X2=0 $Y2=0
cc_344 N_X_c_439_n N_VPWR_c_628_n 0.00240527f $X=1.55 $Y=1.69 $X2=0 $Y2=0
cc_345 N_X_c_445_n N_VPWR_c_628_n 0.00240527f $X=2.41 $Y=1.69 $X2=0 $Y2=0
cc_346 N_X_c_451_n N_VPWR_c_628_n 0.00240527f $X=3.27 $Y=1.69 $X2=0 $Y2=0
cc_347 X N_VPWR_c_628_n 0.00240527f $X=3.825 $Y=1.445 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dfbbn_2.spice.SKY130_FD_SC_HD__DFBBN_2.pxi
* Created: Thu Aug 27 14:14:05 2020
* 
x_PM_SKY130_FD_SC_HD__DFBBN_2%CLK_N N_CLK_N_c_268_n N_CLK_N_c_263_n
+ N_CLK_N_M1038_g N_CLK_N_c_269_n N_CLK_N_M1023_g N_CLK_N_c_264_n
+ N_CLK_N_c_270_n CLK_N CLK_N N_CLK_N_c_266_n N_CLK_N_c_267_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%CLK_N
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_27_47# N_A_27_47#_M1038_s N_A_27_47#_M1023_s
+ N_A_27_47#_M1025_g N_A_27_47#_M1000_g N_A_27_47#_M1018_g N_A_27_47#_c_309_n
+ N_A_27_47#_c_310_n N_A_27_47#_M1006_g N_A_27_47#_c_312_n N_A_27_47#_c_313_n
+ N_A_27_47#_M1007_g N_A_27_47#_M1019_g N_A_27_47#_c_314_n N_A_27_47#_c_315_n
+ N_A_27_47#_c_316_n N_A_27_47#_c_336_n N_A_27_47#_c_317_n N_A_27_47#_c_318_n
+ N_A_27_47#_c_319_n N_A_27_47#_c_337_n N_A_27_47#_c_338_n N_A_27_47#_c_339_n
+ N_A_27_47#_c_320_n N_A_27_47#_c_321_n N_A_27_47#_c_322_n N_A_27_47#_c_323_n
+ N_A_27_47#_c_324_n N_A_27_47#_c_325_n N_A_27_47#_c_326_n N_A_27_47#_c_327_n
+ N_A_27_47#_c_328_n N_A_27_47#_c_329_n N_A_27_47#_c_330_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%D N_D_M1011_g N_D_M1029_g D D N_D_c_570_n
+ N_D_c_571_n PM_SKY130_FD_SC_HD__DFBBN_2%D
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_193_47# N_A_193_47#_M1025_d N_A_193_47#_M1000_d
+ N_A_193_47#_c_610_n N_A_193_47#_M1036_g N_A_193_47#_M1009_g
+ N_A_193_47#_M1031_g N_A_193_47#_c_611_n N_A_193_47#_c_612_n
+ N_A_193_47#_M1004_g N_A_193_47#_c_614_n N_A_193_47#_c_615_n
+ N_A_193_47#_c_622_n N_A_193_47#_c_623_n N_A_193_47#_c_624_n
+ N_A_193_47#_c_625_n N_A_193_47#_c_626_n N_A_193_47#_c_627_n
+ N_A_193_47#_c_628_n N_A_193_47#_c_629_n N_A_193_47#_c_630_n
+ N_A_193_47#_c_631_n N_A_193_47#_c_616_n PM_SKY130_FD_SC_HD__DFBBN_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_650_21# N_A_650_21#_M1035_d N_A_650_21#_M1041_d
+ N_A_650_21#_M1012_g N_A_650_21#_M1015_g N_A_650_21#_M1028_g
+ N_A_650_21#_c_813_n N_A_650_21#_M1021_g N_A_650_21#_c_822_n
+ N_A_650_21#_c_869_p N_A_650_21#_c_834_n N_A_650_21#_c_814_n
+ N_A_650_21#_c_815_n N_A_650_21#_c_816_n N_A_650_21#_c_824_n
+ N_A_650_21#_c_825_n N_A_650_21#_c_839_n N_A_650_21#_c_817_n
+ N_A_650_21#_c_818_n PM_SKY130_FD_SC_HD__DFBBN_2%A_650_21#
x_PM_SKY130_FD_SC_HD__DFBBN_2%SET_B N_SET_B_c_957_n N_SET_B_M1041_g
+ N_SET_B_M1037_g N_SET_B_M1005_g N_SET_B_M1013_g SET_B N_SET_B_c_963_n
+ N_SET_B_c_964_n N_SET_B_c_965_n N_SET_B_c_966_n N_SET_B_c_967_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%SET_B
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_476_47# N_A_476_47#_M1036_d N_A_476_47#_M1018_d
+ N_A_476_47#_M1035_g N_A_476_47#_M1020_g N_A_476_47#_c_1099_n
+ N_A_476_47#_c_1100_n N_A_476_47#_c_1094_n N_A_476_47#_c_1089_n
+ N_A_476_47#_c_1090_n N_A_476_47#_c_1091_n N_A_476_47#_c_1092_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_476_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_944_21# N_A_944_21#_M1027_s N_A_944_21#_M1001_s
+ N_A_944_21#_M1042_g N_A_944_21#_M1032_g N_A_944_21#_M1043_g
+ N_A_944_21#_M1016_g N_A_944_21#_c_1195_n N_A_944_21#_c_1196_n
+ N_A_944_21#_c_1204_n N_A_944_21#_c_1205_n N_A_944_21#_c_1197_n
+ N_A_944_21#_c_1198_n N_A_944_21#_c_1199_n N_A_944_21#_c_1208_n
+ N_A_944_21#_c_1209_n N_A_944_21#_c_1210_n N_A_944_21#_c_1211_n
+ N_A_944_21#_c_1200_n N_A_944_21#_c_1201_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_944_21#
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_1431_21# N_A_1431_21#_M1008_d
+ N_A_1431_21#_M1013_d N_A_1431_21#_M1024_g N_A_1431_21#_M1034_g
+ N_A_1431_21#_c_1352_n N_A_1431_21#_M1003_g N_A_1431_21#_M1014_g
+ N_A_1431_21#_M1022_g N_A_1431_21#_M1030_g N_A_1431_21#_c_1355_n
+ N_A_1431_21#_c_1356_n N_A_1431_21#_c_1357_n N_A_1431_21#_c_1358_n
+ N_A_1431_21#_c_1359_n N_A_1431_21#_M1017_g N_A_1431_21#_c_1370_n
+ N_A_1431_21#_M1026_g N_A_1431_21#_c_1360_n N_A_1431_21#_c_1361_n
+ N_A_1431_21#_c_1371_n N_A_1431_21#_c_1372_n N_A_1431_21#_c_1373_n
+ N_A_1431_21#_c_1374_n N_A_1431_21#_c_1429_p N_A_1431_21#_c_1483_p
+ N_A_1431_21#_c_1400_n N_A_1431_21#_c_1362_n N_A_1431_21#_c_1376_n
+ N_A_1431_21#_c_1377_n N_A_1431_21#_c_1417_n N_A_1431_21#_c_1393_n
+ N_A_1431_21#_c_1420_n N_A_1431_21#_c_1363_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_1431_21#
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_1257_47# N_A_1257_47#_M1007_d
+ N_A_1257_47#_M1031_d N_A_1257_47#_M1008_g N_A_1257_47#_M1039_g
+ N_A_1257_47#_c_1559_n N_A_1257_47#_c_1562_n N_A_1257_47#_c_1548_n
+ N_A_1257_47#_c_1554_n N_A_1257_47#_c_1549_n N_A_1257_47#_c_1550_n
+ N_A_1257_47#_c_1551_n N_A_1257_47#_c_1552_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_1257_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%RESET_B N_RESET_B_M1027_g N_RESET_B_M1001_g
+ RESET_B N_RESET_B_c_1648_n PM_SKY130_FD_SC_HD__DFBBN_2%RESET_B
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_2236_47# N_A_2236_47#_M1017_s
+ N_A_2236_47#_M1026_s N_A_2236_47#_c_1682_n N_A_2236_47#_M1033_g
+ N_A_2236_47#_M1002_g N_A_2236_47#_c_1683_n N_A_2236_47#_M1040_g
+ N_A_2236_47#_M1010_g N_A_2236_47#_c_1684_n N_A_2236_47#_c_1690_n
+ N_A_2236_47#_c_1685_n N_A_2236_47#_c_1686_n N_A_2236_47#_c_1687_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_2236_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%VPWR N_VPWR_M1023_d N_VPWR_M1029_s N_VPWR_M1015_d
+ N_VPWR_M1032_d N_VPWR_M1034_d N_VPWR_M1043_d N_VPWR_M1001_d N_VPWR_M1030_s
+ N_VPWR_M1026_d N_VPWR_M1010_d N_VPWR_c_1755_n N_VPWR_c_1756_n N_VPWR_c_1757_n
+ N_VPWR_c_1758_n N_VPWR_c_1759_n N_VPWR_c_1760_n N_VPWR_c_1761_n
+ N_VPWR_c_1762_n N_VPWR_c_1763_n N_VPWR_c_1764_n N_VPWR_c_1765_n
+ N_VPWR_c_1766_n N_VPWR_c_1767_n VPWR VPWR N_VPWR_c_1768_n N_VPWR_c_1769_n
+ N_VPWR_c_1770_n N_VPWR_c_1771_n N_VPWR_c_1772_n N_VPWR_c_1773_n
+ N_VPWR_c_1774_n N_VPWR_c_1775_n N_VPWR_c_1776_n N_VPWR_c_1777_n
+ N_VPWR_c_1778_n N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n
+ N_VPWR_c_1754_n VPWR PM_SKY130_FD_SC_HD__DFBBN_2%VPWR
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_381_47# N_A_381_47#_M1011_d N_A_381_47#_M1029_d
+ N_A_381_47#_c_1955_n N_A_381_47#_c_1956_n N_A_381_47#_c_1957_n
+ N_A_381_47#_c_1959_n N_A_381_47#_c_1960_n N_A_381_47#_c_1990_n
+ N_A_381_47#_c_1961_n PM_SKY130_FD_SC_HD__DFBBN_2%A_381_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%Q_N N_Q_N_M1003_s N_Q_N_M1014_d N_Q_N_c_2032_n
+ N_Q_N_c_2030_n Q_N Q_N Q_N N_Q_N_c_2043_n Q_N PM_SKY130_FD_SC_HD__DFBBN_2%Q_N
x_PM_SKY130_FD_SC_HD__DFBBN_2%Q N_Q_M1033_d N_Q_M1002_s N_Q_c_2056_n
+ N_Q_c_2054_n N_Q_c_2053_n Q Q Q PM_SKY130_FD_SC_HD__DFBBN_2%Q
x_PM_SKY130_FD_SC_HD__DFBBN_2%VGND N_VGND_M1038_d N_VGND_M1011_s N_VGND_M1012_d
+ N_VGND_M1021_s N_VGND_M1024_d N_VGND_M1027_d N_VGND_M1022_d N_VGND_M1017_d
+ N_VGND_M1040_s N_VGND_c_2075_n N_VGND_c_2076_n N_VGND_c_2077_n N_VGND_c_2078_n
+ N_VGND_c_2079_n N_VGND_c_2080_n N_VGND_c_2081_n N_VGND_c_2082_n
+ N_VGND_c_2083_n N_VGND_c_2084_n N_VGND_c_2085_n N_VGND_c_2086_n
+ N_VGND_c_2087_n N_VGND_c_2088_n N_VGND_c_2089_n N_VGND_c_2090_n
+ N_VGND_c_2091_n VGND VGND N_VGND_c_2092_n VGND N_VGND_c_2093_n N_VGND_c_2094_n
+ N_VGND_c_2095_n N_VGND_c_2096_n N_VGND_c_2097_n N_VGND_c_2098_n
+ N_VGND_c_2099_n N_VGND_c_2100_n N_VGND_c_2101_n N_VGND_c_2102_n VGND
+ PM_SKY130_FD_SC_HD__DFBBN_2%VGND
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_790_47# N_A_790_47#_M1037_d N_A_790_47#_M1042_d
+ N_A_790_47#_c_2285_n N_A_790_47#_c_2286_n N_A_790_47#_c_2297_n
+ PM_SKY130_FD_SC_HD__DFBBN_2%A_790_47#
x_PM_SKY130_FD_SC_HD__DFBBN_2%A_1547_47# N_A_1547_47#_M1005_d
+ N_A_1547_47#_M1016_d N_A_1547_47#_c_2322_n N_A_1547_47#_c_2318_n
+ N_A_1547_47#_c_2323_n PM_SKY130_FD_SC_HD__DFBBN_2%A_1547_47#
cc_1 VNB N_CLK_N_c_263_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_N_c_264_n 0.0229857f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK_N 0.0161955f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_CLK_N_c_266_n 0.0197972f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_CLK_N_c_267_n 0.0141141f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1025_g 0.0382529f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_309_n 0.0133502f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_c_310_n 0.00435992f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_9 VNB N_A_27_47#_M1006_g 0.0198711f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_10 VNB N_A_27_47#_c_312_n 0.00878653f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_11 VNB N_A_27_47#_c_313_n 0.018063f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_12 VNB N_A_27_47#_c_314_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_315_n 9.27212e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_316_n 0.00789919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_317_n 0.00302353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_318_n 0.0315468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_319_n 0.00458399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_320_n 0.0249608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_321_n 0.00430479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_322_n 0.00124359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_323_n 0.0216332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_324_n 0.00235584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_325_n 0.00292248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_326_n 0.00201153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_327_n 0.00493055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_328_n 0.00147534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_329_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_330_n 0.0249207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_D_M1011_g 0.0338938f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_30 VNB N_D_c_570_n 0.0258509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_D_c_571_n 0.00430425f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_32 VNB N_A_193_47#_c_610_n 0.0179685f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_33 VNB N_A_193_47#_c_611_n 0.0124337f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_34 VNB N_A_193_47#_c_612_n 0.00338665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_M1004_g 0.0470935f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_36 VNB N_A_193_47#_c_614_n 0.00432857f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.19
cc_37 VNB N_A_193_47#_c_615_n 0.0315548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_616_n 0.0164942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_650_21#_M1012_g 0.0393082f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_40 VNB N_A_650_21#_c_813_n 0.0192786f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_41 VNB N_A_650_21#_c_814_n 0.00190301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_650_21#_c_815_n 0.00419895f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_43 VNB N_A_650_21#_c_816_n 0.0109044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_650_21#_c_817_n 0.00589338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_650_21#_c_818_n 0.0321818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_SET_B_c_957_n 0.031114f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_47 VNB N_SET_B_M1041_g 0.00696335f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_48 VNB N_SET_B_M1037_g 0.0204338f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_49 VNB N_SET_B_M1005_g 0.0200444f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_50 VNB N_SET_B_M1013_g 0.00793898f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_51 VNB SET_B 0.00769431f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_52 VNB N_SET_B_c_963_n 0.0150191f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_53 VNB N_SET_B_c_964_n 0.00178135f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_54 VNB N_SET_B_c_965_n 0.00209085f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_55 VNB N_SET_B_c_966_n 0.00538514f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_56 VNB N_SET_B_c_967_n 0.0316983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_476_47#_M1035_g 0.0259951f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_58 VNB N_A_476_47#_c_1089_n 0.00755759f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_59 VNB N_A_476_47#_c_1090_n 0.00778508f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_60 VNB N_A_476_47#_c_1091_n 0.0040045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_476_47#_c_1092_n 0.0141708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_944_21#_M1042_g 0.0293266f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_63 VNB N_A_944_21#_M1016_g 0.0279621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_944_21#_c_1195_n 0.0113702f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_65 VNB N_A_944_21#_c_1196_n 0.00176384f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_66 VNB N_A_944_21#_c_1197_n 0.00662861f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_67 VNB N_A_944_21#_c_1198_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_944_21#_c_1199_n 0.0213679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_944_21#_c_1200_n 0.0193899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_944_21#_c_1201_n 0.00516932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1431_21#_M1024_g 0.0441996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_72 VNB N_A_1431_21#_c_1352_n 0.0165362f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_73 VNB N_A_1431_21#_M1022_g 0.021473f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_74 VNB N_A_1431_21#_M1030_g 5.33203e-19 $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.19
cc_75 VNB N_A_1431_21#_c_1355_n 0.0607006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1431_21#_c_1356_n 0.0331492f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_77 VNB N_A_1431_21#_c_1357_n 0.00814182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1431_21#_c_1358_n 4.88264e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1431_21#_c_1359_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1431_21#_c_1360_n 0.0184739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1431_21#_c_1361_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1431_21#_c_1362_n 0.00321658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1431_21#_c_1363_n 0.00365923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1257_47#_M1008_g 0.0224258f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_85 VNB N_A_1257_47#_c_1548_n 0.0117849f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_86 VNB N_A_1257_47#_c_1549_n 0.0114143f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_87 VNB N_A_1257_47#_c_1550_n 4.91252e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1257_47#_c_1551_n 0.00186712f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_89 VNB N_A_1257_47#_c_1552_n 0.017672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_RESET_B_M1027_g 0.0350169f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_91 VNB RESET_B 0.00385601f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_92 VNB N_RESET_B_c_1648_n 0.0299154f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_93 VNB N_A_2236_47#_c_1682_n 0.0168966f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_94 VNB N_A_2236_47#_c_1683_n 0.0215106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2236_47#_c_1684_n 0.00521072f $X=-0.19 $Y=-0.24 $X2=0.242
+ $Y2=1.235
cc_96 VNB N_A_2236_47#_c_1685_n 0.0051319f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_97 VNB N_A_2236_47#_c_1686_n 6.65975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_2236_47#_c_1687_n 0.0519216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VPWR_c_1754_n 0.535415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_381_47#_c_1955_n 0.00964401f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_101 VNB N_A_381_47#_c_1956_n 0.0042849f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_102 VNB N_A_381_47#_c_1957_n 0.00297622f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_103 VNB N_Q_N_c_2030_n 0.00127808f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_104 VNB N_Q_c_2053_n 0.00102326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_2075_n 4.10922e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_2076_n 0.00510315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2077_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2078_n 0.00541886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2079_n 0.0024154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2080_n 0.00550287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2081_n 0.00678097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2082_n 0.020975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2083_n 0.00254068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2084_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2085_n 0.0335145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2086_n 0.0443619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2087_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2088_n 0.0384102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2089_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2090_n 0.0404697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2091_n 0.00372951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2092_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2093_n 0.0161167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2094_n 0.0547685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2095_n 0.015741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2096_n 0.0147637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2097_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2098_n 0.00526381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2099_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2100_n 0.00442399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2101_n 0.00440331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2102_n 0.600481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_A_790_47#_c_2285_n 0.00181668f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_134 VNB N_A_790_47#_c_2286_n 0.00425766f $X=-0.19 $Y=-0.24 $X2=0.305
+ $Y2=0.805
cc_135 VPB N_CLK_N_c_268_n 0.0118724f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_136 VPB N_CLK_N_c_269_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_137 VPB N_CLK_N_c_270_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_138 VPB CLK_N 0.0152683f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_139 VPB N_CLK_N_c_266_n 0.0102819f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_140 VPB N_A_27_47#_M1000_g 0.0362832f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_141 VPB N_A_27_47#_M1018_g 0.046414f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_142 VPB N_A_27_47#_c_309_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_143 VPB N_A_27_47#_c_310_n 0.00326624f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_144 VPB N_A_27_47#_M1019_g 0.0222026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_336_n 0.00205657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_337_n 0.00384216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_338_n 0.0287783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_27_47#_c_339_n 0.0299356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_325_n 0.00320885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_27_47#_c_328_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_27_47#_c_329_n 0.0115872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_D_M1029_g 0.0544931f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_153 VPB N_D_c_570_n 0.00539635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_D_c_571_n 0.00442628f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_155 VPB N_A_193_47#_M1009_g 0.0215879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_193_47#_M1031_g 0.020906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_193_47#_c_611_n 0.0178865f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_158 VPB N_A_193_47#_c_612_n 0.00403646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_193_47#_c_614_n 0.00245106f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.19
cc_160 VPB N_A_193_47#_c_622_n 0.00948586f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.53
cc_161 VPB N_A_193_47#_c_623_n 0.00448953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_193_47#_c_624_n 0.00875464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_193_47#_c_625_n 0.00166689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_193_47#_c_626_n 0.00361706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_193_47#_c_627_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_193_47#_c_628_n 0.00575214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_193_47#_c_629_n 0.0282388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_193_47#_c_630_n 0.00514398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_193_47#_c_631_n 0.0125285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_193_47#_c_616_n 0.0179362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_650_21#_M1012_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_172 VPB N_A_650_21#_M1015_g 0.0210587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_173 VPB N_A_650_21#_M1028_g 0.0318679f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_174 VPB N_A_650_21#_c_822_n 0.0055347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_650_21#_c_815_n 0.00618914f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.53
cc_176 VPB N_A_650_21#_c_824_n 0.00575673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_650_21#_c_825_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_650_21#_c_818_n 0.00659461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_SET_B_M1041_g 0.0508831f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_180 VPB N_SET_B_M1013_g 0.0496547f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_181 VPB N_A_476_47#_M1020_g 0.0201414f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_182 VPB N_A_476_47#_c_1094_n 0.0121994f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_183 VPB N_A_476_47#_c_1090_n 0.00799914f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_184 VPB N_A_476_47#_c_1091_n 0.00260739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_476_47#_c_1092_n 0.0165426f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_944_21#_M1032_g 0.0212617f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_187 VPB N_A_944_21#_M1043_g 0.0210664f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_188 VPB N_A_944_21#_c_1204_n 0.00188964f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_189 VPB N_A_944_21#_c_1205_n 0.00545735f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_190 VPB N_A_944_21#_c_1198_n 0.00255288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_944_21#_c_1199_n 0.0226279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_944_21#_c_1208_n 0.0329117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_944_21#_c_1209_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_944_21#_c_1210_n 0.00738232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_944_21#_c_1211_n 0.00334233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_944_21#_c_1200_n 0.0260777f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_944_21#_c_1201_n 0.00362741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1431_21#_M1024_g 0.0159543f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_199 VPB N_A_1431_21#_M1034_g 0.021027f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_200 VPB N_A_1431_21#_M1014_g 0.0200318f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_201 VPB N_A_1431_21#_M1030_g 0.0238663f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.19
cc_202 VPB N_A_1431_21#_c_1356_n 0.00453783f $X=-0.19 $Y=1.305 $X2=0.262
+ $Y2=1.53
cc_203 VPB N_A_1431_21#_c_1358_n 0.0133375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1431_21#_c_1370_n 0.0186731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1431_21#_c_1371_n 0.0185133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1431_21#_c_1372_n 0.00421617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_1431_21#_c_1373_n 0.0324865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_1431_21#_c_1374_n 0.00304218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_1431_21#_c_1362_n 0.00331499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_1431_21#_c_1376_n 0.00752745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_A_1431_21#_c_1377_n 0.0015533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1257_47#_M1039_g 0.021833f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_213 VPB N_A_1257_47#_c_1554_n 0.0118251f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_214 VPB N_A_1257_47#_c_1549_n 0.00584496f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_215 VPB N_A_1257_47#_c_1550_n 7.62954e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1257_47#_c_1551_n 0.00126723f $X=-0.19 $Y=1.305 $X2=0.262
+ $Y2=1.53
cc_217 VPB N_A_1257_47#_c_1552_n 0.00899175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_RESET_B_M1001_g 0.0249643f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_219 VPB RESET_B 9.54549e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_220 VPB N_RESET_B_c_1648_n 0.00997209f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_221 VPB N_A_2236_47#_M1002_g 0.02086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_2236_47#_M1010_g 0.0247731f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_223 VPB N_A_2236_47#_c_1690_n 0.00930606f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_224 VPB N_A_2236_47#_c_1685_n 0.00518989f $X=-0.19 $Y=1.305 $X2=0.262
+ $Y2=1.53
cc_225 VPB N_A_2236_47#_c_1686_n 3.32987e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_2236_47#_c_1687_n 0.00966347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1755_n 0.00105975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1756_n 0.00598362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1757_n 0.00313724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1758_n 0.00562936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1759_n 0.00726169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1760_n 0.0213133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1761_n 0.00353439f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1762_n 0.0102689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1763_n 0.0483911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1764_n 0.0292737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1765_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1766_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1767_n 0.022998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1768_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1769_n 0.015989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1770_n 0.0413206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1771_n 0.0591311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1772_n 0.0317596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1773_n 0.0157351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1774_n 0.0147637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1775_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1776_n 0.00527066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1777_n 0.00609488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1778_n 0.00928062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1779_n 0.00456774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1780_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1781_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1754_n 0.0691573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_A_381_47#_c_1955_n 0.00981434f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_256 VPB N_A_381_47#_c_1959_n 0.00962247f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=0.805
cc_257 VPB N_A_381_47#_c_1960_n 0.00326874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_A_381_47#_c_1961_n 0.00183453f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_259 VPB N_Q_N_c_2030_n 0.00118602f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_260 VPB N_Q_c_2054_n 9.72879e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_261 VPB N_Q_c_2053_n 0.00110698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 N_CLK_N_c_263_n N_A_27_47#_M1025_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_263 CLK_N N_A_27_47#_M1025_g 3.10561e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_264 N_CLK_N_c_267_n N_A_27_47#_M1025_g 0.00508036f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_265 N_CLK_N_c_270_n N_A_27_47#_M1000_g 0.0275602f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_266 CLK_N N_A_27_47#_M1000_g 5.74563e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_267 N_CLK_N_c_266_n N_A_27_47#_M1000_g 0.00530931f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_268 N_CLK_N_c_263_n N_A_27_47#_c_315_n 0.00695828f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_269 N_CLK_N_c_264_n N_A_27_47#_c_315_n 0.00787672f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_270 CLK_N N_A_27_47#_c_315_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_271 N_CLK_N_c_264_n N_A_27_47#_c_316_n 0.00615556f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_272 CLK_N N_A_27_47#_c_316_n 0.0224836f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_273 N_CLK_N_c_266_n N_A_27_47#_c_316_n 7.46966e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_274 N_CLK_N_c_269_n N_A_27_47#_c_336_n 0.0128417f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_275 N_CLK_N_c_270_n N_A_27_47#_c_336_n 0.0013816f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_276 CLK_N N_A_27_47#_c_336_n 0.00728212f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_277 N_CLK_N_c_269_n N_A_27_47#_c_339_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_278 N_CLK_N_c_270_n N_A_27_47#_c_339_n 0.00358837f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_279 CLK_N N_A_27_47#_c_339_n 0.0236377f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_280 N_CLK_N_c_266_n N_A_27_47#_c_339_n 5.90345e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_281 N_CLK_N_c_264_n N_A_27_47#_c_321_n 0.00170897f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_282 N_CLK_N_c_267_n N_A_27_47#_c_321_n 0.00154636f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_283 N_CLK_N_c_264_n N_A_27_47#_c_325_n 0.001616f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_284 N_CLK_N_c_270_n N_A_27_47#_c_325_n 0.00454961f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_285 CLK_N N_A_27_47#_c_325_n 0.0517716f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_286 N_CLK_N_c_266_n N_A_27_47#_c_325_n 9.99163e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_287 N_CLK_N_c_267_n N_A_27_47#_c_325_n 0.00207113f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_288 CLK_N N_A_27_47#_c_329_n 0.00162113f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_289 N_CLK_N_c_266_n N_A_27_47#_c_329_n 0.0169711f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_290 N_CLK_N_c_269_n N_VPWR_c_1755_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_291 N_CLK_N_c_269_n N_VPWR_c_1768_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_292 N_CLK_N_c_269_n N_VPWR_c_1754_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_293 N_CLK_N_c_263_n N_VGND_c_2075_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_294 N_CLK_N_c_263_n N_VGND_c_2092_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_295 N_CLK_N_c_264_n N_VGND_c_2092_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_296 N_CLK_N_c_263_n N_VGND_c_2102_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_320_n N_D_M1011_g 0.00365815f $X=2.84 $Y=0.85 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_310_n N_D_M1029_g 0.0317155f $X=2.38 $Y=1.32 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_310_n N_D_c_570_n 0.00467503f $X=2.38 $Y=1.32 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_320_n N_D_c_570_n 0.00114217f $X=2.84 $Y=0.85 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_310_n N_D_c_571_n 0.00326853f $X=2.38 $Y=1.32 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_320_n N_D_c_571_n 0.012399f $X=2.84 $Y=0.85 $X2=0 $Y2=0
cc_303 N_A_27_47#_M1006_g N_A_193_47#_c_610_n 0.013193f $X=2.845 $Y=0.415 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_327_n N_A_193_47#_c_610_n 5.17882e-19 $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1018_g N_A_193_47#_M1009_g 0.0190768f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_319_n N_A_193_47#_c_611_n 0.0110561f $X=6.652 $Y=1.305 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_337_n N_A_193_47#_c_611_n 0.00853911f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_338_n N_A_193_47#_c_611_n 0.0216716f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_328_n N_A_193_47#_c_611_n 3.23054e-19 $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_317_n N_A_193_47#_c_612_n 2.62384e-19 $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_318_n N_A_193_47#_c_612_n 0.0209335f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_319_n N_A_193_47#_c_612_n 0.00356667f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_328_n N_A_193_47#_c_612_n 9.01357e-19 $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_313_n N_A_193_47#_M1004_g 0.0129153f $X=6.21 $Y=0.705 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_317_n N_A_193_47#_M1004_g 0.00307377f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_318_n N_A_193_47#_M1004_g 0.021369f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_319_n N_A_193_47#_M1004_g 0.00622479f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_M1018_g N_A_193_47#_c_614_n 0.00534118f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_309_n N_A_193_47#_c_614_n 0.010154f $X=2.77 $Y=1.32 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_310_n N_A_193_47#_c_614_n 0.00204083f $X=2.38 $Y=1.32 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1006_g N_A_193_47#_c_614_n 4.48322e-19 $X=2.845 $Y=0.415
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_320_n N_A_193_47#_c_614_n 0.0173204f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_322_n N_A_193_47#_c_614_n 0.00927819f $X=3.032 $Y=1.12 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_326_n N_A_193_47#_c_614_n 4.97018e-19 $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_327_n N_A_193_47#_c_614_n 0.020859f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_330_n N_A_193_47#_c_614_n 0.00673428f $X=2.905 $Y=0.93 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_310_n N_A_193_47#_c_615_n 0.0232695f $X=2.38 $Y=1.32 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_M1006_g N_A_193_47#_c_615_n 0.0213778f $X=2.845 $Y=0.415 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_320_n N_A_193_47#_c_615_n 0.00539068f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_327_n N_A_193_47#_c_615_n 0.00153923f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_M1018_g N_A_193_47#_c_622_n 0.00700258f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_M1000_g N_A_193_47#_c_623_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_336_n N_A_193_47#_c_623_n 0.00560035f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_325_n N_A_193_47#_c_623_n 0.00113282f $X=0.695 $Y=0.85 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_309_n N_A_193_47#_c_624_n 3.83457e-19 $X=2.77 $Y=1.32 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_324_n N_A_193_47#_c_624_n 0.111194f $X=3.13 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_M1018_g N_A_193_47#_c_625_n 5.24592e-19 $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_M1019_g N_A_193_47#_c_626_n 0.00133927f $X=6.64 $Y=2.275 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_337_n N_A_193_47#_c_626_n 0.00483121f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_338_n N_A_193_47#_c_626_n 0.00219663f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_M1018_g N_A_193_47#_c_627_n 0.0174486f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_309_n N_A_193_47#_c_627_n 0.0212215f $X=2.77 $Y=1.32 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_327_n N_A_193_47#_c_627_n 3.19045e-19 $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_M1018_g N_A_193_47#_c_628_n 0.0103939f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_309_n N_A_193_47#_c_628_n 0.00655916f $X=2.77 $Y=1.32 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_327_n N_A_193_47#_c_628_n 0.00336529f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_M1019_g N_A_193_47#_c_629_n 0.0192968f $X=6.64 $Y=2.275 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_337_n N_A_193_47#_c_629_n 5.88448e-19 $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_338_n N_A_193_47#_c_629_n 0.0169266f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_323_n N_A_193_47#_c_629_n 2.37019e-19 $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_M1019_g N_A_193_47#_c_630_n 6.52047e-19 $X=6.64 $Y=2.275 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_319_n N_A_193_47#_c_630_n 0.00682571f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_337_n N_A_193_47#_c_630_n 0.0168759f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_338_n N_A_193_47#_c_630_n 0.00153059f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_328_n N_A_193_47#_c_630_n 0.00149027f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_337_n N_A_193_47#_c_631_n 0.00347329f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_M1025_g N_A_193_47#_c_616_n 0.0270874f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_315_n N_A_193_47#_c_616_n 0.0116735f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_336_n N_A_193_47#_c_616_n 0.00890309f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_320_n N_A_193_47#_c_616_n 0.0242694f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_321_n N_A_193_47#_c_616_n 0.0014643f $X=0.84 $Y=0.85 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_325_n N_A_193_47#_c_616_n 0.0705599f $X=0.695 $Y=0.85 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_M1006_g N_A_650_21#_M1012_g 0.0243315f $X=2.845 $Y=0.415 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_312_n N_A_650_21#_M1012_g 0.0102862f $X=2.845 $Y=1.245 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_327_n N_A_650_21#_M1012_g 0.0010488f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_330_n N_A_650_21#_M1012_g 0.021533f $X=2.905 $Y=0.93 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_313_n N_A_650_21#_c_813_n 0.0187265f $X=6.21 $Y=0.705 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_317_n N_A_650_21#_c_813_n 0.001702f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_323_n N_A_650_21#_c_822_n 0.00196084f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_323_n N_A_650_21#_c_834_n 0.00348372f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_323_n N_A_650_21#_c_814_n 0.00165548f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_323_n N_A_650_21#_c_815_n 0.016449f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_323_n N_A_650_21#_c_816_n 0.00907541f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_323_n N_A_650_21#_c_824_n 8.24776e-19 $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_323_n N_A_650_21#_c_839_n 6.83984e-19 $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_317_n N_A_650_21#_c_817_n 0.0111636f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_318_n N_A_650_21#_c_817_n 9.14426e-19 $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_319_n N_A_650_21#_c_817_n 0.00462764f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_323_n N_A_650_21#_c_817_n 0.0153364f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_328_n N_A_650_21#_c_817_n 0.00129536f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_317_n N_A_650_21#_c_818_n 5.13187e-19 $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_318_n N_A_650_21#_c_818_n 0.0187265f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_319_n N_A_650_21#_c_818_n 0.00174717f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_323_n N_A_650_21#_c_818_n 0.00365485f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_328_n N_A_650_21#_c_818_n 6.8647e-19 $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_323_n N_SET_B_c_957_n 0.00392015f $X=6.08 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_387 N_A_27_47#_c_323_n N_SET_B_M1041_g 0.0011704f $X=6.08 $Y=1.19 $X2=0 $Y2=0
cc_388 N_A_27_47#_c_323_n SET_B 0.00590244f $X=6.08 $Y=1.19 $X2=0 $Y2=0
cc_389 N_A_27_47#_c_317_n N_SET_B_c_963_n 0.0194369f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_318_n N_SET_B_c_963_n 0.0023282f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_319_n N_SET_B_c_963_n 0.0053562f $X=6.652 $Y=1.305 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_323_n N_SET_B_c_963_n 0.158115f $X=6.08 $Y=1.19 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_328_n N_SET_B_c_963_n 0.0254944f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_323_n N_SET_B_c_964_n 0.0265121f $X=6.08 $Y=1.19 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_323_n N_A_476_47#_M1035_g 0.00188875f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1018_g N_A_476_47#_c_1099_n 0.00281679f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_M1006_g N_A_476_47#_c_1100_n 0.00882839f $X=2.845 $Y=0.415
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_320_n N_A_476_47#_c_1100_n 0.00575474f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_326_n N_A_476_47#_c_1100_n 0.00258895f $X=2.985 $Y=0.85
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_327_n N_A_476_47#_c_1100_n 0.0182033f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_330_n N_A_476_47#_c_1100_n 5.24271e-19 $X=2.905 $Y=0.93
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_M1018_g N_A_476_47#_c_1094_n 8.73767e-19 $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_324_n N_A_476_47#_c_1094_n 3.06883e-19 $X=3.13 $Y=1.19 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_M1006_g N_A_476_47#_c_1089_n 2.58936e-19 $X=2.845 $Y=0.415
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_312_n N_A_476_47#_c_1089_n 0.00144384f $X=2.845 $Y=1.245
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_323_n N_A_476_47#_c_1089_n 0.0152458f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_326_n N_A_476_47#_c_1089_n 0.0143395f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_327_n N_A_476_47#_c_1089_n 0.0251282f $X=2.985 $Y=0.85 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_330_n N_A_476_47#_c_1089_n 0.00218717f $X=2.905 $Y=0.93
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_323_n N_A_476_47#_c_1090_n 0.0384689f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_312_n N_A_476_47#_c_1091_n 0.00268821f $X=2.845 $Y=1.245
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_323_n N_A_476_47#_c_1091_n 0.0110554f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_324_n N_A_476_47#_c_1091_n 0.0060147f $X=3.13 $Y=1.19 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_327_n N_A_476_47#_c_1091_n 0.00391072f $X=2.985 $Y=0.85
+ $X2=0 $Y2=0
cc_415 N_A_27_47#_c_330_n N_A_476_47#_c_1091_n 5.70501e-19 $X=2.905 $Y=0.93
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_323_n N_A_476_47#_c_1092_n 0.00386813f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_323_n N_A_944_21#_M1042_g 0.00150073f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_323_n N_A_944_21#_c_1198_n 0.0122826f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_323_n N_A_944_21#_c_1199_n 0.00611237f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_319_n N_A_944_21#_c_1208_n 0.00715591f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_337_n N_A_944_21#_c_1208_n 0.0157692f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_338_n N_A_944_21#_c_1208_n 0.00184742f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_323_n N_A_944_21#_c_1208_n 0.014133f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_328_n N_A_944_21#_c_1208_n 0.027417f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_323_n N_A_944_21#_c_1209_n 0.0276968f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_337_n N_A_944_21#_c_1210_n 0.00264766f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_323_n N_A_944_21#_c_1210_n 0.00618009f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_337_n N_A_1431_21#_M1024_g 3.51933e-19 $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_M1019_g N_A_1431_21#_c_1373_n 0.0162278f $X=6.64 $Y=2.275
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_338_n N_A_1431_21#_c_1373_n 0.00879184f $X=6.67 $Y=1.74
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_M1019_g N_A_1257_47#_c_1559_n 0.00935459f $X=6.64 $Y=2.275
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_337_n N_A_1257_47#_c_1559_n 0.00669245f $X=6.67 $Y=1.74
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_338_n N_A_1257_47#_c_1559_n 0.0028948f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_317_n N_A_1257_47#_c_1562_n 0.00390894f $X=6.335 $Y=0.87
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_318_n N_A_1257_47#_c_1562_n 0.00184507f $X=6.335 $Y=0.87
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_319_n N_A_1257_47#_c_1562_n 0.00315233f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_317_n N_A_1257_47#_c_1548_n 0.0117718f $X=6.335 $Y=0.87
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_319_n N_A_1257_47#_c_1548_n 0.00837612f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_328_n N_A_1257_47#_c_1548_n 6.65017e-19 $X=6.225 $Y=1.19
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_M1019_g N_A_1257_47#_c_1554_n 0.00655877f $X=6.64 $Y=2.275
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_337_n N_A_1257_47#_c_1554_n 0.0359925f $X=6.67 $Y=1.74 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_338_n N_A_1257_47#_c_1554_n 0.00212049f $X=6.67 $Y=1.74
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_319_n N_A_1257_47#_c_1550_n 0.00588724f $X=6.652 $Y=1.305
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_337_n N_A_1257_47#_c_1550_n 0.00820578f $X=6.67 $Y=1.74
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_328_n N_A_1257_47#_c_1550_n 2.68785e-19 $X=6.225 $Y=1.19
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_336_n N_VPWR_M1023_d 0.00167655f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_447 N_A_27_47#_M1000_g N_VPWR_c_1755_n 0.00827522f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_336_n N_VPWR_c_1755_n 0.0175536f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_339_n N_VPWR_c_1755_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_450 N_A_27_47#_M1000_g N_VPWR_c_1756_n 0.00191302f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_M1018_g N_VPWR_c_1756_n 0.00110623f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_336_n N_VPWR_c_1768_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_453 N_A_27_47#_c_339_n N_VPWR_c_1768_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_454 N_A_27_47#_M1000_g N_VPWR_c_1769_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_M1018_g N_VPWR_c_1770_n 0.00541732f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_M1019_g N_VPWR_c_1771_n 0.00367119f $X=6.64 $Y=2.275 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_M1000_g N_VPWR_c_1754_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_M1018_g N_VPWR_c_1754_n 0.00624914f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_M1019_g N_VPWR_c_1754_n 0.00567418f $X=6.64 $Y=2.275 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_336_n N_VPWR_c_1754_n 0.00507261f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_339_n N_VPWR_c_1754_n 0.00993215f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_320_n N_A_381_47#_c_1955_n 0.0149439f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_320_n N_A_381_47#_c_1956_n 0.0203199f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_327_n N_A_381_47#_c_1956_n 0.00212753f $X=2.985 $Y=0.85
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_c_320_n N_A_381_47#_c_1957_n 0.00433679f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_M1018_g N_A_381_47#_c_1959_n 0.00142476f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_M1018_g N_A_381_47#_c_1961_n 0.00730615f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_468 N_A_27_47#_c_315_n N_VGND_M1038_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_469 N_A_27_47#_M1025_g N_VGND_c_2075_n 0.00783511f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_315_n N_VGND_c_2075_n 0.0158742f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_471 N_A_27_47#_c_321_n N_VGND_c_2075_n 0.00116283f $X=0.84 $Y=0.85 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_329_n N_VGND_c_2075_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_M1025_g N_VGND_c_2076_n 0.00299798f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_320_n N_VGND_c_2076_n 0.00126774f $X=2.84 $Y=0.85 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_323_n N_VGND_c_2077_n 9.89759e-19 $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_313_n N_VGND_c_2078_n 0.00174046f $X=6.21 $Y=0.705 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_M1006_g N_VGND_c_2086_n 0.00359964f $X=2.845 $Y=0.415 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_313_n N_VGND_c_2090_n 0.00435972f $X=6.21 $Y=0.705 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_317_n N_VGND_c_2090_n 0.00288727f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_318_n N_VGND_c_2090_n 2.15978e-19 $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_314_n N_VGND_c_2092_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_482 N_A_27_47#_c_315_n N_VGND_c_2092_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_M1025_g N_VGND_c_2093_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_M1038_s N_VGND_c_2102_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_M1025_g N_VGND_c_2102_n 0.00581646f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_M1006_g N_VGND_c_2102_n 0.00561651f $X=2.845 $Y=0.415 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_313_n N_VGND_c_2102_n 0.00616197f $X=6.21 $Y=0.705 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_314_n N_VGND_c_2102_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_315_n N_VGND_c_2102_n 0.00526087f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_317_n N_VGND_c_2102_n 0.00224883f $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_c_320_n N_VGND_c_2102_n 0.0940283f $X=2.84 $Y=0.85 $X2=0 $Y2=0
cc_492 N_A_27_47#_c_321_n N_VGND_c_2102_n 0.0131302f $X=0.84 $Y=0.85 $X2=0 $Y2=0
cc_493 N_A_27_47#_c_326_n N_VGND_c_2102_n 0.015297f $X=2.985 $Y=0.85 $X2=0 $Y2=0
cc_494 N_A_27_47#_c_327_n A_584_47# 8.80342e-19 $X=2.985 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_495 N_D_M1011_g N_A_193_47#_c_610_n 0.0212588f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_496 N_D_M1011_g N_A_193_47#_c_614_n 0.0012229f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_497 N_D_c_570_n N_A_193_47#_c_614_n 0.0010617f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_498 N_D_c_571_n N_A_193_47#_c_614_n 0.0453933f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_499 N_D_c_570_n N_A_193_47#_c_615_n 0.0014765f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_500 N_D_c_571_n N_A_193_47#_c_615_n 2.3625e-19 $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_501 N_D_c_571_n N_A_193_47#_c_622_n 0.0053193f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_502 N_D_M1029_g N_A_193_47#_c_623_n 4.12204e-19 $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_503 N_D_M1029_g N_A_193_47#_c_628_n 0.00106128f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_504 N_D_c_571_n N_A_193_47#_c_628_n 0.00408526f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_505 N_D_M1011_g N_A_193_47#_c_616_n 0.00375157f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_506 N_D_M1029_g N_A_193_47#_c_616_n 0.00498234f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_507 N_D_M1029_g N_VPWR_c_1756_n 0.0117009f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_508 N_D_M1029_g N_VPWR_c_1770_n 0.0035268f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_509 N_D_M1029_g N_VPWR_c_1754_n 0.00400653f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_510 N_D_M1011_g N_A_381_47#_c_1955_n 0.00549247f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_511 N_D_M1029_g N_A_381_47#_c_1955_n 0.0113867f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_512 N_D_c_570_n N_A_381_47#_c_1955_n 0.00753248f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_513 N_D_c_571_n N_A_381_47#_c_1955_n 0.0473422f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_514 N_D_M1011_g N_A_381_47#_c_1956_n 0.0126207f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_515 N_D_c_570_n N_A_381_47#_c_1956_n 0.00200368f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_516 N_D_c_571_n N_A_381_47#_c_1956_n 0.023609f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_517 N_D_M1029_g N_A_381_47#_c_1959_n 0.0131516f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_518 N_D_c_570_n N_A_381_47#_c_1959_n 0.00153518f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_519 N_D_c_571_n N_A_381_47#_c_1959_n 0.0278526f $X=1.845 $Y=1.17 $X2=0 $Y2=0
cc_520 N_D_M1029_g N_A_381_47#_c_1961_n 0.00261491f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_521 N_D_M1011_g N_VGND_c_2076_n 0.00943841f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_522 N_D_M1011_g N_VGND_c_2086_n 0.00339367f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_523 N_D_M1011_g N_VGND_c_2102_n 0.00393034f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_524 N_A_193_47#_c_614_n N_A_650_21#_M1012_g 5.35023e-19 $X=2.425 $Y=0.87
+ $X2=0 $Y2=0
cc_525 N_A_193_47#_c_624_n N_A_650_21#_M1015_g 0.00197541f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_526 N_A_193_47#_M1031_g N_A_650_21#_M1028_g 0.0164618f $X=6.22 $Y=2.275 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_c_612_n N_A_650_21#_M1028_g 0.00557961f $X=6.295 $Y=1.32
+ $X2=0 $Y2=0
cc_528 N_A_193_47#_c_624_n N_A_650_21#_M1028_g 0.00753824f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_c_629_n N_A_650_21#_M1028_g 0.00910409f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_530 N_A_193_47#_c_630_n N_A_650_21#_M1028_g 0.00264318f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_531 N_A_193_47#_c_624_n N_A_650_21#_c_822_n 0.0240118f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_532 N_A_193_47#_c_624_n N_A_650_21#_c_834_n 0.0279846f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_533 N_A_193_47#_c_624_n N_A_650_21#_c_824_n 0.0141612f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_534 N_A_193_47#_M1009_g N_A_650_21#_c_825_n 0.0161827f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_535 N_A_193_47#_c_624_n N_A_650_21#_c_825_n 0.00193898f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_536 N_A_193_47#_c_627_n N_A_650_21#_c_825_n 0.00927772f $X=2.755 $Y=1.74
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_c_624_n N_A_650_21#_c_839_n 0.00959465f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_538 N_A_193_47#_c_612_n N_A_650_21#_c_818_n 0.00272432f $X=6.295 $Y=1.32
+ $X2=0 $Y2=0
cc_539 N_A_193_47#_M1004_g N_SET_B_c_963_n 0.00574501f $X=6.755 $Y=0.415 $X2=0
+ $Y2=0
cc_540 N_A_193_47#_M1009_g N_A_476_47#_c_1099_n 0.0091014f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_541 N_A_193_47#_c_622_n N_A_476_47#_c_1099_n 2.09728e-19 $X=2.4 $Y=1.87 $X2=0
+ $Y2=0
cc_542 N_A_193_47#_c_624_n N_A_476_47#_c_1099_n 0.00506942f $X=6.08 $Y=1.87
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_c_625_n N_A_476_47#_c_1099_n 0.00303545f $X=2.69 $Y=1.87
+ $X2=0 $Y2=0
cc_544 N_A_193_47#_c_627_n N_A_476_47#_c_1099_n 0.00186639f $X=2.755 $Y=1.74
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_628_n N_A_476_47#_c_1099_n 0.0152514f $X=2.755 $Y=1.74
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_614_n N_A_476_47#_c_1100_n 0.00653862f $X=2.425 $Y=0.87
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_c_615_n N_A_476_47#_c_1100_n 8.98642e-19 $X=2.425 $Y=0.87
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_M1009_g N_A_476_47#_c_1094_n 0.00650943f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_614_n N_A_476_47#_c_1094_n 0.00666284f $X=2.425 $Y=0.87
+ $X2=0 $Y2=0
cc_550 N_A_193_47#_c_624_n N_A_476_47#_c_1094_n 0.013911f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_551 N_A_193_47#_c_625_n N_A_476_47#_c_1094_n 0.00149623f $X=2.69 $Y=1.87
+ $X2=0 $Y2=0
cc_552 N_A_193_47#_c_627_n N_A_476_47#_c_1094_n 0.00203066f $X=2.755 $Y=1.74
+ $X2=0 $Y2=0
cc_553 N_A_193_47#_c_628_n N_A_476_47#_c_1094_n 0.0282877f $X=2.755 $Y=1.74
+ $X2=0 $Y2=0
cc_554 N_A_193_47#_c_624_n N_A_476_47#_c_1090_n 0.00350894f $X=6.08 $Y=1.87
+ $X2=0 $Y2=0
cc_555 N_A_193_47#_c_614_n N_A_476_47#_c_1091_n 0.00728836f $X=2.425 $Y=0.87
+ $X2=0 $Y2=0
cc_556 N_A_193_47#_c_624_n N_A_476_47#_c_1091_n 0.00456412f $X=6.08 $Y=1.87
+ $X2=0 $Y2=0
cc_557 N_A_193_47#_c_624_n N_A_944_21#_M1032_g 0.00583916f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_558 N_A_193_47#_c_624_n N_A_944_21#_c_1198_n 0.00487283f $X=6.08 $Y=1.87
+ $X2=0 $Y2=0
cc_559 N_A_193_47#_c_611_n N_A_944_21#_c_1208_n 0.00389341f $X=6.68 $Y=1.32
+ $X2=0 $Y2=0
cc_560 N_A_193_47#_c_624_n N_A_944_21#_c_1208_n 0.0139809f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_561 N_A_193_47#_c_626_n N_A_944_21#_c_1208_n 0.0255925f $X=6.225 $Y=1.87
+ $X2=0 $Y2=0
cc_562 N_A_193_47#_c_629_n N_A_944_21#_c_1208_n 0.00176885f $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_563 N_A_193_47#_c_630_n N_A_944_21#_c_1208_n 0.00661378f $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_564 N_A_193_47#_c_631_n N_A_944_21#_c_1208_n 0.00371524f $X=6.16 $Y=1.575
+ $X2=0 $Y2=0
cc_565 N_A_193_47#_c_624_n N_A_944_21#_c_1209_n 0.0264578f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_566 N_A_193_47#_c_629_n N_A_944_21#_c_1209_n 7.96394e-19 $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_567 N_A_193_47#_c_630_n N_A_944_21#_c_1209_n 0.00130051f $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_568 N_A_193_47#_c_631_n N_A_944_21#_c_1209_n 7.27878e-19 $X=6.16 $Y=1.575
+ $X2=0 $Y2=0
cc_569 N_A_193_47#_c_624_n N_A_944_21#_c_1210_n 0.020032f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_570 N_A_193_47#_c_629_n N_A_944_21#_c_1210_n 6.45403e-19 $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_571 N_A_193_47#_c_630_n N_A_944_21#_c_1210_n 0.00461622f $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_572 N_A_193_47#_c_631_n N_A_944_21#_c_1210_n 0.00148716f $X=6.16 $Y=1.575
+ $X2=0 $Y2=0
cc_573 N_A_193_47#_M1004_g N_A_1431_21#_M1024_g 0.0428045f $X=6.755 $Y=0.415
+ $X2=0 $Y2=0
cc_574 N_A_193_47#_M1031_g N_A_1257_47#_c_1559_n 0.00496872f $X=6.22 $Y=2.275
+ $X2=0 $Y2=0
cc_575 N_A_193_47#_c_626_n N_A_1257_47#_c_1559_n 0.00187313f $X=6.225 $Y=1.87
+ $X2=0 $Y2=0
cc_576 N_A_193_47#_c_630_n N_A_1257_47#_c_1559_n 0.00141396f $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_577 N_A_193_47#_M1004_g N_A_1257_47#_c_1562_n 0.0096406f $X=6.755 $Y=0.415
+ $X2=0 $Y2=0
cc_578 N_A_193_47#_M1004_g N_A_1257_47#_c_1548_n 0.010696f $X=6.755 $Y=0.415
+ $X2=0 $Y2=0
cc_579 N_A_193_47#_c_626_n N_A_1257_47#_c_1554_n 0.00214622f $X=6.225 $Y=1.87
+ $X2=0 $Y2=0
cc_580 N_A_193_47#_c_630_n N_A_1257_47#_c_1554_n 0.0013353f $X=6.16 $Y=1.74
+ $X2=0 $Y2=0
cc_581 N_A_193_47#_M1004_g N_A_1257_47#_c_1550_n 0.00156831f $X=6.755 $Y=0.415
+ $X2=0 $Y2=0
cc_582 N_A_193_47#_c_624_n N_VPWR_M1032_d 0.00710211f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_583 N_A_193_47#_c_616_n N_VPWR_c_1755_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_584 N_A_193_47#_c_622_n N_VPWR_c_1756_n 0.00172075f $X=2.4 $Y=1.87 $X2=0
+ $Y2=0
cc_585 N_A_193_47#_c_616_n N_VPWR_c_1756_n 0.0234727f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_586 N_A_193_47#_c_624_n N_VPWR_c_1757_n 0.00160449f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_587 N_A_193_47#_c_624_n N_VPWR_c_1758_n 0.0137334f $X=6.08 $Y=1.87 $X2=0
+ $Y2=0
cc_588 N_A_193_47#_c_616_n N_VPWR_c_1769_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_589 N_A_193_47#_M1009_g N_VPWR_c_1770_n 0.00367119f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_590 N_A_193_47#_M1031_g N_VPWR_c_1771_n 0.00424681f $X=6.22 $Y=2.275 $X2=0
+ $Y2=0
cc_591 N_A_193_47#_c_630_n N_VPWR_c_1771_n 0.00254851f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_592 N_A_193_47#_M1009_g N_VPWR_c_1754_n 0.00562272f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_593 N_A_193_47#_M1031_g N_VPWR_c_1754_n 0.0061745f $X=6.22 $Y=2.275 $X2=0
+ $Y2=0
cc_594 N_A_193_47#_c_622_n N_VPWR_c_1754_n 0.0505224f $X=2.4 $Y=1.87 $X2=0 $Y2=0
cc_595 N_A_193_47#_c_623_n N_VPWR_c_1754_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_596 N_A_193_47#_c_624_n N_VPWR_c_1754_n 0.159053f $X=6.08 $Y=1.87 $X2=0 $Y2=0
cc_597 N_A_193_47#_c_625_n N_VPWR_c_1754_n 0.0160117f $X=2.69 $Y=1.87 $X2=0
+ $Y2=0
cc_598 N_A_193_47#_c_626_n N_VPWR_c_1754_n 0.0148451f $X=6.225 $Y=1.87 $X2=0
+ $Y2=0
cc_599 N_A_193_47#_c_628_n N_VPWR_c_1754_n 3.19863e-19 $X=2.755 $Y=1.74 $X2=0
+ $Y2=0
cc_600 N_A_193_47#_c_629_n N_VPWR_c_1754_n 3.05853e-19 $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_601 N_A_193_47#_c_630_n N_VPWR_c_1754_n 0.00131252f $X=6.16 $Y=1.74 $X2=0
+ $Y2=0
cc_602 N_A_193_47#_c_616_n N_VPWR_c_1754_n 0.00389918f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_603 N_A_193_47#_c_623_n N_A_381_47#_c_1955_n 0.00121388f $X=1.3 $Y=1.87 $X2=0
+ $Y2=0
cc_604 N_A_193_47#_c_616_n N_A_381_47#_c_1955_n 0.0703675f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_605 N_A_193_47#_c_610_n N_A_381_47#_c_1956_n 0.00221174f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_606 N_A_193_47#_c_614_n N_A_381_47#_c_1956_n 0.0076355f $X=2.425 $Y=0.87
+ $X2=0 $Y2=0
cc_607 N_A_193_47#_c_616_n N_A_381_47#_c_1957_n 0.0149979f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_608 N_A_193_47#_c_622_n N_A_381_47#_c_1959_n 0.030474f $X=2.4 $Y=1.87 $X2=0
+ $Y2=0
cc_609 N_A_193_47#_c_625_n N_A_381_47#_c_1959_n 6.96814e-19 $X=2.69 $Y=1.87
+ $X2=0 $Y2=0
cc_610 N_A_193_47#_c_628_n N_A_381_47#_c_1959_n 0.00893286f $X=2.755 $Y=1.74
+ $X2=0 $Y2=0
cc_611 N_A_193_47#_c_622_n N_A_381_47#_c_1960_n 0.0156655f $X=2.4 $Y=1.87 $X2=0
+ $Y2=0
cc_612 N_A_193_47#_c_623_n N_A_381_47#_c_1960_n 9.4615e-19 $X=1.3 $Y=1.87 $X2=0
+ $Y2=0
cc_613 N_A_193_47#_c_616_n N_A_381_47#_c_1960_n 0.0117002f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_614 N_A_193_47#_c_610_n N_A_381_47#_c_1990_n 0.00397815f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_615 N_A_193_47#_c_625_n N_A_381_47#_c_1961_n 8.58786e-19 $X=2.69 $Y=1.87
+ $X2=0 $Y2=0
cc_616 N_A_193_47#_c_624_n A_894_329# 5.39371e-19 $X=6.08 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_617 N_A_193_47#_c_624_n A_1115_329# 0.00532504f $X=6.08 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_618 N_A_193_47#_c_610_n N_VGND_c_2076_n 0.00121072f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_619 N_A_193_47#_c_616_n N_VGND_c_2076_n 0.00853554f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_620 N_A_193_47#_M1004_g N_VGND_c_2079_n 0.00126137f $X=6.755 $Y=0.415 $X2=0
+ $Y2=0
cc_621 N_A_193_47#_c_610_n N_VGND_c_2086_n 0.00546277f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_622 N_A_193_47#_c_614_n N_VGND_c_2086_n 0.00113905f $X=2.425 $Y=0.87 $X2=0
+ $Y2=0
cc_623 N_A_193_47#_c_615_n N_VGND_c_2086_n 2.1168e-19 $X=2.425 $Y=0.87 $X2=0
+ $Y2=0
cc_624 N_A_193_47#_M1004_g N_VGND_c_2090_n 0.00359964f $X=6.755 $Y=0.415 $X2=0
+ $Y2=0
cc_625 N_A_193_47#_c_616_n N_VGND_c_2093_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_626 N_A_193_47#_M1025_d N_VGND_c_2102_n 0.00217251f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_627 N_A_193_47#_c_610_n N_VGND_c_2102_n 0.00671269f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_628 N_A_193_47#_M1004_g N_VGND_c_2102_n 0.00564067f $X=6.755 $Y=0.415 $X2=0
+ $Y2=0
cc_629 N_A_193_47#_c_614_n N_VGND_c_2102_n 0.00121387f $X=2.425 $Y=0.87 $X2=0
+ $Y2=0
cc_630 N_A_193_47#_c_616_n N_VGND_c_2102_n 0.00389166f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_631 N_A_650_21#_M1012_g N_SET_B_c_957_n 0.0190011f $X=3.325 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_632 N_A_650_21#_M1012_g N_SET_B_M1041_g 0.0137896f $X=3.325 $Y=0.445 $X2=0
+ $Y2=0
cc_633 N_A_650_21#_M1015_g N_SET_B_M1041_g 0.0101628f $X=3.325 $Y=2.275 $X2=0
+ $Y2=0
cc_634 N_A_650_21#_c_822_n N_SET_B_M1041_g 0.0159332f $X=4.1 $Y=1.91 $X2=0 $Y2=0
cc_635 N_A_650_21#_c_869_p N_SET_B_M1041_g 0.00507112f $X=4.185 $Y=2.21 $X2=0
+ $Y2=0
cc_636 N_A_650_21#_c_824_n N_SET_B_M1041_g 0.00473578f $X=3.435 $Y=1.74 $X2=0
+ $Y2=0
cc_637 N_A_650_21#_c_825_n N_SET_B_M1041_g 0.020182f $X=3.435 $Y=1.74 $X2=0
+ $Y2=0
cc_638 N_A_650_21#_M1012_g N_SET_B_M1037_g 0.0156014f $X=3.325 $Y=0.445 $X2=0
+ $Y2=0
cc_639 N_A_650_21#_c_814_n N_SET_B_M1037_g 5.56585e-19 $X=4.615 $Y=1.065 $X2=0
+ $Y2=0
cc_640 N_A_650_21#_M1012_g SET_B 0.00118793f $X=3.325 $Y=0.445 $X2=0 $Y2=0
cc_641 N_A_650_21#_c_814_n SET_B 0.00825406f $X=4.615 $Y=1.065 $X2=0 $Y2=0
cc_642 N_A_650_21#_M1035_d N_SET_B_c_963_n 5.1491e-19 $X=4.45 $Y=0.235 $X2=0
+ $Y2=0
cc_643 N_A_650_21#_c_813_n N_SET_B_c_963_n 0.00507207f $X=5.735 $Y=0.985 $X2=0
+ $Y2=0
cc_644 N_A_650_21#_c_814_n N_SET_B_c_963_n 0.0208059f $X=4.615 $Y=1.065 $X2=0
+ $Y2=0
cc_645 N_A_650_21#_c_816_n N_SET_B_c_963_n 0.0198998f $X=5.51 $Y=0.98 $X2=0
+ $Y2=0
cc_646 N_A_650_21#_c_817_n N_SET_B_c_963_n 0.0108883f $X=5.675 $Y=0.98 $X2=0
+ $Y2=0
cc_647 N_A_650_21#_c_814_n N_SET_B_c_964_n 0.00230334f $X=4.615 $Y=1.065 $X2=0
+ $Y2=0
cc_648 N_A_650_21#_c_814_n N_A_476_47#_M1035_g 0.00722888f $X=4.615 $Y=1.065
+ $X2=0 $Y2=0
cc_649 N_A_650_21#_c_815_n N_A_476_47#_M1035_g 0.00191659f $X=4.615 $Y=1.785
+ $X2=0 $Y2=0
cc_650 N_A_650_21#_c_834_n N_A_476_47#_M1020_g 0.012508f $X=4.53 $Y=1.91 $X2=0
+ $Y2=0
cc_651 N_A_650_21#_M1015_g N_A_476_47#_c_1099_n 0.00191115f $X=3.325 $Y=2.275
+ $X2=0 $Y2=0
cc_652 N_A_650_21#_M1012_g N_A_476_47#_c_1100_n 0.00797698f $X=3.325 $Y=0.445
+ $X2=0 $Y2=0
cc_653 N_A_650_21#_M1012_g N_A_476_47#_c_1094_n 0.0154362f $X=3.325 $Y=0.445
+ $X2=0 $Y2=0
cc_654 N_A_650_21#_c_824_n N_A_476_47#_c_1094_n 0.0330453f $X=3.435 $Y=1.74
+ $X2=0 $Y2=0
cc_655 N_A_650_21#_M1012_g N_A_476_47#_c_1089_n 0.0153158f $X=3.325 $Y=0.445
+ $X2=0 $Y2=0
cc_656 N_A_650_21#_c_822_n N_A_476_47#_c_1090_n 0.0141289f $X=4.1 $Y=1.91 $X2=0
+ $Y2=0
cc_657 N_A_650_21#_c_834_n N_A_476_47#_c_1090_n 0.00218253f $X=4.53 $Y=1.91
+ $X2=0 $Y2=0
cc_658 N_A_650_21#_c_815_n N_A_476_47#_c_1090_n 0.0246731f $X=4.615 $Y=1.785
+ $X2=0 $Y2=0
cc_659 N_A_650_21#_c_839_n N_A_476_47#_c_1090_n 0.00650509f $X=4.185 $Y=1.87
+ $X2=0 $Y2=0
cc_660 N_A_650_21#_M1012_g N_A_476_47#_c_1091_n 0.0106244f $X=3.325 $Y=0.445
+ $X2=0 $Y2=0
cc_661 N_A_650_21#_c_824_n N_A_476_47#_c_1091_n 0.0169621f $X=3.435 $Y=1.74
+ $X2=0 $Y2=0
cc_662 N_A_650_21#_c_825_n N_A_476_47#_c_1091_n 0.00119732f $X=3.435 $Y=1.74
+ $X2=0 $Y2=0
cc_663 N_A_650_21#_c_815_n N_A_476_47#_c_1092_n 0.00921796f $X=4.615 $Y=1.785
+ $X2=0 $Y2=0
cc_664 N_A_650_21#_c_839_n N_A_476_47#_c_1092_n 9.09922e-19 $X=4.185 $Y=1.87
+ $X2=0 $Y2=0
cc_665 N_A_650_21#_c_814_n N_A_944_21#_M1042_g 0.00957438f $X=4.615 $Y=1.065
+ $X2=0 $Y2=0
cc_666 N_A_650_21#_c_815_n N_A_944_21#_M1042_g 0.00757744f $X=4.615 $Y=1.785
+ $X2=0 $Y2=0
cc_667 N_A_650_21#_c_816_n N_A_944_21#_M1042_g 0.00930678f $X=5.51 $Y=0.98 $X2=0
+ $Y2=0
cc_668 N_A_650_21#_c_817_n N_A_944_21#_M1042_g 0.00136887f $X=5.675 $Y=0.98
+ $X2=0 $Y2=0
cc_669 N_A_650_21#_c_818_n N_A_944_21#_M1042_g 0.00197459f $X=5.675 $Y=1.15
+ $X2=0 $Y2=0
cc_670 N_A_650_21#_M1028_g N_A_944_21#_M1032_g 0.0142344f $X=5.5 $Y=2.065 $X2=0
+ $Y2=0
cc_671 N_A_650_21#_c_834_n N_A_944_21#_M1032_g 0.00222516f $X=4.53 $Y=1.91 $X2=0
+ $Y2=0
cc_672 N_A_650_21#_M1028_g N_A_944_21#_c_1198_n 2.9354e-19 $X=5.5 $Y=2.065 $X2=0
+ $Y2=0
cc_673 N_A_650_21#_c_815_n N_A_944_21#_c_1198_n 0.0312021f $X=4.615 $Y=1.785
+ $X2=0 $Y2=0
cc_674 N_A_650_21#_c_816_n N_A_944_21#_c_1198_n 0.0205705f $X=5.51 $Y=0.98 $X2=0
+ $Y2=0
cc_675 N_A_650_21#_c_818_n N_A_944_21#_c_1198_n 0.00382982f $X=5.675 $Y=1.15
+ $X2=0 $Y2=0
cc_676 N_A_650_21#_c_816_n N_A_944_21#_c_1199_n 0.00590751f $X=5.51 $Y=0.98
+ $X2=0 $Y2=0
cc_677 N_A_650_21#_c_817_n N_A_944_21#_c_1199_n 7.54142e-19 $X=5.675 $Y=0.98
+ $X2=0 $Y2=0
cc_678 N_A_650_21#_c_818_n N_A_944_21#_c_1199_n 0.0166765f $X=5.675 $Y=1.15
+ $X2=0 $Y2=0
cc_679 N_A_650_21#_c_817_n N_A_944_21#_c_1209_n 9.59092e-19 $X=5.675 $Y=0.98
+ $X2=0 $Y2=0
cc_680 N_A_650_21#_c_818_n N_A_944_21#_c_1209_n 0.00358318f $X=5.675 $Y=1.15
+ $X2=0 $Y2=0
cc_681 N_A_650_21#_M1028_g N_A_944_21#_c_1210_n 0.0143513f $X=5.5 $Y=2.065 $X2=0
+ $Y2=0
cc_682 N_A_650_21#_c_816_n N_A_944_21#_c_1210_n 0.00760725f $X=5.51 $Y=0.98
+ $X2=0 $Y2=0
cc_683 N_A_650_21#_c_817_n N_A_944_21#_c_1210_n 0.0207118f $X=5.675 $Y=0.98
+ $X2=0 $Y2=0
cc_684 N_A_650_21#_c_818_n N_A_944_21#_c_1210_n 0.00632961f $X=5.675 $Y=1.15
+ $X2=0 $Y2=0
cc_685 N_A_650_21#_M1028_g N_A_1257_47#_c_1559_n 7.04843e-19 $X=5.5 $Y=2.065
+ $X2=0 $Y2=0
cc_686 N_A_650_21#_M1015_g N_VPWR_c_1757_n 0.00326498f $X=3.325 $Y=2.275 $X2=0
+ $Y2=0
cc_687 N_A_650_21#_c_822_n N_VPWR_c_1757_n 0.0124698f $X=4.1 $Y=1.91 $X2=0 $Y2=0
cc_688 N_A_650_21#_c_869_p N_VPWR_c_1757_n 0.00820313f $X=4.185 $Y=2.21 $X2=0
+ $Y2=0
cc_689 N_A_650_21#_c_824_n N_VPWR_c_1757_n 0.0125544f $X=3.435 $Y=1.74 $X2=0
+ $Y2=0
cc_690 N_A_650_21#_c_825_n N_VPWR_c_1757_n 7.62241e-19 $X=3.435 $Y=1.74 $X2=0
+ $Y2=0
cc_691 N_A_650_21#_M1028_g N_VPWR_c_1758_n 0.0164544f $X=5.5 $Y=2.065 $X2=0
+ $Y2=0
cc_692 N_A_650_21#_c_834_n N_VPWR_c_1758_n 8.19852e-19 $X=4.53 $Y=1.91 $X2=0
+ $Y2=0
cc_693 N_A_650_21#_c_822_n N_VPWR_c_1764_n 0.00474052f $X=4.1 $Y=1.91 $X2=0
+ $Y2=0
cc_694 N_A_650_21#_c_869_p N_VPWR_c_1764_n 0.00725778f $X=4.185 $Y=2.21 $X2=0
+ $Y2=0
cc_695 N_A_650_21#_c_834_n N_VPWR_c_1764_n 0.00580887f $X=4.53 $Y=1.91 $X2=0
+ $Y2=0
cc_696 N_A_650_21#_M1015_g N_VPWR_c_1770_n 0.00535335f $X=3.325 $Y=2.275 $X2=0
+ $Y2=0
cc_697 N_A_650_21#_c_824_n N_VPWR_c_1770_n 0.00111392f $X=3.435 $Y=1.74 $X2=0
+ $Y2=0
cc_698 N_A_650_21#_M1028_g N_VPWR_c_1771_n 0.00585385f $X=5.5 $Y=2.065 $X2=0
+ $Y2=0
cc_699 N_A_650_21#_M1041_d N_VPWR_c_1754_n 0.0031612f $X=3.93 $Y=2.065 $X2=0
+ $Y2=0
cc_700 N_A_650_21#_M1015_g N_VPWR_c_1754_n 0.00664368f $X=3.325 $Y=2.275 $X2=0
+ $Y2=0
cc_701 N_A_650_21#_M1028_g N_VPWR_c_1754_n 0.00765939f $X=5.5 $Y=2.065 $X2=0
+ $Y2=0
cc_702 N_A_650_21#_c_822_n N_VPWR_c_1754_n 0.00386836f $X=4.1 $Y=1.91 $X2=0
+ $Y2=0
cc_703 N_A_650_21#_c_869_p N_VPWR_c_1754_n 0.0029026f $X=4.185 $Y=2.21 $X2=0
+ $Y2=0
cc_704 N_A_650_21#_c_834_n N_VPWR_c_1754_n 0.00505387f $X=4.53 $Y=1.91 $X2=0
+ $Y2=0
cc_705 N_A_650_21#_c_824_n N_VPWR_c_1754_n 0.00128163f $X=3.435 $Y=1.74 $X2=0
+ $Y2=0
cc_706 N_A_650_21#_c_834_n A_894_329# 0.00273228f $X=4.53 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_707 N_A_650_21#_c_815_n A_894_329# 0.00162899f $X=4.615 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_708 N_A_650_21#_M1012_g N_VGND_c_2077_n 0.00372247f $X=3.325 $Y=0.445 $X2=0
+ $Y2=0
cc_709 N_A_650_21#_c_813_n N_VGND_c_2078_n 0.0111314f $X=5.735 $Y=0.985 $X2=0
+ $Y2=0
cc_710 N_A_650_21#_c_816_n N_VGND_c_2078_n 0.00387395f $X=5.51 $Y=0.98 $X2=0
+ $Y2=0
cc_711 N_A_650_21#_c_817_n N_VGND_c_2078_n 0.00379129f $X=5.675 $Y=0.98 $X2=0
+ $Y2=0
cc_712 N_A_650_21#_c_818_n N_VGND_c_2078_n 8.52393e-19 $X=5.675 $Y=1.15 $X2=0
+ $Y2=0
cc_713 N_A_650_21#_M1012_g N_VGND_c_2086_n 0.00359757f $X=3.325 $Y=0.445 $X2=0
+ $Y2=0
cc_714 N_A_650_21#_c_813_n N_VGND_c_2090_n 0.0046653f $X=5.735 $Y=0.985 $X2=0
+ $Y2=0
cc_715 N_A_650_21#_M1035_d N_VGND_c_2102_n 0.00178362f $X=4.45 $Y=0.235 $X2=0
+ $Y2=0
cc_716 N_A_650_21#_M1012_g N_VGND_c_2102_n 0.00576589f $X=3.325 $Y=0.445 $X2=0
+ $Y2=0
cc_717 N_A_650_21#_c_813_n N_VGND_c_2102_n 0.00460207f $X=5.735 $Y=0.985 $X2=0
+ $Y2=0
cc_718 N_A_650_21#_M1035_d N_A_790_47#_c_2285_n 0.0030477f $X=4.45 $Y=0.235
+ $X2=0 $Y2=0
cc_719 N_A_650_21#_c_814_n N_A_790_47#_c_2285_n 0.0147704f $X=4.615 $Y=1.065
+ $X2=0 $Y2=0
cc_720 N_A_650_21#_c_816_n N_A_790_47#_c_2285_n 0.00259503f $X=5.51 $Y=0.98
+ $X2=0 $Y2=0
cc_721 N_A_650_21#_c_813_n N_A_790_47#_c_2286_n 0.00507683f $X=5.735 $Y=0.985
+ $X2=0 $Y2=0
cc_722 N_A_650_21#_c_816_n N_A_790_47#_c_2286_n 0.0158487f $X=5.51 $Y=0.98 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_957_n N_A_476_47#_M1035_g 0.00619508f $X=3.855 $Y=1.145 $X2=0
+ $Y2=0
cc_724 N_SET_B_M1037_g N_A_476_47#_M1035_g 0.0234092f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_725 SET_B N_A_476_47#_M1035_g 0.0018678f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_726 N_SET_B_c_963_n N_A_476_47#_M1035_g 0.00496613f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_727 N_SET_B_c_964_n N_A_476_47#_M1035_g 0.00135305f $X=4.07 $Y=0.85 $X2=0
+ $Y2=0
cc_728 N_SET_B_M1041_g N_A_476_47#_M1020_g 0.0228864f $X=3.855 $Y=2.275 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_957_n N_A_476_47#_c_1089_n 0.00214594f $X=3.855 $Y=1.145 $X2=0
+ $Y2=0
cc_730 N_SET_B_M1041_g N_A_476_47#_c_1089_n 5.82142e-19 $X=3.855 $Y=2.275 $X2=0
+ $Y2=0
cc_731 N_SET_B_M1037_g N_A_476_47#_c_1089_n 0.0018137f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_732 SET_B N_A_476_47#_c_1089_n 0.0221461f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_733 N_SET_B_c_964_n N_A_476_47#_c_1089_n 0.00112047f $X=4.07 $Y=0.85 $X2=0
+ $Y2=0
cc_734 N_SET_B_c_957_n N_A_476_47#_c_1090_n 0.00299221f $X=3.855 $Y=1.145 $X2=0
+ $Y2=0
cc_735 N_SET_B_M1041_g N_A_476_47#_c_1090_n 0.0131452f $X=3.855 $Y=2.275 $X2=0
+ $Y2=0
cc_736 SET_B N_A_476_47#_c_1090_n 0.024648f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_737 N_SET_B_c_963_n N_A_476_47#_c_1090_n 0.00284271f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_738 N_SET_B_c_964_n N_A_476_47#_c_1090_n 6.67689e-19 $X=4.07 $Y=0.85 $X2=0
+ $Y2=0
cc_739 N_SET_B_M1041_g N_A_476_47#_c_1091_n 4.98733e-19 $X=3.855 $Y=2.275 $X2=0
+ $Y2=0
cc_740 N_SET_B_M1041_g N_A_476_47#_c_1092_n 0.021088f $X=3.855 $Y=2.275 $X2=0
+ $Y2=0
cc_741 N_SET_B_c_963_n N_A_944_21#_M1042_g 0.00317213f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_742 N_SET_B_c_963_n N_A_944_21#_c_1198_n 5.29205e-19 $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_743 N_SET_B_M1013_g N_A_944_21#_c_1208_n 0.00583258f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_744 N_SET_B_c_963_n N_A_944_21#_c_1208_n 0.0486538f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_745 N_SET_B_c_965_n N_A_944_21#_c_1208_n 0.0135087f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_746 N_SET_B_M1005_g N_A_1431_21#_M1024_g 0.0180201f $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_747 N_SET_B_M1013_g N_A_1431_21#_M1024_g 0.0136409f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_748 N_SET_B_c_963_n N_A_1431_21#_M1024_g 0.00627116f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_749 N_SET_B_c_965_n N_A_1431_21#_M1024_g 0.00136404f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_750 N_SET_B_c_966_n N_A_1431_21#_M1024_g 0.00227945f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_751 N_SET_B_c_967_n N_A_1431_21#_M1024_g 0.020875f $X=7.65 $Y=0.98 $X2=0
+ $Y2=0
cc_752 N_SET_B_M1013_g N_A_1431_21#_M1034_g 0.0109753f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_753 N_SET_B_M1013_g N_A_1431_21#_c_1372_n 0.00710111f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_754 N_SET_B_M1013_g N_A_1431_21#_c_1373_n 0.019738f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_755 N_SET_B_M1013_g N_A_1431_21#_c_1374_n 0.0136222f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_756 N_SET_B_c_966_n N_A_1431_21#_c_1362_n 0.00828511f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_757 N_SET_B_M1005_g N_A_1431_21#_c_1393_n 6.74813e-19 $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_758 N_SET_B_c_965_n N_A_1431_21#_c_1393_n 2.37563e-19 $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_759 N_SET_B_c_966_n N_A_1431_21#_c_1393_n 0.00144717f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_760 N_SET_B_M1005_g N_A_1257_47#_M1008_g 0.0175593f $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_761 N_SET_B_c_966_n N_A_1257_47#_M1008_g 0.00170408f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_762 N_SET_B_c_967_n N_A_1257_47#_M1008_g 0.009306f $X=7.65 $Y=0.98 $X2=0
+ $Y2=0
cc_763 N_SET_B_M1013_g N_A_1257_47#_M1039_g 0.0325064f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_764 N_SET_B_c_963_n N_A_1257_47#_c_1562_n 0.00883541f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_765 N_SET_B_c_963_n N_A_1257_47#_c_1548_n 0.017797f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_766 N_SET_B_c_965_n N_A_1257_47#_c_1548_n 0.0022902f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_767 N_SET_B_c_966_n N_A_1257_47#_c_1548_n 0.0118231f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_768 N_SET_B_M1013_g N_A_1257_47#_c_1549_n 0.0117331f $X=7.77 $Y=2.275 $X2=0
+ $Y2=0
cc_769 N_SET_B_c_963_n N_A_1257_47#_c_1549_n 0.00876649f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_770 N_SET_B_c_965_n N_A_1257_47#_c_1549_n 0.00124273f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_771 N_SET_B_c_966_n N_A_1257_47#_c_1549_n 0.0248283f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_772 N_SET_B_c_967_n N_A_1257_47#_c_1549_n 0.00490678f $X=7.65 $Y=0.98 $X2=0
+ $Y2=0
cc_773 N_SET_B_c_967_n N_A_1257_47#_c_1551_n 0.00111089f $X=7.65 $Y=0.98 $X2=0
+ $Y2=0
cc_774 N_SET_B_c_967_n N_A_1257_47#_c_1552_n 0.0212822f $X=7.65 $Y=0.98 $X2=0
+ $Y2=0
cc_775 N_SET_B_M1041_g N_VPWR_c_1757_n 0.0094739f $X=3.855 $Y=2.275 $X2=0 $Y2=0
cc_776 N_SET_B_M1041_g N_VPWR_c_1764_n 0.00373914f $X=3.855 $Y=2.275 $X2=0 $Y2=0
cc_777 N_SET_B_M1013_g N_VPWR_c_1767_n 0.00368415f $X=7.77 $Y=2.275 $X2=0 $Y2=0
cc_778 N_SET_B_M1013_g N_VPWR_c_1778_n 0.00857728f $X=7.77 $Y=2.275 $X2=0 $Y2=0
cc_779 N_SET_B_M1041_g N_VPWR_c_1754_n 0.00439789f $X=3.855 $Y=2.275 $X2=0 $Y2=0
cc_780 N_SET_B_M1013_g N_VPWR_c_1754_n 0.00444663f $X=7.77 $Y=2.275 $X2=0 $Y2=0
cc_781 N_SET_B_c_963_n N_VGND_M1021_s 0.00213341f $X=7.46 $Y=0.85 $X2=0 $Y2=0
cc_782 N_SET_B_c_957_n N_VGND_c_2077_n 7.32772e-19 $X=3.855 $Y=1.145 $X2=0 $Y2=0
cc_783 N_SET_B_M1037_g N_VGND_c_2077_n 0.00287306f $X=3.875 $Y=0.445 $X2=0 $Y2=0
cc_784 SET_B N_VGND_c_2077_n 0.00971383f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_785 N_SET_B_c_963_n N_VGND_c_2078_n 0.00404506f $X=7.46 $Y=0.85 $X2=0 $Y2=0
cc_786 N_SET_B_M1005_g N_VGND_c_2079_n 0.00282278f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_787 N_SET_B_c_963_n N_VGND_c_2079_n 0.00604269f $X=7.46 $Y=0.85 $X2=0 $Y2=0
cc_788 N_SET_B_c_965_n N_VGND_c_2079_n 7.41662e-19 $X=7.605 $Y=0.85 $X2=0 $Y2=0
cc_789 N_SET_B_c_966_n N_VGND_c_2079_n 0.00350326f $X=7.605 $Y=0.85 $X2=0 $Y2=0
cc_790 N_SET_B_M1037_g N_VGND_c_2088_n 0.00423333f $X=3.875 $Y=0.445 $X2=0 $Y2=0
cc_791 SET_B N_VGND_c_2088_n 0.00223437f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_792 N_SET_B_M1005_g N_VGND_c_2094_n 0.00439071f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_793 N_SET_B_c_966_n N_VGND_c_2094_n 0.00352663f $X=7.605 $Y=0.85 $X2=0 $Y2=0
cc_794 N_SET_B_M1037_g N_VGND_c_2102_n 0.00593301f $X=3.875 $Y=0.445 $X2=0 $Y2=0
cc_795 N_SET_B_M1005_g N_VGND_c_2102_n 0.00595177f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_796 SET_B N_VGND_c_2102_n 0.00248323f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_797 N_SET_B_c_963_n N_VGND_c_2102_n 0.165266f $X=7.46 $Y=0.85 $X2=0 $Y2=0
cc_798 N_SET_B_c_964_n N_VGND_c_2102_n 0.014763f $X=4.07 $Y=0.85 $X2=0 $Y2=0
cc_799 N_SET_B_c_965_n N_VGND_c_2102_n 0.0141642f $X=7.605 $Y=0.85 $X2=0 $Y2=0
cc_800 N_SET_B_c_966_n N_VGND_c_2102_n 0.00284893f $X=7.605 $Y=0.85 $X2=0 $Y2=0
cc_801 N_SET_B_c_963_n N_A_790_47#_M1037_d 0.00177886f $X=7.46 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_802 N_SET_B_c_964_n N_A_790_47#_M1037_d 6.34838e-19 $X=4.07 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_803 N_SET_B_c_963_n N_A_790_47#_M1042_d 0.00184007f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_804 N_SET_B_c_963_n N_A_790_47#_c_2285_n 0.00611167f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_805 N_SET_B_c_963_n N_A_790_47#_c_2286_n 0.00346721f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_806 N_SET_B_M1037_g N_A_790_47#_c_2297_n 0.0039841f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_807 SET_B N_A_790_47#_c_2297_n 0.00361223f $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_808 N_SET_B_c_963_n N_A_790_47#_c_2297_n 0.00386944f $X=7.46 $Y=0.85 $X2=0
+ $Y2=0
cc_809 N_SET_B_c_964_n N_A_790_47#_c_2297_n 0.00238177f $X=4.07 $Y=0.85 $X2=0
+ $Y2=0
cc_810 N_SET_B_c_963_n A_1162_47# 0.00369541f $X=7.46 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_811 N_SET_B_M1005_g N_A_1547_47#_c_2318_n 0.00349862f $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_812 N_SET_B_c_966_n N_A_1547_47#_c_2318_n 0.00344477f $X=7.605 $Y=0.85 $X2=0
+ $Y2=0
cc_813 N_SET_B_c_967_n N_A_1547_47#_c_2318_n 2.8008e-19 $X=7.65 $Y=0.98 $X2=0
+ $Y2=0
cc_814 N_A_476_47#_M1035_g N_A_944_21#_M1042_g 0.0306362f $X=4.375 $Y=0.555
+ $X2=0 $Y2=0
cc_815 N_A_476_47#_M1020_g N_A_944_21#_M1032_g 0.0354948f $X=4.395 $Y=2.065
+ $X2=0 $Y2=0
cc_816 N_A_476_47#_c_1092_n N_A_944_21#_c_1199_n 0.0354948f $X=4.275 $Y=1.32
+ $X2=0 $Y2=0
cc_817 N_A_476_47#_M1020_g N_VPWR_c_1757_n 0.00136797f $X=4.395 $Y=2.065 $X2=0
+ $Y2=0
cc_818 N_A_476_47#_M1020_g N_VPWR_c_1764_n 0.00432313f $X=4.395 $Y=2.065 $X2=0
+ $Y2=0
cc_819 N_A_476_47#_c_1099_n N_VPWR_c_1770_n 0.0377433f $X=3.01 $Y=2.335 $X2=0
+ $Y2=0
cc_820 N_A_476_47#_M1018_d N_VPWR_c_1754_n 0.00173085f $X=2.38 $Y=2.065 $X2=0
+ $Y2=0
cc_821 N_A_476_47#_M1020_g N_VPWR_c_1754_n 0.0059524f $X=4.395 $Y=2.065 $X2=0
+ $Y2=0
cc_822 N_A_476_47#_c_1099_n N_VPWR_c_1754_n 0.0132511f $X=3.01 $Y=2.335 $X2=0
+ $Y2=0
cc_823 N_A_476_47#_c_1099_n N_A_381_47#_c_1961_n 0.010625f $X=3.01 $Y=2.335
+ $X2=0 $Y2=0
cc_824 N_A_476_47#_c_1099_n A_560_413# 0.00858887f $X=3.01 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_825 N_A_476_47#_c_1094_n A_560_413# 0.00579571f $X=3.095 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_826 N_A_476_47#_c_1100_n N_VGND_c_2086_n 0.0547511f $X=3.24 $Y=0.365 $X2=0
+ $Y2=0
cc_827 N_A_476_47#_M1035_g N_VGND_c_2088_n 0.00357877f $X=4.375 $Y=0.555 $X2=0
+ $Y2=0
cc_828 N_A_476_47#_M1036_d N_VGND_c_2102_n 0.00266057f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_829 N_A_476_47#_M1035_g N_VGND_c_2102_n 0.00545888f $X=4.375 $Y=0.555 $X2=0
+ $Y2=0
cc_830 N_A_476_47#_c_1100_n N_VGND_c_2102_n 0.021542f $X=3.24 $Y=0.365 $X2=0
+ $Y2=0
cc_831 N_A_476_47#_c_1100_n A_584_47# 0.00625863f $X=3.24 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_832 N_A_476_47#_M1035_g N_A_790_47#_c_2285_n 0.00927812f $X=4.375 $Y=0.555
+ $X2=0 $Y2=0
cc_833 N_A_476_47#_c_1090_n N_A_790_47#_c_2297_n 0.00119392f $X=4.11 $Y=1.32
+ $X2=0 $Y2=0
cc_834 N_A_476_47#_c_1092_n N_A_790_47#_c_2297_n 5.73033e-19 $X=4.275 $Y=1.32
+ $X2=0 $Y2=0
cc_835 N_A_944_21#_c_1208_n N_A_1431_21#_M1024_g 0.00413345f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_836 N_A_944_21#_c_1208_n N_A_1431_21#_c_1372_n 0.015309f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_837 N_A_944_21#_c_1208_n N_A_1431_21#_c_1373_n 0.00677286f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_838 N_A_944_21#_c_1208_n N_A_1431_21#_c_1374_n 0.010417f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_839 N_A_944_21#_c_1208_n N_A_1431_21#_c_1400_n 0.00964432f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_840 N_A_944_21#_M1043_g N_A_1431_21#_c_1362_n 0.0128951f $X=8.61 $Y=2.065
+ $X2=0 $Y2=0
cc_841 N_A_944_21#_M1016_g N_A_1431_21#_c_1362_n 0.00626744f $X=8.67 $Y=0.555
+ $X2=0 $Y2=0
cc_842 N_A_944_21#_c_1196_n N_A_1431_21#_c_1362_n 0.00727786f $X=9.07 $Y=0.84
+ $X2=0 $Y2=0
cc_843 N_A_944_21#_c_1204_n N_A_1431_21#_c_1362_n 0.0130479f $X=9.07 $Y=1.66
+ $X2=0 $Y2=0
cc_844 N_A_944_21#_c_1208_n N_A_1431_21#_c_1362_n 0.0270698f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_845 N_A_944_21#_c_1211_n N_A_1431_21#_c_1362_n 5.62937e-19 $X=8.985 $Y=1.53
+ $X2=0 $Y2=0
cc_846 N_A_944_21#_c_1200_n N_A_1431_21#_c_1362_n 0.00930156f $X=8.67 $Y=1.32
+ $X2=0 $Y2=0
cc_847 N_A_944_21#_c_1201_n N_A_1431_21#_c_1362_n 0.046128f $X=8.88 $Y=1.32
+ $X2=0 $Y2=0
cc_848 N_A_944_21#_M1001_s N_A_1431_21#_c_1376_n 0.00522551f $X=9.28 $Y=1.505
+ $X2=0 $Y2=0
cc_849 N_A_944_21#_M1043_g N_A_1431_21#_c_1376_n 0.00712539f $X=8.61 $Y=2.065
+ $X2=0 $Y2=0
cc_850 N_A_944_21#_c_1204_n N_A_1431_21#_c_1376_n 0.0212381f $X=9.07 $Y=1.66
+ $X2=0 $Y2=0
cc_851 N_A_944_21#_c_1205_n N_A_1431_21#_c_1376_n 0.0322551f $X=9.405 $Y=1.66
+ $X2=0 $Y2=0
cc_852 N_A_944_21#_c_1208_n N_A_1431_21#_c_1376_n 0.00648571f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_853 N_A_944_21#_c_1211_n N_A_1431_21#_c_1376_n 0.00170504f $X=8.985 $Y=1.53
+ $X2=0 $Y2=0
cc_854 N_A_944_21#_c_1200_n N_A_1431_21#_c_1376_n 0.0026574f $X=8.67 $Y=1.32
+ $X2=0 $Y2=0
cc_855 N_A_944_21#_c_1205_n N_A_1431_21#_c_1377_n 0.00790422f $X=9.405 $Y=1.66
+ $X2=0 $Y2=0
cc_856 N_A_944_21#_c_1208_n N_A_1431_21#_c_1417_n 0.00453864f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_857 N_A_944_21#_M1016_g N_A_1431_21#_c_1393_n 0.00431602f $X=8.67 $Y=0.555
+ $X2=0 $Y2=0
cc_858 N_A_944_21#_c_1197_n N_A_1431_21#_c_1393_n 0.00435313f $X=9.415 $Y=0.43
+ $X2=0 $Y2=0
cc_859 N_A_944_21#_M1043_g N_A_1431_21#_c_1420_n 0.00499743f $X=8.61 $Y=2.065
+ $X2=0 $Y2=0
cc_860 N_A_944_21#_M1016_g N_A_1257_47#_M1008_g 0.0191895f $X=8.67 $Y=0.555
+ $X2=0 $Y2=0
cc_861 N_A_944_21#_M1043_g N_A_1257_47#_M1039_g 0.039703f $X=8.61 $Y=2.065 $X2=0
+ $Y2=0
cc_862 N_A_944_21#_c_1208_n N_A_1257_47#_M1039_g 0.00713863f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_863 N_A_944_21#_c_1208_n N_A_1257_47#_c_1554_n 0.0219541f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_864 N_A_944_21#_c_1208_n N_A_1257_47#_c_1549_n 0.0228947f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_865 N_A_944_21#_M1016_g N_A_1257_47#_c_1551_n 2.36981e-19 $X=8.67 $Y=0.555
+ $X2=0 $Y2=0
cc_866 N_A_944_21#_c_1208_n N_A_1257_47#_c_1551_n 0.00714757f $X=8.84 $Y=1.53
+ $X2=0 $Y2=0
cc_867 N_A_944_21#_c_1200_n N_A_1257_47#_c_1552_n 0.0588925f $X=8.67 $Y=1.32
+ $X2=0 $Y2=0
cc_868 N_A_944_21#_c_1195_n N_RESET_B_M1027_g 0.00679798f $X=9.28 $Y=0.84 $X2=0
+ $Y2=0
cc_869 N_A_944_21#_c_1197_n N_RESET_B_M1027_g 0.0028847f $X=9.415 $Y=0.43 $X2=0
+ $Y2=0
cc_870 N_A_944_21#_c_1201_n N_RESET_B_M1027_g 0.00231874f $X=8.88 $Y=1.32 $X2=0
+ $Y2=0
cc_871 N_A_944_21#_c_1205_n N_RESET_B_M1001_g 0.00264716f $X=9.405 $Y=1.66 $X2=0
+ $Y2=0
cc_872 N_A_944_21#_c_1211_n N_RESET_B_M1001_g 0.00261411f $X=8.985 $Y=1.53 $X2=0
+ $Y2=0
cc_873 N_A_944_21#_c_1200_n N_RESET_B_M1001_g 0.00233488f $X=8.67 $Y=1.32 $X2=0
+ $Y2=0
cc_874 N_A_944_21#_c_1201_n N_RESET_B_M1001_g 0.00300666f $X=8.88 $Y=1.32 $X2=0
+ $Y2=0
cc_875 N_A_944_21#_c_1195_n RESET_B 0.0203337f $X=9.28 $Y=0.84 $X2=0 $Y2=0
cc_876 N_A_944_21#_c_1205_n RESET_B 0.0156391f $X=9.405 $Y=1.66 $X2=0 $Y2=0
cc_877 N_A_944_21#_c_1200_n RESET_B 5.55669e-19 $X=8.67 $Y=1.32 $X2=0 $Y2=0
cc_878 N_A_944_21#_c_1201_n RESET_B 0.0185921f $X=8.88 $Y=1.32 $X2=0 $Y2=0
cc_879 N_A_944_21#_M1016_g N_RESET_B_c_1648_n 0.00205043f $X=8.67 $Y=0.555 $X2=0
+ $Y2=0
cc_880 N_A_944_21#_c_1195_n N_RESET_B_c_1648_n 0.00563333f $X=9.28 $Y=0.84 $X2=0
+ $Y2=0
cc_881 N_A_944_21#_c_1205_n N_RESET_B_c_1648_n 0.00581996f $X=9.405 $Y=1.66
+ $X2=0 $Y2=0
cc_882 N_A_944_21#_c_1200_n N_RESET_B_c_1648_n 0.00924079f $X=8.67 $Y=1.32 $X2=0
+ $Y2=0
cc_883 N_A_944_21#_c_1201_n N_RESET_B_c_1648_n 0.00328056f $X=8.88 $Y=1.32 $X2=0
+ $Y2=0
cc_884 N_A_944_21#_c_1198_n N_VPWR_M1032_d 0.00320447f $X=5.035 $Y=1.32 $X2=0
+ $Y2=0
cc_885 N_A_944_21#_c_1210_n N_VPWR_M1032_d 0.00221031f $X=5.765 $Y=1.53 $X2=0
+ $Y2=0
cc_886 N_A_944_21#_c_1204_n N_VPWR_M1043_d 0.00311394f $X=9.07 $Y=1.66 $X2=0
+ $Y2=0
cc_887 N_A_944_21#_M1032_g N_VPWR_c_1758_n 0.0034982f $X=4.795 $Y=2.065 $X2=0
+ $Y2=0
cc_888 N_A_944_21#_c_1198_n N_VPWR_c_1758_n 0.0121469f $X=5.035 $Y=1.32 $X2=0
+ $Y2=0
cc_889 N_A_944_21#_c_1199_n N_VPWR_c_1758_n 0.00112967f $X=5.035 $Y=1.32 $X2=0
+ $Y2=0
cc_890 N_A_944_21#_c_1210_n N_VPWR_c_1758_n 7.83548e-19 $X=5.765 $Y=1.53 $X2=0
+ $Y2=0
cc_891 N_A_944_21#_M1032_g N_VPWR_c_1764_n 0.00585385f $X=4.795 $Y=2.065 $X2=0
+ $Y2=0
cc_892 N_A_944_21#_M1043_g N_VPWR_c_1766_n 0.0111257f $X=8.61 $Y=2.065 $X2=0
+ $Y2=0
cc_893 N_A_944_21#_M1043_g N_VPWR_c_1767_n 0.00339278f $X=8.61 $Y=2.065 $X2=0
+ $Y2=0
cc_894 N_A_944_21#_M1032_g N_VPWR_c_1754_n 0.00674623f $X=4.795 $Y=2.065 $X2=0
+ $Y2=0
cc_895 N_A_944_21#_M1043_g N_VPWR_c_1754_n 0.0038354f $X=8.61 $Y=2.065 $X2=0
+ $Y2=0
cc_896 N_A_944_21#_c_1210_n A_1115_329# 0.00272182f $X=5.765 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_897 N_A_944_21#_M1042_g N_VGND_c_2078_n 0.00307943f $X=4.795 $Y=0.555 $X2=0
+ $Y2=0
cc_898 N_A_944_21#_c_1195_n N_VGND_c_2080_n 0.00347746f $X=9.28 $Y=0.84 $X2=0
+ $Y2=0
cc_899 N_A_944_21#_c_1197_n N_VGND_c_2080_n 0.00624747f $X=9.415 $Y=0.43 $X2=0
+ $Y2=0
cc_900 N_A_944_21#_M1042_g N_VGND_c_2088_n 0.00357877f $X=4.795 $Y=0.555 $X2=0
+ $Y2=0
cc_901 N_A_944_21#_M1016_g N_VGND_c_2094_n 0.00357877f $X=8.67 $Y=0.555 $X2=0
+ $Y2=0
cc_902 N_A_944_21#_c_1195_n N_VGND_c_2094_n 0.00300947f $X=9.28 $Y=0.84 $X2=0
+ $Y2=0
cc_903 N_A_944_21#_c_1196_n N_VGND_c_2094_n 0.00166179f $X=9.07 $Y=0.84 $X2=0
+ $Y2=0
cc_904 N_A_944_21#_c_1197_n N_VGND_c_2094_n 0.0143536f $X=9.415 $Y=0.43 $X2=0
+ $Y2=0
cc_905 N_A_944_21#_M1027_s N_VGND_c_2102_n 0.00404615f $X=9.29 $Y=0.235 $X2=0
+ $Y2=0
cc_906 N_A_944_21#_M1042_g N_VGND_c_2102_n 0.00661646f $X=4.795 $Y=0.555 $X2=0
+ $Y2=0
cc_907 N_A_944_21#_M1016_g N_VGND_c_2102_n 0.00657041f $X=8.67 $Y=0.555 $X2=0
+ $Y2=0
cc_908 N_A_944_21#_c_1195_n N_VGND_c_2102_n 0.00541125f $X=9.28 $Y=0.84 $X2=0
+ $Y2=0
cc_909 N_A_944_21#_c_1196_n N_VGND_c_2102_n 0.00329575f $X=9.07 $Y=0.84 $X2=0
+ $Y2=0
cc_910 N_A_944_21#_c_1197_n N_VGND_c_2102_n 0.00834371f $X=9.415 $Y=0.43 $X2=0
+ $Y2=0
cc_911 N_A_944_21#_M1042_g N_A_790_47#_c_2285_n 0.0106822f $X=4.795 $Y=0.555
+ $X2=0 $Y2=0
cc_912 N_A_944_21#_c_1196_n N_A_1547_47#_M1016_d 0.0043454f $X=9.07 $Y=0.84
+ $X2=0 $Y2=0
cc_913 N_A_944_21#_M1016_g N_A_1547_47#_c_2322_n 0.0112006f $X=8.67 $Y=0.555
+ $X2=0 $Y2=0
cc_914 N_A_944_21#_c_1196_n N_A_1547_47#_c_2323_n 0.0133877f $X=9.07 $Y=0.84
+ $X2=0 $Y2=0
cc_915 N_A_944_21#_c_1197_n N_A_1547_47#_c_2323_n 0.0155579f $X=9.415 $Y=0.43
+ $X2=0 $Y2=0
cc_916 N_A_944_21#_c_1200_n N_A_1547_47#_c_2323_n 5.38954e-19 $X=8.67 $Y=1.32
+ $X2=0 $Y2=0
cc_917 N_A_1431_21#_c_1362_n N_A_1257_47#_M1008_g 0.0153921f $X=8.535 $Y=1.915
+ $X2=0 $Y2=0
cc_918 N_A_1431_21#_c_1393_n N_A_1257_47#_M1008_g 0.00536261f $X=8.535 $Y=0.687
+ $X2=0 $Y2=0
cc_919 N_A_1431_21#_c_1400_n N_A_1257_47#_M1039_g 0.0118664f $X=8.445 $Y=2 $X2=0
+ $Y2=0
cc_920 N_A_1431_21#_M1034_g N_A_1257_47#_c_1559_n 0.00204127f $X=7.23 $Y=2.275
+ $X2=0 $Y2=0
cc_921 N_A_1431_21#_M1024_g N_A_1257_47#_c_1562_n 0.0017558f $X=7.23 $Y=0.445
+ $X2=0 $Y2=0
cc_922 N_A_1431_21#_M1024_g N_A_1257_47#_c_1548_n 0.0128435f $X=7.23 $Y=0.445
+ $X2=0 $Y2=0
cc_923 N_A_1431_21#_M1024_g N_A_1257_47#_c_1554_n 0.0148682f $X=7.23 $Y=0.445
+ $X2=0 $Y2=0
cc_924 N_A_1431_21#_c_1372_n N_A_1257_47#_c_1554_n 0.0248026f $X=7.35 $Y=1.74
+ $X2=0 $Y2=0
cc_925 N_A_1431_21#_c_1429_p N_A_1257_47#_c_1554_n 0.0135579f $X=7.515 $Y=2
+ $X2=0 $Y2=0
cc_926 N_A_1431_21#_M1024_g N_A_1257_47#_c_1549_n 0.0115171f $X=7.23 $Y=0.445
+ $X2=0 $Y2=0
cc_927 N_A_1431_21#_c_1372_n N_A_1257_47#_c_1549_n 0.0154844f $X=7.35 $Y=1.74
+ $X2=0 $Y2=0
cc_928 N_A_1431_21#_c_1373_n N_A_1257_47#_c_1549_n 0.00126891f $X=7.35 $Y=1.74
+ $X2=0 $Y2=0
cc_929 N_A_1431_21#_c_1374_n N_A_1257_47#_c_1549_n 0.00635717f $X=7.955 $Y=2
+ $X2=0 $Y2=0
cc_930 N_A_1431_21#_c_1417_n N_A_1257_47#_c_1549_n 0.00162703f $X=8.04 $Y=2
+ $X2=0 $Y2=0
cc_931 N_A_1431_21#_c_1400_n N_A_1257_47#_c_1551_n 0.00158774f $X=8.445 $Y=2
+ $X2=0 $Y2=0
cc_932 N_A_1431_21#_c_1362_n N_A_1257_47#_c_1551_n 0.0241621f $X=8.535 $Y=1.915
+ $X2=0 $Y2=0
cc_933 N_A_1431_21#_c_1417_n N_A_1257_47#_c_1551_n 9.97507e-19 $X=8.04 $Y=2
+ $X2=0 $Y2=0
cc_934 N_A_1431_21#_c_1417_n N_A_1257_47#_c_1552_n 4.0151e-19 $X=8.04 $Y=2 $X2=0
+ $Y2=0
cc_935 N_A_1431_21#_c_1352_n N_RESET_B_M1027_g 0.0181841f $X=10.115 $Y=0.995
+ $X2=0 $Y2=0
cc_936 N_A_1431_21#_c_1356_n N_RESET_B_M1027_g 0.0206659f $X=10.61 $Y=1.16 $X2=0
+ $Y2=0
cc_937 N_A_1431_21#_c_1363_n N_RESET_B_M1027_g 0.00215032f $X=10.055 $Y=1.16
+ $X2=0 $Y2=0
cc_938 N_A_1431_21#_c_1376_n N_RESET_B_M1001_g 0.0145711f $X=9.9 $Y=2 $X2=0
+ $Y2=0
cc_939 N_A_1431_21#_c_1377_n N_RESET_B_M1001_g 0.00498182f $X=9.985 $Y=1.915
+ $X2=0 $Y2=0
cc_940 N_A_1431_21#_c_1356_n RESET_B 7.65575e-19 $X=10.61 $Y=1.16 $X2=0 $Y2=0
cc_941 N_A_1431_21#_c_1376_n RESET_B 0.00376763f $X=9.9 $Y=2 $X2=0 $Y2=0
cc_942 N_A_1431_21#_c_1363_n RESET_B 0.0191707f $X=10.055 $Y=1.16 $X2=0 $Y2=0
cc_943 N_A_1431_21#_M1014_g N_RESET_B_c_1648_n 0.0294515f $X=10.115 $Y=1.985
+ $X2=0 $Y2=0
cc_944 N_A_1431_21#_c_1363_n N_RESET_B_c_1648_n 0.00564908f $X=10.055 $Y=1.16
+ $X2=0 $Y2=0
cc_945 N_A_1431_21#_c_1357_n N_A_2236_47#_c_1682_n 0.00248624f $X=11.385
+ $Y=1.025 $X2=0 $Y2=0
cc_946 N_A_1431_21#_c_1359_n N_A_2236_47#_c_1682_n 0.0159717f $X=11.515 $Y=0.73
+ $X2=0 $Y2=0
cc_947 N_A_1431_21#_c_1358_n N_A_2236_47#_M1002_g 0.00455389f $X=11.385 $Y=1.535
+ $X2=0 $Y2=0
cc_948 N_A_1431_21#_c_1371_n N_A_2236_47#_M1002_g 0.0111821f $X=11.515 $Y=1.61
+ $X2=0 $Y2=0
cc_949 N_A_1431_21#_M1022_g N_A_2236_47#_c_1684_n 0.00289093f $X=10.535 $Y=0.56
+ $X2=0 $Y2=0
cc_950 N_A_1431_21#_c_1357_n N_A_2236_47#_c_1684_n 0.00371526f $X=11.385
+ $Y=1.025 $X2=0 $Y2=0
cc_951 N_A_1431_21#_c_1359_n N_A_2236_47#_c_1684_n 0.00952994f $X=11.515 $Y=0.73
+ $X2=0 $Y2=0
cc_952 N_A_1431_21#_c_1360_n N_A_2236_47#_c_1684_n 0.00973927f $X=11.515
+ $Y=0.805 $X2=0 $Y2=0
cc_953 N_A_1431_21#_M1030_g N_A_2236_47#_c_1690_n 0.00396263f $X=10.535 $Y=1.985
+ $X2=0 $Y2=0
cc_954 N_A_1431_21#_c_1358_n N_A_2236_47#_c_1690_n 0.00693146f $X=11.385
+ $Y=1.535 $X2=0 $Y2=0
cc_955 N_A_1431_21#_c_1370_n N_A_2236_47#_c_1690_n 0.0104643f $X=11.515 $Y=1.685
+ $X2=0 $Y2=0
cc_956 N_A_1431_21#_c_1371_n N_A_2236_47#_c_1690_n 0.0101644f $X=11.515 $Y=1.61
+ $X2=0 $Y2=0
cc_957 N_A_1431_21#_c_1360_n N_A_2236_47#_c_1685_n 0.00384385f $X=11.515
+ $Y=0.805 $X2=0 $Y2=0
cc_958 N_A_1431_21#_c_1371_n N_A_2236_47#_c_1685_n 0.0033881f $X=11.515 $Y=1.61
+ $X2=0 $Y2=0
cc_959 N_A_1431_21#_M1022_g N_A_2236_47#_c_1686_n 5.62277e-19 $X=10.535 $Y=0.56
+ $X2=0 $Y2=0
cc_960 N_A_1431_21#_M1030_g N_A_2236_47#_c_1686_n 5.62277e-19 $X=10.535 $Y=1.985
+ $X2=0 $Y2=0
cc_961 N_A_1431_21#_c_1355_n N_A_2236_47#_c_1686_n 0.0166518f $X=11.31 $Y=1.16
+ $X2=0 $Y2=0
cc_962 N_A_1431_21#_c_1357_n N_A_2236_47#_c_1686_n 0.00114357f $X=11.385
+ $Y=1.025 $X2=0 $Y2=0
cc_963 N_A_1431_21#_c_1358_n N_A_2236_47#_c_1686_n 0.00114357f $X=11.385
+ $Y=1.535 $X2=0 $Y2=0
cc_964 N_A_1431_21#_c_1361_n N_A_2236_47#_c_1686_n 0.00732445f $X=11.385 $Y=1.16
+ $X2=0 $Y2=0
cc_965 N_A_1431_21#_c_1357_n N_A_2236_47#_c_1687_n 0.0132039f $X=11.385 $Y=1.025
+ $X2=0 $Y2=0
cc_966 N_A_1431_21#_c_1374_n N_VPWR_M1034_d 0.00124767f $X=7.955 $Y=2 $X2=0
+ $Y2=0
cc_967 N_A_1431_21#_c_1429_p N_VPWR_M1034_d 0.00160397f $X=7.515 $Y=2 $X2=0
+ $Y2=0
cc_968 N_A_1431_21#_c_1376_n N_VPWR_M1043_d 0.0044189f $X=9.9 $Y=2 $X2=0 $Y2=0
cc_969 N_A_1431_21#_c_1376_n N_VPWR_M1001_d 0.00750664f $X=9.9 $Y=2 $X2=0 $Y2=0
cc_970 N_A_1431_21#_c_1377_n N_VPWR_M1001_d 0.00494076f $X=9.985 $Y=1.915 $X2=0
+ $Y2=0
cc_971 N_A_1431_21#_M1030_g N_VPWR_c_1759_n 0.00636974f $X=10.535 $Y=1.985 $X2=0
+ $Y2=0
cc_972 N_A_1431_21#_c_1355_n N_VPWR_c_1759_n 0.00589606f $X=11.31 $Y=1.16 $X2=0
+ $Y2=0
cc_973 N_A_1431_21#_c_1358_n N_VPWR_c_1759_n 7.93027e-19 $X=11.385 $Y=1.535
+ $X2=0 $Y2=0
cc_974 N_A_1431_21#_c_1370_n N_VPWR_c_1759_n 0.00410891f $X=11.515 $Y=1.685
+ $X2=0 $Y2=0
cc_975 N_A_1431_21#_c_1370_n N_VPWR_c_1760_n 0.00471278f $X=11.515 $Y=1.685
+ $X2=0 $Y2=0
cc_976 N_A_1431_21#_c_1370_n N_VPWR_c_1761_n 0.00513511f $X=11.515 $Y=1.685
+ $X2=0 $Y2=0
cc_977 N_A_1431_21#_c_1376_n N_VPWR_c_1766_n 0.0863621f $X=9.9 $Y=2 $X2=0 $Y2=0
cc_978 N_A_1431_21#_c_1374_n N_VPWR_c_1767_n 0.00359839f $X=7.955 $Y=2 $X2=0
+ $Y2=0
cc_979 N_A_1431_21#_c_1483_p N_VPWR_c_1767_n 0.00713694f $X=8.04 $Y=2.21 $X2=0
+ $Y2=0
cc_980 N_A_1431_21#_c_1400_n N_VPWR_c_1767_n 0.00458994f $X=8.445 $Y=2 $X2=0
+ $Y2=0
cc_981 N_A_1431_21#_c_1376_n N_VPWR_c_1767_n 4.74543e-19 $X=9.9 $Y=2 $X2=0 $Y2=0
cc_982 N_A_1431_21#_c_1420_n N_VPWR_c_1767_n 0.00279601f $X=8.535 $Y=2 $X2=0
+ $Y2=0
cc_983 N_A_1431_21#_M1034_g N_VPWR_c_1771_n 0.00542601f $X=7.23 $Y=2.275 $X2=0
+ $Y2=0
cc_984 N_A_1431_21#_c_1429_p N_VPWR_c_1771_n 9.91118e-19 $X=7.515 $Y=2 $X2=0
+ $Y2=0
cc_985 N_A_1431_21#_M1014_g N_VPWR_c_1773_n 0.0046653f $X=10.115 $Y=1.985 $X2=0
+ $Y2=0
cc_986 N_A_1431_21#_M1030_g N_VPWR_c_1773_n 0.00526178f $X=10.535 $Y=1.985 $X2=0
+ $Y2=0
cc_987 N_A_1431_21#_M1034_g N_VPWR_c_1778_n 0.00321606f $X=7.23 $Y=2.275 $X2=0
+ $Y2=0
cc_988 N_A_1431_21#_c_1373_n N_VPWR_c_1778_n 7.01948e-19 $X=7.35 $Y=1.74 $X2=0
+ $Y2=0
cc_989 N_A_1431_21#_c_1374_n N_VPWR_c_1778_n 0.0106677f $X=7.955 $Y=2 $X2=0
+ $Y2=0
cc_990 N_A_1431_21#_c_1429_p N_VPWR_c_1778_n 0.0126362f $X=7.515 $Y=2 $X2=0
+ $Y2=0
cc_991 N_A_1431_21#_c_1483_p N_VPWR_c_1778_n 0.00687131f $X=8.04 $Y=2.21 $X2=0
+ $Y2=0
cc_992 N_A_1431_21#_M1014_g N_VPWR_c_1779_n 0.00851349f $X=10.115 $Y=1.985 $X2=0
+ $Y2=0
cc_993 N_A_1431_21#_M1030_g N_VPWR_c_1779_n 6.62288e-19 $X=10.535 $Y=1.985 $X2=0
+ $Y2=0
cc_994 N_A_1431_21#_c_1376_n N_VPWR_c_1779_n 0.00915613f $X=9.9 $Y=2 $X2=0 $Y2=0
cc_995 N_A_1431_21#_M1013_d N_VPWR_c_1754_n 0.00327257f $X=7.845 $Y=2.065 $X2=0
+ $Y2=0
cc_996 N_A_1431_21#_M1034_g N_VPWR_c_1754_n 0.00997697f $X=7.23 $Y=2.275 $X2=0
+ $Y2=0
cc_997 N_A_1431_21#_M1014_g N_VPWR_c_1754_n 0.00791913f $X=10.115 $Y=1.985 $X2=0
+ $Y2=0
cc_998 N_A_1431_21#_M1030_g N_VPWR_c_1754_n 0.0105468f $X=10.535 $Y=1.985 $X2=0
+ $Y2=0
cc_999 N_A_1431_21#_c_1370_n N_VPWR_c_1754_n 0.00941266f $X=11.515 $Y=1.685
+ $X2=0 $Y2=0
cc_1000 N_A_1431_21#_c_1374_n N_VPWR_c_1754_n 0.00704318f $X=7.955 $Y=2 $X2=0
+ $Y2=0
cc_1001 N_A_1431_21#_c_1429_p N_VPWR_c_1754_n 0.00270501f $X=7.515 $Y=2 $X2=0
+ $Y2=0
cc_1002 N_A_1431_21#_c_1483_p N_VPWR_c_1754_n 0.00608739f $X=8.04 $Y=2.21 $X2=0
+ $Y2=0
cc_1003 N_A_1431_21#_c_1400_n N_VPWR_c_1754_n 0.00829558f $X=8.445 $Y=2 $X2=0
+ $Y2=0
cc_1004 N_A_1431_21#_c_1376_n N_VPWR_c_1754_n 0.00700558f $X=9.9 $Y=2 $X2=0
+ $Y2=0
cc_1005 N_A_1431_21#_c_1420_n N_VPWR_c_1754_n 0.0049407f $X=8.535 $Y=2 $X2=0
+ $Y2=0
cc_1006 N_A_1431_21#_c_1400_n A_1665_329# 0.00202121f $X=8.445 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1007 N_A_1431_21#_c_1362_n A_1665_329# 0.00305059f $X=8.535 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1008 N_A_1431_21#_c_1420_n A_1665_329# 5.84995e-19 $X=8.535 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1009 N_A_1431_21#_M1030_g N_Q_N_c_2032_n 0.00155132f $X=10.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1010 N_A_1431_21#_c_1356_n N_Q_N_c_2032_n 0.00146072f $X=10.61 $Y=1.16 $X2=0
+ $Y2=0
cc_1011 N_A_1431_21#_c_1352_n N_Q_N_c_2030_n 0.00485794f $X=10.115 $Y=0.995
+ $X2=0 $Y2=0
cc_1012 N_A_1431_21#_M1022_g N_Q_N_c_2030_n 0.00977427f $X=10.535 $Y=0.56 $X2=0
+ $Y2=0
cc_1013 N_A_1431_21#_M1030_g N_Q_N_c_2030_n 0.0112823f $X=10.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1014 N_A_1431_21#_c_1356_n N_Q_N_c_2030_n 0.0249052f $X=10.61 $Y=1.16 $X2=0
+ $Y2=0
cc_1015 N_A_1431_21#_c_1377_n N_Q_N_c_2030_n 0.0161779f $X=9.985 $Y=1.915 $X2=0
+ $Y2=0
cc_1016 N_A_1431_21#_c_1363_n N_Q_N_c_2030_n 0.0222693f $X=10.055 $Y=1.16 $X2=0
+ $Y2=0
cc_1017 N_A_1431_21#_M1022_g Q_N 0.00155132f $X=10.535 $Y=0.56 $X2=0 $Y2=0
cc_1018 N_A_1431_21#_c_1356_n Q_N 0.00141867f $X=10.61 $Y=1.16 $X2=0 $Y2=0
cc_1019 N_A_1431_21#_M1030_g Q_N 0.00974836f $X=10.535 $Y=1.985 $X2=0 $Y2=0
cc_1020 N_A_1431_21#_M1022_g N_Q_N_c_2043_n 0.00514122f $X=10.535 $Y=0.56 $X2=0
+ $Y2=0
cc_1021 N_A_1431_21#_M1024_g N_VGND_c_2079_n 0.00846638f $X=7.23 $Y=0.445 $X2=0
+ $Y2=0
cc_1022 N_A_1431_21#_c_1352_n N_VGND_c_2080_n 0.0106158f $X=10.115 $Y=0.995
+ $X2=0 $Y2=0
cc_1023 N_A_1431_21#_M1022_g N_VGND_c_2080_n 7.74e-19 $X=10.535 $Y=0.56 $X2=0
+ $Y2=0
cc_1024 N_A_1431_21#_c_1356_n N_VGND_c_2080_n 7.52163e-19 $X=10.61 $Y=1.16 $X2=0
+ $Y2=0
cc_1025 N_A_1431_21#_c_1363_n N_VGND_c_2080_n 0.0110684f $X=10.055 $Y=1.16 $X2=0
+ $Y2=0
cc_1026 N_A_1431_21#_M1022_g N_VGND_c_2081_n 0.00507375f $X=10.535 $Y=0.56 $X2=0
+ $Y2=0
cc_1027 N_A_1431_21#_c_1355_n N_VGND_c_2081_n 0.0061362f $X=11.31 $Y=1.16 $X2=0
+ $Y2=0
cc_1028 N_A_1431_21#_c_1359_n N_VGND_c_2081_n 0.00363002f $X=11.515 $Y=0.73
+ $X2=0 $Y2=0
cc_1029 N_A_1431_21#_c_1360_n N_VGND_c_2081_n 5.57729e-19 $X=11.515 $Y=0.805
+ $X2=0 $Y2=0
cc_1030 N_A_1431_21#_c_1359_n N_VGND_c_2082_n 0.00541359f $X=11.515 $Y=0.73
+ $X2=0 $Y2=0
cc_1031 N_A_1431_21#_c_1360_n N_VGND_c_2082_n 2.96334e-19 $X=11.515 $Y=0.805
+ $X2=0 $Y2=0
cc_1032 N_A_1431_21#_c_1359_n N_VGND_c_2083_n 0.00420958f $X=11.515 $Y=0.73
+ $X2=0 $Y2=0
cc_1033 N_A_1431_21#_M1024_g N_VGND_c_2090_n 0.0046653f $X=7.23 $Y=0.445 $X2=0
+ $Y2=0
cc_1034 N_A_1431_21#_c_1352_n N_VGND_c_2095_n 0.0046653f $X=10.115 $Y=0.995
+ $X2=0 $Y2=0
cc_1035 N_A_1431_21#_M1022_g N_VGND_c_2095_n 0.00526178f $X=10.535 $Y=0.56 $X2=0
+ $Y2=0
cc_1036 N_A_1431_21#_M1008_d N_VGND_c_2102_n 0.00216833f $X=8.325 $Y=0.235 $X2=0
+ $Y2=0
cc_1037 N_A_1431_21#_M1024_g N_VGND_c_2102_n 0.00460207f $X=7.23 $Y=0.445 $X2=0
+ $Y2=0
cc_1038 N_A_1431_21#_c_1352_n N_VGND_c_2102_n 0.00796766f $X=10.115 $Y=0.995
+ $X2=0 $Y2=0
cc_1039 N_A_1431_21#_M1022_g N_VGND_c_2102_n 0.0105468f $X=10.535 $Y=0.56 $X2=0
+ $Y2=0
cc_1040 N_A_1431_21#_c_1359_n N_VGND_c_2102_n 0.0110992f $X=11.515 $Y=0.73 $X2=0
+ $Y2=0
cc_1041 N_A_1431_21#_M1008_d N_A_1547_47#_c_2322_n 0.00312752f $X=8.325 $Y=0.235
+ $X2=0 $Y2=0
cc_1042 N_A_1431_21#_c_1393_n N_A_1547_47#_c_2322_n 0.0145304f $X=8.535 $Y=0.687
+ $X2=0 $Y2=0
cc_1043 N_A_1257_47#_M1039_g N_VPWR_c_1766_n 0.00209073f $X=8.25 $Y=2.065 $X2=0
+ $Y2=0
cc_1044 N_A_1257_47#_M1039_g N_VPWR_c_1767_n 0.00425094f $X=8.25 $Y=2.065 $X2=0
+ $Y2=0
cc_1045 N_A_1257_47#_c_1559_n N_VPWR_c_1771_n 0.0377433f $X=6.925 $Y=2.335 $X2=0
+ $Y2=0
cc_1046 N_A_1257_47#_M1039_g N_VPWR_c_1778_n 0.00144209f $X=8.25 $Y=2.065 $X2=0
+ $Y2=0
cc_1047 N_A_1257_47#_M1031_d N_VPWR_c_1754_n 0.00205544f $X=6.295 $Y=2.065 $X2=0
+ $Y2=0
cc_1048 N_A_1257_47#_M1039_g N_VPWR_c_1754_n 0.00591666f $X=8.25 $Y=2.065 $X2=0
+ $Y2=0
cc_1049 N_A_1257_47#_c_1559_n N_VPWR_c_1754_n 0.0272797f $X=6.925 $Y=2.335 $X2=0
+ $Y2=0
cc_1050 N_A_1257_47#_c_1559_n A_1343_413# 0.0111731f $X=6.925 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1051 N_A_1257_47#_c_1554_n A_1343_413# 0.00577347f $X=7.01 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1052 N_A_1257_47#_c_1562_n N_VGND_c_2079_n 0.0155419f $X=6.925 $Y=0.365 $X2=0
+ $Y2=0
cc_1053 N_A_1257_47#_c_1548_n N_VGND_c_2079_n 0.00412668f $X=7.01 $Y=1.235 $X2=0
+ $Y2=0
cc_1054 N_A_1257_47#_c_1562_n N_VGND_c_2090_n 0.0433655f $X=6.925 $Y=0.365 $X2=0
+ $Y2=0
cc_1055 N_A_1257_47#_M1008_g N_VGND_c_2094_n 0.00357877f $X=8.25 $Y=0.555 $X2=0
+ $Y2=0
cc_1056 N_A_1257_47#_M1007_d N_VGND_c_2102_n 0.00272713f $X=6.285 $Y=0.235 $X2=0
+ $Y2=0
cc_1057 N_A_1257_47#_M1008_g N_VGND_c_2102_n 0.00569618f $X=8.25 $Y=0.555 $X2=0
+ $Y2=0
cc_1058 N_A_1257_47#_c_1562_n N_VGND_c_2102_n 0.0129183f $X=6.925 $Y=0.365 $X2=0
+ $Y2=0
cc_1059 N_A_1257_47#_c_1562_n A_1366_47# 0.0053026f $X=6.925 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1060 N_A_1257_47#_c_1548_n A_1366_47# 0.00495481f $X=7.01 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_1061 N_A_1257_47#_M1008_g N_A_1547_47#_c_2322_n 0.0110234f $X=8.25 $Y=0.555
+ $X2=0 $Y2=0
cc_1062 N_A_1257_47#_c_1551_n N_A_1547_47#_c_2322_n 0.00293167f $X=8.19 $Y=1.24
+ $X2=0 $Y2=0
cc_1063 N_A_1257_47#_c_1551_n N_A_1547_47#_c_2318_n 0.00206243f $X=8.19 $Y=1.24
+ $X2=0 $Y2=0
cc_1064 N_A_1257_47#_c_1552_n N_A_1547_47#_c_2318_n 3.6952e-19 $X=8.19 $Y=1.24
+ $X2=0 $Y2=0
cc_1065 N_RESET_B_M1001_g N_VPWR_c_1772_n 0.00655753f $X=9.63 $Y=1.825 $X2=0
+ $Y2=0
cc_1066 N_RESET_B_M1027_g N_VGND_c_2080_n 0.00666592f $X=9.63 $Y=0.445 $X2=0
+ $Y2=0
cc_1067 N_RESET_B_M1027_g N_VGND_c_2094_n 0.00585385f $X=9.63 $Y=0.445 $X2=0
+ $Y2=0
cc_1068 N_RESET_B_M1027_g N_VGND_c_2102_n 0.0120869f $X=9.63 $Y=0.445 $X2=0
+ $Y2=0
cc_1069 N_A_2236_47#_c_1690_n N_VPWR_c_1759_n 0.0478695f $X=11.305 $Y=1.91 $X2=0
+ $Y2=0
cc_1070 N_A_2236_47#_c_1690_n N_VPWR_c_1760_n 0.0136791f $X=11.305 $Y=1.91 $X2=0
+ $Y2=0
cc_1071 N_A_2236_47#_M1002_g N_VPWR_c_1761_n 0.0129007f $X=11.99 $Y=1.985 $X2=0
+ $Y2=0
cc_1072 N_A_2236_47#_M1010_g N_VPWR_c_1761_n 7.65813e-19 $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_1073 N_A_2236_47#_c_1690_n N_VPWR_c_1761_n 0.0469761f $X=11.305 $Y=1.91 $X2=0
+ $Y2=0
cc_1074 N_A_2236_47#_c_1685_n N_VPWR_c_1761_n 0.010742f $X=11.905 $Y=1.16 $X2=0
+ $Y2=0
cc_1075 N_A_2236_47#_c_1687_n N_VPWR_c_1761_n 0.00259291f $X=12.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1076 N_A_2236_47#_M1010_g N_VPWR_c_1763_n 0.00369093f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_1077 N_A_2236_47#_M1002_g N_VPWR_c_1774_n 0.0046653f $X=11.99 $Y=1.985 $X2=0
+ $Y2=0
cc_1078 N_A_2236_47#_M1010_g N_VPWR_c_1774_n 0.00571722f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_1079 N_A_2236_47#_M1002_g N_VPWR_c_1754_n 0.00796766f $X=11.99 $Y=1.985 $X2=0
+ $Y2=0
cc_1080 N_A_2236_47#_M1010_g N_VPWR_c_1754_n 0.0111841f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_1081 N_A_2236_47#_c_1690_n N_VPWR_c_1754_n 0.00936305f $X=11.305 $Y=1.91
+ $X2=0 $Y2=0
cc_1082 N_A_2236_47#_c_1683_n N_Q_c_2056_n 0.00172265f $X=12.41 $Y=0.995 $X2=0
+ $Y2=0
cc_1083 N_A_2236_47#_M1002_g N_Q_c_2054_n 0.00155635f $X=11.99 $Y=1.985 $X2=0
+ $Y2=0
cc_1084 N_A_2236_47#_M1010_g N_Q_c_2054_n 0.00273509f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_1085 N_A_2236_47#_c_1690_n N_Q_c_2054_n 0.00473041f $X=11.305 $Y=1.91 $X2=0
+ $Y2=0
cc_1086 N_A_2236_47#_c_1682_n N_Q_c_2053_n 0.00387645f $X=11.99 $Y=0.995 $X2=0
+ $Y2=0
cc_1087 N_A_2236_47#_M1002_g N_Q_c_2053_n 0.00272957f $X=11.99 $Y=1.985 $X2=0
+ $Y2=0
cc_1088 N_A_2236_47#_c_1683_n N_Q_c_2053_n 0.00618256f $X=12.41 $Y=0.995 $X2=0
+ $Y2=0
cc_1089 N_A_2236_47#_M1010_g N_Q_c_2053_n 0.00557758f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_1090 N_A_2236_47#_c_1685_n N_Q_c_2053_n 0.0251318f $X=11.905 $Y=1.16 $X2=0
+ $Y2=0
cc_1091 N_A_2236_47#_c_1687_n N_Q_c_2053_n 0.0270739f $X=12.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1092 N_A_2236_47#_c_1683_n Q 0.00541215f $X=12.41 $Y=0.995 $X2=0 $Y2=0
cc_1093 N_A_2236_47#_M1010_g Q 0.0103034f $X=12.41 $Y=1.985 $X2=0 $Y2=0
cc_1094 N_A_2236_47#_c_1684_n N_VGND_c_2081_n 0.0317632f $X=11.305 $Y=0.51 $X2=0
+ $Y2=0
cc_1095 N_A_2236_47#_c_1684_n N_VGND_c_2082_n 0.0157432f $X=11.305 $Y=0.51 $X2=0
+ $Y2=0
cc_1096 N_A_2236_47#_c_1682_n N_VGND_c_2083_n 0.0078127f $X=11.99 $Y=0.995 $X2=0
+ $Y2=0
cc_1097 N_A_2236_47#_c_1683_n N_VGND_c_2083_n 6.44631e-19 $X=12.41 $Y=0.995
+ $X2=0 $Y2=0
cc_1098 N_A_2236_47#_c_1684_n N_VGND_c_2083_n 0.0209519f $X=11.305 $Y=0.51 $X2=0
+ $Y2=0
cc_1099 N_A_2236_47#_c_1685_n N_VGND_c_2083_n 0.0104995f $X=11.905 $Y=1.16 $X2=0
+ $Y2=0
cc_1100 N_A_2236_47#_c_1687_n N_VGND_c_2083_n 0.00255976f $X=12.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1101 N_A_2236_47#_c_1683_n N_VGND_c_2085_n 0.00323465f $X=12.41 $Y=0.995
+ $X2=0 $Y2=0
cc_1102 N_A_2236_47#_c_1682_n N_VGND_c_2096_n 0.0046653f $X=11.99 $Y=0.995 $X2=0
+ $Y2=0
cc_1103 N_A_2236_47#_c_1683_n N_VGND_c_2096_n 0.00571722f $X=12.41 $Y=0.995
+ $X2=0 $Y2=0
cc_1104 N_A_2236_47#_M1017_s N_VGND_c_2102_n 0.00335098f $X=11.18 $Y=0.235 $X2=0
+ $Y2=0
cc_1105 N_A_2236_47#_c_1682_n N_VGND_c_2102_n 0.00796766f $X=11.99 $Y=0.995
+ $X2=0 $Y2=0
cc_1106 N_A_2236_47#_c_1683_n N_VGND_c_2102_n 0.0111841f $X=12.41 $Y=0.995 $X2=0
+ $Y2=0
cc_1107 N_A_2236_47#_c_1684_n N_VGND_c_2102_n 0.00961085f $X=11.305 $Y=0.51
+ $X2=0 $Y2=0
cc_1108 N_VPWR_c_1754_n N_A_381_47#_M1029_d 0.00309406f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1109 N_VPWR_c_1756_n N_A_381_47#_c_1959_n 0.011655f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_1110 N_VPWR_c_1770_n N_A_381_47#_c_1959_n 0.00221328f $X=3.42 $Y=2.72 $X2=0
+ $Y2=0
cc_1111 N_VPWR_c_1754_n N_A_381_47#_c_1959_n 0.00201225f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1112 N_VPWR_c_1756_n N_A_381_47#_c_1960_n 0.0116681f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_1113 N_VPWR_c_1769_n N_A_381_47#_c_1960_n 3.86777e-19 $X=1.445 $Y=2.72 $X2=0
+ $Y2=0
cc_1114 N_VPWR_c_1754_n N_A_381_47#_c_1960_n 7.1462e-19 $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1115 N_VPWR_c_1770_n N_A_381_47#_c_1961_n 0.0115924f $X=3.42 $Y=2.72 $X2=0
+ $Y2=0
cc_1116 N_VPWR_c_1754_n N_A_381_47#_c_1961_n 0.00307944f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1117 N_VPWR_c_1754_n A_560_413# 0.00355877f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1118 N_VPWR_c_1754_n A_894_329# 0.00239341f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1119 N_VPWR_c_1754_n A_1115_329# 0.00777501f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1120 N_VPWR_c_1754_n A_1343_413# 0.00566996f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1121 N_VPWR_c_1754_n A_1665_329# 0.00245111f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1122 N_VPWR_c_1754_n N_Q_N_M1014_d 0.00393857f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1123 N_VPWR_c_1759_n N_Q_N_c_2030_n 0.0706187f $X=10.785 $Y=1.63 $X2=0 $Y2=0
cc_1124 N_VPWR_c_1773_n Q_N 0.0158644f $X=10.68 $Y=2.72 $X2=0 $Y2=0
cc_1125 N_VPWR_c_1754_n Q_N 0.00975768f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1126 N_VPWR_c_1754_n N_Q_M1002_s 0.00393857f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1127 N_VPWR_c_1763_n N_Q_c_2054_n 0.0362378f $X=12.62 $Y=1.63 $X2=0 $Y2=0
cc_1128 N_VPWR_c_1774_n Q 0.013819f $X=12.515 $Y=2.72 $X2=0 $Y2=0
cc_1129 N_VPWR_c_1754_n Q 0.00873952f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1130 N_VPWR_c_1759_n N_VGND_c_2081_n 0.0085478f $X=10.785 $Y=1.63 $X2=0 $Y2=0
cc_1131 N_VPWR_c_1763_n N_VGND_c_2085_n 0.0101366f $X=12.62 $Y=1.63 $X2=0 $Y2=0
cc_1132 N_A_381_47#_c_1956_n N_VGND_M1011_s 0.00109803f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1133 N_A_381_47#_c_1957_n N_VGND_M1011_s 0.00109988f $X=1.59 $Y=0.73 $X2=0
+ $Y2=0
cc_1134 N_A_381_47#_c_1956_n N_VGND_c_2076_n 0.00955176f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1135 N_A_381_47#_c_1957_n N_VGND_c_2076_n 0.0114768f $X=1.59 $Y=0.73 $X2=0
+ $Y2=0
cc_1136 N_A_381_47#_c_1956_n N_VGND_c_2086_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1137 N_A_381_47#_c_1990_n N_VGND_c_2086_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1138 N_A_381_47#_c_1957_n N_VGND_c_2093_n 4.97798e-19 $X=1.59 $Y=0.73 $X2=0
+ $Y2=0
cc_1139 N_A_381_47#_M1011_d N_VGND_c_2102_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1140 N_A_381_47#_c_1956_n N_VGND_c_2102_n 0.0023552f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1141 N_A_381_47#_c_1957_n N_VGND_c_2102_n 8.52239e-19 $X=1.59 $Y=0.73 $X2=0
+ $Y2=0
cc_1142 N_A_381_47#_c_1990_n N_VGND_c_2102_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1143 N_Q_N_c_2030_n N_VGND_c_2080_n 0.00493434f $X=10.37 $Y=1.63 $X2=0 $Y2=0
cc_1144 N_Q_N_c_2043_n N_VGND_c_2081_n 0.0443217f $X=10.37 $Y=0.585 $X2=0 $Y2=0
cc_1145 N_Q_N_c_2043_n N_VGND_c_2095_n 0.0157211f $X=10.37 $Y=0.585 $X2=0 $Y2=0
cc_1146 N_Q_N_M1003_s N_VGND_c_2102_n 0.00393857f $X=10.19 $Y=0.235 $X2=0 $Y2=0
cc_1147 N_Q_N_c_2043_n N_VGND_c_2102_n 0.00972746f $X=10.37 $Y=0.585 $X2=0 $Y2=0
cc_1148 Q N_VGND_c_2096_n 0.0137848f $X=12.14 $Y=0.425 $X2=0 $Y2=0
cc_1149 N_Q_M1033_d N_VGND_c_2102_n 0.00393857f $X=12.065 $Y=0.235 $X2=0 $Y2=0
cc_1150 Q N_VGND_c_2102_n 0.00873176f $X=12.14 $Y=0.425 $X2=0 $Y2=0
cc_1151 N_VGND_c_2102_n A_584_47# 0.00230551f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1152 N_VGND_c_2102_n N_A_790_47#_M1037_d 0.00227745f $X=12.65 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1153 N_VGND_c_2102_n N_A_790_47#_M1042_d 0.00173088f $X=12.65 $Y=0 $X2=0
+ $Y2=0
cc_1154 N_VGND_c_2078_n N_A_790_47#_c_2285_n 0.0139f $X=5.525 $Y=0.38 $X2=0
+ $Y2=0
cc_1155 N_VGND_c_2088_n N_A_790_47#_c_2285_n 0.0528039f $X=5.36 $Y=0 $X2=0 $Y2=0
cc_1156 N_VGND_c_2102_n N_A_790_47#_c_2285_n 0.015297f $X=12.65 $Y=0 $X2=0 $Y2=0
cc_1157 N_VGND_c_2078_n N_A_790_47#_c_2286_n 0.00297978f $X=5.525 $Y=0.38 $X2=0
+ $Y2=0
cc_1158 N_VGND_c_2088_n N_A_790_47#_c_2297_n 0.0197166f $X=5.36 $Y=0 $X2=0 $Y2=0
cc_1159 N_VGND_c_2102_n N_A_790_47#_c_2297_n 0.00556798f $X=12.65 $Y=0 $X2=0
+ $Y2=0
cc_1160 N_VGND_c_2102_n A_1162_47# 0.00467499f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1161 N_VGND_c_2102_n A_1366_47# 0.00261578f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1162 N_VGND_c_2102_n N_A_1547_47#_M1005_d 0.00378249f $X=12.65 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1163 N_VGND_c_2102_n N_A_1547_47#_M1016_d 0.00251082f $X=12.65 $Y=0 $X2=0
+ $Y2=0
cc_1164 N_VGND_c_2094_n N_A_1547_47#_c_2322_n 0.0358653f $X=9.74 $Y=0 $X2=0
+ $Y2=0
cc_1165 N_VGND_c_2102_n N_A_1547_47#_c_2322_n 0.0235203f $X=12.65 $Y=0 $X2=0
+ $Y2=0
cc_1166 N_VGND_c_2094_n N_A_1547_47#_c_2318_n 0.0215241f $X=9.74 $Y=0 $X2=0
+ $Y2=0
cc_1167 N_VGND_c_2102_n N_A_1547_47#_c_2318_n 0.01237f $X=12.65 $Y=0 $X2=0 $Y2=0
cc_1168 N_VGND_c_2094_n N_A_1547_47#_c_2323_n 0.0110309f $X=9.74 $Y=0 $X2=0
+ $Y2=0
cc_1169 N_VGND_c_2102_n N_A_1547_47#_c_2323_n 0.0063548f $X=12.65 $Y=0 $X2=0
+ $Y2=0

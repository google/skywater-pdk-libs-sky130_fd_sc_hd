* File: sky130_fd_sc_hd__o221a_1.pex.spice
* Created: Tue Sep  1 19:22:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O221A_1%C1 1 3 6 8 9 10
c29 9 0 8.85515e-21 $X=0.67 $Y=1.16
r30 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r31 8 13 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.25 $Y2=1.16
r32 8 9 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.595 $Y=1.16 $X2=0.67
+ $Y2=1.16
r33 4 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.325
+ $X2=0.67 $Y2=1.16
r34 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.67 $Y=1.325 $X2=0.67
+ $Y2=1.985
r35 1 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=0.995
+ $X2=0.67 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.67 $Y=0.995 $X2=0.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%B1 3 6 8 11 13
r37 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.16
+ $X2=1.09 $Y2=1.325
r38 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.16
+ $X2=1.09 $Y2=0.995
r39 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.16 $X2=1.09 $Y2=1.16
r40 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.15 $Y=1.985
+ $X2=1.15 $Y2=1.325
r41 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.125 $Y=0.56
+ $X2=1.125 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%B2 3 7 8 9 13 15
c41 8 0 1.49676e-19 $X=1.61 $Y=1.19
r42 13 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.61 $Y2=1.325
r43 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.61 $Y2=0.995
r44 9 24 7.38284 $w=3.18e-07 $l=2.05e-07 $layer=LI1_cond $X=1.655 $Y=1.53
+ $X2=1.655 $Y2=1.325
r45 8 24 5.32494 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=1.16
+ $X2=1.625 $Y2=1.325
r46 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.16 $X2=1.65 $Y2=1.16
r47 7 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.545 $Y=0.56
+ $X2=1.545 $Y2=0.995
r48 3 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.51 $Y=1.985
+ $X2=1.51 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%A2 3 6 8 9 13 14 15
c35 14 0 1.96039e-19 $X=2.325 $Y=1.16
c36 9 0 3.0922e-19 $X=2.07 $Y=1.53
r37 13 16 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.16
+ $X2=2.375 $Y2=1.325
r38 13 15 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.16
+ $X2=2.375 $Y2=0.995
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.16 $X2=2.325 $Y2=1.16
r40 9 25 7.52929 $w=3.73e-07 $l=2.45e-07 $layer=LI1_cond $X=2.192 $Y=1.53
+ $X2=2.192 $Y2=1.285
r41 8 25 2.98932 $w=4.83e-07 $l=9.5e-08 $layer=LI1_cond $X=2.247 $Y=1.19
+ $X2=2.247 $Y2=1.285
r42 8 14 0.739842 $w=4.83e-07 $l=3e-08 $layer=LI1_cond $X=2.247 $Y=1.19
+ $X2=2.247 $Y2=1.16
r43 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.485 $Y=1.985
+ $X2=2.485 $Y2=1.325
r44 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.485 $Y=0.56
+ $X2=2.485 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%A1 3 5 7 8 11
c34 11 0 3.82587e-19 $X=2.905 $Y=1.16
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.16
+ $X2=2.905 $Y2=1.325
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.16 $X2=2.905 $Y2=1.16
r37 8 12 5.54545 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=3.01 $Y=1.18
+ $X2=2.905 $Y2=1.18
r38 5 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=0.995
+ $X2=2.905 $Y2=1.16
r39 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.905 $Y=0.995
+ $X2=2.905 $Y2=0.56
r40 3 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.845 $Y=1.985
+ $X2=2.845 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%A_51_297# 1 2 3 12 15 19 23 26 27 28 30 31
+ 32 34 35 36 38 46 49 54 55 58
r119 55 59 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.427 $Y=1.16
+ $X2=3.427 $Y2=1.325
r120 55 58 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.427 $Y=1.16
+ $X2=3.427 $Y2=0.995
r121 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.16 $X2=3.47 $Y2=1.16
r122 51 54 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=1.18
+ $X2=3.47 $Y2=1.18
r123 37 51 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.385 $Y=1.285
+ $X2=3.385 $Y2=1.18
r124 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.385 $Y=1.285
+ $X2=3.385 $Y2=1.455
r125 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.3 $Y=1.54
+ $X2=3.385 $Y2=1.455
r126 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.3 $Y=1.54
+ $X2=2.72 $Y2=1.54
r127 34 49 9.44516 $w=4.65e-07 $l=4.85592e-07 $layer=LI1_cond $X=2.635 $Y=1.875
+ $X2=2.275 $Y2=2.17
r128 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.635 $Y=1.625
+ $X2=2.72 $Y2=1.54
r129 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.635 $Y=1.625
+ $X2=2.635 $Y2=1.875
r130 31 49 23.5314 $w=4.65e-07 $l=7.98123e-07 $layer=LI1_cond $X=1.575 $Y=1.96
+ $X2=2.275 $Y2=2.17
r131 31 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.575 $Y=1.96
+ $X2=1.325 $Y2=1.96
r132 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.24 $Y=1.875
+ $X2=1.325 $Y2=1.96
r133 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.24 $Y=1.625
+ $X2=1.24 $Y2=1.875
r134 28 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=1.54
+ $X2=0.67 $Y2=1.54
r135 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.155 $Y=1.54
+ $X2=1.24 $Y2=1.625
r136 27 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.155 $Y=1.54
+ $X2=0.755 $Y2=1.54
r137 26 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.455
+ $X2=0.67 $Y2=1.54
r138 25 46 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.67 $Y=0.825 $X2=0.67
+ $Y2=0.735
r139 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.67 $Y=0.825
+ $X2=0.67 $Y2=1.455
r140 21 46 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=0.41 $Y=0.735
+ $X2=0.67 $Y2=0.735
r141 21 23 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.41 $Y=0.645
+ $X2=0.41 $Y2=0.39
r142 17 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.39 $Y=1.54
+ $X2=0.67 $Y2=1.54
r143 17 19 25.93 $w=2.98e-07 $l=6.75e-07 $layer=LI1_cond $X=0.39 $Y=1.625
+ $X2=0.39 $Y2=2.3
r144 15 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.325 $Y=1.985
+ $X2=3.325 $Y2=1.325
r145 12 58 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.325 $Y=0.56
+ $X2=3.325 $Y2=0.995
r146 3 49 150 $w=1.7e-07 $l=8.96577e-07 $layer=licon1_PDIFF $count=4 $X=1.585
+ $Y=1.485 $X2=2.275 $Y2=1.96
r147 2 17 400 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=1.485 $X2=0.455 $Y2=1.62
r148 2 19 400 $w=1.7e-07 $l=9.09519e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=1.485 $X2=0.455 $Y2=2.3
r149 1 21 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.235 $X2=0.41 $Y2=0.73
r150 1 23 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.235 $X2=0.41 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%VPWR 1 2 9 13 16 17 18 24 33 34 37
r48 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r49 34 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r51 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=2.72
+ $X2=3.055 $Y2=2.72
r52 31 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.22 $Y=2.72 $X2=3.91
+ $Y2=2.72
r53 30 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=2.72
+ $X2=3.055 $Y2=2.72
r59 24 29 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.89 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 22 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 16 21 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.735 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.735 $Y=2.72
+ $X2=0.86 $Y2=2.72
r65 15 26 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=0.86 $Y2=2.72
r67 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=2.635
+ $X2=3.055 $Y2=2.72
r68 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.055 $Y=2.635
+ $X2=3.055 $Y2=1.96
r69 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=2.635
+ $X2=0.86 $Y2=2.72
r70 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.86 $Y=2.635 $X2=0.86
+ $Y2=1.96
r71 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.92
+ $Y=1.485 $X2=3.055 $Y2=1.96
r72 1 9 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=0.745
+ $Y=1.485 $X2=0.9 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%X 1 2 10 13 19 24
r25 16 24 5.79663 $w=2.5e-07 $l=2.95e-07 $layer=LI1_cond $X=3.93 $Y=1.875
+ $X2=3.93 $Y2=2.17
r26 16 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.93 $Y=1.875
+ $X2=3.93 $Y2=1.87
r27 13 24 0.40545 $w=5.88e-07 $l=2e-08 $layer=LI1_cond $X=3.91 $Y=2.17 $X2=3.93
+ $Y2=2.17
r28 13 21 7.19674 $w=5.88e-07 $l=3.55e-07 $layer=LI1_cond $X=3.91 $Y=2.17
+ $X2=3.555 $Y2=2.17
r29 13 19 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.93 $Y=1.83 $X2=3.93
+ $Y2=1.87
r30 11 13 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=3.93 $Y=0.905
+ $X2=3.93 $Y2=1.83
r31 10 11 6.29411 $w=2.5e-07 $l=3.2e-07 $layer=LI1_cond $X=3.93 $Y=0.585
+ $X2=3.93 $Y2=0.905
r32 8 10 7.38205 $w=6.38e-07 $l=3.95e-07 $layer=LI1_cond $X=3.535 $Y=0.585
+ $X2=3.93 $Y2=0.585
r33 2 21 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=3.4
+ $Y=1.485 $X2=3.555 $Y2=1.96
r34 1 8 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.4
+ $Y=0.235 $X2=3.535 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%A_149_47# 1 2 11
r14 8 11 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.91 $Y=0.39
+ $X2=1.755 $Y2=0.39
r15 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.62
+ $Y=0.235 $X2=1.755 $Y2=0.39
r16 1 8 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=0.745
+ $Y=0.235 $X2=0.91 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%A_240_47# 1 2 7 11 16
r36 14 16 10.6882 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.335 $Y=0.775
+ $X2=1.545 $Y2=0.775
r37 9 11 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.695 $Y=0.735
+ $X2=2.695 $Y2=0.39
r38 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=2.695 $Y2=0.735
r39 7 16 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=1.545 $Y2=0.82
r40 2 11 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.56
+ $Y=0.235 $X2=2.695 $Y2=0.39
r41 1 14 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.235 $X2=1.335 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r51 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r52 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r53 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r54 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r55 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r56 24 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r57 21 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r58 21 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r59 19 31 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.99
+ $Y2=0
r60 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.115
+ $Y2=0
r61 18 34 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.91
+ $Y2=0
r62 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.115
+ $Y2=0
r63 16 28 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.07
+ $Y2=0
r64 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.275
+ $Y2=0
r65 15 31 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.99
+ $Y2=0
r66 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.275
+ $Y2=0
r67 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0
r68 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0.39
r69 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0.085
+ $X2=2.275 $Y2=0
r70 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.275 $Y=0.085
+ $X2=2.275 $Y2=0.39
r71 2 13 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.98
+ $Y=0.235 $X2=3.115 $Y2=0.39
r72 1 9 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.235 $X2=2.275 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__dlxbp_1.pxi.spice
* Created: Tue Sep  1 19:06:01 2020
* 
x_PM_SKY130_FD_SC_HD__DLXBP_1%GATE N_GATE_c_156_n N_GATE_c_151_n N_GATE_M1018_g
+ N_GATE_c_157_n N_GATE_M1008_g N_GATE_c_152_n N_GATE_c_158_n GATE GATE
+ N_GATE_c_154_n N_GATE_c_155_n PM_SKY130_FD_SC_HD__DLXBP_1%GATE
x_PM_SKY130_FD_SC_HD__DLXBP_1%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1008_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_M1021_g N_A_27_47#_c_195_n
+ N_A_27_47#_M1012_g N_A_27_47#_c_196_n N_A_27_47#_c_331_p N_A_27_47#_c_197_n
+ N_A_27_47#_c_198_n N_A_27_47#_c_205_n N_A_27_47#_c_206_n N_A_27_47#_c_199_n
+ N_A_27_47#_c_200_n N_A_27_47#_c_208_n N_A_27_47#_c_209_n N_A_27_47#_c_210_n
+ N_A_27_47#_c_255_p N_A_27_47#_c_211_n N_A_27_47#_c_201_n N_A_27_47#_c_202_n
+ PM_SKY130_FD_SC_HD__DLXBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLXBP_1%D N_D_c_340_n N_D_c_341_n N_D_M1002_g N_D_M1009_g
+ N_D_c_342_n N_D_c_343_n N_D_c_348_n D N_D_c_344_n N_D_c_345_n
+ PM_SKY130_FD_SC_HD__DLXBP_1%D
x_PM_SKY130_FD_SC_HD__DLXBP_1%A_299_47# N_A_299_47#_M1002_s N_A_299_47#_M1009_s
+ N_A_299_47#_M1006_g N_A_299_47#_M1005_g N_A_299_47#_c_395_n
+ N_A_299_47#_c_391_n N_A_299_47#_c_392_n N_A_299_47#_c_393_n
+ PM_SKY130_FD_SC_HD__DLXBP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLXBP_1%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_c_464_n N_A_193_47#_M1016_g N_A_193_47#_c_469_n
+ N_A_193_47#_M1013_g N_A_193_47#_c_466_n N_A_193_47#_c_467_n
+ N_A_193_47#_c_468_n N_A_193_47#_c_473_n N_A_193_47#_c_474_n
+ N_A_193_47#_c_475_n N_A_193_47#_c_476_n N_A_193_47#_c_477_n
+ N_A_193_47#_c_478_n PM_SKY130_FD_SC_HD__DLXBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLXBP_1%A_716_21# N_A_716_21#_M1020_s N_A_716_21#_M1019_s
+ N_A_716_21#_M1004_g N_A_716_21#_M1001_g N_A_716_21#_c_591_n
+ N_A_716_21#_M1017_g N_A_716_21#_M1007_g N_A_716_21#_c_592_n
+ N_A_716_21#_c_593_n N_A_716_21#_c_594_n N_A_716_21#_M1003_g
+ N_A_716_21#_M1014_g N_A_716_21#_c_603_n N_A_716_21#_c_604_n
+ N_A_716_21#_c_605_n N_A_716_21#_c_606_n N_A_716_21#_c_636_p
+ N_A_716_21#_c_595_n N_A_716_21#_c_607_n N_A_716_21#_c_596_n
+ N_A_716_21#_c_597_n N_A_716_21#_c_619_p N_A_716_21#_c_627_p
+ N_A_716_21#_c_628_p PM_SKY130_FD_SC_HD__DLXBP_1%A_716_21#
x_PM_SKY130_FD_SC_HD__DLXBP_1%A_560_47# N_A_560_47#_M1016_d N_A_560_47#_M1021_d
+ N_A_560_47#_c_706_n N_A_560_47#_M1020_g N_A_560_47#_M1019_g
+ N_A_560_47#_c_707_n N_A_560_47#_c_708_n N_A_560_47#_c_717_n
+ N_A_560_47#_c_719_n N_A_560_47#_c_709_n N_A_560_47#_c_732_n
+ N_A_560_47#_c_715_n N_A_560_47#_c_710_n N_A_560_47#_c_711_n
+ PM_SKY130_FD_SC_HD__DLXBP_1%A_560_47#
x_PM_SKY130_FD_SC_HD__DLXBP_1%A_1124_47# N_A_1124_47#_M1003_s
+ N_A_1124_47#_M1014_s N_A_1124_47#_M1015_g N_A_1124_47#_M1011_g
+ N_A_1124_47#_c_797_n N_A_1124_47#_c_802_n N_A_1124_47#_c_798_n
+ N_A_1124_47#_c_799_n N_A_1124_47#_c_816_n N_A_1124_47#_c_800_n
+ PM_SKY130_FD_SC_HD__DLXBP_1%A_1124_47#
x_PM_SKY130_FD_SC_HD__DLXBP_1%VPWR N_VPWR_M1008_d N_VPWR_M1009_d N_VPWR_M1001_d
+ N_VPWR_M1019_d N_VPWR_M1014_d N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_848_n
+ N_VPWR_c_849_n N_VPWR_c_850_n N_VPWR_c_851_n N_VPWR_c_852_n VPWR
+ N_VPWR_c_853_n N_VPWR_c_854_n N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n
+ N_VPWR_c_845_n N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n
+ PM_SKY130_FD_SC_HD__DLXBP_1%VPWR
x_PM_SKY130_FD_SC_HD__DLXBP_1%Q N_Q_M1017_d N_Q_M1007_d N_Q_c_956_n Q Q Q
+ N_Q_c_957_n Q N_Q_c_958_n PM_SKY130_FD_SC_HD__DLXBP_1%Q
x_PM_SKY130_FD_SC_HD__DLXBP_1%Q_N N_Q_N_M1015_d N_Q_N_M1011_d N_Q_N_c_984_n
+ N_Q_N_c_987_n N_Q_N_c_985_n Q_N Q_N Q_N PM_SKY130_FD_SC_HD__DLXBP_1%Q_N
x_PM_SKY130_FD_SC_HD__DLXBP_1%VGND N_VGND_M1018_d N_VGND_M1002_d N_VGND_M1004_d
+ N_VGND_M1020_d N_VGND_M1003_d N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n
+ N_VGND_c_1003_n N_VGND_c_1004_n VGND N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n
+ N_VGND_c_1015_n N_VGND_c_1016_n PM_SKY130_FD_SC_HD__DLXBP_1%VGND
cc_1 VNB N_GATE_c_151_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_152_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_c_154_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_c_155_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0398895f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_195_n 0.0228812f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_c_196_n 0.0206274f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_9 VNB N_A_27_47#_c_197_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_198_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_11 VNB N_A_27_47#_c_199_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_200_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_201_n 0.0231477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_202_n 0.021629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_D_c_340_n 0.00566197f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.07
cc_16 VNB N_D_c_341_n 0.017236f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_c_342_n 0.0315818f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_18 VNB N_D_c_343_n 0.0122081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_D_c_344_n 0.0111024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_c_345_n 0.00609199f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_21 VNB N_A_299_47#_M1006_g 0.0239837f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_22 VNB N_A_299_47#_M1005_g 0.00433259f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_23 VNB N_A_299_47#_c_391_n 0.00838199f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB N_A_299_47#_c_392_n 0.00121169f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_25 VNB N_A_299_47#_c_393_n 0.0318617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_464_n 0.0299719f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_27 VNB N_A_193_47#_M1016_g 0.0184062f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_28 VNB N_A_193_47#_c_466_n 0.0130942f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_29 VNB N_A_193_47#_c_467_n 0.00884872f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_30 VNB N_A_193_47#_c_468_n 0.00296442f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_31 VNB N_A_716_21#_M1004_g 0.0475314f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_716_21#_c_591_n 0.0193358f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_33 VNB N_A_716_21#_c_592_n 0.0447184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_716_21#_c_593_n 0.0275964f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_35 VNB N_A_716_21#_c_594_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_36 VNB N_A_716_21#_c_595_n 0.00158082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_716_21#_c_596_n 0.00424373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_716_21#_c_597_n 0.00937387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_560_47#_c_706_n 0.0201814f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_40 VNB N_A_560_47#_c_707_n 0.0433679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_560_47#_c_708_n 0.00878515f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_42 VNB N_A_560_47#_c_709_n 0.0070098f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_560_47#_c_710_n 0.011498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_560_47#_c_711_n 0.00318788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_1124_47#_c_797_n 0.00257988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1124_47#_c_798_n 0.00423483f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_47 VNB N_A_1124_47#_c_799_n 0.0242779f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_48 VNB N_A_1124_47#_c_800_n 0.0197732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_845_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Q_c_956_n 0.00206234f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_51 VNB N_Q_c_957_n 0.00567627f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_52 VNB N_Q_c_958_n 0.00226957f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_53 VNB N_Q_N_c_984_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_54 VNB N_Q_N_c_985_n 0.0230748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB Q_N 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_56 VNB N_VGND_c_1000_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1001_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1002_n 0.00639151f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_59 VNB N_VGND_c_1003_n 0.0018397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1004_n 0.00262354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1005_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1006_n 0.0269729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1007_n 0.0394538f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1008_n 0.0196078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1009_n 0.0287938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1010_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1011_n 0.359087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1012_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1013_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1014_n 0.00536381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1015_n 0.00356594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1016_n 0.00440331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VPB N_GATE_c_156_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_74 VPB N_GATE_c_157_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_75 VPB N_GATE_c_158_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_76 VPB GATE 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_77 VPB N_GATE_c_154_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_78 VPB N_A_27_47#_M1000_g 0.0387186f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_79 VPB N_A_27_47#_M1021_g 0.0302557f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_80 VPB N_A_27_47#_c_205_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_206_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_199_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_208_n 0.0214251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_209_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_210_n 0.0054554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_211_n 0.0062278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_201_n 0.0118328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_202_n 0.0465512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_D_c_340_n 0.0132141f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_90 VPB N_D_M1009_g 0.0227921f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_91 VPB N_D_c_348_n 0.0253967f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_92 VPB N_D_c_345_n 0.00184345f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_93 VPB N_A_299_47#_M1005_g 0.0394961f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_94 VPB N_A_299_47#_c_395_n 0.00712846f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_95 VPB N_A_299_47#_c_392_n 0.0100201f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_96 VPB N_A_193_47#_c_469_n 0.0271083f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_97 VPB N_A_193_47#_M1013_g 0.0205692f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_98 VPB N_A_193_47#_c_466_n 0.00733188f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_99 VPB N_A_193_47#_c_468_n 0.00228174f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_100 VPB N_A_193_47#_c_473_n 0.00289677f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_101 VPB N_A_193_47#_c_474_n 0.00832819f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_102 VPB N_A_193_47#_c_475_n 0.00237077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_193_47#_c_476_n 0.00692284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_47#_c_477_n 0.00258762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_193_47#_c_478_n 0.00824469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_716_21#_M1004_g 0.0149439f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_107 VPB N_A_716_21#_M1001_g 0.0256586f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_108 VPB N_A_716_21#_M1007_g 0.0222272f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_109 VPB N_A_716_21#_c_592_n 0.021816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_716_21#_c_593_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_111 VPB N_A_716_21#_c_603_n 0.0194583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_716_21#_c_604_n 0.0303904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_716_21#_c_605_n 0.00647507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_716_21#_c_606_n 0.0439608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_716_21#_c_607_n 0.00367821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_716_21#_c_596_n 0.00318503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_716_21#_c_597_n 8.29733e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_560_47#_M1019_g 0.0221883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_560_47#_c_707_n 0.0152272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_560_47#_c_708_n 5.55128e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_121 VPB N_A_560_47#_c_715_n 0.00664709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_560_47#_c_711_n 0.00185821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_1124_47#_M1011_g 0.0227239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_1124_47#_c_802_n 0.00398137f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_125 VPB N_A_1124_47#_c_798_n 0.00438424f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_126 VPB N_A_1124_47#_c_799_n 0.00574638f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_127 VPB N_VPWR_c_846_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_847_n 0.00348418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_848_n 0.00485902f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_130 VPB N_VPWR_c_849_n 0.00255346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_850_n 0.00289402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_851_n 0.0400902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_852_n 0.0038195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_853_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_854_n 0.0295328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_855_n 0.0203481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_856_n 0.0288571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_857_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_845_n 0.0662682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_859_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_860_n 0.00393955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_861_n 0.00421326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_862_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB Q 0.00208691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB Q 0.00833228f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_146 VPB N_Q_c_958_n 0.00474547f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_147 VPB N_Q_N_c_987_n 0.00617439f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_148 VPB N_Q_N_c_985_n 0.00721226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB Q_N 0.0341455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 N_GATE_c_151_n N_A_27_47#_M1010_g 0.0187834f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_151 N_GATE_c_155_n N_A_27_47#_M1010_g 0.0041981f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_152 N_GATE_c_158_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_153 N_GATE_c_154_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_154 N_GATE_c_151_n N_A_27_47#_c_197_n 0.00663556f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_155 N_GATE_c_152_n N_A_27_47#_c_197_n 0.0105293f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_156 N_GATE_c_152_n N_A_27_47#_c_198_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_157 GATE N_A_27_47#_c_198_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_158 N_GATE_c_154_n N_A_27_47#_c_198_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_159 N_GATE_c_157_n N_A_27_47#_c_205_n 0.0135489f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_160 N_GATE_c_158_n N_A_27_47#_c_205_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_161 N_GATE_c_157_n N_A_27_47#_c_206_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_162 N_GATE_c_158_n N_A_27_47#_c_206_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_163 GATE N_A_27_47#_c_206_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_164 N_GATE_c_154_n N_A_27_47#_c_206_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_165 N_GATE_c_154_n N_A_27_47#_c_199_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_166 N_GATE_c_152_n N_A_27_47#_c_200_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_167 GATE N_A_27_47#_c_200_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_168 N_GATE_c_155_n N_A_27_47#_c_200_n 0.0015185f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_169 N_GATE_c_156_n N_A_27_47#_c_209_n 0.0033897f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_170 N_GATE_c_158_n N_A_27_47#_c_209_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_171 GATE N_A_27_47#_c_209_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_172 N_GATE_c_156_n N_A_27_47#_c_210_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_173 N_GATE_c_158_n N_A_27_47#_c_210_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_174 GATE N_A_27_47#_c_201_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_175 N_GATE_c_154_n N_A_27_47#_c_201_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_176 N_GATE_c_157_n N_VPWR_c_846_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_177 N_GATE_c_157_n N_VPWR_c_853_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_178 N_GATE_c_157_n N_VPWR_c_845_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_179 N_GATE_c_151_n N_VGND_c_1000_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_180 N_GATE_c_151_n N_VGND_c_1005_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_181 N_GATE_c_152_n N_VGND_c_1005_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_182 N_GATE_c_151_n N_VGND_c_1011_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_208_n N_D_c_340_n 0.00166885f $X=2.495 $Y=1.53 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_201_n N_D_c_340_n 0.00398519f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1010_g N_D_c_342_n 0.00594648f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_208_n N_D_c_342_n 0.00202509f $X=2.495 $Y=1.53 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1000_g N_D_c_348_n 0.00398519f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_201_n N_D_c_344_n 0.00374568f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_208_n N_D_c_345_n 0.00994501f $X=2.495 $Y=1.53 $X2=0 $Y2=0
cc_190 N_A_27_47#_M1021_g N_A_299_47#_M1005_g 0.0362042f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_208_n N_A_299_47#_M1005_g 0.00578627f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_211_n N_A_299_47#_M1005_g 0.00249161f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_202_n N_A_299_47#_M1005_g 0.025438f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_208_n N_A_299_47#_c_395_n 5.38705e-19 $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_211_n N_A_299_47#_c_395_n 5.28447e-19 $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_208_n N_A_299_47#_c_391_n 0.00707632f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_208_n N_A_299_47#_c_392_n 0.0352966f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_255_p N_A_299_47#_c_392_n 6.56874e-19 $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_211_n N_A_299_47#_c_392_n 0.0127261f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_208_n N_A_299_47#_c_393_n 4.67313e-19 $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_202_n N_A_299_47#_c_393_n 6.94876e-19 $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_195_n N_A_193_47#_c_464_n 0.00210217f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_196_n N_A_193_47#_c_464_n 0.0137281f $X=3.215 $Y=1.175 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_211_n N_A_193_47#_c_464_n 3.34828e-19 $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_202_n N_A_193_47#_c_464_n 0.0208787f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_195_n N_A_193_47#_M1016_g 0.0129164f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1021_g N_A_193_47#_c_469_n 0.0108369f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_202_n N_A_193_47#_c_469_n 0.0205499f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1021_g N_A_193_47#_M1013_g 0.0187214f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_M1010_g N_A_193_47#_c_466_n 0.00508307f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_197_n N_A_193_47#_c_466_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_199_n N_A_193_47#_c_466_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_200_n N_A_193_47#_c_466_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_208_n N_A_193_47#_c_466_n 0.0180404f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_209_n N_A_193_47#_c_466_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_210_n N_A_193_47#_c_466_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_195_n N_A_193_47#_c_467_n 0.00255901f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_196_n N_A_193_47#_c_467_n 0.00254458f $X=3.215 $Y=1.175
+ $X2=0 $Y2=0
cc_219 N_A_27_47#_c_255_p N_A_193_47#_c_467_n 0.00140771f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_211_n N_A_193_47#_c_467_n 0.00982389f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_202_n N_A_193_47#_c_467_n 0.00618484f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_196_n N_A_193_47#_c_468_n 0.00256585f $X=3.215 $Y=1.175
+ $X2=0 $Y2=0
cc_223 N_A_27_47#_c_255_p N_A_193_47#_c_468_n 0.00114357f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_211_n N_A_193_47#_c_468_n 0.0151775f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_202_n N_A_193_47#_c_468_n 0.0186948f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_205_n N_A_193_47#_c_473_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_208_n N_A_193_47#_c_473_n 0.00195186f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_201_n N_A_193_47#_c_473_n 0.00508307f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1021_g N_A_193_47#_c_474_n 0.00615873f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_230 N_A_27_47#_c_208_n N_A_193_47#_c_474_n 0.093966f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_255_p N_A_193_47#_c_474_n 0.026178f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_211_n N_A_193_47#_c_474_n 0.00861087f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_202_n N_A_193_47#_c_474_n 0.00378075f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_M1000_g N_A_193_47#_c_475_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_205_n N_A_193_47#_c_475_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_208_n N_A_193_47#_c_475_n 0.0259095f $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_210_n N_A_193_47#_c_475_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1000_g N_A_193_47#_c_476_n 0.00508307f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1021_g N_A_193_47#_c_477_n 0.00143061f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_240 N_A_27_47#_c_202_n N_A_193_47#_c_477_n 0.00128779f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1021_g N_A_193_47#_c_478_n 0.00594922f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_242 N_A_27_47#_c_255_p N_A_193_47#_c_478_n 5.35887e-19 $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_211_n N_A_193_47#_c_478_n 0.00816604f $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_202_n N_A_193_47#_c_478_n 0.00500321f $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_195_n N_A_716_21#_M1004_g 0.0469991f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_202_n N_A_716_21#_M1004_g 8.19949e-19 $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_M1021_g N_A_560_47#_c_717_n 0.00528621f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_248 N_A_27_47#_c_211_n N_A_560_47#_c_717_n 4.9211e-19 $X=2.64 $Y=1.53 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_195_n N_A_560_47#_c_719_n 0.0115399f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_195_n N_A_560_47#_c_709_n 0.00522274f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_202_n N_A_560_47#_c_715_n 7.10824e-19 $X=2.735 $Y=1.43 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_196_n N_A_560_47#_c_710_n 0.00307428f $X=3.215 $Y=1.175
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_205_n N_VPWR_M1008_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_254 N_A_27_47#_M1000_g N_VPWR_c_846_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_205_n N_VPWR_c_846_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_206_n N_VPWR_c_846_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_209_n N_VPWR_c_846_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_258 N_A_27_47#_M1021_g N_VPWR_c_847_n 0.00427372f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_208_n N_VPWR_c_847_n 8.71018e-19 $X=2.495 $Y=1.53 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1021_g N_VPWR_c_851_n 0.00497675f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_205_n N_VPWR_c_853_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_206_n N_VPWR_c_853_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_263 N_A_27_47#_M1000_g N_VPWR_c_854_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1000_g N_VPWR_c_845_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1021_g N_VPWR_c_845_n 0.00612727f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_205_n N_VPWR_c_845_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_206_n N_VPWR_c_845_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_197_n N_VGND_M1018_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_269 N_A_27_47#_M1010_g N_VGND_c_1000_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_197_n N_VGND_c_1000_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_199_n N_VGND_c_1000_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_201_n N_VGND_c_1000_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_195_n N_VGND_c_1002_n 0.00172915f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_331_p N_VGND_c_1005_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_197_n N_VGND_c_1005_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1010_g N_VGND_c_1006_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_195_n N_VGND_c_1007_n 0.00378965f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1018_s N_VGND_c_1011_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1010_g N_VGND_c_1011_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_195_n N_VGND_c_1011_n 0.00558598f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_331_p N_VGND_c_1011_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_197_n N_VGND_c_1011_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_283 N_D_c_341_n N_A_299_47#_M1006_g 0.0161281f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_284 N_D_c_342_n N_A_299_47#_M1006_g 0.00339235f $X=1.52 $Y=0.88 $X2=0 $Y2=0
cc_285 N_D_c_340_n N_A_299_47#_M1005_g 0.00304642f $X=1.58 $Y=1.54 $X2=0 $Y2=0
cc_286 N_D_c_348_n N_A_299_47#_M1005_g 0.0209394f $X=1.84 $Y=1.615 $X2=0 $Y2=0
cc_287 N_D_M1009_g N_A_299_47#_c_395_n 0.0119836f $X=1.84 $Y=2.165 $X2=0 $Y2=0
cc_288 N_D_c_348_n N_A_299_47#_c_395_n 0.00866293f $X=1.84 $Y=1.615 $X2=0 $Y2=0
cc_289 N_D_c_341_n N_A_299_47#_c_391_n 0.00708994f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_290 N_D_c_342_n N_A_299_47#_c_391_n 0.0209069f $X=1.52 $Y=0.88 $X2=0 $Y2=0
cc_291 N_D_c_344_n N_A_299_47#_c_391_n 0.00102253f $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_c_345_n N_A_299_47#_c_391_n 0.037824f $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_293 N_D_c_340_n N_A_299_47#_c_392_n 0.00411666f $X=1.58 $Y=1.54 $X2=0 $Y2=0
cc_294 N_D_c_342_n N_A_299_47#_c_392_n 0.00180773f $X=1.52 $Y=0.88 $X2=0 $Y2=0
cc_295 N_D_c_343_n N_A_299_47#_c_392_n 3.54152e-19 $X=1.52 $Y=1.205 $X2=0 $Y2=0
cc_296 N_D_c_348_n N_A_299_47#_c_392_n 0.0131272f $X=1.84 $Y=1.615 $X2=0 $Y2=0
cc_297 N_D_c_345_n N_A_299_47#_c_392_n 0.0240586f $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_298 N_D_c_344_n N_A_299_47#_c_393_n 0.00656842f $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_299 N_D_c_345_n N_A_299_47#_c_393_n 6.7858e-19 $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_300 N_D_c_340_n N_A_193_47#_c_466_n 0.00244425f $X=1.58 $Y=1.54 $X2=0 $Y2=0
cc_301 N_D_c_341_n N_A_193_47#_c_466_n 3.74107e-19 $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_302 N_D_c_342_n N_A_193_47#_c_466_n 0.00251305f $X=1.52 $Y=0.88 $X2=0 $Y2=0
cc_303 N_D_c_344_n N_A_193_47#_c_466_n 8.19938e-19 $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_304 N_D_c_345_n N_A_193_47#_c_466_n 0.0293308f $X=1.52 $Y=1.04 $X2=0 $Y2=0
cc_305 N_D_M1009_g N_A_193_47#_c_473_n 0.00119622f $X=1.84 $Y=2.165 $X2=0 $Y2=0
cc_306 N_D_M1009_g N_A_193_47#_c_474_n 0.00297192f $X=1.84 $Y=2.165 $X2=0 $Y2=0
cc_307 N_D_M1009_g N_VPWR_c_847_n 0.00301012f $X=1.84 $Y=2.165 $X2=0 $Y2=0
cc_308 N_D_M1009_g N_VPWR_c_854_n 0.00543342f $X=1.84 $Y=2.165 $X2=0 $Y2=0
cc_309 N_D_M1009_g N_VPWR_c_845_n 0.00734866f $X=1.84 $Y=2.165 $X2=0 $Y2=0
cc_310 N_D_c_341_n N_VGND_c_1001_n 0.0110368f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_311 N_D_c_341_n N_VGND_c_1006_n 0.00336882f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_312 N_D_c_342_n N_VGND_c_1006_n 9.59663e-19 $X=1.52 $Y=0.88 $X2=0 $Y2=0
cc_313 N_D_c_341_n N_VGND_c_1011_n 0.00532348f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_314 N_D_c_342_n N_VGND_c_1011_n 0.00281935f $X=1.52 $Y=0.88 $X2=0 $Y2=0
cc_315 N_A_299_47#_M1006_g N_A_193_47#_c_464_n 0.00895289f $X=2.25 $Y=0.445
+ $X2=0 $Y2=0
cc_316 N_A_299_47#_c_391_n N_A_193_47#_c_464_n 6.80619e-19 $X=1.985 $Y=1.235
+ $X2=0 $Y2=0
cc_317 N_A_299_47#_c_393_n N_A_193_47#_c_464_n 0.00848951f $X=2.22 $Y=1.07 $X2=0
+ $Y2=0
cc_318 N_A_299_47#_M1006_g N_A_193_47#_M1016_g 0.0248806f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_319 N_A_299_47#_c_395_n N_A_193_47#_c_466_n 0.00120958f $X=1.63 $Y=1.99 $X2=0
+ $Y2=0
cc_320 N_A_299_47#_c_391_n N_A_193_47#_c_466_n 0.0259409f $X=1.985 $Y=1.235
+ $X2=0 $Y2=0
cc_321 N_A_299_47#_c_392_n N_A_193_47#_c_466_n 0.0137392f $X=1.985 $Y=1.495
+ $X2=0 $Y2=0
cc_322 N_A_299_47#_M1006_g N_A_193_47#_c_467_n 7.60915e-19 $X=2.25 $Y=0.445
+ $X2=0 $Y2=0
cc_323 N_A_299_47#_c_391_n N_A_193_47#_c_467_n 0.0186413f $X=1.985 $Y=1.235
+ $X2=0 $Y2=0
cc_324 N_A_299_47#_c_393_n N_A_193_47#_c_467_n 8.80463e-19 $X=2.22 $Y=1.07 $X2=0
+ $Y2=0
cc_325 N_A_299_47#_M1005_g N_A_193_47#_c_468_n 5.84459e-19 $X=2.26 $Y=2.165
+ $X2=0 $Y2=0
cc_326 N_A_299_47#_c_391_n N_A_193_47#_c_468_n 0.00483521f $X=1.985 $Y=1.235
+ $X2=0 $Y2=0
cc_327 N_A_299_47#_c_393_n N_A_193_47#_c_468_n 0.00212443f $X=2.22 $Y=1.07 $X2=0
+ $Y2=0
cc_328 N_A_299_47#_c_395_n N_A_193_47#_c_473_n 0.0522135f $X=1.63 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_299_47#_M1005_g N_A_193_47#_c_474_n 0.00391501f $X=2.26 $Y=2.165
+ $X2=0 $Y2=0
cc_330 N_A_299_47#_c_395_n N_A_193_47#_c_474_n 0.0225182f $X=1.63 $Y=1.99 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_c_392_n N_A_193_47#_c_474_n 0.00548892f $X=1.985 $Y=1.495
+ $X2=0 $Y2=0
cc_332 N_A_299_47#_c_395_n N_A_193_47#_c_475_n 0.00277433f $X=1.63 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_M1005_g N_A_560_47#_c_717_n 5.29815e-19 $X=2.26 $Y=2.165
+ $X2=0 $Y2=0
cc_334 N_A_299_47#_M1005_g N_VPWR_c_847_n 0.0203828f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_395_n N_VPWR_c_847_n 0.0235712f $X=1.63 $Y=1.99 $X2=0 $Y2=0
cc_336 N_A_299_47#_c_391_n N_VPWR_c_847_n 0.00165706f $X=1.985 $Y=1.235 $X2=0
+ $Y2=0
cc_337 N_A_299_47#_c_392_n N_VPWR_c_847_n 0.0100007f $X=1.985 $Y=1.495 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_393_n N_VPWR_c_847_n 2.89143e-19 $X=2.22 $Y=1.07 $X2=0
+ $Y2=0
cc_339 N_A_299_47#_M1005_g N_VPWR_c_851_n 0.00349454f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_c_395_n N_VPWR_c_854_n 0.0178472f $X=1.63 $Y=1.99 $X2=0 $Y2=0
cc_341 N_A_299_47#_M1009_s N_VPWR_c_845_n 0.00174533f $X=1.505 $Y=1.845 $X2=0
+ $Y2=0
cc_342 N_A_299_47#_M1005_g N_VPWR_c_845_n 0.00365666f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_343 N_A_299_47#_c_395_n N_VPWR_c_845_n 0.00639203f $X=1.63 $Y=1.99 $X2=0
+ $Y2=0
cc_344 N_A_299_47#_c_391_n N_VGND_M1002_d 0.0016772f $X=1.985 $Y=1.235 $X2=0
+ $Y2=0
cc_345 N_A_299_47#_M1006_g N_VGND_c_1001_n 0.0095526f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_c_391_n N_VGND_c_1001_n 0.0172492f $X=1.985 $Y=1.235 $X2=0
+ $Y2=0
cc_347 N_A_299_47#_c_393_n N_VGND_c_1001_n 2.75008e-19 $X=2.22 $Y=1.07 $X2=0
+ $Y2=0
cc_348 N_A_299_47#_c_391_n N_VGND_c_1006_n 0.0108554f $X=1.985 $Y=1.235 $X2=0
+ $Y2=0
cc_349 N_A_299_47#_M1006_g N_VGND_c_1007_n 0.0046653f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_350 N_A_299_47#_M1002_s N_VGND_c_1011_n 0.002505f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_351 N_A_299_47#_M1006_g N_VGND_c_1011_n 0.00813035f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_352 N_A_299_47#_c_391_n N_VGND_c_1011_n 0.0127569f $X=1.985 $Y=1.235 $X2=0
+ $Y2=0
cc_353 N_A_193_47#_c_468_n N_A_716_21#_M1004_g 9.32151e-19 $X=3.05 $Y=1.575
+ $X2=0 $Y2=0
cc_354 N_A_193_47#_M1013_g N_A_716_21#_M1001_g 0.0253162f $X=3.165 $Y=2.275
+ $X2=0 $Y2=0
cc_355 N_A_193_47#_c_478_n N_A_716_21#_M1001_g 2.13425e-19 $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_356 N_A_193_47#_c_469_n N_A_716_21#_c_606_n 0.0167028f $X=3.165 $Y=1.88 $X2=0
+ $Y2=0
cc_357 N_A_193_47#_c_478_n N_A_716_21#_c_606_n 4.26054e-19 $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_358 N_A_193_47#_c_469_n N_A_560_47#_c_717_n 0.00226187f $X=3.165 $Y=1.88
+ $X2=0 $Y2=0
cc_359 N_A_193_47#_M1013_g N_A_560_47#_c_717_n 0.00882514f $X=3.165 $Y=2.275
+ $X2=0 $Y2=0
cc_360 N_A_193_47#_c_474_n N_A_560_47#_c_717_n 0.00321126f $X=2.905 $Y=1.87
+ $X2=0 $Y2=0
cc_361 N_A_193_47#_c_477_n N_A_560_47#_c_717_n 0.00264142f $X=3.05 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_193_47#_c_478_n N_A_560_47#_c_717_n 0.0116912f $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_363 N_A_193_47#_c_464_n N_A_560_47#_c_719_n 5.71128e-19 $X=2.725 $Y=0.73
+ $X2=0 $Y2=0
cc_364 N_A_193_47#_c_467_n N_A_560_47#_c_719_n 0.0214775f $X=2.965 $Y=0.885
+ $X2=0 $Y2=0
cc_365 N_A_193_47#_c_467_n N_A_560_47#_c_709_n 0.0236825f $X=2.965 $Y=0.885
+ $X2=0 $Y2=0
cc_366 N_A_193_47#_M1013_g N_A_560_47#_c_732_n 0.0034713f $X=3.165 $Y=2.275
+ $X2=0 $Y2=0
cc_367 N_A_193_47#_c_469_n N_A_560_47#_c_715_n 0.00168822f $X=3.165 $Y=1.88
+ $X2=0 $Y2=0
cc_368 N_A_193_47#_M1013_g N_A_560_47#_c_715_n 0.00272415f $X=3.165 $Y=2.275
+ $X2=0 $Y2=0
cc_369 N_A_193_47#_c_468_n N_A_560_47#_c_715_n 0.0117785f $X=3.05 $Y=1.575 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_477_n N_A_560_47#_c_715_n 0.00143506f $X=3.05 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_478_n N_A_560_47#_c_715_n 0.0283386f $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_372 N_A_193_47#_c_469_n N_A_560_47#_c_710_n 0.00211754f $X=3.165 $Y=1.88
+ $X2=0 $Y2=0
cc_373 N_A_193_47#_c_467_n N_A_560_47#_c_710_n 0.00645692f $X=2.965 $Y=0.885
+ $X2=0 $Y2=0
cc_374 N_A_193_47#_c_468_n N_A_560_47#_c_710_n 0.0164566f $X=3.05 $Y=1.575 $X2=0
+ $Y2=0
cc_375 N_A_193_47#_c_474_n N_VPWR_M1009_d 6.81311e-19 $X=2.905 $Y=1.87 $X2=0
+ $Y2=0
cc_376 N_A_193_47#_c_476_n N_VPWR_c_846_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_474_n N_VPWR_c_847_n 0.0168221f $X=2.905 $Y=1.87 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_M1013_g N_VPWR_c_851_n 0.00366111f $X=3.165 $Y=2.275 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_476_n N_VPWR_c_854_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_380 N_A_193_47#_M1013_g N_VPWR_c_845_n 0.00541551f $X=3.165 $Y=2.275 $X2=0
+ $Y2=0
cc_381 N_A_193_47#_c_474_n N_VPWR_c_845_n 0.0768976f $X=2.905 $Y=1.87 $X2=0
+ $Y2=0
cc_382 N_A_193_47#_c_475_n N_VPWR_c_845_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_383 N_A_193_47#_c_476_n N_VPWR_c_845_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_c_477_n N_VPWR_c_845_n 0.0147476f $X=3.05 $Y=1.87 $X2=0 $Y2=0
cc_385 N_A_193_47#_c_474_n A_467_369# 0.00398287f $X=2.905 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_386 N_A_193_47#_M1016_g N_VGND_c_1001_n 0.00184148f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_387 N_A_193_47#_c_466_n N_VGND_c_1006_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_c_464_n N_VGND_c_1007_n 5.15715e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_389 N_A_193_47#_M1016_g N_VGND_c_1007_n 0.00435108f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_390 N_A_193_47#_c_467_n N_VGND_c_1007_n 0.00337743f $X=2.965 $Y=0.885 $X2=0
+ $Y2=0
cc_391 N_A_193_47#_M1010_d N_VGND_c_1011_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_392 N_A_193_47#_c_464_n N_VGND_c_1011_n 3.58005e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_393 N_A_193_47#_M1016_g N_VGND_c_1011_n 0.00632668f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_394 N_A_193_47#_c_466_n N_VGND_c_1011_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_395 N_A_193_47#_c_467_n N_VGND_c_1011_n 0.0056644f $X=2.965 $Y=0.885 $X2=0
+ $Y2=0
cc_396 N_A_716_21#_c_591_n N_A_560_47#_c_706_n 0.0226161f $X=5.015 $Y=0.995
+ $X2=0 $Y2=0
cc_397 N_A_716_21#_c_595_n N_A_560_47#_c_706_n 0.00838476f $X=4.447 $Y=0.995
+ $X2=0 $Y2=0
cc_398 N_A_716_21#_c_619_p N_A_560_47#_c_706_n 0.0041185f $X=4.385 $Y=0.58 $X2=0
+ $Y2=0
cc_399 N_A_716_21#_M1007_g N_A_560_47#_M1019_g 0.0248218f $X=5.015 $Y=1.985
+ $X2=0 $Y2=0
cc_400 N_A_716_21#_c_606_n N_A_560_47#_M1019_g 0.00365118f $X=3.905 $Y=1.7 $X2=0
+ $Y2=0
cc_401 N_A_716_21#_c_607_n N_A_560_47#_M1019_g 0.00751288f $X=4.43 $Y=1.535
+ $X2=0 $Y2=0
cc_402 N_A_716_21#_M1004_g N_A_560_47#_c_707_n 0.0196777f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_716_21#_c_605_n N_A_560_47#_c_707_n 0.00753869f $X=4.285 $Y=1.7 $X2=0
+ $Y2=0
cc_404 N_A_716_21#_c_606_n N_A_560_47#_c_707_n 0.00517995f $X=3.905 $Y=1.7 $X2=0
+ $Y2=0
cc_405 N_A_716_21#_c_619_p N_A_560_47#_c_707_n 0.00219273f $X=4.385 $Y=0.58
+ $X2=0 $Y2=0
cc_406 N_A_716_21#_c_627_p N_A_560_47#_c_707_n 0.00255404f $X=4.385 $Y=1.755
+ $X2=0 $Y2=0
cc_407 N_A_716_21#_c_628_p N_A_560_47#_c_707_n 0.0181886f $X=4.447 $Y=1.16 $X2=0
+ $Y2=0
cc_408 N_A_716_21#_c_596_n N_A_560_47#_c_708_n 0.018719f $X=5.065 $Y=1.16 $X2=0
+ $Y2=0
cc_409 N_A_716_21#_c_597_n N_A_560_47#_c_708_n 0.0166057f $X=5.065 $Y=1.16 $X2=0
+ $Y2=0
cc_410 N_A_716_21#_c_628_p N_A_560_47#_c_708_n 0.00248969f $X=4.447 $Y=1.16
+ $X2=0 $Y2=0
cc_411 N_A_716_21#_M1001_g N_A_560_47#_c_717_n 0.0045197f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_412 N_A_716_21#_M1004_g N_A_560_47#_c_719_n 0.00159662f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_413 N_A_716_21#_M1004_g N_A_560_47#_c_709_n 0.0103959f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_414 N_A_716_21#_M1001_g N_A_560_47#_c_732_n 0.00423932f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_415 N_A_716_21#_c_636_p N_A_560_47#_c_732_n 0.00205148f $X=4.385 $Y=2.27
+ $X2=0 $Y2=0
cc_416 N_A_716_21#_M1004_g N_A_560_47#_c_715_n 0.0117131f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_716_21#_M1001_g N_A_560_47#_c_715_n 0.00823168f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_418 N_A_716_21#_c_605_n N_A_560_47#_c_715_n 0.0252243f $X=4.285 $Y=1.7 $X2=0
+ $Y2=0
cc_419 N_A_716_21#_c_606_n N_A_560_47#_c_715_n 0.00913418f $X=3.905 $Y=1.7 $X2=0
+ $Y2=0
cc_420 N_A_716_21#_c_636_p N_A_560_47#_c_715_n 0.00574382f $X=4.385 $Y=2.27
+ $X2=0 $Y2=0
cc_421 N_A_716_21#_M1004_g N_A_560_47#_c_710_n 0.00864866f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_422 N_A_716_21#_M1004_g N_A_560_47#_c_711_n 0.0124531f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_423 N_A_716_21#_c_605_n N_A_560_47#_c_711_n 0.0236312f $X=4.285 $Y=1.7 $X2=0
+ $Y2=0
cc_424 N_A_716_21#_c_606_n N_A_560_47#_c_711_n 0.00678362f $X=3.905 $Y=1.7 $X2=0
+ $Y2=0
cc_425 N_A_716_21#_c_628_p N_A_560_47#_c_711_n 0.0278171f $X=4.447 $Y=1.16 $X2=0
+ $Y2=0
cc_426 N_A_716_21#_c_603_n N_A_1124_47#_M1011_g 0.00909592f $X=5.94 $Y=1.62
+ $X2=0 $Y2=0
cc_427 N_A_716_21#_c_604_n N_A_1124_47#_M1011_g 0.0122907f $X=5.94 $Y=1.77 $X2=0
+ $Y2=0
cc_428 N_A_716_21#_c_591_n N_A_1124_47#_c_797_n 0.00141284f $X=5.015 $Y=0.995
+ $X2=0 $Y2=0
cc_429 N_A_716_21#_c_593_n N_A_1124_47#_c_797_n 0.0112708f $X=5.925 $Y=1.325
+ $X2=0 $Y2=0
cc_430 N_A_716_21#_c_594_n N_A_1124_47#_c_797_n 0.00951761f $X=5.955 $Y=0.73
+ $X2=0 $Y2=0
cc_431 N_A_716_21#_M1007_g N_A_1124_47#_c_802_n 0.00165518f $X=5.015 $Y=1.985
+ $X2=0 $Y2=0
cc_432 N_A_716_21#_c_603_n N_A_1124_47#_c_802_n 0.0117262f $X=5.94 $Y=1.62 $X2=0
+ $Y2=0
cc_433 N_A_716_21#_c_604_n N_A_1124_47#_c_802_n 0.0208659f $X=5.94 $Y=1.77 $X2=0
+ $Y2=0
cc_434 N_A_716_21#_c_593_n N_A_1124_47#_c_798_n 0.0156725f $X=5.925 $Y=1.325
+ $X2=0 $Y2=0
cc_435 N_A_716_21#_c_604_n N_A_1124_47#_c_798_n 0.00116449f $X=5.94 $Y=1.77
+ $X2=0 $Y2=0
cc_436 N_A_716_21#_c_593_n N_A_1124_47#_c_799_n 0.0215069f $X=5.925 $Y=1.325
+ $X2=0 $Y2=0
cc_437 N_A_716_21#_c_592_n N_A_1124_47#_c_816_n 0.0155499f $X=5.85 $Y=1.16 $X2=0
+ $Y2=0
cc_438 N_A_716_21#_c_593_n N_A_1124_47#_c_816_n 0.00186446f $X=5.925 $Y=1.325
+ $X2=0 $Y2=0
cc_439 N_A_716_21#_c_593_n N_A_1124_47#_c_800_n 0.00357247f $X=5.925 $Y=1.325
+ $X2=0 $Y2=0
cc_440 N_A_716_21#_c_594_n N_A_1124_47#_c_800_n 0.0157829f $X=5.955 $Y=0.73
+ $X2=0 $Y2=0
cc_441 N_A_716_21#_M1001_g N_VPWR_c_848_n 0.00443168f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_442 N_A_716_21#_c_605_n N_VPWR_c_848_n 0.00755153f $X=4.285 $Y=1.7 $X2=0
+ $Y2=0
cc_443 N_A_716_21#_c_606_n N_VPWR_c_848_n 0.00474199f $X=3.905 $Y=1.7 $X2=0
+ $Y2=0
cc_444 N_A_716_21#_c_636_p N_VPWR_c_848_n 0.0127245f $X=4.385 $Y=2.27 $X2=0
+ $Y2=0
cc_445 N_A_716_21#_M1007_g N_VPWR_c_849_n 0.0198221f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_446 N_A_716_21#_c_596_n N_VPWR_c_849_n 0.0152127f $X=5.065 $Y=1.16 $X2=0
+ $Y2=0
cc_447 N_A_716_21#_c_604_n N_VPWR_c_850_n 0.00537515f $X=5.94 $Y=1.77 $X2=0
+ $Y2=0
cc_448 N_A_716_21#_M1001_g N_VPWR_c_851_n 0.00498998f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_449 N_A_716_21#_c_636_p N_VPWR_c_855_n 0.0119709f $X=4.385 $Y=2.27 $X2=0
+ $Y2=0
cc_450 N_A_716_21#_M1007_g N_VPWR_c_856_n 0.0046653f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_451 N_A_716_21#_c_604_n N_VPWR_c_856_n 0.00541359f $X=5.94 $Y=1.77 $X2=0
+ $Y2=0
cc_452 N_A_716_21#_M1019_s N_VPWR_c_845_n 0.00248707f $X=4.26 $Y=1.485 $X2=0
+ $Y2=0
cc_453 N_A_716_21#_M1001_g N_VPWR_c_845_n 0.00971782f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_454 N_A_716_21#_M1007_g N_VPWR_c_845_n 0.00921786f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_716_21#_c_604_n N_VPWR_c_845_n 0.0110992f $X=5.94 $Y=1.77 $X2=0 $Y2=0
cc_456 N_A_716_21#_c_605_n N_VPWR_c_845_n 0.0113987f $X=4.285 $Y=1.7 $X2=0 $Y2=0
cc_457 N_A_716_21#_c_606_n N_VPWR_c_845_n 0.00246751f $X=3.905 $Y=1.7 $X2=0
+ $Y2=0
cc_458 N_A_716_21#_c_636_p N_VPWR_c_845_n 0.0086523f $X=4.385 $Y=2.27 $X2=0
+ $Y2=0
cc_459 N_A_716_21#_c_592_n N_Q_c_956_n 0.00600702f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_460 N_A_716_21#_c_593_n N_Q_c_956_n 0.00127001f $X=5.925 $Y=1.325 $X2=0 $Y2=0
cc_461 N_A_716_21#_c_596_n N_Q_c_956_n 4.59641e-19 $X=5.065 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_716_21#_c_592_n Q 0.0051645f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_463 N_A_716_21#_c_604_n Q 0.00304572f $X=5.94 $Y=1.77 $X2=0 $Y2=0
cc_464 N_A_716_21#_c_596_n Q 2.71773e-19 $X=5.065 $Y=1.16 $X2=0 $Y2=0
cc_465 N_A_716_21#_c_594_n N_Q_c_957_n 0.00119211f $X=5.955 $Y=0.73 $X2=0 $Y2=0
cc_466 N_A_716_21#_c_591_n N_Q_c_958_n 0.00399642f $X=5.015 $Y=0.995 $X2=0 $Y2=0
cc_467 N_A_716_21#_M1007_g N_Q_c_958_n 0.00882731f $X=5.015 $Y=1.985 $X2=0 $Y2=0
cc_468 N_A_716_21#_c_592_n N_Q_c_958_n 0.0223494f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_716_21#_c_603_n N_Q_c_958_n 0.0010384f $X=5.94 $Y=1.62 $X2=0 $Y2=0
cc_470 N_A_716_21#_c_596_n N_Q_c_958_n 0.0249855f $X=5.065 $Y=1.16 $X2=0 $Y2=0
cc_471 N_A_716_21#_M1004_g N_VGND_c_1002_n 0.0115017f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_472 N_A_716_21#_c_619_p N_VGND_c_1002_n 0.00725053f $X=4.385 $Y=0.58 $X2=0
+ $Y2=0
cc_473 N_A_716_21#_c_591_n N_VGND_c_1003_n 0.0119032f $X=5.015 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_716_21#_c_596_n N_VGND_c_1003_n 0.0127851f $X=5.065 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_716_21#_c_594_n N_VGND_c_1004_n 0.00420958f $X=5.955 $Y=0.73 $X2=0
+ $Y2=0
cc_476 N_A_716_21#_M1004_g N_VGND_c_1007_n 0.0046653f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_477 N_A_716_21#_c_619_p N_VGND_c_1008_n 0.00795251f $X=4.385 $Y=0.58 $X2=0
+ $Y2=0
cc_478 N_A_716_21#_c_591_n N_VGND_c_1009_n 0.0046653f $X=5.015 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_A_716_21#_c_594_n N_VGND_c_1009_n 0.00541359f $X=5.955 $Y=0.73 $X2=0
+ $Y2=0
cc_480 N_A_716_21#_M1020_s N_VGND_c_1011_n 0.00321007f $X=4.26 $Y=0.235 $X2=0
+ $Y2=0
cc_481 N_A_716_21#_M1004_g N_VGND_c_1011_n 0.00813035f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_482 N_A_716_21#_c_591_n N_VGND_c_1011_n 0.00921786f $X=5.015 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_716_21#_c_594_n N_VGND_c_1011_n 0.0110992f $X=5.955 $Y=0.73 $X2=0
+ $Y2=0
cc_484 N_A_716_21#_c_619_p N_VGND_c_1011_n 0.00902972f $X=4.385 $Y=0.58 $X2=0
+ $Y2=0
cc_485 N_A_560_47#_c_717_n N_VPWR_c_847_n 0.00543374f $X=3.425 $Y=2.34 $X2=0
+ $Y2=0
cc_486 N_A_560_47#_M1019_g N_VPWR_c_848_n 0.00316529f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_487 N_A_560_47#_M1019_g N_VPWR_c_849_n 0.00396306f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_A_560_47#_c_717_n N_VPWR_c_851_n 0.0386273f $X=3.425 $Y=2.34 $X2=0
+ $Y2=0
cc_489 N_A_560_47#_c_715_n N_VPWR_c_851_n 6.98957e-19 $X=3.555 $Y=1.995 $X2=0
+ $Y2=0
cc_490 N_A_560_47#_M1019_g N_VPWR_c_855_n 0.00585385f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_A_560_47#_M1021_d N_VPWR_c_845_n 0.00180969f $X=2.81 $Y=2.065 $X2=0
+ $Y2=0
cc_492 N_A_560_47#_M1019_g N_VPWR_c_845_n 0.0119294f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_560_47#_c_717_n N_VPWR_c_845_n 0.0217052f $X=3.425 $Y=2.34 $X2=0
+ $Y2=0
cc_494 N_A_560_47#_c_715_n N_VPWR_c_845_n 9.85588e-19 $X=3.555 $Y=1.995 $X2=0
+ $Y2=0
cc_495 N_A_560_47#_c_717_n A_648_413# 0.0054034f $X=3.425 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_496 N_A_560_47#_c_732_n A_648_413# 0.00192965f $X=3.517 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_497 N_A_560_47#_c_715_n A_648_413# 2.998e-19 $X=3.555 $Y=1.995 $X2=-0.19
+ $Y2=-0.24
cc_498 N_A_560_47#_c_719_n N_VGND_c_1001_n 0.00258705f $X=3.305 $Y=0.45 $X2=0
+ $Y2=0
cc_499 N_A_560_47#_c_706_n N_VGND_c_1002_n 0.00410674f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_500 N_A_560_47#_c_707_n N_VGND_c_1002_n 0.00169847f $X=4.52 $Y=1.16 $X2=0
+ $Y2=0
cc_501 N_A_560_47#_c_719_n N_VGND_c_1002_n 0.011006f $X=3.305 $Y=0.45 $X2=0
+ $Y2=0
cc_502 N_A_560_47#_c_711_n N_VGND_c_1002_n 0.012642f $X=4.09 $Y=1.16 $X2=0 $Y2=0
cc_503 N_A_560_47#_c_706_n N_VGND_c_1003_n 0.0020107f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_560_47#_c_719_n N_VGND_c_1007_n 0.0228254f $X=3.305 $Y=0.45 $X2=0
+ $Y2=0
cc_505 N_A_560_47#_c_706_n N_VGND_c_1008_n 0.00547395f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_560_47#_M1016_d N_VGND_c_1011_n 0.00259228f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_507 N_A_560_47#_c_706_n N_VGND_c_1011_n 0.0110501f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_508 N_A_560_47#_c_719_n N_VGND_c_1011_n 0.0229382f $X=3.305 $Y=0.45 $X2=0
+ $Y2=0
cc_509 N_A_560_47#_c_719_n A_651_47# 0.00393298f $X=3.305 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_510 N_A_560_47#_c_709_n A_651_47# 0.00158748f $X=3.39 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_511 N_A_1124_47#_M1011_g N_VPWR_c_850_n 0.0132029f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_A_1124_47#_c_802_n N_VPWR_c_850_n 0.0454653f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_513 N_A_1124_47#_c_798_n N_VPWR_c_850_n 0.00959603f $X=6.345 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_A_1124_47#_c_799_n N_VPWR_c_850_n 0.00244466f $X=6.345 $Y=1.16 $X2=0
+ $Y2=0
cc_515 N_A_1124_47#_c_802_n N_VPWR_c_856_n 0.0153916f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_516 N_A_1124_47#_M1011_g N_VPWR_c_857_n 0.0046653f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_517 N_A_1124_47#_M1014_s N_VPWR_c_845_n 0.00352456f $X=5.62 $Y=1.845 $X2=0
+ $Y2=0
cc_518 N_A_1124_47#_M1011_g N_VPWR_c_845_n 0.00895857f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_519 N_A_1124_47#_c_802_n N_VPWR_c_845_n 0.00941829f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_520 N_A_1124_47#_c_797_n N_Q_c_957_n 0.0595964f $X=5.745 $Y=0.51 $X2=0 $Y2=0
cc_521 N_A_1124_47#_c_802_n N_Q_c_958_n 0.0905032f $X=5.745 $Y=2.165 $X2=0 $Y2=0
cc_522 N_A_1124_47#_c_816_n N_Q_c_958_n 0.0251378f $X=5.785 $Y=1.16 $X2=0 $Y2=0
cc_523 N_A_1124_47#_M1011_g N_Q_N_c_987_n 0.00595806f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_524 N_A_1124_47#_c_802_n N_Q_N_c_987_n 0.00519826f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_525 N_A_1124_47#_c_798_n N_Q_N_c_985_n 0.0266603f $X=6.345 $Y=1.16 $X2=0
+ $Y2=0
cc_526 N_A_1124_47#_c_800_n N_Q_N_c_985_n 0.0189779f $X=6.357 $Y=0.995 $X2=0
+ $Y2=0
cc_527 N_A_1124_47#_c_797_n N_VGND_c_1004_n 0.0209216f $X=5.745 $Y=0.51 $X2=0
+ $Y2=0
cc_528 N_A_1124_47#_c_798_n N_VGND_c_1004_n 0.0104995f $X=6.345 $Y=1.16 $X2=0
+ $Y2=0
cc_529 N_A_1124_47#_c_799_n N_VGND_c_1004_n 0.00255976f $X=6.345 $Y=1.16 $X2=0
+ $Y2=0
cc_530 N_A_1124_47#_c_800_n N_VGND_c_1004_n 0.00941229f $X=6.357 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_1124_47#_c_797_n N_VGND_c_1009_n 0.0153916f $X=5.745 $Y=0.51 $X2=0
+ $Y2=0
cc_532 N_A_1124_47#_c_800_n N_VGND_c_1010_n 0.0046653f $X=6.357 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_A_1124_47#_M1003_s N_VGND_c_1011_n 0.00352456f $X=5.62 $Y=0.235 $X2=0
+ $Y2=0
cc_534 N_A_1124_47#_c_797_n N_VGND_c_1011_n 0.00941829f $X=5.745 $Y=0.51 $X2=0
+ $Y2=0
cc_535 N_A_1124_47#_c_800_n N_VGND_c_1011_n 0.00895857f $X=6.357 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_845_n A_467_369# 0.00469785f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_537 N_VPWR_c_845_n A_648_413# 0.00276026f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_538 N_VPWR_c_845_n N_Q_M1007_d 0.00383158f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_c_856_n Q 0.0229891f $X=6.09 $Y=2.72 $X2=0 $Y2=0
cc_540 N_VPWR_c_845_n Q 0.0133387f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_541 N_VPWR_c_849_n N_Q_c_958_n 0.0020953f $X=4.805 $Y=1.735 $X2=0 $Y2=0
cc_542 N_VPWR_c_845_n N_Q_N_M1011_d 0.00387172f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_543 N_VPWR_c_857_n Q_N 0.018001f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_544 N_VPWR_c_845_n Q_N 0.00993603f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_545 N_Q_c_957_n N_VGND_c_1009_n 0.0242903f $X=5.225 $Y=0.42 $X2=0 $Y2=0
cc_546 N_Q_M1017_d N_VGND_c_1011_n 0.00382897f $X=5.09 $Y=0.235 $X2=0 $Y2=0
cc_547 N_Q_c_957_n N_VGND_c_1011_n 0.013369f $X=5.225 $Y=0.42 $X2=0 $Y2=0
cc_548 Q_N N_VGND_c_1010_n 0.0179668f $X=6.595 $Y=0.425 $X2=0 $Y2=0
cc_549 N_Q_N_M1015_d N_VGND_c_1011_n 0.00387172f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_550 Q_N N_VGND_c_1011_n 0.00992828f $X=6.595 $Y=0.425 $X2=0 $Y2=0
cc_551 N_VGND_c_1011_n A_465_47# 0.0114412f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_552 N_VGND_c_1011_n A_651_47# 0.00635689f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__nand4_2.spice.pex
* Created: Thu Aug 27 14:30:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4_2%D 3 7 9 11 15 17 18
c47 18 0 1.6164e-19 $X=0.695 $Y=1.19
c48 11 0 8.56806e-20 $X=0.89 $Y=0.56
r49 21 23 36.15 $w=2.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.68
+ $Y2=1.16
r50 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.68
+ $Y=1.16 $X2=0.68 $Y2=1.16
r51 17 18 24.6773 $w=1.98e-07 $l=4.45e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.68 $Y2=1.175
r52 9 23 36.15 $w=2.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=0.68
+ $Y2=1.16
r53 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r54 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r55 5 21 17.3521 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r56 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r57 1 21 17.3521 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r58 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%C 3 7 11 15 17 18 26
c48 26 0 1.6164e-19 $X=1.73 $Y=1.16
c49 3 0 1.79953e-19 $X=1.31 $Y=0.56
r50 24 26 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.73 $Y2=1.16
r51 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r52 21 24 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r53 18 25 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.52 $Y2=1.175
r54 17 25 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.52 $Y2=1.175
r55 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r56 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r57 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r58 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r59 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r60 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295 $X2=1.31
+ $Y2=1.985
r61 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r62 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%B 3 7 11 15 17 18 28
c48 18 0 1.78369e-19 $X=2.995 $Y=1.19
r49 26 28 53.3217 $w=2.7e-07 $l=2.4e-07 $layer=POLY_cond $X=2.89 $Y=1.16
+ $X2=3.13 $Y2=1.16
r50 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.89
+ $Y=1.16 $X2=2.89 $Y2=1.16
r51 24 26 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=2.89 $Y2=1.16
r52 23 24 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=2.71 $Y=1.16 $X2=2.73
+ $Y2=1.16
r53 21 23 88.8695 $w=2.7e-07 $l=4e-07 $layer=POLY_cond $X=2.31 $Y=1.16 $X2=2.71
+ $Y2=1.16
r54 18 27 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=2.89 $Y2=1.175
r55 17 27 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.89 $Y2=1.175
r56 13 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.13 $Y=1.025
+ $X2=3.13 $Y2=1.16
r57 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.13 $Y=1.025
+ $X2=3.13 $Y2=0.56
r58 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.73 $Y=1.295
+ $X2=2.73 $Y2=1.16
r59 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.73 $Y=1.295
+ $X2=2.73 $Y2=1.985
r60 5 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.71 $Y=1.025
+ $X2=2.71 $Y2=1.16
r61 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.71 $Y=1.025
+ $X2=2.71 $Y2=0.56
r62 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.31 $Y=1.295
+ $X2=2.31 $Y2=1.16
r63 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.31 $Y=1.295 $X2=2.31
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%A 3 7 11 15 17 20 23
c40 17 0 1.78369e-19 $X=4.045 $Y=1.16
c41 3 0 1.27323e-19 $X=3.55 $Y=0.56
r42 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.33
+ $Y=1.16 $X2=4.33 $Y2=1.16
r43 17 23 58.9526 $w=2.9e-07 $l=2.85e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=4.33 $Y2=1.16
r44 17 19 12.6442 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=3.97 $Y2=1.16
r45 13 19 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.97 $Y=1.305
+ $X2=3.97 $Y2=1.16
r46 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.97 $Y=1.305
+ $X2=3.97 $Y2=1.985
r47 9 19 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.97 $Y=1.015
+ $X2=3.97 $Y2=1.16
r48 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.97 $Y=1.015
+ $X2=3.97 $Y2=0.56
r49 1 19 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=3.55 $Y=1.16
+ $X2=3.97 $Y2=1.16
r50 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.55 $Y=1.295 $X2=3.55
+ $Y2=1.985
r51 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.55 $Y=1.025
+ $X2=3.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%VPWR 1 2 3 4 5 16 18 24 28 32 34 36 41 42 44
+ 45 46 52 60 68 72
r68 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r69 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r70 63 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r71 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 60 71 4.61575 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=4.347 $Y2=2.72
r73 60 62 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 59 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 56 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=2.72
+ $X2=2.02 $Y2=2.72
r78 56 58 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.185 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 55 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 52 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=2.02 $Y2=2.72
r82 52 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r83 51 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r84 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r85 48 65 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r86 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r87 46 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 46 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 44 58 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r90 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.16 $Y2=2.72
r91 43 62 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.91 $Y2=2.72
r92 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.16 $Y2=2.72
r93 41 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72 $X2=1.1
+ $Y2=2.72
r95 40 54 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r96 40 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72 $X2=1.1
+ $Y2=2.72
r97 36 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.26 $Y=1.66
+ $X2=4.26 $Y2=2.34
r98 34 71 3.15043 $w=3.3e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.26 $Y=2.635
+ $X2=4.347 $Y2=2.72
r99 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.26 $Y=2.635
+ $X2=4.26 $Y2=2.34
r100 30 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=2.635
+ $X2=3.16 $Y2=2.72
r101 30 32 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.16 $Y=2.635
+ $X2=3.16 $Y2=2
r102 26 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=2.635
+ $X2=2.02 $Y2=2.72
r103 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.02 $Y=2.635
+ $X2=2.02 $Y2=2
r104 22 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r105 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r106 18 21 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r107 16 65 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r108 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r109 5 39 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.485 $X2=4.26 $Y2=2.34
r110 5 36 400 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.485 $X2=4.26 $Y2=1.66
r111 4 32 300 $w=1.7e-07 $l=6.69365e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=3.16 $Y2=2
r112 3 28 300 $w=1.7e-07 $l=6.13148e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=2.02 $Y2=2
r113 2 24 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r114 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r115 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%Y 1 2 3 4 5 16 18 20 24 26 30 34 38 43 44 45
+ 46 47
c86 47 0 1.57533e-19 $X=3.455 $Y=1.53
r87 68 69 2.05776 $w=5.53e-07 $l=5e-09 $layer=LI1_cond $X=3.647 $Y=1.66
+ $X2=3.647 $Y2=1.665
r88 47 68 2.26285 $w=5.53e-07 $l=1.05e-07 $layer=LI1_cond $X=3.647 $Y=1.555
+ $X2=3.647 $Y2=1.66
r89 46 47 7.32733 $w=5.53e-07 $l=3.4e-07 $layer=LI1_cond $X=3.647 $Y=1.19
+ $X2=3.647 $Y2=1.53
r90 46 62 4.85939 $w=5.53e-07 $l=1.35e-07 $layer=LI1_cond $X=3.647 $Y=1.19
+ $X2=3.647 $Y2=1.055
r91 45 47 13.253 $w=3.88e-07 $l=3.75e-07 $layer=LI1_cond $X=2.995 $Y=1.555
+ $X2=3.37 $Y2=1.555
r92 45 54 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=2.995 $Y=1.555
+ $X2=2.685 $Y2=1.555
r93 44 54 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.52 $Y=1.555
+ $X2=2.685 $Y2=1.555
r94 38 69 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.76 $Y=2.34
+ $X2=3.76 $Y2=1.665
r95 34 62 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.76 $Y=0.72
+ $X2=3.76 $Y2=1.055
r96 28 44 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.52 $Y=1.665
+ $X2=2.52 $Y2=1.555
r97 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.52 $Y=1.665
+ $X2=2.52 $Y2=2.34
r98 27 43 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.555
+ $X2=1.52 $Y2=1.555
r99 26 44 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=1.555
+ $X2=2.52 $Y2=1.555
r100 26 27 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.355 $Y=1.555
+ $X2=1.685 $Y2=1.555
r101 22 43 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.555
r102 22 24 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r103 21 41 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.555
+ $X2=0.68 $Y2=1.555
r104 20 43 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=1.52 $Y2=1.555
r105 20 21 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=0.845 $Y2=1.555
r106 16 41 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.555
r107 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r108 5 68 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.485 $X2=3.76 $Y2=1.66
r109 5 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.485 $X2=3.76 $Y2=2.34
r110 4 44 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.485 $X2=2.52 $Y2=1.66
r111 4 30 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.485 $X2=2.52 $Y2=2.34
r112 3 43 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r113 3 24 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r114 2 41 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r115 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r116 1 34 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.76 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%A_27_47# 1 2 3 12 14 15 16 19 22
c41 14 0 1.79953e-19 $X=0.935 $Y=0.82
r42 20 25 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.185 $Y=0.36
+ $X2=1.06 $Y2=0.36
r43 20 22 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=1.185 $Y=0.36
+ $X2=1.96 $Y2=0.36
r44 17 19 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.06 $Y=0.735
+ $X2=1.06 $Y2=0.72
r45 16 25 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.06 $Y=0.465
+ $X2=1.06 $Y2=0.36
r46 16 19 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.06 $Y=0.465
+ $X2=1.06 $Y2=0.72
r47 14 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=1.06 $Y2=0.735
r48 14 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=0.425 $Y2=0.82
r49 10 15 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r50 10 12 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.38
r51 3 22 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.96 $Y2=0.38
r52 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r53 2 19 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.72
r54 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%VGND 1 6 8 10 17 18 21
r53 21 22 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r54 18 22 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=0.69
+ $Y2=0
r55 17 18 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r56 15 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r57 15 17 235.193 $w=1.68e-07 $l=3.605e-06 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=4.37 $Y2=0
r58 10 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r59 10 12 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r60 8 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 4 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r63 4 6 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0.38
r64 1 6 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%A_277_47# 1 2 11
c22 11 0 3.70537e-19 $X=2.92 $Y=0.72
r23 8 11 59.7563 $w=2.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.52 $Y=0.77 $X2=2.92
+ $Y2=0.77
r24 2 11 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.235 $X2=2.92 $Y2=0.72
r25 1 8 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_2%A_471_47# 1 2 3 10 16 18 20 22 25
r34 20 27 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=4.26 $Y=0.465
+ $X2=4.26 $Y2=0.36
r35 20 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.26 $Y=0.465
+ $X2=4.26 $Y2=0.72
r36 19 25 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=0.36 $X2=3.34
+ $Y2=0.36
r37 18 27 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0.36
+ $X2=4.26 $Y2=0.36
r38 18 19 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=4.095 $Y=0.36
+ $X2=3.425 $Y2=0.36
r39 14 25 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.34 $Y=0.465
+ $X2=3.34 $Y2=0.36
r40 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.34 $Y=0.465
+ $X2=3.34 $Y2=0.72
r41 10 25 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.255 $Y=0.36 $X2=3.34
+ $Y2=0.36
r42 10 12 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=3.255 $Y=0.36
+ $X2=2.48 $Y2=0.36
r43 3 27 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=4.045
+ $Y=0.235 $X2=4.26 $Y2=0.38
r44 3 22 182 $w=1.7e-07 $l=5.82666e-07 $layer=licon1_NDIFF $count=1 $X=4.045
+ $Y=0.235 $X2=4.26 $Y2=0.72
r45 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.34 $Y2=0.38
r46 2 16 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.34 $Y2=0.72
r47 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.48 $Y2=0.38
.ends


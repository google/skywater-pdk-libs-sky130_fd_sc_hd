* File: sky130_fd_sc_hd__clkinv_2.pxi.spice
* Created: Thu Aug 27 14:12:35 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINV_2%A N_A_M1000_g N_A_M1001_g N_A_M1002_g N_A_c_39_n
+ N_A_M1003_g N_A_M1004_g A A A PM_SKY130_FD_SC_HD__CLKINV_2%A
x_PM_SKY130_FD_SC_HD__CLKINV_2%Y N_Y_M1002_d N_Y_M1000_s N_Y_M1001_s N_Y_c_122_p
+ N_Y_c_91_n N_Y_c_92_n N_Y_c_123_p N_Y_c_86_n N_Y_c_87_n N_Y_c_88_n N_Y_c_93_n
+ N_Y_c_94_n Y Y Y N_Y_c_90_n N_Y_c_96_n PM_SKY130_FD_SC_HD__CLKINV_2%Y
x_PM_SKY130_FD_SC_HD__CLKINV_2%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_c_137_n
+ N_VPWR_c_138_n N_VPWR_c_139_n VPWR N_VPWR_c_140_n N_VPWR_c_141_n
+ N_VPWR_c_142_n N_VPWR_c_136_n PM_SKY130_FD_SC_HD__CLKINV_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKINV_2%VGND N_VGND_M1002_s N_VGND_M1004_s N_VGND_c_163_n
+ N_VGND_c_164_n N_VGND_c_165_n VGND N_VGND_c_166_n N_VGND_c_167_n
+ N_VGND_c_168_n N_VGND_c_169_n PM_SKY130_FD_SC_HD__CLKINV_2%VGND
cc_1 VNB N_A_M1001_g 4.57292e-19 $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_2 VNB N_A_M1002_g 0.0421156f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.445
cc_3 VNB N_A_c_39_n 0.0934495f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.295
cc_4 VNB N_A_M1003_g 4.91581e-19 $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.985
cc_5 VNB N_A_M1004_g 0.0349086f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=0.445
cc_6 VNB A 0.0140604f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_7 VNB N_Y_c_86_n 0.00149799f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_8 VNB N_Y_c_87_n 0.00167495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_Y_c_88_n 0.00410962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB Y 0.0210583f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_11 VNB N_Y_c_90_n 0.0101921f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.16
cc_12 VNB N_VPWR_c_136_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_13 VNB N_VGND_c_163_n 0.0193788f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.015
cc_14 VNB N_VGND_c_164_n 0.0101596f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.445
cc_15 VNB N_VGND_c_165_n 0.0154987f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.295
cc_16 VNB N_VGND_c_166_n 0.0199636f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.025
cc_17 VNB N_VGND_c_167_n 0.0142308f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_18 VNB N_VGND_c_168_n 0.00564902f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_19 VNB N_VGND_c_169_n 0.141662f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_20 VPB N_A_M1000_g 0.0271137f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_21 VPB N_A_M1001_g 0.0195484f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_22 VPB N_A_c_39_n 0.00626485f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.295
cc_23 VPB N_A_M1003_g 0.0231397f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_24 VPB N_Y_c_91_n 0.00238943f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_25 VPB N_Y_c_92_n 0.00852947f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_26 VPB N_Y_c_93_n 6.00816e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_Y_c_94_n 0.0021151f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_28 VPB Y 0.00792875f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_29 VPB N_Y_c_96_n 0.00978245f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.177
cc_30 VPB N_VPWR_c_137_n 0.00461568f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.015
cc_31 VPB N_VPWR_c_138_n 0.0117052f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.445
cc_32 VPB N_VPWR_c_139_n 0.00460237f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.295
cc_33 VPB N_VPWR_c_140_n 0.0183554f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.025
cc_34 VPB N_VPWR_c_141_n 0.0167406f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_35 VPB N_VPWR_c_142_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_36 VPB N_VPWR_c_136_n 0.0475378f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_37 N_A_M1000_g N_Y_c_91_n 0.0163534f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_38 N_A_M1001_g N_Y_c_91_n 0.0150272f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_39 N_A_c_39_n N_Y_c_91_n 0.00240036f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_40 A N_Y_c_91_n 0.0426147f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_41 N_A_c_39_n N_Y_c_92_n 0.00589614f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_42 A N_Y_c_92_n 0.0209563f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_43 N_A_M1002_g N_Y_c_86_n 0.00189162f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_44 N_A_M1004_g N_Y_c_86_n 0.00180689f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_45 N_A_M1004_g N_Y_c_87_n 0.0146405f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_46 A N_Y_c_87_n 0.00394157f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A_M1002_g N_Y_c_88_n 0.00568793f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_48 N_A_c_39_n N_Y_c_88_n 0.00241459f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_49 A N_Y_c_88_n 0.0183373f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A_c_39_n N_Y_c_93_n 4.58912e-19 $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_51 N_A_M1003_g N_Y_c_93_n 0.0180233f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_52 A N_Y_c_93_n 0.0024245f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_53 N_A_c_39_n N_Y_c_94_n 0.00232565f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_54 A N_Y_c_94_n 0.0213708f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A_M1003_g Y 0.00683246f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_56 N_A_M1004_g Y 0.0148622f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_57 A Y 0.0184815f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_M1000_g N_VPWR_c_137_n 0.00304967f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_137_n 0.00161372f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_60 N_A_M1003_g N_VPWR_c_139_n 0.00339731f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_M1000_g N_VPWR_c_140_n 0.00585385f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1001_g N_VPWR_c_141_n 0.00585385f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_M1003_g N_VPWR_c_141_n 0.00585385f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_VPWR_c_136_n 0.011554f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_VPWR_c_136_n 0.0105664f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_VPWR_c_136_n 0.0115083f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_VGND_c_163_n 0.00365907f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_39_n N_VGND_c_163_n 0.00633207f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_69 A N_VGND_c_163_n 0.0101104f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_M1002_g N_VGND_c_165_n 5.86108e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_VGND_c_165_n 0.00871096f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_VGND_c_167_n 0.00585385f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_VGND_c_167_n 0.00364083f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1002_g N_VGND_c_169_n 0.0119927f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_VGND_c_169_n 0.00434306f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_76 N_Y_c_91_n N_VPWR_M1000_d 0.00176461f $X=1.01 $Y=1.545 $X2=-0.19 $Y2=-0.24
cc_77 N_Y_c_96_n N_VPWR_M1003_d 0.0029729f $X=1.615 $Y=1.46 $X2=0 $Y2=0
cc_78 N_Y_c_91_n N_VPWR_c_137_n 0.0135055f $X=1.01 $Y=1.545 $X2=0 $Y2=0
cc_79 N_Y_c_96_n N_VPWR_c_139_n 0.0186635f $X=1.615 $Y=1.46 $X2=0 $Y2=0
cc_80 N_Y_c_122_p N_VPWR_c_140_n 0.0135879f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_81 N_Y_c_123_p N_VPWR_c_141_n 0.0125603f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_82 N_Y_M1000_s N_VPWR_c_136_n 0.00253019f $X=0.155 $Y=1.485 $X2=0 $Y2=0
cc_83 N_Y_M1001_s N_VPWR_c_136_n 0.00302653f $X=1 $Y=1.485 $X2=0 $Y2=0
cc_84 N_Y_c_122_p N_VPWR_c_136_n 0.00960102f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_85 N_Y_c_123_p N_VPWR_c_136_n 0.00979076f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_86 N_Y_c_87_n N_VGND_c_165_n 0.0027328f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_87 N_Y_c_90_n N_VGND_c_165_n 0.0230152f $X=1.615 $Y=0.895 $X2=0 $Y2=0
cc_88 N_Y_c_86_n N_VGND_c_167_n 0.0117468f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_89 N_Y_c_87_n N_VGND_c_167_n 0.0023442f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_90 N_Y_M1002_d N_VGND_c_169_n 0.00285545f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_91 N_Y_c_86_n N_VGND_c_169_n 0.00845997f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_92 N_Y_c_87_n N_VGND_c_169_n 0.00409036f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_93 N_Y_c_90_n N_VGND_c_169_n 0.00136789f $X=1.615 $Y=0.895 $X2=0 $Y2=0

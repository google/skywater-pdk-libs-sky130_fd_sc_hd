* File: sky130_fd_sc_hd__a21oi_2.spice
* Created: Thu Aug 27 14:01:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21oi_2.pex.spice"
.subckt sky130_fd_sc_hd__a21oi_2  VNB VPB A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1001 A_285_47# N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.18525 PD=0.925 PS=1.87 NRD=15.228 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_285_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.089375 PD=0.93 PS=0.925 NRD=0 NRS=15.228 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1000_d N_A1_M1009_g A_114_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.06825 PD=0.93 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.1 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1003 A_114_47# N_A2_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.10725 PD=0.86 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.4 SB=75001.2
+ A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1004_d N_B1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.26 PD=0.92 PS=2.1 NRD=0 NRS=24.912 M=1 R=4.33333 SA=75002.3
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_297#_M1002_d N_A2_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1002_s N_A1_M1006_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.14 PD=1.27 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 N_A_27_297#_M1005_d N_A2_M1005_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1010 N_A_27_297#_M1005_d N_B1_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_297#_M1011_d N_B1_M1011_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.36 AS=0.135 PD=2.72 PS=1.27 NRD=18.715 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a21oi_2.pxi.spice"
*
.ends
*
*

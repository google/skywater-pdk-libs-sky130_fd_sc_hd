* File: sky130_fd_sc_hd__bufbuf_8.pex.spice
* Created: Tue Sep  1 18:59:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%A 3 7 9 15
c30 9 0 1.54613e-19 $X=0.235 $Y=1.19
r31 12 15 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r32 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r33 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r34 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.805
r35 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r36 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%A_27_47# 1 2 9 12 16 20 22 23 24 25 28 29
+ 32
c68 29 0 1.54613e-19 $X=0.955 $Y=1.16
c69 24 0 7.44113e-20 $X=0.61 $Y=1.53
r70 29 33 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.947 $Y=1.16
+ $X2=0.947 $Y2=1.325
r71 29 32 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.947 $Y=1.16
+ $X2=0.947 $Y2=0.995
r72 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=1.16 $X2=0.955 $Y2=1.16
r73 24 28 16.9064 $w=2.67e-07 $l=4.65242e-07 $layer=LI1_cond $X=0.61 $Y=1.53
+ $X2=0.825 $Y2=1.16
r74 24 25 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.61 $Y=1.53
+ $X2=0.425 $Y2=1.53
r75 22 28 15.5356 $w=2.67e-07 $l=4.34396e-07 $layer=LI1_cond $X=0.61 $Y=0.82
+ $X2=0.825 $Y2=1.16
r76 22 23 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.61 $Y=0.82
+ $X2=0.425 $Y2=0.82
r77 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r78 18 20 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r79 14 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.425 $Y2=0.82
r80 14 16 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.47
r81 12 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.985
+ $X2=0.955 $Y2=1.325
r82 9 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.56
+ $X2=0.955 $Y2=0.995
r83 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r84 1 16 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%A_206_47# 1 2 9 13 17 21 25 29 33 36 41 45
+ 49 50 51 56
c104 41 0 1.44067e-19 $X=2.475 $Y=1.16
c105 29 0 1.25206e-19 $X=2.765 $Y=1.985
c106 25 0 1.25206e-19 $X=2.765 $Y=0.56
r107 52 54 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.925 $Y=1.16
+ $X2=2.345 $Y2=1.16
r108 49 50 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=1.63 $X2=1.19
+ $Y2=1.545
r109 45 47 16.4563 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=1.19 $Y=0.4
+ $X2=1.19 $Y2=0.825
r110 42 56 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.475 $Y=1.16
+ $X2=2.765 $Y2=1.16
r111 42 54 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=2.475 $Y=1.16
+ $X2=2.345 $Y2=1.16
r112 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.475
+ $Y=1.16 $X2=2.475 $Y2=1.16
r113 39 51 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=1.175
+ $X2=1.295 $Y2=1.175
r114 39 41 60.7227 $w=1.98e-07 $l=1.095e-06 $layer=LI1_cond $X=1.38 $Y=1.175
+ $X2=2.475 $Y2=1.175
r115 37 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.295 $Y=1.275
+ $X2=1.295 $Y2=1.175
r116 37 50 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.295 $Y=1.275
+ $X2=1.295 $Y2=1.545
r117 36 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.295 $Y=1.075
+ $X2=1.295 $Y2=1.175
r118 36 47 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.295 $Y=1.075
+ $X2=1.295 $Y2=0.825
r119 31 49 3.18438 $w=3.78e-07 $l=1.05e-07 $layer=LI1_cond $X=1.19 $Y=1.735
+ $X2=1.19 $Y2=1.63
r120 31 33 17.4383 $w=3.78e-07 $l=5.75e-07 $layer=LI1_cond $X=1.19 $Y=1.735
+ $X2=1.19 $Y2=2.31
r121 27 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.295
+ $X2=2.765 $Y2=1.16
r122 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.765 $Y=1.295
+ $X2=2.765 $Y2=1.985
r123 23 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.025
+ $X2=2.765 $Y2=1.16
r124 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.765 $Y=1.025
+ $X2=2.765 $Y2=0.56
r125 19 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.345 $Y=1.295
+ $X2=2.345 $Y2=1.16
r126 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.345 $Y=1.295
+ $X2=2.345 $Y2=1.985
r127 15 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.345 $Y=1.025
+ $X2=2.345 $Y2=1.16
r128 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.345 $Y=1.025
+ $X2=2.345 $Y2=0.56
r129 11 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.925 $Y=1.295
+ $X2=1.925 $Y2=1.16
r130 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.925 $Y=1.295
+ $X2=1.925 $Y2=1.985
r131 7 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.925 $Y=1.025
+ $X2=1.925 $Y2=1.16
r132 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.925 $Y=1.025
+ $X2=1.925 $Y2=0.56
r133 2 49 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.63
r134 2 33 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=2.31
r135 1 45 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.235 $X2=1.165 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%A_318_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 83 87 88 89 90 93 97 102 104 110 114 117 119 130
c238 130 0 1.44067e-19 $X=6.125 $Y=1.16
r239 129 130 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.705 $Y=1.16
+ $X2=6.125 $Y2=1.16
r240 128 129 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.285 $Y=1.16
+ $X2=5.705 $Y2=1.16
r241 125 126 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.445 $Y=1.16
+ $X2=4.865 $Y2=1.16
r242 124 125 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.025 $Y=1.16
+ $X2=4.445 $Y2=1.16
r243 123 124 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.605 $Y=1.16
+ $X2=4.025 $Y2=1.16
r244 111 128 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=5.015 $Y=1.16
+ $X2=5.285 $Y2=1.16
r245 111 126 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=5.015 $Y=1.16
+ $X2=4.865 $Y2=1.16
r246 110 111 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=5.015
+ $Y=1.16 $X2=5.015 $Y2=1.16
r247 108 123 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=3.315 $Y=1.16
+ $X2=3.605 $Y2=1.16
r248 108 120 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=3.315 $Y=1.16
+ $X2=3.185 $Y2=1.16
r249 107 110 94.2727 $w=1.98e-07 $l=1.7e-06 $layer=LI1_cond $X=3.315 $Y=1.175
+ $X2=5.015 $Y2=1.175
r250 107 108 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.315
+ $Y=1.16 $X2=3.315 $Y2=1.16
r251 105 119 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=1.175
+ $X2=2.975 $Y2=1.175
r252 105 107 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.06 $Y=1.175
+ $X2=3.315 $Y2=1.175
r253 104 117 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=1.445
+ $X2=2.975 $Y2=1.53
r254 103 119 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.975 $Y=1.275
+ $X2=2.975 $Y2=1.175
r255 103 104 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.975 $Y=1.275
+ $X2=2.975 $Y2=1.445
r256 102 119 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.975 $Y=1.075
+ $X2=2.975 $Y2=1.175
r257 101 114 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=0.905
+ $X2=2.975 $Y2=0.82
r258 101 102 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.975 $Y=0.905
+ $X2=2.975 $Y2=1.075
r259 97 99 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.555 $Y=1.63
+ $X2=2.555 $Y2=2.31
r260 95 117 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.555 $Y=1.53
+ $X2=2.975 $Y2=1.53
r261 95 97 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.555 $Y=1.615
+ $X2=2.555 $Y2=1.63
r262 91 114 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.555 $Y=0.82
+ $X2=2.975 $Y2=0.82
r263 91 93 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.555 $Y=0.735
+ $X2=2.555 $Y2=0.4
r264 89 95 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=1.53
+ $X2=2.555 $Y2=1.53
r265 89 90 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.39 $Y=1.53
+ $X2=1.88 $Y2=1.53
r266 87 91 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=0.82
+ $X2=2.555 $Y2=0.82
r267 87 88 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.39 $Y=0.82
+ $X2=1.88 $Y2=0.82
r268 83 85 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.715 $Y=1.63
+ $X2=1.715 $Y2=2.31
r269 81 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.715 $Y=1.615
+ $X2=1.88 $Y2=1.53
r270 81 83 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.715 $Y=1.615
+ $X2=1.715 $Y2=1.63
r271 77 88 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.715 $Y=0.735
+ $X2=1.88 $Y2=0.82
r272 77 79 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.715 $Y=0.735
+ $X2=1.715 $Y2=0.4
r273 73 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.125 $Y=1.295
+ $X2=6.125 $Y2=1.16
r274 73 75 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.125 $Y=1.295
+ $X2=6.125 $Y2=1.985
r275 69 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.125 $Y=1.025
+ $X2=6.125 $Y2=1.16
r276 69 71 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.125 $Y=1.025
+ $X2=6.125 $Y2=0.56
r277 65 129 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.705 $Y=1.295
+ $X2=5.705 $Y2=1.16
r278 65 67 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.705 $Y=1.295
+ $X2=5.705 $Y2=1.985
r279 61 129 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.705 $Y=1.025
+ $X2=5.705 $Y2=1.16
r280 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.705 $Y=1.025
+ $X2=5.705 $Y2=0.56
r281 57 128 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.285 $Y=1.295
+ $X2=5.285 $Y2=1.16
r282 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.285 $Y=1.295
+ $X2=5.285 $Y2=1.985
r283 53 128 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.285 $Y=1.025
+ $X2=5.285 $Y2=1.16
r284 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.285 $Y=1.025
+ $X2=5.285 $Y2=0.56
r285 49 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.865 $Y=1.295
+ $X2=4.865 $Y2=1.16
r286 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.865 $Y=1.295
+ $X2=4.865 $Y2=1.985
r287 45 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.865 $Y=1.025
+ $X2=4.865 $Y2=1.16
r288 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.865 $Y=1.025
+ $X2=4.865 $Y2=0.56
r289 41 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.445 $Y=1.295
+ $X2=4.445 $Y2=1.16
r290 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.445 $Y=1.295
+ $X2=4.445 $Y2=1.985
r291 37 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.445 $Y=1.025
+ $X2=4.445 $Y2=1.16
r292 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.445 $Y=1.025
+ $X2=4.445 $Y2=0.56
r293 33 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.025 $Y=1.295
+ $X2=4.025 $Y2=1.16
r294 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.025 $Y=1.295
+ $X2=4.025 $Y2=1.985
r295 29 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.025 $Y=1.025
+ $X2=4.025 $Y2=1.16
r296 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.025 $Y=1.025
+ $X2=4.025 $Y2=0.56
r297 25 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.605 $Y=1.295
+ $X2=3.605 $Y2=1.16
r298 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.605 $Y=1.295
+ $X2=3.605 $Y2=1.985
r299 21 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.605 $Y=1.025
+ $X2=3.605 $Y2=1.16
r300 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.605 $Y=1.025
+ $X2=3.605 $Y2=0.56
r301 17 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.185 $Y=1.295
+ $X2=3.185 $Y2=1.16
r302 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.185 $Y=1.295
+ $X2=3.185 $Y2=1.985
r303 13 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.185 $Y=1.025
+ $X2=3.185 $Y2=1.16
r304 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.185 $Y=1.025
+ $X2=3.185 $Y2=0.56
r305 4 99 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.485 $X2=2.555 $Y2=2.31
r306 4 97 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.485 $X2=2.555 $Y2=1.63
r307 3 85 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.715 $Y2=2.31
r308 3 83 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.715 $Y2=1.63
r309 2 93 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.42
+ $Y=0.235 $X2=2.555 $Y2=0.4
r310 1 79 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.235 $X2=1.715 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%VPWR 1 2 3 4 5 6 7 24 26 30 34 38 42 46 50
+ 53 54 56 57 59 60 62 63 65 66 67 69 91 92 95 98
c104 1 0 7.44113e-20 $X=0.545 $Y=1.485
r105 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r106 96 99 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r107 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r108 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r109 89 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r110 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r112 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r113 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r114 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r116 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r117 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 77 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 74 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.135 $Y2=2.72
r121 74 76 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 69 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r123 69 71 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 67 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 67 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 65 88 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.25 $Y=2.72 $X2=6.21
+ $Y2=2.72
r127 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.25 $Y=2.72
+ $X2=6.335 $Y2=2.72
r128 64 91 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.42 $Y=2.72
+ $X2=6.67 $Y2=2.72
r129 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.72
+ $X2=6.335 $Y2=2.72
r130 62 85 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.41 $Y=2.72
+ $X2=5.29 $Y2=2.72
r131 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=2.72
+ $X2=5.495 $Y2=2.72
r132 61 88 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.58 $Y=2.72
+ $X2=6.21 $Y2=2.72
r133 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=2.72
+ $X2=5.495 $Y2=2.72
r134 59 82 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.57 $Y=2.72 $X2=4.37
+ $Y2=2.72
r135 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=2.72
+ $X2=4.655 $Y2=2.72
r136 58 85 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.74 $Y=2.72
+ $X2=5.29 $Y2=2.72
r137 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=2.72
+ $X2=4.655 $Y2=2.72
r138 56 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.815 $Y2=2.72
r140 55 82 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.9 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=2.72
+ $X2=3.815 $Y2=2.72
r142 53 76 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.89 $Y=2.72
+ $X2=2.53 $Y2=2.72
r143 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=2.72
+ $X2=2.975 $Y2=2.72
r144 52 79 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=3.45 $Y2=2.72
r145 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=2.975 $Y2=2.72
r146 48 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=2.635
+ $X2=6.335 $Y2=2.72
r147 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.335 $Y=2.635
+ $X2=6.335 $Y2=2
r148 44 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.72
r149 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2
r150 40 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=2.635
+ $X2=4.655 $Y2=2.72
r151 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.655 $Y=2.635
+ $X2=4.655 $Y2=2
r152 36 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=2.635
+ $X2=3.815 $Y2=2.72
r153 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.815 $Y=2.635
+ $X2=3.815 $Y2=2
r154 32 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.72
r155 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2
r156 28 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.635
+ $X2=2.135 $Y2=2.72
r157 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.135 $Y=2.635
+ $X2=2.135 $Y2=2
r158 27 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r159 26 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.72
+ $X2=2.135 $Y2=2.72
r160 26 27 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=2.05 $Y=2.72
+ $X2=0.765 $Y2=2.72
r161 22 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r162 22 24 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=1.95
r163 7 50 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.2
+ $Y=1.485 $X2=6.335 $Y2=2
r164 6 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.36
+ $Y=1.485 $X2=5.495 $Y2=2
r165 5 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.52
+ $Y=1.485 $X2=4.655 $Y2=2
r166 4 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=1.485 $X2=3.815 $Y2=2
r167 3 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.84
+ $Y=1.485 $X2=2.975 $Y2=2
r168 2 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.485 $X2=2.135 $Y2=2
r169 1 24 600 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 79 81 82 83 84 85 86 88 89
c163 38 0 1.25206e-19 $X=3.56 $Y=1.53
c164 36 0 1.25206e-19 $X=3.56 $Y=0.82
r165 88 89 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.625 $Y=1.19
+ $X2=6.625 $Y2=1.445
r166 87 88 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=6.625 $Y=0.905
+ $X2=6.625 $Y2=1.19
r167 80 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=1.53
+ $X2=5.915 $Y2=1.53
r168 79 89 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.435 $Y=1.53
+ $X2=6.625 $Y2=1.53
r169 79 80 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.435 $Y=1.53
+ $X2=6.08 $Y2=1.53
r170 78 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0.82
+ $X2=5.915 $Y2=0.82
r171 77 87 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=6.435 $Y=0.82
+ $X2=6.625 $Y2=0.905
r172 77 78 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.435 $Y=0.82
+ $X2=6.08 $Y2=0.82
r173 73 75 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.915 $Y=1.63
+ $X2=5.915 $Y2=2.31
r174 71 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=1.615
+ $X2=5.915 $Y2=1.53
r175 71 73 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.915 $Y=1.615
+ $X2=5.915 $Y2=1.63
r176 67 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=0.735
+ $X2=5.915 $Y2=0.82
r177 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.915 $Y=0.735
+ $X2=5.915 $Y2=0.4
r178 66 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.24 $Y=1.53
+ $X2=5.075 $Y2=1.53
r179 65 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=1.53
+ $X2=5.915 $Y2=1.53
r180 65 66 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.75 $Y=1.53
+ $X2=5.24 $Y2=1.53
r181 64 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.24 $Y=0.82
+ $X2=5.075 $Y2=0.82
r182 63 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=0.82
+ $X2=5.915 $Y2=0.82
r183 63 64 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.75 $Y=0.82
+ $X2=5.24 $Y2=0.82
r184 59 61 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.075 $Y=1.63
+ $X2=5.075 $Y2=2.31
r185 57 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=1.615
+ $X2=5.075 $Y2=1.53
r186 57 59 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.075 $Y=1.615
+ $X2=5.075 $Y2=1.63
r187 53 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=0.735
+ $X2=5.075 $Y2=0.82
r188 53 55 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.075 $Y=0.735
+ $X2=5.075 $Y2=0.4
r189 52 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=1.53
+ $X2=4.235 $Y2=1.53
r190 51 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.91 $Y=1.53
+ $X2=5.075 $Y2=1.53
r191 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.91 $Y=1.53
+ $X2=4.4 $Y2=1.53
r192 50 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=0.82
+ $X2=4.235 $Y2=0.82
r193 49 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.91 $Y=0.82
+ $X2=5.075 $Y2=0.82
r194 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.91 $Y=0.82
+ $X2=4.4 $Y2=0.82
r195 45 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.235 $Y=1.63
+ $X2=4.235 $Y2=2.31
r196 43 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.235 $Y=1.615
+ $X2=4.235 $Y2=1.53
r197 43 45 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.235 $Y=1.615
+ $X2=4.235 $Y2=1.63
r198 39 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.235 $Y=0.735
+ $X2=4.235 $Y2=0.82
r199 39 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.235 $Y=0.735
+ $X2=4.235 $Y2=0.4
r200 37 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=1.53
+ $X2=4.235 $Y2=1.53
r201 37 38 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.07 $Y=1.53
+ $X2=3.56 $Y2=1.53
r202 35 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0.82
+ $X2=4.235 $Y2=0.82
r203 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.07 $Y=0.82
+ $X2=3.56 $Y2=0.82
r204 31 33 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.395 $Y=1.63
+ $X2=3.395 $Y2=2.31
r205 29 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=1.615
+ $X2=3.56 $Y2=1.53
r206 29 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.395 $Y=1.615
+ $X2=3.395 $Y2=1.63
r207 25 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=0.735
+ $X2=3.56 $Y2=0.82
r208 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.395 $Y=0.735
+ $X2=3.395 $Y2=0.4
r209 8 75 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=1.485 $X2=5.915 $Y2=2.31
r210 8 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=1.485 $X2=5.915 $Y2=1.63
r211 7 61 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=4.94
+ $Y=1.485 $X2=5.075 $Y2=2.31
r212 7 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.94
+ $Y=1.485 $X2=5.075 $Y2=1.63
r213 6 47 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=4.1
+ $Y=1.485 $X2=4.235 $Y2=2.31
r214 6 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.1
+ $Y=1.485 $X2=4.235 $Y2=1.63
r215 5 33 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.485 $X2=3.395 $Y2=2.31
r216 5 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.485 $X2=3.395 $Y2=1.63
r217 4 69 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.78
+ $Y=0.235 $X2=5.915 $Y2=0.4
r218 3 55 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.94
+ $Y=0.235 $X2=5.075 $Y2=0.4
r219 2 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.1
+ $Y=0.235 $X2=4.235 $Y2=0.4
r220 1 27 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.26
+ $Y=0.235 $X2=3.395 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_8%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 50
+ 53 54 56 57 59 60 62 63 65 66 67 69 91 92 95 98
r122 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r123 96 99 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r124 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r125 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r126 89 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r127 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r128 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r129 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r130 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r131 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r132 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r133 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r134 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r135 77 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r136 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r137 74 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.135
+ $Y2=0
r138 74 76 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.53
+ $Y2=0
r139 69 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r140 69 71 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r141 67 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r142 67 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r143 65 88 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.25 $Y=0 $X2=6.21
+ $Y2=0
r144 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.25 $Y=0 $X2=6.335
+ $Y2=0
r145 64 91 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.42 $Y=0 $X2=6.67
+ $Y2=0
r146 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0 $X2=6.335
+ $Y2=0
r147 62 85 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.29
+ $Y2=0
r148 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.495
+ $Y2=0
r149 61 88 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.58 $Y=0 $X2=6.21
+ $Y2=0
r150 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=0 $X2=5.495
+ $Y2=0
r151 59 82 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.57 $Y=0 $X2=4.37
+ $Y2=0
r152 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=0 $X2=4.655
+ $Y2=0
r153 58 85 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=5.29
+ $Y2=0
r154 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.655
+ $Y2=0
r155 56 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=0 $X2=3.45
+ $Y2=0
r156 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=0 $X2=3.815
+ $Y2=0
r157 55 82 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.9 $Y=0 $X2=4.37
+ $Y2=0
r158 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=0 $X2=3.815
+ $Y2=0
r159 53 76 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.53
+ $Y2=0
r160 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.975
+ $Y2=0
r161 52 79 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.06 $Y=0 $X2=3.45
+ $Y2=0
r162 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=0 $X2=2.975
+ $Y2=0
r163 48 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0.085
+ $X2=6.335 $Y2=0
r164 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.335 $Y=0.085
+ $X2=6.335 $Y2=0.4
r165 44 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=0.085
+ $X2=5.495 $Y2=0
r166 44 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.495 $Y=0.085
+ $X2=5.495 $Y2=0.4
r167 40 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0
r168 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0.4
r169 36 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r170 36 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.4
r171 32 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=0.085
+ $X2=2.975 $Y2=0
r172 32 34 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.975 $Y=0.085
+ $X2=2.975 $Y2=0.4
r173 28 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.135 $Y2=0
r174 28 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.135 $Y2=0.4
r175 27 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r176 26 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.135
+ $Y2=0
r177 26 27 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=2.05 $Y=0
+ $X2=0.765 $Y2=0
r178 22 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r179 22 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r180 7 50 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.235 $X2=6.335 $Y2=0.4
r181 6 46 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.36
+ $Y=0.235 $X2=5.495 $Y2=0.4
r182 5 42 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.52
+ $Y=0.235 $X2=4.655 $Y2=0.4
r183 4 38 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.68
+ $Y=0.235 $X2=3.815 $Y2=0.4
r184 3 34 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.235 $X2=2.975 $Y2=0.4
r185 2 30 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.235 $X2=2.135 $Y2=0.4
r186 1 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends


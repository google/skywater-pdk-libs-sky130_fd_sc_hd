* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
M1000 a_455_47# a_301_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.7485e+12p pd=1.708e+07u as=1.1245e+12p ps=1.126e+07u
M1001 Z a_116_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=0p ps=0u
M1002 a_407_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=2.8613e+12p pd=2.338e+07u as=1.6652e+12p ps=1.498e+07u
M1003 a_407_309# a_116_47# Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.08e+12p ps=1.016e+07u
M1004 VGND A a_116_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1005 a_455_47# a_301_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_455_47# a_116_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_301_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR TE_B a_407_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z a_116_47# a_407_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_301_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR TE_B a_407_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_301_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_407_309# a_116_47# Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_301_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_455_47# a_301_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_407_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_407_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_407_309# a_116_47# Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_116_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1020 a_116_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_455_47# a_301_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR TE_B a_407_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z a_116_47# a_407_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Z a_116_47# a_407_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_301_47# TE_B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1026 Z a_116_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_455_47# a_116_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR TE_B a_407_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Z a_116_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_407_309# a_116_47# Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_301_47# TE_B VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1032 a_455_47# a_116_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_455_47# a_116_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Z a_116_47# a_455_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Z a_116_47# a_407_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_116_47# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_407_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__a21boi_0.pex.spice
* Created: Thu Aug 27 14:00:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BOI_0%B1_N 3 6 9 11 12 15 16
c35 3 0 4.73589e-20 $X=0.475 $Y=0.445
r36 15 17 41.4854 $w=3.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.575 $Y=1.4
+ $X2=0.575 $Y2=1.265
r37 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.4 $X2=0.585 $Y2=1.4
r38 12 16 12.7447 $w=4.23e-07 $l=4.7e-07 $layer=LI1_cond $X=0.682 $Y=1.87
+ $X2=0.682 $Y2=1.4
r39 9 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.475 $Y=2.275
+ $X2=0.475 $Y2=1.885
r40 6 11 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.575 $Y=1.71
+ $X2=0.575 $Y2=1.885
r41 5 15 6.59477 $w=3.5e-07 $l=4e-08 $layer=POLY_cond $X=0.575 $Y=1.44 $X2=0.575
+ $Y2=1.4
r42 5 6 44.5147 $w=3.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.575 $Y=1.44
+ $X2=0.575 $Y2=1.71
r43 3 17 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.265
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%A_27_47# 1 2 7 8 9 11 14 16 19 25 28 30 31
c59 9 0 1.11678e-19 $X=1.245 $Y=0.77
r60 30 31 10.0776 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.225 $Y=2.3
+ $X2=0.225 $Y2=2.085
r61 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=0.93 $X2=0.98 $Y2=0.93
r62 23 28 1.26991 $w=2.5e-07 $l=1.43e-07 $layer=LI1_cond $X=0.38 $Y=0.905
+ $X2=0.237 $Y2=0.905
r63 23 25 27.6586 $w=2.48e-07 $l=6e-07 $layer=LI1_cond $X=0.38 $Y=0.905 $X2=0.98
+ $Y2=0.905
r64 21 28 5.25345 $w=2.45e-07 $l=1.43614e-07 $layer=LI1_cond $X=0.197 $Y=1.03
+ $X2=0.237 $Y2=0.905
r65 21 31 57.0776 $w=2.03e-07 $l=1.055e-06 $layer=LI1_cond $X=0.197 $Y=1.03
+ $X2=0.197 $Y2=2.085
r66 17 28 5.25345 $w=2.45e-07 $l=1.25e-07 $layer=LI1_cond $X=0.237 $Y=0.78
+ $X2=0.237 $Y2=0.905
r67 17 19 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=0.237 $Y=0.78
+ $X2=0.237 $Y2=0.445
r68 14 16 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.425 $Y=2.165
+ $X2=1.425 $Y2=1.68
r69 9 26 45.6624 $w=6.54e-07 $l=1.99198e-07 $layer=POLY_cond $X=1.245 $Y=0.77
+ $X2=1.157 $Y2=0.93
r70 9 11 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.245 $Y=0.77
+ $X2=1.245 $Y2=0.445
r71 8 16 54.9885 $w=4.9e-07 $l=2.45e-07 $layer=POLY_cond $X=1.255 $Y=1.435
+ $X2=1.255 $Y2=1.68
r72 7 26 13.088 $w=6.54e-07 $l=1.77356e-07 $layer=POLY_cond $X=1.255 $Y=1.065
+ $X2=1.157 $Y2=0.93
r73 7 8 40.4002 $w=4.9e-07 $l=3.7e-07 $layer=POLY_cond $X=1.255 $Y=1.065
+ $X2=1.255 $Y2=1.435
r74 2 30 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r75 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%A1 3 7 8 9 11 12 15 16
c44 16 0 3.43796e-21 $X=1.865 $Y=0.93
c45 8 0 1.0824e-19 $X=1.865 $Y=0.9
c46 3 0 1.07878e-19 $X=1.855 $Y=2.165
r47 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.865
+ $Y=0.93 $X2=1.865 $Y2=0.93
r48 12 16 17.7299 $w=3.88e-07 $l=6e-07 $layer=LI1_cond $X=1.975 $Y=1.53
+ $X2=1.975 $Y2=0.93
r49 10 15 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=1.865 $Y=1.3
+ $X2=1.865 $Y2=0.93
r50 10 11 36.4065 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.865 $Y=1.3
+ $X2=1.865 $Y2=1.435
r51 8 15 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=1.865 $Y=0.9 $X2=1.865
+ $Y2=0.93
r52 8 9 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.865 $Y=0.9
+ $X2=1.865 $Y2=0.765
r53 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=0.445
+ $X2=1.925 $Y2=0.765
r54 3 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.855 $Y=2.165
+ $X2=1.855 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%A2 3 5 8 10 11 14 16
r30 14 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=0.93
+ $X2=2.39 $Y2=0.765
r31 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.435
+ $Y=0.93 $X2=2.435 $Y2=0.93
r32 11 15 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=2.477 $Y=0.85
+ $X2=2.477 $Y2=0.93
r33 8 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.285 $Y=2.165
+ $X2=2.285 $Y2=1.435
r34 5 10 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.39 $Y=1.255 $X2=2.39
+ $Y2=1.435
r35 4 14 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.39 $Y=0.945
+ $X2=2.39 $Y2=0.93
r36 4 5 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=2.39 $Y=0.945 $X2=2.39
+ $Y2=1.255
r37 3 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.285 $Y=0.445
+ $X2=2.285 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%VPWR 1 2 9 13 15 17 22 29 30 33 36
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 27 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r49 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 23 25 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 22 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r59 11 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.635
+ $X2=2.07 $Y2=2.72
r60 11 13 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.07 $Y=2.635
+ $X2=2.07 $Y2=2.34
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635 $X2=0.69
+ $Y2=2.72
r62 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=2.635 $X2=0.69
+ $Y2=2.3
r63 2 13 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.845 $X2=2.07 $Y2=2.34
r64 1 9 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.065 $X2=0.69 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%Y 1 2 7 9 16
c33 16 0 1.07878e-19 $X=1.15 $Y=2.21
c34 7 0 4.73589e-20 $X=1.462 $Y=1.2
r35 12 16 24.4894 $w=2.38e-07 $l=5.1e-07 $layer=LI1_cond $X=1.185 $Y=1.655
+ $X2=1.185 $Y2=2.165
r36 11 12 4.4837 $w=2.4e-07 $l=2.28e-07 $layer=LI1_cond $X=1.185 $Y=1.427
+ $X2=1.185 $Y2=1.655
r37 7 11 7.28162 $w=4.53e-07 $l=2.77e-07 $layer=LI1_cond $X=1.462 $Y=1.427
+ $X2=1.185 $Y2=1.427
r38 7 9 29.4947 $w=2.93e-07 $l=7.55e-07 $layer=LI1_cond $X=1.462 $Y=1.2
+ $X2=1.462 $Y2=0.445
r39 2 16 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.845 $X2=1.21 $Y2=2.165
r40 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.32
+ $Y=0.235 $X2=1.46 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%A_300_369# 1 2 9 14 16
r29 10 14 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=1.915
+ $X2=1.64 $Y2=1.915
r30 9 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=1.915
+ $X2=2.5 $Y2=1.915
r31 9 10 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=2.335 $Y=1.915
+ $X2=1.805 $Y2=1.915
r32 2 16 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=1.845 $X2=2.5 $Y2=1.99
r33 1 14 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.845 $X2=1.64 $Y2=1.97
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_0%VGND 1 2 7 9 11 13 18 35
r34 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r35 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r36 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r37 22 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r38 22 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r39 21 24 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r40 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r41 19 21 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.145 $Y=0 $X2=1.15
+ $Y2=0
r42 18 34 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.547
+ $Y2=0
r43 18 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.07
+ $Y2=0
r44 13 31 8.94546 $w=5.93e-07 $l=4.45e-07 $layer=LI1_cond $X=0.847 $Y=0
+ $X2=0.847 $Y2=0.445
r45 13 19 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.847 $Y=0 $X2=1.145
+ $Y2=0
r46 13 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 13 15 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.23
+ $Y2=0
r48 11 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r49 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r50 7 34 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.5 $Y=0.085
+ $X2=2.547 $Y2=0
r51 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.5 $Y=0.085 $X2=2.5
+ $Y2=0.43
r52 2 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.235 $X2=2.5 $Y2=0.43
r53 1 31 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.03 $Y2=0.445
.ends


* File: sky130_fd_sc_hd__fa_1.spice.SKY130_FD_SC_HD__FA_1.pxi
* Created: Thu Aug 27 14:21:04 2020
* 
x_PM_SKY130_FD_SC_HD__FA_1%A_76_199# N_A_76_199#_M1025_d N_A_76_199#_M1018_d
+ N_A_76_199#_M1024_g N_A_76_199#_M1017_g N_A_76_199#_M1007_g
+ N_A_76_199#_M1010_g N_A_76_199#_c_191_n N_A_76_199#_c_178_n
+ N_A_76_199#_c_309_p N_A_76_199#_c_242_p N_A_76_199#_c_179_n
+ N_A_76_199#_c_180_n N_A_76_199#_c_181_n N_A_76_199#_c_182_n
+ N_A_76_199#_c_183_n N_A_76_199#_c_184_n N_A_76_199#_c_185_n
+ N_A_76_199#_c_186_n N_A_76_199#_c_187_n N_A_76_199#_c_188_n
+ PM_SKY130_FD_SC_HD__FA_1%A_76_199#
x_PM_SKY130_FD_SC_HD__FA_1%A N_A_M1020_g N_A_M1011_g N_A_M1001_g N_A_M1009_g
+ N_A_M1019_g N_A_M1003_g N_A_M1013_g N_A_M1015_g A N_A_c_351_n N_A_c_352_n
+ N_A_c_353_n N_A_c_354_n N_A_c_355_n N_A_c_356_n N_A_c_357_n N_A_c_358_n
+ N_A_c_359_n N_A_c_360_n N_A_c_361_n N_A_c_362_n N_A_c_363_n N_A_c_364_n
+ PM_SKY130_FD_SC_HD__FA_1%A
x_PM_SKY130_FD_SC_HD__FA_1%B N_B_M1025_g N_B_M1018_g N_B_c_587_n N_B_M1000_g
+ N_B_c_595_n N_B_M1005_g N_B_c_588_n N_B_c_589_n N_B_c_596_n N_B_c_597_n
+ N_B_M1026_g N_B_c_598_n N_B_M1022_g N_B_M1004_g N_B_M1027_g N_B_c_601_n
+ N_B_c_591_n N_B_c_603_n N_B_c_592_n B N_B_c_605_n N_B_c_606_n N_B_c_607_n
+ N_B_c_608_n N_B_c_609_n N_B_c_610_n N_B_c_611_n N_B_c_612_n N_B_c_613_n
+ N_B_c_614_n PM_SKY130_FD_SC_HD__FA_1%B
x_PM_SKY130_FD_SC_HD__FA_1%CIN N_CIN_M1023_g N_CIN_M1012_g N_CIN_M1014_g
+ N_CIN_M1008_g N_CIN_M1002_g N_CIN_M1021_g N_CIN_c_811_n N_CIN_c_812_n
+ N_CIN_c_813_n N_CIN_c_826_n N_CIN_c_827_n N_CIN_c_814_n N_CIN_c_815_n
+ N_CIN_c_816_n N_CIN_c_817_n N_CIN_c_830_n N_CIN_c_831_n N_CIN_c_832_n
+ N_CIN_c_818_n N_CIN_c_819_n CIN N_CIN_c_820_n N_CIN_c_835_n N_CIN_c_836_n
+ PM_SKY130_FD_SC_HD__FA_1%CIN
x_PM_SKY130_FD_SC_HD__FA_1%A_995_47# N_A_995_47#_M1007_d N_A_995_47#_M1010_d
+ N_A_995_47#_M1016_g N_A_995_47#_M1006_g N_A_995_47#_c_1052_n
+ N_A_995_47#_c_1034_n N_A_995_47#_c_1035_n N_A_995_47#_c_1041_n
+ N_A_995_47#_c_1042_n N_A_995_47#_c_1048_n N_A_995_47#_c_1043_n
+ N_A_995_47#_c_1036_n N_A_995_47#_c_1037_n N_A_995_47#_c_1038_n
+ N_A_995_47#_c_1039_n PM_SKY130_FD_SC_HD__FA_1%A_995_47#
x_PM_SKY130_FD_SC_HD__FA_1%COUT N_COUT_M1024_s N_COUT_M1017_s N_COUT_c_1129_n
+ N_COUT_c_1132_n N_COUT_c_1130_n COUT COUT COUT N_COUT_c_1134_n
+ PM_SKY130_FD_SC_HD__FA_1%COUT
x_PM_SKY130_FD_SC_HD__FA_1%VPWR N_VPWR_M1017_d N_VPWR_M1009_d N_VPWR_M1022_s
+ N_VPWR_M1008_d N_VPWR_M1015_d N_VPWR_c_1148_n N_VPWR_c_1149_n N_VPWR_c_1150_n
+ N_VPWR_c_1151_n N_VPWR_c_1152_n N_VPWR_c_1153_n N_VPWR_c_1154_n VPWR VPWR
+ N_VPWR_c_1155_n VPWR N_VPWR_c_1156_n N_VPWR_c_1157_n N_VPWR_c_1158_n
+ N_VPWR_c_1159_n N_VPWR_c_1147_n N_VPWR_c_1161_n N_VPWR_c_1162_n
+ N_VPWR_c_1163_n N_VPWR_c_1164_n PM_SKY130_FD_SC_HD__FA_1%VPWR
x_PM_SKY130_FD_SC_HD__FA_1%A_382_413# N_A_382_413#_M1012_d N_A_382_413#_M1005_d
+ N_A_382_413#_c_1281_n N_A_382_413#_c_1264_n N_A_382_413#_c_1265_n
+ N_A_382_413#_c_1266_n PM_SKY130_FD_SC_HD__FA_1%A_382_413#
x_PM_SKY130_FD_SC_HD__FA_1%A_738_413# N_A_738_413#_M1022_d N_A_738_413#_M1003_d
+ N_A_738_413#_c_1308_n N_A_738_413#_c_1291_n N_A_738_413#_c_1292_n
+ N_A_738_413#_c_1305_n PM_SKY130_FD_SC_HD__FA_1%A_738_413#
x_PM_SKY130_FD_SC_HD__FA_1%SUM N_SUM_M1016_d N_SUM_M1006_d SUM SUM SUM SUM SUM
+ SUM SUM N_SUM_c_1325_n SUM PM_SKY130_FD_SC_HD__FA_1%SUM
x_PM_SKY130_FD_SC_HD__FA_1%VGND N_VGND_M1024_d N_VGND_M1001_d N_VGND_M1026_s
+ N_VGND_M1014_d N_VGND_M1013_d N_VGND_c_1337_n N_VGND_c_1338_n N_VGND_c_1339_n
+ N_VGND_c_1340_n N_VGND_c_1341_n N_VGND_c_1342_n N_VGND_c_1343_n VGND VGND
+ N_VGND_c_1344_n VGND N_VGND_c_1345_n N_VGND_c_1346_n N_VGND_c_1347_n
+ N_VGND_c_1348_n N_VGND_c_1349_n N_VGND_c_1350_n N_VGND_c_1351_n
+ N_VGND_c_1352_n N_VGND_c_1353_n PM_SKY130_FD_SC_HD__FA_1%VGND
x_PM_SKY130_FD_SC_HD__FA_1%A_382_47# N_A_382_47#_M1023_d N_A_382_47#_M1000_d
+ N_A_382_47#_c_1492_n N_A_382_47#_c_1467_n N_A_382_47#_c_1468_n
+ N_A_382_47#_c_1484_n PM_SKY130_FD_SC_HD__FA_1%A_382_47#
x_PM_SKY130_FD_SC_HD__FA_1%A_738_47# N_A_738_47#_M1026_d N_A_738_47#_M1019_d
+ N_A_738_47#_c_1524_n N_A_738_47#_c_1502_n N_A_738_47#_c_1503_n
+ N_A_738_47#_c_1521_n PM_SKY130_FD_SC_HD__FA_1%A_738_47#
cc_1 VNB N_A_76_199#_M1007_g 0.0223326f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=0.445
cc_2 VNB N_A_76_199#_M1010_g 0.00503421f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=2.275
cc_3 VNB N_A_76_199#_c_178_n 0.00254803f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=0.72
cc_4 VNB N_A_76_199#_c_179_n 0.00184612f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_5 VNB N_A_76_199#_c_180_n 0.0229624f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_6 VNB N_A_76_199#_c_181_n 0.00107287f $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=0.995
cc_7 VNB N_A_76_199#_c_182_n 0.0121497f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.85
cc_8 VNB N_A_76_199#_c_183_n 0.00176616f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=0.85
cc_9 VNB N_A_76_199#_c_184_n 0.0070582f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=0.85
cc_10 VNB N_A_76_199#_c_185_n 0.00440688f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=0.85
cc_11 VNB N_A_76_199#_c_186_n 0.0192349f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_12 VNB N_A_76_199#_c_187_n 0.024338f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=1.04
cc_13 VNB N_A_76_199#_c_188_n 0.0102777f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=1.04
cc_14 VNB N_A_M1020_g 0.0287646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_M1001_g 0.0299029f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_16 VNB N_A_M1019_g 0.0198556f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=2.275
cc_17 VNB N_A_M1003_g 0.00424732f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.995
cc_18 VNB N_A_M1013_g 0.0269376f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.72
cc_19 VNB N_A_M1015_g 8.20116e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB A 0.00573968f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_21 VNB N_A_c_351_n 0.00312666f $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=0.995
cc_22 VNB N_A_c_352_n 0.00156436f $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=1.325
cc_23 VNB N_A_c_353_n 0.00605362f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=2.265
cc_24 VNB N_A_c_354_n 8.64789e-19 $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.85
cc_25 VNB N_A_c_355_n 0.00817331f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=0.85
cc_26 VNB N_A_c_356_n 0.00123023f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=0.85
cc_27 VNB N_A_c_357_n 0.00253456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_c_358_n 0.00243525f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=1.04
cc_29 VNB N_A_c_359_n 0.0204657f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=0.595
cc_30 VNB N_A_c_360_n 0.0224949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_c_361_n 0.0244928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_c_362_n 0.0070021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_c_363_n 0.0243451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_c_364_n 0.00687449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_B_M1025_g 0.0402388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_B_c_587_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_37 VNB N_B_c_588_n 0.0642743f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=0.445
cc_38 VNB N_B_c_589_n 0.00947258f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=0.445
cc_39 VNB N_B_M1004_g 0.0420425f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=2.265
cc_40 VNB N_B_c_591_n 0.0213839f $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=1.325
cc_41 VNB N_B_c_592_n 0.0171497f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=0.85
cc_42 VNB N_CIN_M1023_g 0.0283504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_CIN_M1002_g 0.0375252f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=2.275
cc_44 VNB N_CIN_c_811_n 0.0134432f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=0.72
cc_45 VNB N_CIN_c_812_n 0.00665379f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.72
cc_46 VNB N_CIN_c_813_n 3.21027e-19 $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=2.265
cc_47 VNB N_CIN_c_814_n 0.00130567f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_48 VNB N_CIN_c_815_n 0.0174754f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_49 VNB N_CIN_c_816_n 0.00451859f $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=0.995
cc_50 VNB N_CIN_c_817_n 7.97928e-19 $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=2.265
cc_51 VNB N_CIN_c_818_n 0.019004f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=0.85
cc_52 VNB N_CIN_c_819_n 0.00314327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_CIN_c_820_n 0.0206121f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=1.04
cc_54 VNB N_A_995_47#_c_1034_n 0.00271197f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=1.205
cc_55 VNB N_A_995_47#_c_1035_n 0.00150869f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=2.275
cc_56 VNB N_A_995_47#_c_1036_n 0.00172275f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=0.85
cc_57 VNB N_A_995_47#_c_1037_n 0.0228508f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=0.85
cc_58 VNB N_A_995_47#_c_1038_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_995_47#_c_1039_n 0.0194896f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=0.85
cc_60 VNB N_COUT_c_1129_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_61 VNB N_COUT_c_1130_n 0.0215722f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_62 VNB COUT 0.0172322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VPWR_c_1147_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB SUM 0.0264328f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_65 VNB SUM 0.0263963f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.325
cc_66 VNB N_VGND_c_1337_n 0.00280508f $X=-0.19 $Y=-0.24 $X2=4.9 $Y2=1.205
cc_67 VNB N_VGND_c_1338_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.805
cc_68 VNB N_VGND_c_1339_n 0.0049662f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=0.72
cc_69 VNB N_VGND_c_1340_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=2.275
cc_70 VNB N_VGND_c_1341_n 0.00280508f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_71 VNB N_VGND_c_1342_n 0.0439664f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=2.265
cc_72 VNB N_VGND_c_1343_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.85
cc_73 VNB N_VGND_c_1344_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1345_n 0.035829f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.325
cc_75 VNB N_VGND_c_1346_n 0.0159136f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=0.445
cc_76 VNB N_VGND_c_1347_n 0.0116974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1348_n 0.0224232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1349_n 0.35695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1350_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1351_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1352_n 0.00507318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1353_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_382_47#_c_1467_n 0.00310751f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_84 VNB N_A_382_47#_c_1468_n 0.00259269f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_85 VNB N_A_738_47#_c_1502_n 0.00560037f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_86 VNB N_A_738_47#_c_1503_n 0.00218712f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_87 VPB N_A_76_199#_M1017_g 0.0219161f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_88 VPB N_A_76_199#_M1010_g 0.0499078f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=2.275
cc_89 VPB N_A_76_199#_c_191_n 0.00946185f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.625
cc_90 VPB N_A_76_199#_c_180_n 0.00500576f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_91 VPB N_A_M1011_g 0.0477743f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_92 VPB N_A_M1009_g 0.0513423f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=0.445
cc_93 VPB N_A_M1003_g 0.0468785f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.995
cc_94 VPB N_A_M1015_g 0.0522983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB A 4.61303e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_96 VPB N_A_c_352_n 0.0052097f $X=-0.19 $Y=1.305 $X2=0.557 $Y2=1.325
cc_97 VPB N_A_c_354_n 2.38594e-19 $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.85
cc_98 VPB N_A_c_356_n 5.14832e-19 $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.85
cc_99 VPB N_A_c_357_n 0.00184442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_c_358_n 0.00521027f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=1.04
cc_101 VPB N_A_c_359_n 0.00510517f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.595
cc_102 VPB N_A_c_360_n 0.00705974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_B_M1025_g 0.0117641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_B_M1018_g 0.0207646f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_105 VPB N_B_c_595_n 0.0172359f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_106 VPB N_B_c_596_n 0.0370539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_B_c_597_n 0.00873481f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=1.205
cc_108 VPB N_B_c_598_n 0.0170553f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_109 VPB N_B_M1004_g 0.00999311f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=2.265
cc_110 VPB N_B_M1027_g 0.0222209f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_111 VPB N_B_c_601_n 0.0158992f $X=-0.19 $Y=1.305 $X2=0.557 $Y2=0.995
cc_112 VPB N_B_c_591_n 0.0085167f $X=-0.19 $Y=1.305 $X2=0.557 $Y2=1.325
cc_113 VPB N_B_c_603_n 0.0144932f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.85
cc_114 VPB B 0.00726369f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.85
cc_115 VPB N_B_c_605_n 0.00754267f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.85
cc_116 VPB N_B_c_606_n 0.00312395f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.85
cc_117 VPB N_B_c_607_n 0.0115214f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.85
cc_118 VPB N_B_c_608_n 7.35744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_B_c_609_n 0.00504967f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=0.875
cc_120 VPB N_B_c_610_n 0.00238729f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.595
cc_121 VPB N_B_c_611_n 0.00894792f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=0.595
cc_122 VPB N_B_c_612_n 0.0215382f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.945
cc_123 VPB N_B_c_613_n 0.0254707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_B_c_614_n 0.0237398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_CIN_M1012_g 0.0444312f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_126 VPB N_CIN_M1008_g 0.0249875f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=0.875
cc_127 VPB N_CIN_M1002_g 0.0105544f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=2.275
cc_128 VPB N_CIN_M1021_g 0.0216681f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_129 VPB N_CIN_c_813_n 0.00299774f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=2.265
cc_130 VPB N_CIN_c_826_n 0.0149956f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=2.275
cc_131 VPB N_CIN_c_827_n 0.00269299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_CIN_c_814_n 0.00743298f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_133 VPB N_CIN_c_817_n 0.00264134f $X=-0.19 $Y=1.305 $X2=1.105 $Y2=2.265
cc_134 VPB N_CIN_c_830_n 0.0176538f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.85
cc_135 VPB N_CIN_c_831_n 0.00211333f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=0.85
cc_136 VPB N_CIN_c_832_n 0.0248509f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.85
cc_137 VPB N_CIN_c_818_n 0.00663712f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.85
cc_138 VPB N_CIN_c_820_n 0.0070998f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=1.04
cc_139 VPB N_CIN_c_835_n 0.024639f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=1.205
cc_140 VPB N_CIN_c_836_n 0.00516339f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=1.04
cc_141 VPB N_A_995_47#_M1006_g 0.0218927f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_142 VPB N_A_995_47#_c_1041_n 0.00238948f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.805
cc_143 VPB N_A_995_47#_c_1042_n 0.00133231f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.72
cc_144 VPB N_A_995_47#_c_1043_n 0.00291829f $X=-0.19 $Y=1.305 $X2=0.557
+ $Y2=1.325
cc_145 VPB N_A_995_47#_c_1036_n 2.05126e-19 $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.85
cc_146 VPB N_A_995_47#_c_1037_n 0.00468357f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=0.85
cc_147 VPB N_COUT_c_1132_n 0.00610764f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_148 VPB N_COUT_c_1130_n 0.00845538f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_149 VPB N_COUT_c_1134_n 0.0326252f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_150 VPB N_VPWR_c_1148_n 0.00232309f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=1.205
cc_151 VPB N_VPWR_c_1149_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.805
cc_152 VPB N_VPWR_c_1150_n 0.00463137f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=0.72
cc_153 VPB N_VPWR_c_1151_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.625 $Y2=2.275
cc_154 VPB N_VPWR_c_1152_n 0.00276129f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_155 VPB N_VPWR_c_1153_n 0.0465801f $X=-0.19 $Y=1.305 $X2=1.105 $Y2=2.265
cc_156 VPB N_VPWR_c_1154_n 0.0050671f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.85
cc_157 VPB N_VPWR_c_1155_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1156_n 0.0377979f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.325
cc_159 VPB N_VPWR_c_1157_n 0.0153021f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=1.205
cc_160 VPB N_VPWR_c_1158_n 0.0116974f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.945
cc_161 VPB N_VPWR_c_1159_n 0.0193094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1147_n 0.0507754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1161_n 0.00353539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1162_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1163_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1164_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_382_413#_c_1264_n 0.0041398f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_168 VPB N_A_382_413#_c_1265_n 0.00291826f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.985
cc_169 VPB N_A_382_413#_c_1266_n 0.00404454f $X=-0.19 $Y=1.305 $X2=4.9 $Y2=0.445
cc_170 VPB N_A_738_413#_c_1291_n 0.00612081f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.985
cc_171 VPB N_A_738_413#_c_1292_n 0.00336306f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.985
cc_172 VPB SUM 0.00997423f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_173 VPB N_SUM_c_1325_n 0.0365457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB SUM 0.00998997f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=0.85
cc_175 N_A_76_199#_c_178_n N_A_M1020_g 0.0129484f $X=1.11 $Y=0.72 $X2=0 $Y2=0
cc_176 N_A_76_199#_c_181_n N_A_M1020_g 0.00384891f $X=0.557 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_76_199#_c_184_n N_A_M1020_g 0.00821975f $X=1.615 $Y=0.85 $X2=0 $Y2=0
cc_178 N_A_76_199#_c_186_n N_A_M1020_g 0.023207f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_76_199#_M1017_g N_A_M1011_g 0.035455f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_76_199#_c_191_n N_A_M1011_g 0.035268f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_181 N_A_76_199#_c_182_n N_A_M1001_g 0.00338905f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_182 N_A_76_199#_M1007_g N_A_M1019_g 0.0165256f $X=4.9 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A_76_199#_c_182_n N_A_M1019_g 0.00113591f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_184 N_A_76_199#_c_188_n N_A_M1019_g 7.03584e-19 $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_185 N_A_76_199#_M1010_g N_A_M1003_g 0.0451521f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_186 N_A_76_199#_c_191_n A 0.008897f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_187 N_A_76_199#_c_178_n A 0.0127285f $X=1.11 $Y=0.72 $X2=0 $Y2=0
cc_188 N_A_76_199#_c_179_n A 0.0191017f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_76_199#_c_180_n A 3.62419e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_76_199#_c_184_n A 0.00931512f $X=1.615 $Y=0.85 $X2=0 $Y2=0
cc_191 N_A_76_199#_c_182_n N_A_c_351_n 0.0499403f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_192 N_A_76_199#_c_183_n N_A_c_351_n 0.0274258f $X=1.76 $Y=0.85 $X2=0 $Y2=0
cc_193 N_A_76_199#_c_184_n N_A_c_351_n 0.00503003f $X=1.615 $Y=0.85 $X2=0 $Y2=0
cc_194 N_A_76_199#_c_191_n N_A_c_352_n 0.00111151f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_195 N_A_76_199#_c_178_n N_A_c_352_n 5.98459e-19 $X=1.11 $Y=0.72 $X2=0 $Y2=0
cc_196 N_A_76_199#_c_179_n N_A_c_352_n 0.00137149f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_76_199#_c_184_n N_A_c_352_n 0.00380863f $X=1.615 $Y=0.85 $X2=0 $Y2=0
cc_198 N_A_76_199#_c_182_n N_A_c_353_n 0.124199f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_199 N_A_76_199#_c_182_n N_A_c_354_n 0.0266325f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_200 N_A_76_199#_M1010_g N_A_c_355_n 0.00194937f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_201 N_A_76_199#_c_182_n N_A_c_355_n 0.0490684f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_202 N_A_76_199#_c_185_n N_A_c_355_n 0.0249445f $X=5.315 $Y=0.85 $X2=0 $Y2=0
cc_203 N_A_76_199#_c_187_n N_A_c_355_n 0.00189249f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_204 N_A_76_199#_c_188_n N_A_c_355_n 0.017351f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_205 N_A_76_199#_M1010_g N_A_c_356_n 4.24426e-19 $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_206 N_A_76_199#_c_182_n N_A_c_356_n 0.0260464f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_207 N_A_76_199#_c_188_n N_A_c_356_n 3.06648e-19 $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_208 N_A_76_199#_c_182_n N_A_c_357_n 0.00306165f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_209 N_A_76_199#_c_191_n N_A_c_359_n 0.00190359f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_210 N_A_76_199#_c_178_n N_A_c_359_n 0.00158237f $X=1.11 $Y=0.72 $X2=0 $Y2=0
cc_211 N_A_76_199#_c_179_n N_A_c_359_n 0.00197416f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_76_199#_c_180_n N_A_c_359_n 0.0203259f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_76_199#_c_182_n N_A_c_360_n 0.00187757f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_214 N_A_76_199#_c_182_n N_A_c_361_n 0.00347599f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_215 N_A_76_199#_c_187_n N_A_c_361_n 0.0196997f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_216 N_A_76_199#_c_188_n N_A_c_361_n 0.0011512f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_217 N_A_76_199#_c_182_n N_A_c_362_n 0.00264956f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_218 N_A_76_199#_c_187_n N_A_c_362_n 0.00313209f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_219 N_A_76_199#_c_188_n N_A_c_362_n 0.0147194f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_220 N_A_76_199#_c_188_n N_A_c_364_n 0.00414166f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_221 N_A_76_199#_c_183_n N_B_M1025_g 0.0032555f $X=1.76 $Y=0.85 $X2=0 $Y2=0
cc_222 N_A_76_199#_c_184_n N_B_M1025_g 0.0240484f $X=1.615 $Y=0.85 $X2=0 $Y2=0
cc_223 N_A_76_199#_c_191_n N_B_M1018_g 0.00392696f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_224 N_A_76_199#_c_242_p N_B_M1018_g 0.0141314f $X=1.625 $Y=2.275 $X2=0 $Y2=0
cc_225 N_A_76_199#_c_182_n N_B_c_588_n 0.0180258f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_226 N_A_76_199#_c_182_n N_B_c_589_n 0.00188483f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_227 N_A_76_199#_c_185_n N_B_M1004_g 4.321e-19 $X=5.315 $Y=0.85 $X2=0 $Y2=0
cc_228 N_A_76_199#_c_188_n N_B_M1004_g 0.00577511f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_229 N_A_76_199#_c_191_n B 0.02463f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_230 N_A_76_199#_c_242_p B 0.0250439f $X=1.625 $Y=2.275 $X2=0 $Y2=0
cc_231 N_A_76_199#_c_184_n B 0.00628162f $X=1.615 $Y=0.85 $X2=0 $Y2=0
cc_232 N_A_76_199#_c_242_p N_B_c_606_n 0.00152729f $X=1.625 $Y=2.275 $X2=0 $Y2=0
cc_233 N_A_76_199#_M1010_g N_B_c_607_n 0.00179768f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_234 N_A_76_199#_c_187_n N_B_c_607_n 5.89663e-19 $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_235 N_A_76_199#_c_188_n N_B_c_607_n 0.00309513f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_236 N_A_76_199#_c_191_n N_B_c_613_n 0.00169219f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_237 N_A_76_199#_c_242_p N_B_c_613_n 0.00247661f $X=1.625 $Y=2.275 $X2=0 $Y2=0
cc_238 N_A_76_199#_c_182_n N_CIN_M1023_g 0.00462124f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_239 N_A_76_199#_c_183_n N_CIN_M1023_g 0.0024037f $X=1.76 $Y=0.85 $X2=0 $Y2=0
cc_240 N_A_76_199#_c_184_n N_CIN_M1023_g 0.00443973f $X=1.615 $Y=0.85 $X2=0
+ $Y2=0
cc_241 N_A_76_199#_M1007_g N_CIN_M1002_g 0.015353f $X=4.9 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_76_199#_M1010_g N_CIN_M1002_g 0.0132203f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_243 N_A_76_199#_c_185_n N_CIN_M1002_g 0.00147214f $X=5.315 $Y=0.85 $X2=0
+ $Y2=0
cc_244 N_A_76_199#_c_187_n N_CIN_M1002_g 0.0217272f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_245 N_A_76_199#_c_188_n N_CIN_M1002_g 0.0136455f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_246 N_A_76_199#_M1010_g N_CIN_M1021_g 0.0149126f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_247 N_A_76_199#_c_182_n N_CIN_c_812_n 0.00117889f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_248 N_A_76_199#_c_182_n N_CIN_c_815_n 0.0209196f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_249 N_A_76_199#_c_182_n N_CIN_c_816_n 0.00158362f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_250 N_A_76_199#_M1010_g N_CIN_c_830_n 0.0144105f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_251 N_A_76_199#_c_187_n N_CIN_c_830_n 0.00169335f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_252 N_A_76_199#_c_188_n N_CIN_c_830_n 0.00955271f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_253 N_A_76_199#_c_182_n N_CIN_c_818_n 9.52651e-19 $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_254 N_A_76_199#_c_183_n N_CIN_c_818_n 9.74524e-19 $X=1.76 $Y=0.85 $X2=0 $Y2=0
cc_255 N_A_76_199#_c_184_n N_CIN_c_818_n 2.46291e-19 $X=1.615 $Y=0.85 $X2=0
+ $Y2=0
cc_256 N_A_76_199#_c_182_n N_CIN_c_819_n 0.00500146f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_257 N_A_76_199#_c_183_n N_CIN_c_819_n 0.0013906f $X=1.76 $Y=0.85 $X2=0 $Y2=0
cc_258 N_A_76_199#_c_184_n N_CIN_c_819_n 0.00266523f $X=1.615 $Y=0.85 $X2=0
+ $Y2=0
cc_259 N_A_76_199#_c_182_n N_CIN_c_820_n 0.00189437f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_260 N_A_76_199#_M1010_g N_CIN_c_835_n 0.0204361f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_261 N_A_76_199#_c_188_n N_CIN_c_835_n 6.09232e-19 $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_262 N_A_76_199#_M1010_g N_CIN_c_836_n 0.00575383f $X=4.9 $Y=2.275 $X2=0 $Y2=0
cc_263 N_A_76_199#_c_188_n N_CIN_c_836_n 0.00657808f $X=4.96 $Y=1.04 $X2=0 $Y2=0
cc_264 N_A_76_199#_c_185_n N_A_995_47#_c_1034_n 0.00325379f $X=5.315 $Y=0.85
+ $X2=0 $Y2=0
cc_265 N_A_76_199#_c_188_n N_A_995_47#_c_1034_n 0.00750162f $X=4.96 $Y=1.04
+ $X2=0 $Y2=0
cc_266 N_A_76_199#_c_182_n N_A_995_47#_c_1048_n 4.08874e-19 $X=5.17 $Y=0.85
+ $X2=0 $Y2=0
cc_267 N_A_76_199#_c_185_n N_A_995_47#_c_1048_n 0.00101125f $X=5.315 $Y=0.85
+ $X2=0 $Y2=0
cc_268 N_A_76_199#_c_188_n N_A_995_47#_c_1048_n 0.0118074f $X=4.96 $Y=1.04 $X2=0
+ $Y2=0
cc_269 N_A_76_199#_M1017_g N_COUT_c_1130_n 0.00333486f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_270 N_A_76_199#_c_191_n N_COUT_c_1130_n 0.00842515f $X=0.6 $Y=1.625 $X2=0
+ $Y2=0
cc_271 N_A_76_199#_c_179_n N_COUT_c_1130_n 0.0243753f $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_76_199#_c_180_n N_COUT_c_1130_n 0.00753785f $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_76_199#_c_181_n N_COUT_c_1130_n 0.00861302f $X=0.557 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_76_199#_c_186_n N_COUT_c_1130_n 0.00343973f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_76_199#_c_191_n N_VPWR_M1017_d 0.00967615f $X=0.6 $Y=1.625 $X2=-0.19
+ $Y2=-0.24
cc_276 N_A_76_199#_M1017_g N_VPWR_c_1148_n 0.0093716f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_277 N_A_76_199#_c_191_n N_VPWR_c_1148_n 0.039151f $X=0.6 $Y=1.625 $X2=0 $Y2=0
cc_278 N_A_76_199#_M1010_g N_VPWR_c_1151_n 0.00114511f $X=4.9 $Y=2.275 $X2=0
+ $Y2=0
cc_279 N_A_76_199#_M1010_g N_VPWR_c_1153_n 0.00585385f $X=4.9 $Y=2.275 $X2=0
+ $Y2=0
cc_280 N_A_76_199#_M1017_g N_VPWR_c_1155_n 0.0046653f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A_76_199#_c_191_n N_VPWR_c_1156_n 0.00974389f $X=0.6 $Y=1.625 $X2=0
+ $Y2=0
cc_282 N_A_76_199#_c_242_p N_VPWR_c_1156_n 0.0364401f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_283 N_A_76_199#_M1018_d N_VPWR_c_1147_n 0.00390407f $X=1.49 $Y=2.065 $X2=0
+ $Y2=0
cc_284 N_A_76_199#_M1017_g N_VPWR_c_1147_n 0.00895857f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_285 N_A_76_199#_M1010_g N_VPWR_c_1147_n 0.0109946f $X=4.9 $Y=2.275 $X2=0
+ $Y2=0
cc_286 N_A_76_199#_c_191_n N_VPWR_c_1147_n 0.0133726f $X=0.6 $Y=1.625 $X2=0
+ $Y2=0
cc_287 N_A_76_199#_c_242_p N_VPWR_c_1147_n 0.022276f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_288 N_A_76_199#_c_242_p A_208_413# 0.00822779f $X=1.625 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_289 N_A_76_199#_M1010_g N_A_738_413#_c_1291_n 0.00479826f $X=4.9 $Y=2.275
+ $X2=0 $Y2=0
cc_290 N_A_76_199#_c_178_n N_VGND_M1024_d 0.00604386f $X=1.11 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_291 N_A_76_199#_c_309_p N_VGND_M1024_d 8.83574e-19 $X=0.685 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_292 N_A_76_199#_c_181_n N_VGND_M1024_d 9.39224e-19 $X=0.557 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_293 N_A_76_199#_c_178_n N_VGND_c_1337_n 0.0112591f $X=1.11 $Y=0.72 $X2=0
+ $Y2=0
cc_294 N_A_76_199#_c_309_p N_VGND_c_1337_n 0.00924733f $X=0.685 $Y=0.72 $X2=0
+ $Y2=0
cc_295 N_A_76_199#_c_180_n N_VGND_c_1337_n 2.98237e-19 $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_296 N_A_76_199#_c_186_n N_VGND_c_1337_n 0.00837852f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_76_199#_c_182_n N_VGND_c_1338_n 0.00115864f $X=5.17 $Y=0.85 $X2=0
+ $Y2=0
cc_298 N_A_76_199#_c_182_n N_VGND_c_1339_n 0.00407154f $X=5.17 $Y=0.85 $X2=0
+ $Y2=0
cc_299 N_A_76_199#_M1007_g N_VGND_c_1340_n 0.00114511f $X=4.9 $Y=0.445 $X2=0
+ $Y2=0
cc_300 N_A_76_199#_c_182_n N_VGND_c_1340_n 0.00115864f $X=5.17 $Y=0.85 $X2=0
+ $Y2=0
cc_301 N_A_76_199#_M1007_g N_VGND_c_1342_n 0.00585385f $X=4.9 $Y=0.445 $X2=0
+ $Y2=0
cc_302 N_A_76_199#_c_186_n N_VGND_c_1344_n 0.0046653f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_76_199#_c_178_n N_VGND_c_1345_n 0.00366264f $X=1.11 $Y=0.72 $X2=0
+ $Y2=0
cc_304 N_A_76_199#_c_184_n N_VGND_c_1345_n 0.0373012f $X=1.615 $Y=0.85 $X2=0
+ $Y2=0
cc_305 N_A_76_199#_M1025_d N_VGND_c_1349_n 0.00208923f $X=1.49 $Y=0.235 $X2=0
+ $Y2=0
cc_306 N_A_76_199#_M1007_g N_VGND_c_1349_n 0.00660978f $X=4.9 $Y=0.445 $X2=0
+ $Y2=0
cc_307 N_A_76_199#_c_178_n N_VGND_c_1349_n 0.00745304f $X=1.11 $Y=0.72 $X2=0
+ $Y2=0
cc_308 N_A_76_199#_c_309_p N_VGND_c_1349_n 8.3983e-19 $X=0.685 $Y=0.72 $X2=0
+ $Y2=0
cc_309 N_A_76_199#_c_182_n N_VGND_c_1349_n 0.156698f $X=5.17 $Y=0.85 $X2=0 $Y2=0
cc_310 N_A_76_199#_c_183_n N_VGND_c_1349_n 0.0149056f $X=1.76 $Y=0.85 $X2=0
+ $Y2=0
cc_311 N_A_76_199#_c_184_n N_VGND_c_1349_n 0.0173394f $X=1.615 $Y=0.85 $X2=0
+ $Y2=0
cc_312 N_A_76_199#_c_185_n N_VGND_c_1349_n 0.0156759f $X=5.315 $Y=0.85 $X2=0
+ $Y2=0
cc_313 N_A_76_199#_c_186_n N_VGND_c_1349_n 0.00895857f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_76_199#_c_188_n N_VGND_c_1349_n 0.00304902f $X=4.96 $Y=1.04 $X2=0
+ $Y2=0
cc_315 N_A_76_199#_c_178_n A_208_47# 2.09292e-19 $X=1.11 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_316 N_A_76_199#_c_184_n A_208_47# 0.00654395f $X=1.615 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_317 N_A_76_199#_c_182_n N_A_382_47#_c_1467_n 0.0271275f $X=5.17 $Y=0.85 $X2=0
+ $Y2=0
cc_318 N_A_76_199#_c_182_n N_A_382_47#_c_1468_n 0.00797006f $X=5.17 $Y=0.85
+ $X2=0 $Y2=0
cc_319 N_A_76_199#_c_183_n N_A_382_47#_c_1468_n 0.00117968f $X=1.76 $Y=0.85
+ $X2=0 $Y2=0
cc_320 N_A_76_199#_c_184_n N_A_382_47#_c_1468_n 0.0081472f $X=1.615 $Y=0.85
+ $X2=0 $Y2=0
cc_321 N_A_76_199#_M1007_g N_A_738_47#_c_1502_n 0.00472067f $X=4.9 $Y=0.445
+ $X2=0 $Y2=0
cc_322 N_A_76_199#_c_182_n N_A_738_47#_c_1502_n 0.0297995f $X=5.17 $Y=0.85 $X2=0
+ $Y2=0
cc_323 N_A_76_199#_c_185_n N_A_738_47#_c_1502_n 0.00140299f $X=5.315 $Y=0.85
+ $X2=0 $Y2=0
cc_324 N_A_76_199#_c_188_n N_A_738_47#_c_1502_n 0.00128001f $X=4.96 $Y=1.04
+ $X2=0 $Y2=0
cc_325 N_A_76_199#_c_182_n N_A_738_47#_c_1503_n 0.00610445f $X=5.17 $Y=0.85
+ $X2=0 $Y2=0
cc_326 N_A_M1020_g N_B_M1025_g 0.035483f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_327 N_A_M1011_g N_B_M1025_g 0.00918325f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_328 A N_B_M1025_g 0.00432518f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_329 N_A_c_351_n N_B_M1025_g 0.00510287f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_330 N_A_c_352_n N_B_M1025_g 0.00145512f $X=1.3 $Y=1.19 $X2=0 $Y2=0
cc_331 N_A_c_359_n N_B_M1025_g 0.0207319f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_M1011_g N_B_M1018_g 0.0303588f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_333 N_A_M1001_g N_B_c_587_n 0.0218633f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_334 N_A_c_353_n N_B_c_589_n 5.6387e-19 $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_335 N_A_c_354_n N_B_c_589_n 3.21623e-19 $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_336 N_A_c_357_n N_B_c_589_n 4.12248e-19 $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_337 N_A_M1009_g N_B_c_597_n 0.0224258f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_338 N_A_M1013_g N_B_M1004_g 0.0289497f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_339 N_A_M1015_g N_B_M1004_g 0.0086241f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_340 N_A_c_355_n N_B_M1004_g 0.00521518f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_341 N_A_c_358_n N_B_M1004_g 3.42408e-19 $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_342 N_A_c_363_n N_B_M1004_g 0.0210546f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_343 N_A_c_364_n N_B_M1004_g 0.0041572f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_344 N_A_M1015_g N_B_M1027_g 0.0283902f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_345 N_A_c_353_n N_B_c_591_n 0.00134601f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_346 N_A_M1011_g B 0.00155484f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_347 N_A_c_351_n B 0.00571869f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_348 N_A_M1009_g N_B_c_605_n 0.00432516f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_349 N_A_c_351_n N_B_c_605_n 0.0492154f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_350 N_A_c_353_n N_B_c_605_n 0.0518715f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_351 N_A_c_354_n N_B_c_605_n 0.0266284f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_352 N_A_c_357_n N_B_c_605_n 0.00305499f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_353 N_A_c_360_n N_B_c_605_n 0.00189048f $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_354 N_A_c_351_n N_B_c_606_n 0.0274262f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_355 N_A_M1003_g N_B_c_607_n 0.00147004f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_356 N_A_c_353_n N_B_c_607_n 0.0504198f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_357 N_A_c_355_n N_B_c_607_n 0.0897573f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_358 N_A_c_356_n N_B_c_607_n 0.0275368f $X=4.54 $Y=1.19 $X2=0 $Y2=0
cc_359 N_A_c_362_n N_B_c_607_n 0.00173442f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_360 N_A_c_353_n N_B_c_608_n 0.0275518f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_361 N_A_c_353_n N_B_c_609_n 0.00183472f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_362 N_A_M1015_g N_B_c_610_n 4.49035e-19 $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_363 N_A_c_355_n N_B_c_610_n 0.0274019f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_364 N_A_c_364_n N_B_c_610_n 2.20027e-19 $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_365 N_A_M1015_g N_B_c_611_n 0.00341368f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_366 N_A_c_355_n N_B_c_611_n 0.00406245f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_367 N_A_c_363_n N_B_c_611_n 6.68519e-19 $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_368 N_A_c_364_n N_B_c_611_n 0.0121738f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_369 N_A_M1011_g N_B_c_613_n 0.0201434f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_370 N_A_c_352_n N_B_c_613_n 0.00123766f $X=1.3 $Y=1.19 $X2=0 $Y2=0
cc_371 N_A_M1015_g N_B_c_614_n 0.0199227f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_372 N_A_c_364_n N_B_c_614_n 3.00025e-19 $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_373 N_A_M1001_g N_CIN_M1023_g 0.0261054f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_374 N_A_c_360_n N_CIN_M1012_g 0.0412054f $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_375 N_A_M1003_g N_CIN_M1008_g 0.0256653f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_376 N_A_c_355_n N_CIN_M1002_g 0.00283992f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_377 N_A_M1019_g N_CIN_c_811_n 0.0141455f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_378 N_A_M1019_g N_CIN_c_812_n 0.00744646f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_379 N_A_c_361_n N_CIN_c_812_n 0.0209196f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_380 N_A_c_351_n N_CIN_c_813_n 6.23037e-19 $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_381 N_A_c_352_n N_CIN_c_813_n 9.00939e-19 $X=1.3 $Y=1.19 $X2=0 $Y2=0
cc_382 N_A_c_357_n N_CIN_c_813_n 0.00575336f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_383 N_A_c_360_n N_CIN_c_813_n 0.00493779f $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_384 N_A_M1009_g N_CIN_c_826_n 0.0124584f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_385 N_A_c_351_n N_CIN_c_826_n 0.00156522f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_386 N_A_c_353_n N_CIN_c_826_n 5.93941e-19 $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_387 N_A_c_354_n N_CIN_c_826_n 5.3606e-19 $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_388 N_A_c_357_n N_CIN_c_826_n 0.0178288f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_389 N_A_c_360_n N_CIN_c_826_n 0.0024982f $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_390 N_A_M1009_g N_CIN_c_814_n 0.00469718f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_391 N_A_c_353_n N_CIN_c_814_n 0.00319513f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_392 N_A_c_354_n N_CIN_c_814_n 0.00137624f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_393 N_A_c_357_n N_CIN_c_814_n 0.00802988f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_394 N_A_c_360_n N_CIN_c_814_n 5.0579e-19 $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_395 N_A_c_353_n N_CIN_c_815_n 0.0361711f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_396 N_A_c_356_n N_CIN_c_815_n 0.00124935f $X=4.54 $Y=1.19 $X2=0 $Y2=0
cc_397 N_A_c_362_n N_CIN_c_815_n 0.0141315f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_398 N_A_M1001_g N_CIN_c_816_n 0.00195651f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_399 N_A_c_353_n N_CIN_c_816_n 0.00560548f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_400 N_A_c_354_n N_CIN_c_816_n 0.00142282f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_401 N_A_c_357_n N_CIN_c_816_n 0.0168914f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_402 N_A_c_360_n N_CIN_c_816_n 0.0010498f $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_403 N_A_M1003_g N_CIN_c_817_n 4.71687e-19 $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_404 N_A_c_353_n N_CIN_c_817_n 0.0032466f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_405 N_A_c_356_n N_CIN_c_817_n 0.00169222f $X=4.54 $Y=1.19 $X2=0 $Y2=0
cc_406 N_A_c_362_n N_CIN_c_817_n 9.71923e-19 $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_407 N_A_M1003_g N_CIN_c_830_n 0.0100247f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_408 N_A_c_353_n N_CIN_c_830_n 0.00331122f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_409 N_A_c_355_n N_CIN_c_830_n 0.00270801f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_410 N_A_c_356_n N_CIN_c_830_n 0.00108059f $X=4.54 $Y=1.19 $X2=0 $Y2=0
cc_411 N_A_c_361_n N_CIN_c_830_n 5.94361e-19 $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_412 N_A_c_362_n N_CIN_c_830_n 0.0178134f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_413 N_A_M1003_g N_CIN_c_832_n 0.021979f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_414 N_A_c_353_n N_CIN_c_832_n 9.61162e-19 $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_415 N_A_M1001_g N_CIN_c_818_n 0.0215001f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_416 N_A_c_357_n N_CIN_c_818_n 7.99315e-19 $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_417 A N_CIN_c_819_n 0.00465896f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_418 N_A_c_351_n N_CIN_c_819_n 0.0145708f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_419 N_A_c_352_n N_CIN_c_819_n 7.45527e-19 $X=1.3 $Y=1.19 $X2=0 $Y2=0
cc_420 N_A_c_357_n N_CIN_c_819_n 0.0106105f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_421 N_A_c_360_n N_CIN_c_819_n 8.25882e-19 $X=2.315 $Y=1.195 $X2=0 $Y2=0
cc_422 N_A_M1003_g N_CIN_c_820_n 0.0112529f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_423 N_A_c_353_n N_CIN_c_820_n 0.0041373f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_424 N_A_c_356_n N_CIN_c_820_n 0.00137864f $X=4.54 $Y=1.19 $X2=0 $Y2=0
cc_425 N_A_c_362_n N_CIN_c_820_n 0.00226131f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_426 N_A_c_355_n N_CIN_c_836_n 0.00134396f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_427 N_A_M1015_g N_A_995_47#_M1006_g 0.0357912f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_428 N_A_M1015_g N_A_995_47#_c_1052_n 4.38095e-19 $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_429 N_A_M1013_g N_A_995_47#_c_1034_n 4.0244e-19 $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_430 N_A_c_355_n N_A_995_47#_c_1034_n 0.0135777f $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_431 N_A_c_363_n N_A_995_47#_c_1034_n 0.00167625f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_432 N_A_c_364_n N_A_995_47#_c_1034_n 0.0103824f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_433 N_A_M1013_g N_A_995_47#_c_1035_n 0.0111548f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_434 N_A_c_358_n N_A_995_47#_c_1035_n 0.00376691f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_435 N_A_c_363_n N_A_995_47#_c_1035_n 0.00116721f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_436 N_A_c_364_n N_A_995_47#_c_1035_n 0.010611f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_437 N_A_M1015_g N_A_995_47#_c_1041_n 0.0111631f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_438 N_A_c_364_n N_A_995_47#_c_1041_n 0.00256722f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_439 N_A_M1015_g N_A_995_47#_c_1042_n 0.00486613f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_440 N_A_M1015_g N_A_995_47#_c_1043_n 0.0116261f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_441 N_A_c_363_n N_A_995_47#_c_1043_n 0.00120219f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_442 N_A_c_364_n N_A_995_47#_c_1043_n 0.00265067f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_443 N_A_c_358_n N_A_995_47#_c_1036_n 0.00844193f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_444 N_A_c_363_n N_A_995_47#_c_1036_n 0.00815335f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_445 N_A_c_364_n N_A_995_47#_c_1036_n 0.0168513f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_446 N_A_c_363_n N_A_995_47#_c_1037_n 0.019446f $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_447 N_A_c_364_n N_A_995_47#_c_1037_n 6.32783e-19 $X=6.16 $Y=1.12 $X2=0 $Y2=0
cc_448 N_A_M1013_g N_A_995_47#_c_1038_n 0.00258793f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_449 N_A_M1013_g N_A_995_47#_c_1039_n 0.0235984f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_450 N_A_M1011_g N_VPWR_c_1148_n 0.00514543f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_451 N_A_M1009_g N_VPWR_c_1149_n 0.00759908f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_452 N_A_M1003_g N_VPWR_c_1151_n 0.00761262f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_453 N_A_M1015_g N_VPWR_c_1152_n 0.00409489f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_454 N_A_M1003_g N_VPWR_c_1153_n 0.00337001f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_455 N_A_M1015_g N_VPWR_c_1153_n 0.0041289f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_456 N_A_M1011_g N_VPWR_c_1156_n 0.00425983f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_457 N_A_M1009_g N_VPWR_c_1156_n 0.00337001f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_458 N_A_M1011_g N_VPWR_c_1147_n 0.0058625f $X=0.965 $Y=2.275 $X2=0 $Y2=0
cc_459 N_A_M1009_g N_VPWR_c_1147_n 0.00397658f $X=2.255 $Y=2.275 $X2=0 $Y2=0
cc_460 N_A_M1003_g N_VPWR_c_1147_n 0.00403935f $X=4.455 $Y=2.275 $X2=0 $Y2=0
cc_461 N_A_M1015_g N_VPWR_c_1147_n 0.00597277f $X=6.22 $Y=2.275 $X2=0 $Y2=0
cc_462 N_A_M1009_g N_A_382_413#_c_1264_n 0.0105731f $X=2.255 $Y=2.275 $X2=0
+ $Y2=0
cc_463 N_A_M1003_g N_A_738_413#_c_1291_n 0.0111197f $X=4.455 $Y=2.275 $X2=0
+ $Y2=0
cc_464 N_A_M1020_g N_VGND_c_1337_n 0.00419788f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_465 N_A_M1001_g N_VGND_c_1338_n 0.00760016f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_466 N_A_M1019_g N_VGND_c_1340_n 0.00760591f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_467 N_A_M1013_g N_VGND_c_1341_n 0.00769722f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_468 N_A_M1019_g N_VGND_c_1342_n 0.00337001f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_469 N_A_M1013_g N_VGND_c_1342_n 0.00337001f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_470 N_A_M1020_g N_VGND_c_1345_n 0.00425094f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_471 N_A_M1001_g N_VGND_c_1345_n 0.00337001f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_472 N_A_M1020_g N_VGND_c_1349_n 0.006053f $X=0.965 $Y=0.445 $X2=0 $Y2=0
cc_473 N_A_M1001_g N_VGND_c_1349_n 0.00377406f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_474 N_A_M1019_g N_VGND_c_1349_n 0.00383683f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_475 N_A_M1013_g N_VGND_c_1349_n 0.00412258f $X=6.22 $Y=0.445 $X2=0 $Y2=0
cc_476 N_A_M1001_g N_A_382_47#_c_1467_n 0.0108136f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_477 N_A_c_351_n N_A_382_47#_c_1467_n 0.00108134f $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_478 N_A_c_353_n N_A_382_47#_c_1467_n 0.00161385f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_479 N_A_c_354_n N_A_382_47#_c_1467_n 9.66928e-19 $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_480 N_A_c_357_n N_A_382_47#_c_1467_n 0.0169746f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_481 N_A_c_360_n N_A_382_47#_c_1467_n 0.00247695f $X=2.315 $Y=1.195 $X2=0
+ $Y2=0
cc_482 N_A_c_351_n N_A_382_47#_c_1468_n 5.45312e-19 $X=2.39 $Y=1.19 $X2=0 $Y2=0
cc_483 N_A_M1019_g N_A_738_47#_c_1502_n 0.00973522f $X=4.455 $Y=0.445 $X2=0
+ $Y2=0
cc_484 N_A_c_353_n N_A_738_47#_c_1502_n 0.0025772f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_485 N_A_c_355_n N_A_738_47#_c_1502_n 7.16872e-19 $X=6.09 $Y=1.19 $X2=0 $Y2=0
cc_486 N_A_c_356_n N_A_738_47#_c_1502_n 3.2424e-19 $X=4.54 $Y=1.19 $X2=0 $Y2=0
cc_487 N_A_c_361_n N_A_738_47#_c_1502_n 0.00230741f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_488 N_A_c_362_n N_A_738_47#_c_1502_n 0.0240755f $X=4.46 $Y=1.04 $X2=0 $Y2=0
cc_489 N_B_M1025_g N_CIN_M1023_g 0.0261105f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_490 N_B_M1025_g N_CIN_M1012_g 0.00958021f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_491 N_B_M1018_g N_CIN_M1012_g 0.0167915f $X=1.415 $Y=2.275 $X2=0 $Y2=0
cc_492 B N_CIN_M1012_g 0.0051403f $X=1.53 $Y=1.445 $X2=0 $Y2=0
cc_493 N_B_c_605_n N_CIN_M1012_g 0.00515121f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_494 N_B_c_606_n N_CIN_M1012_g 0.0023625f $X=1.76 $Y=1.53 $X2=0 $Y2=0
cc_495 N_B_c_613_n N_CIN_M1012_g 0.0170014f $X=1.385 $Y=1.715 $X2=0 $Y2=0
cc_496 N_B_c_603_n N_CIN_M1008_g 0.0194852f $X=3.502 $Y=1.915 $X2=0 $Y2=0
cc_497 N_B_c_612_n N_CIN_M1008_g 0.00348516f $X=3.45 $Y=1.6 $X2=0 $Y2=0
cc_498 N_B_M1004_g N_CIN_M1002_g 0.0534949f $X=5.74 $Y=0.445 $X2=0 $Y2=0
cc_499 N_B_c_607_n N_CIN_M1002_g 0.00168706f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_500 N_B_c_610_n N_CIN_M1002_g 6.61635e-19 $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_501 N_B_c_611_n N_CIN_M1002_g 0.00259458f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_502 N_B_M1027_g N_CIN_M1021_g 0.0534949f $X=5.74 $Y=2.275 $X2=0 $Y2=0
cc_503 N_B_c_592_n N_CIN_c_811_n 0.00946436f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_504 N_B_c_588_n N_CIN_c_812_n 0.00946436f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_505 N_B_M1025_g N_CIN_c_813_n 9.20834e-19 $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_506 B N_CIN_c_813_n 0.0101863f $X=1.53 $Y=1.445 $X2=0 $Y2=0
cc_507 N_B_c_605_n N_CIN_c_813_n 0.0101343f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_508 N_B_c_606_n N_CIN_c_813_n 0.00173655f $X=1.76 $Y=1.53 $X2=0 $Y2=0
cc_509 N_B_c_596_n N_CIN_c_826_n 0.00421109f $X=3.315 $Y=1.915 $X2=0 $Y2=0
cc_510 N_B_c_597_n N_CIN_c_826_n 0.00556877f $X=2.75 $Y=1.915 $X2=0 $Y2=0
cc_511 N_B_c_605_n N_CIN_c_826_n 0.0247638f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_512 N_B_c_608_n N_CIN_c_826_n 2.87707e-19 $X=3.62 $Y=1.53 $X2=0 $Y2=0
cc_513 N_B_c_609_n N_CIN_c_826_n 0.0114491f $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_514 N_B_c_612_n N_CIN_c_826_n 0.00100465f $X=3.45 $Y=1.6 $X2=0 $Y2=0
cc_515 B N_CIN_c_827_n 0.0137791f $X=1.53 $Y=1.445 $X2=0 $Y2=0
cc_516 N_B_c_605_n N_CIN_c_827_n 0.00525602f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_517 N_B_c_606_n N_CIN_c_827_n 0.00122285f $X=1.76 $Y=1.53 $X2=0 $Y2=0
cc_518 N_B_c_601_n N_CIN_c_814_n 7.30597e-19 $X=3.475 $Y=1.595 $X2=0 $Y2=0
cc_519 N_B_c_591_n N_CIN_c_814_n 0.00417439f $X=3.475 $Y=1.435 $X2=0 $Y2=0
cc_520 N_B_c_605_n N_CIN_c_814_n 0.0115031f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_521 N_B_c_608_n N_CIN_c_814_n 9.40906e-19 $X=3.62 $Y=1.53 $X2=0 $Y2=0
cc_522 N_B_c_609_n N_CIN_c_814_n 0.00826368f $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_523 N_B_c_588_n N_CIN_c_815_n 0.0170405f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_524 N_B_c_596_n N_CIN_c_815_n 0.00437579f $X=3.315 $Y=1.915 $X2=0 $Y2=0
cc_525 N_B_c_601_n N_CIN_c_815_n 5.9469e-19 $X=3.475 $Y=1.595 $X2=0 $Y2=0
cc_526 N_B_c_591_n N_CIN_c_815_n 0.0193458f $X=3.475 $Y=1.435 $X2=0 $Y2=0
cc_527 N_B_c_603_n N_CIN_c_815_n 0.00124084f $X=3.502 $Y=1.915 $X2=0 $Y2=0
cc_528 N_B_c_605_n N_CIN_c_815_n 0.00184797f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_529 N_B_c_607_n N_CIN_c_815_n 0.00127868f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_530 N_B_c_608_n N_CIN_c_815_n 0.00181285f $X=3.62 $Y=1.53 $X2=0 $Y2=0
cc_531 N_B_c_609_n N_CIN_c_815_n 0.022414f $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_532 N_B_c_588_n N_CIN_c_816_n 0.00347447f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_533 N_B_c_591_n N_CIN_c_817_n 0.0044194f $X=3.475 $Y=1.435 $X2=0 $Y2=0
cc_534 N_B_c_607_n N_CIN_c_817_n 0.00577857f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_535 N_B_c_608_n N_CIN_c_817_n 0.00152525f $X=3.62 $Y=1.53 $X2=0 $Y2=0
cc_536 N_B_c_609_n N_CIN_c_817_n 0.00391111f $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_537 N_B_c_607_n N_CIN_c_830_n 0.0508593f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_538 N_B_c_601_n N_CIN_c_831_n 0.00116908f $X=3.475 $Y=1.595 $X2=0 $Y2=0
cc_539 N_B_c_607_n N_CIN_c_831_n 0.00496173f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_540 N_B_c_608_n N_CIN_c_831_n 0.00121328f $X=3.62 $Y=1.53 $X2=0 $Y2=0
cc_541 N_B_c_609_n N_CIN_c_831_n 0.00949903f $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_542 N_B_c_601_n N_CIN_c_832_n 0.0164961f $X=3.475 $Y=1.595 $X2=0 $Y2=0
cc_543 N_B_c_607_n N_CIN_c_832_n 0.00208441f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_544 N_B_c_609_n N_CIN_c_832_n 8.17579e-19 $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_545 N_B_M1025_g N_CIN_c_818_n 0.0214502f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_546 N_B_c_606_n N_CIN_c_818_n 9.74524e-19 $X=1.76 $Y=1.53 $X2=0 $Y2=0
cc_547 N_B_M1025_g N_CIN_c_819_n 0.00110487f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_548 B N_CIN_c_819_n 0.00199359f $X=1.53 $Y=1.445 $X2=0 $Y2=0
cc_549 N_B_c_605_n N_CIN_c_819_n 0.0025168f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_550 N_B_c_606_n N_CIN_c_819_n 0.00156579f $X=1.76 $Y=1.53 $X2=0 $Y2=0
cc_551 N_B_c_588_n N_CIN_c_820_n 0.00388837f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_552 N_B_c_591_n N_CIN_c_820_n 0.0156686f $X=3.475 $Y=1.435 $X2=0 $Y2=0
cc_553 N_B_c_607_n N_CIN_c_835_n 0.00218391f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_554 N_B_c_610_n N_CIN_c_835_n 6.76137e-19 $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_555 N_B_c_614_n N_CIN_c_835_n 0.0534949f $X=5.8 $Y=1.68 $X2=0 $Y2=0
cc_556 N_B_c_607_n N_CIN_c_836_n 0.00989817f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_557 N_B_c_610_n N_CIN_c_836_n 0.00123607f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_558 N_B_c_611_n N_CIN_c_836_n 0.0139966f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_559 N_B_c_614_n N_CIN_c_836_n 0.00142939f $X=5.8 $Y=1.68 $X2=0 $Y2=0
cc_560 N_B_M1027_g N_A_995_47#_c_1052_n 0.0153915f $X=5.74 $Y=2.275 $X2=0 $Y2=0
cc_561 N_B_c_607_n N_A_995_47#_c_1052_n 0.00888491f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_562 N_B_c_610_n N_A_995_47#_c_1052_n 0.00185453f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_563 N_B_c_611_n N_A_995_47#_c_1052_n 0.0127074f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_564 N_B_c_614_n N_A_995_47#_c_1052_n 0.00241517f $X=5.8 $Y=1.68 $X2=0 $Y2=0
cc_565 N_B_M1004_g N_A_995_47#_c_1034_n 0.0183218f $X=5.74 $Y=0.445 $X2=0 $Y2=0
cc_566 N_B_c_610_n N_A_995_47#_c_1042_n 0.00206268f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_567 N_B_c_611_n N_A_995_47#_c_1042_n 0.0117542f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_568 N_B_M1027_g N_A_995_47#_c_1043_n 0.00412533f $X=5.74 $Y=2.275 $X2=0 $Y2=0
cc_569 N_B_c_611_n N_A_995_47#_c_1043_n 0.00460861f $X=5.775 $Y=1.53 $X2=0 $Y2=0
cc_570 N_B_c_595_n N_VPWR_c_1149_n 0.00677587f $X=2.675 $Y=1.99 $X2=0 $Y2=0
cc_571 N_B_c_595_n N_VPWR_c_1150_n 0.00192382f $X=2.675 $Y=1.99 $X2=0 $Y2=0
cc_572 N_B_c_596_n N_VPWR_c_1150_n 0.00517219f $X=3.315 $Y=1.915 $X2=0 $Y2=0
cc_573 N_B_c_598_n N_VPWR_c_1150_n 0.00808089f $X=3.615 $Y=1.99 $X2=0 $Y2=0
cc_574 N_B_c_608_n N_VPWR_c_1150_n 0.00172657f $X=3.62 $Y=1.53 $X2=0 $Y2=0
cc_575 N_B_c_609_n N_VPWR_c_1150_n 0.00938786f $X=3.475 $Y=1.53 $X2=0 $Y2=0
cc_576 N_B_c_598_n N_VPWR_c_1151_n 5.31689e-19 $X=3.615 $Y=1.99 $X2=0 $Y2=0
cc_577 N_B_M1027_g N_VPWR_c_1153_n 0.00357877f $X=5.74 $Y=2.275 $X2=0 $Y2=0
cc_578 N_B_M1018_g N_VPWR_c_1156_n 0.00357877f $X=1.415 $Y=2.275 $X2=0 $Y2=0
cc_579 N_B_c_595_n N_VPWR_c_1157_n 0.00337001f $X=2.675 $Y=1.99 $X2=0 $Y2=0
cc_580 N_B_c_596_n N_VPWR_c_1157_n 0.00378947f $X=3.315 $Y=1.915 $X2=0 $Y2=0
cc_581 N_B_c_598_n N_VPWR_c_1158_n 0.0046653f $X=3.615 $Y=1.99 $X2=0 $Y2=0
cc_582 N_B_M1018_g N_VPWR_c_1147_n 0.00539554f $X=1.415 $Y=2.275 $X2=0 $Y2=0
cc_583 N_B_c_595_n N_VPWR_c_1147_n 0.0053254f $X=2.675 $Y=1.99 $X2=0 $Y2=0
cc_584 N_B_c_596_n N_VPWR_c_1147_n 0.00445861f $X=3.315 $Y=1.915 $X2=0 $Y2=0
cc_585 N_B_c_598_n N_VPWR_c_1147_n 0.00799591f $X=3.615 $Y=1.99 $X2=0 $Y2=0
cc_586 N_B_M1027_g N_VPWR_c_1147_n 0.00530375f $X=5.74 $Y=2.275 $X2=0 $Y2=0
cc_587 N_B_c_595_n N_A_382_413#_c_1264_n 0.00768486f $X=2.675 $Y=1.99 $X2=0
+ $Y2=0
cc_588 N_B_c_596_n N_A_382_413#_c_1264_n 0.0114259f $X=3.315 $Y=1.915 $X2=0
+ $Y2=0
cc_589 N_B_c_597_n N_A_382_413#_c_1264_n 0.00252322f $X=2.75 $Y=1.915 $X2=0
+ $Y2=0
cc_590 N_B_c_598_n N_A_382_413#_c_1264_n 0.0033156f $X=3.615 $Y=1.99 $X2=0 $Y2=0
cc_591 N_B_c_605_n N_A_382_413#_c_1264_n 0.00719178f $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_592 N_B_c_605_n N_A_382_413#_c_1265_n 9.79325e-19 $X=3.33 $Y=1.53 $X2=0 $Y2=0
cc_593 N_B_c_598_n N_A_382_413#_c_1266_n 0.0024353f $X=3.615 $Y=1.99 $X2=0 $Y2=0
cc_594 N_B_c_607_n N_A_738_413#_c_1291_n 0.00513362f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_595 N_B_c_603_n N_A_738_413#_c_1292_n 0.00424941f $X=3.502 $Y=1.915 $X2=0
+ $Y2=0
cc_596 N_B_c_607_n N_A_738_413#_c_1292_n 0.00282827f $X=5.63 $Y=1.53 $X2=0 $Y2=0
cc_597 N_B_c_587_n N_VGND_c_1338_n 0.00676915f $X=2.675 $Y=0.73 $X2=0 $Y2=0
cc_598 N_B_c_587_n N_VGND_c_1339_n 0.00208038f $X=2.675 $Y=0.73 $X2=0 $Y2=0
cc_599 N_B_c_588_n N_VGND_c_1339_n 0.0045972f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_600 N_B_c_592_n N_VGND_c_1339_n 0.00827538f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_601 N_B_c_592_n N_VGND_c_1340_n 5.31689e-19 $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_602 N_B_M1004_g N_VGND_c_1341_n 0.00105809f $X=5.74 $Y=0.445 $X2=0 $Y2=0
cc_603 N_B_M1004_g N_VGND_c_1342_n 0.00357877f $X=5.74 $Y=0.445 $X2=0 $Y2=0
cc_604 N_B_M1025_g N_VGND_c_1345_n 0.00357668f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_605 N_B_c_587_n N_VGND_c_1346_n 0.00337001f $X=2.675 $Y=0.73 $X2=0 $Y2=0
cc_606 N_B_c_588_n N_VGND_c_1346_n 0.00469312f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_607 N_B_c_592_n N_VGND_c_1347_n 0.0046653f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_608 N_B_M1025_g N_VGND_c_1349_n 0.00538188f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_609 N_B_c_587_n N_VGND_c_1349_n 0.00512288f $X=2.675 $Y=0.73 $X2=0 $Y2=0
cc_610 N_B_c_588_n N_VGND_c_1349_n 0.00336079f $X=3.485 $Y=0.805 $X2=0 $Y2=0
cc_611 N_B_M1004_g N_VGND_c_1349_n 0.00530375f $X=5.74 $Y=0.445 $X2=0 $Y2=0
cc_612 N_B_c_592_n N_VGND_c_1349_n 0.00446764f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_613 N_B_c_587_n N_A_382_47#_c_1467_n 0.00758462f $X=2.675 $Y=0.73 $X2=0 $Y2=0
cc_614 N_B_c_588_n N_A_382_47#_c_1467_n 0.00812182f $X=3.485 $Y=0.805 $X2=0
+ $Y2=0
cc_615 N_B_c_589_n N_A_382_47#_c_1467_n 0.00392189f $X=2.75 $Y=0.805 $X2=0 $Y2=0
cc_616 N_B_c_592_n N_A_382_47#_c_1467_n 0.00310565f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_617 N_B_c_592_n N_A_382_47#_c_1484_n 0.00158481f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_618 N_B_c_592_n N_A_738_47#_c_1503_n 0.00420459f $X=3.587 $Y=0.73 $X2=0 $Y2=0
cc_619 N_CIN_M1021_g N_A_995_47#_c_1052_n 0.0116755f $X=5.38 $Y=2.275 $X2=0
+ $Y2=0
cc_620 N_CIN_c_830_n N_A_995_47#_c_1052_n 0.00228311f $X=5.155 $Y=1.6 $X2=0
+ $Y2=0
cc_621 N_CIN_c_835_n N_A_995_47#_c_1052_n 5.57228e-19 $X=5.32 $Y=1.68 $X2=0
+ $Y2=0
cc_622 N_CIN_c_836_n N_A_995_47#_c_1052_n 0.0167105f $X=5.28 $Y=1.6 $X2=0 $Y2=0
cc_623 N_CIN_M1002_g N_A_995_47#_c_1034_n 0.00947783f $X=5.38 $Y=0.445 $X2=0
+ $Y2=0
cc_624 N_CIN_c_836_n N_A_995_47#_c_1043_n 5.66439e-19 $X=5.28 $Y=1.6 $X2=0 $Y2=0
cc_625 N_CIN_M1012_g N_VPWR_c_1149_n 0.00118455f $X=1.835 $Y=2.275 $X2=0 $Y2=0
cc_626 N_CIN_M1008_g N_VPWR_c_1150_n 5.37584e-19 $X=4.035 $Y=2.275 $X2=0 $Y2=0
cc_627 N_CIN_M1008_g N_VPWR_c_1151_n 0.00640108f $X=4.035 $Y=2.275 $X2=0 $Y2=0
cc_628 N_CIN_M1021_g N_VPWR_c_1153_n 0.00357877f $X=5.38 $Y=2.275 $X2=0 $Y2=0
cc_629 N_CIN_M1012_g N_VPWR_c_1156_n 0.00585385f $X=1.835 $Y=2.275 $X2=0 $Y2=0
cc_630 N_CIN_M1008_g N_VPWR_c_1158_n 0.00337001f $X=4.035 $Y=2.275 $X2=0 $Y2=0
cc_631 N_CIN_M1012_g N_VPWR_c_1147_n 0.0108681f $X=1.835 $Y=2.275 $X2=0 $Y2=0
cc_632 N_CIN_M1008_g N_VPWR_c_1147_n 0.00397658f $X=4.035 $Y=2.275 $X2=0 $Y2=0
cc_633 N_CIN_M1021_g N_VPWR_c_1147_n 0.00525841f $X=5.38 $Y=2.275 $X2=0 $Y2=0
cc_634 N_CIN_c_826_n N_A_382_413#_c_1264_n 0.058703f $X=2.79 $Y=1.68 $X2=0 $Y2=0
cc_635 N_CIN_M1012_g N_A_382_413#_c_1265_n 0.00415589f $X=1.835 $Y=2.275 $X2=0
+ $Y2=0
cc_636 N_CIN_c_826_n N_A_382_413#_c_1265_n 0.00691538f $X=2.79 $Y=1.68 $X2=0
+ $Y2=0
cc_637 N_CIN_c_827_n N_A_382_413#_c_1265_n 0.00669798f $X=2.04 $Y=1.68 $X2=0
+ $Y2=0
cc_638 N_CIN_M1008_g N_A_738_413#_c_1291_n 0.0110354f $X=4.035 $Y=2.275 $X2=0
+ $Y2=0
cc_639 N_CIN_c_830_n N_A_738_413#_c_1291_n 0.038655f $X=5.155 $Y=1.6 $X2=0 $Y2=0
cc_640 N_CIN_c_831_n N_A_738_413#_c_1291_n 0.00233744f $X=3.955 $Y=1.6 $X2=0
+ $Y2=0
cc_641 N_CIN_c_832_n N_A_738_413#_c_1291_n 0.00258394f $X=4.035 $Y=1.6 $X2=0
+ $Y2=0
cc_642 N_CIN_c_836_n N_A_738_413#_c_1291_n 9.45372e-19 $X=5.28 $Y=1.6 $X2=0
+ $Y2=0
cc_643 N_CIN_c_831_n N_A_738_413#_c_1292_n 0.00769662f $X=3.955 $Y=1.6 $X2=0
+ $Y2=0
cc_644 N_CIN_c_832_n N_A_738_413#_c_1292_n 2.43081e-19 $X=4.035 $Y=1.6 $X2=0
+ $Y2=0
cc_645 N_CIN_M1023_g N_VGND_c_1338_n 0.00118455f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_646 N_CIN_c_811_n N_VGND_c_1339_n 5.44952e-19 $X=4.037 $Y=0.73 $X2=0 $Y2=0
cc_647 N_CIN_c_815_n N_VGND_c_1339_n 0.00537741f $X=3.785 $Y=1.107 $X2=0 $Y2=0
cc_648 N_CIN_c_811_n N_VGND_c_1340_n 0.00639437f $X=4.037 $Y=0.73 $X2=0 $Y2=0
cc_649 N_CIN_M1002_g N_VGND_c_1342_n 0.00357877f $X=5.38 $Y=0.445 $X2=0 $Y2=0
cc_650 N_CIN_M1023_g N_VGND_c_1345_n 0.00585385f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_651 N_CIN_c_811_n N_VGND_c_1347_n 0.00337001f $X=4.037 $Y=0.73 $X2=0 $Y2=0
cc_652 N_CIN_M1023_g N_VGND_c_1349_n 0.00649423f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_653 N_CIN_M1002_g N_VGND_c_1349_n 0.00515781f $X=5.38 $Y=0.445 $X2=0 $Y2=0
cc_654 N_CIN_c_811_n N_VGND_c_1349_n 0.00377406f $X=4.037 $Y=0.73 $X2=0 $Y2=0
cc_655 N_CIN_c_815_n N_A_382_47#_c_1467_n 5.77639e-19 $X=3.785 $Y=1.107 $X2=0
+ $Y2=0
cc_656 N_CIN_c_816_n N_A_382_47#_c_1467_n 0.0110711f $X=2.96 $Y=1.107 $X2=0
+ $Y2=0
cc_657 N_CIN_M1023_g N_A_382_47#_c_1468_n 0.00129924f $X=1.835 $Y=0.445 $X2=0
+ $Y2=0
cc_658 N_CIN_c_818_n N_A_382_47#_c_1468_n 2.17239e-19 $X=1.835 $Y=1.19 $X2=0
+ $Y2=0
cc_659 N_CIN_c_819_n N_A_382_47#_c_1468_n 0.00270907f $X=1.955 $Y=1.19 $X2=0
+ $Y2=0
cc_660 N_CIN_c_811_n N_A_738_47#_c_1502_n 0.00669222f $X=4.037 $Y=0.73 $X2=0
+ $Y2=0
cc_661 N_CIN_c_812_n N_A_738_47#_c_1502_n 0.00564483f $X=4.037 $Y=0.88 $X2=0
+ $Y2=0
cc_662 N_CIN_c_815_n N_A_738_47#_c_1502_n 0.00301863f $X=3.785 $Y=1.107 $X2=0
+ $Y2=0
cc_663 N_CIN_c_832_n N_A_738_47#_c_1502_n 0.00124331f $X=4.035 $Y=1.6 $X2=0
+ $Y2=0
cc_664 N_CIN_c_815_n N_A_738_47#_c_1503_n 0.0115587f $X=3.785 $Y=1.107 $X2=0
+ $Y2=0
cc_665 N_A_995_47#_c_1041_n N_VPWR_M1015_d 0.00671884f $X=6.495 $Y=2.02 $X2=0
+ $Y2=0
cc_666 N_A_995_47#_c_1042_n N_VPWR_M1015_d 0.00546326f $X=6.58 $Y=1.935 $X2=0
+ $Y2=0
cc_667 N_A_995_47#_M1006_g N_VPWR_c_1152_n 0.00808649f $X=6.715 $Y=1.985 $X2=0
+ $Y2=0
cc_668 N_A_995_47#_c_1041_n N_VPWR_c_1152_n 0.0200213f $X=6.495 $Y=2.02 $X2=0
+ $Y2=0
cc_669 N_A_995_47#_c_1052_n N_VPWR_c_1153_n 0.0530726f $X=6 $Y=2.295 $X2=0 $Y2=0
cc_670 N_A_995_47#_c_1041_n N_VPWR_c_1153_n 0.00259773f $X=6.495 $Y=2.02 $X2=0
+ $Y2=0
cc_671 N_A_995_47#_c_1043_n N_VPWR_c_1153_n 0.00963745f $X=6.085 $Y=2.02 $X2=0
+ $Y2=0
cc_672 N_A_995_47#_M1006_g N_VPWR_c_1159_n 0.0046653f $X=6.715 $Y=1.985 $X2=0
+ $Y2=0
cc_673 N_A_995_47#_M1010_d N_VPWR_c_1147_n 0.00641803f $X=4.975 $Y=2.065 $X2=0
+ $Y2=0
cc_674 N_A_995_47#_M1006_g N_VPWR_c_1147_n 0.0090943f $X=6.715 $Y=1.985 $X2=0
+ $Y2=0
cc_675 N_A_995_47#_c_1052_n N_VPWR_c_1147_n 0.0331712f $X=6 $Y=2.295 $X2=0 $Y2=0
cc_676 N_A_995_47#_c_1041_n N_VPWR_c_1147_n 0.00584423f $X=6.495 $Y=2.02 $X2=0
+ $Y2=0
cc_677 N_A_995_47#_c_1043_n N_VPWR_c_1147_n 0.00631874f $X=6.085 $Y=2.02 $X2=0
+ $Y2=0
cc_678 N_A_995_47#_c_1052_n N_A_738_413#_c_1305_n 0.016651f $X=6 $Y=2.295 $X2=0
+ $Y2=0
cc_679 N_A_995_47#_c_1052_n A_1091_413# 0.00289261f $X=6 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_680 N_A_995_47#_c_1052_n A_1163_413# 0.00379213f $X=6 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_681 N_A_995_47#_c_1043_n A_1163_413# 0.00237999f $X=6.085 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_682 N_A_995_47#_c_1042_n SUM 0.00914827f $X=6.58 $Y=1.935 $X2=0 $Y2=0
cc_683 N_A_995_47#_c_1036_n SUM 0.0249546f $X=6.655 $Y=1.16 $X2=0 $Y2=0
cc_684 N_A_995_47#_c_1038_n SUM 0.010468f $X=6.617 $Y=0.995 $X2=0 $Y2=0
cc_685 N_A_995_47#_c_1039_n SUM 0.0151345f $X=6.655 $Y=0.995 $X2=0 $Y2=0
cc_686 N_A_995_47#_c_1035_n N_VGND_M1013_d 0.00672944f $X=6.495 $Y=0.7 $X2=0
+ $Y2=0
cc_687 N_A_995_47#_c_1038_n N_VGND_M1013_d 0.00117264f $X=6.617 $Y=0.995 $X2=0
+ $Y2=0
cc_688 N_A_995_47#_c_1035_n N_VGND_c_1341_n 0.0201928f $X=6.495 $Y=0.7 $X2=0
+ $Y2=0
cc_689 N_A_995_47#_c_1037_n N_VGND_c_1341_n 2.43955e-19 $X=6.655 $Y=1.16 $X2=0
+ $Y2=0
cc_690 N_A_995_47#_c_1039_n N_VGND_c_1341_n 0.00409489f $X=6.655 $Y=0.995 $X2=0
+ $Y2=0
cc_691 N_A_995_47#_c_1034_n N_VGND_c_1342_n 0.0114f $X=5.925 $Y=0.38 $X2=0 $Y2=0
cc_692 N_A_995_47#_c_1035_n N_VGND_c_1342_n 0.00256355f $X=6.495 $Y=0.7 $X2=0
+ $Y2=0
cc_693 N_A_995_47#_c_1048_n N_VGND_c_1342_n 0.0474775f $X=5.255 $Y=0.425 $X2=0
+ $Y2=0
cc_694 N_A_995_47#_c_1035_n N_VGND_c_1348_n 9.25461e-19 $X=6.495 $Y=0.7 $X2=0
+ $Y2=0
cc_695 N_A_995_47#_c_1039_n N_VGND_c_1348_n 0.00558147f $X=6.655 $Y=0.995 $X2=0
+ $Y2=0
cc_696 N_A_995_47#_M1007_d N_VGND_c_1349_n 0.0024769f $X=4.975 $Y=0.235 $X2=0
+ $Y2=0
cc_697 N_A_995_47#_c_1034_n N_VGND_c_1349_n 0.00642843f $X=5.925 $Y=0.38 $X2=0
+ $Y2=0
cc_698 N_A_995_47#_c_1035_n N_VGND_c_1349_n 0.00789204f $X=6.495 $Y=0.7 $X2=0
+ $Y2=0
cc_699 N_A_995_47#_c_1048_n N_VGND_c_1349_n 0.0227627f $X=5.255 $Y=0.425 $X2=0
+ $Y2=0
cc_700 N_A_995_47#_c_1039_n N_VGND_c_1349_n 0.0111802f $X=6.655 $Y=0.995 $X2=0
+ $Y2=0
cc_701 N_A_995_47#_c_1048_n N_A_738_47#_c_1521_n 0.0162015f $X=5.255 $Y=0.425
+ $X2=0 $Y2=0
cc_702 N_A_995_47#_c_1034_n A_1091_47# 0.00296887f $X=5.925 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_703 N_A_995_47#_c_1034_n A_1163_47# 0.00709994f $X=5.925 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_704 N_COUT_c_1134_n N_VPWR_c_1155_n 0.018001f $X=0.26 $Y=1.775 $X2=0 $Y2=0
cc_705 N_COUT_M1017_s N_VPWR_c_1147_n 0.00387172f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_706 N_COUT_c_1134_n N_VPWR_c_1147_n 0.00993603f $X=0.26 $Y=1.775 $X2=0 $Y2=0
cc_707 COUT N_VGND_c_1344_n 0.0179343f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_708 N_COUT_M1024_s N_VGND_c_1349_n 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_709 COUT N_VGND_c_1349_n 0.00992194f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_710 N_VPWR_c_1147_n A_208_413# 0.00240919f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_711 N_VPWR_c_1147_n N_A_382_413#_M1012_d 0.00409863f $X=7.13 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_712 N_VPWR_c_1147_n N_A_382_413#_M1005_d 0.00226128f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_713 N_VPWR_c_1156_n N_A_382_413#_c_1281_n 0.0111986f $X=2.3 $Y=2.72 $X2=0
+ $Y2=0
cc_714 N_VPWR_c_1147_n N_A_382_413#_c_1281_n 0.00642843f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_715 N_VPWR_M1009_d N_A_382_413#_c_1264_n 0.00158918f $X=2.33 $Y=2.065 $X2=0
+ $Y2=0
cc_716 N_VPWR_c_1149_n N_A_382_413#_c_1264_n 0.0158599f $X=2.465 $Y=2.36 $X2=0
+ $Y2=0
cc_717 N_VPWR_c_1156_n N_A_382_413#_c_1264_n 0.00255672f $X=2.3 $Y=2.72 $X2=0
+ $Y2=0
cc_718 N_VPWR_c_1157_n N_A_382_413#_c_1264_n 0.00255672f $X=3.24 $Y=2.72 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_1147_n N_A_382_413#_c_1264_n 0.0101119f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_1150_n N_A_382_413#_c_1266_n 0.0149504f $X=3.405 $Y=2.34 $X2=0
+ $Y2=0
cc_721 N_VPWR_c_1157_n N_A_382_413#_c_1266_n 0.0159201f $X=3.24 $Y=2.72 $X2=0
+ $Y2=0
cc_722 N_VPWR_c_1147_n N_A_382_413#_c_1266_n 0.00891562f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_723 N_VPWR_c_1147_n N_A_738_413#_M1022_d 0.00409863f $X=7.13 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_724 N_VPWR_c_1147_n N_A_738_413#_M1003_d 0.00516727f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_725 N_VPWR_c_1158_n N_A_738_413#_c_1308_n 0.0111986f $X=4.08 $Y=2.72 $X2=0
+ $Y2=0
cc_726 N_VPWR_c_1147_n N_A_738_413#_c_1308_n 0.00642843f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_727 N_VPWR_M1008_d N_A_738_413#_c_1291_n 0.00158918f $X=4.11 $Y=2.065 $X2=0
+ $Y2=0
cc_728 N_VPWR_c_1151_n N_A_738_413#_c_1291_n 0.0158599f $X=4.245 $Y=2.36 $X2=0
+ $Y2=0
cc_729 N_VPWR_c_1153_n N_A_738_413#_c_1291_n 0.00255672f $X=6.34 $Y=2.72 $X2=0
+ $Y2=0
cc_730 N_VPWR_c_1158_n N_A_738_413#_c_1291_n 0.00255672f $X=4.08 $Y=2.72 $X2=0
+ $Y2=0
cc_731 N_VPWR_c_1147_n N_A_738_413#_c_1291_n 0.0101119f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_732 N_VPWR_c_1153_n N_A_738_413#_c_1305_n 0.0114f $X=6.34 $Y=2.72 $X2=0 $Y2=0
cc_733 N_VPWR_c_1147_n N_A_738_413#_c_1305_n 0.00642843f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_734 N_VPWR_c_1147_n A_1091_413# 0.00168648f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_735 N_VPWR_c_1147_n A_1163_413# 0.00264201f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_736 N_VPWR_c_1147_n N_SUM_M1006_d 0.00387172f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_737 N_VPWR_c_1159_n N_SUM_c_1325_n 0.0280384f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_738 N_VPWR_c_1147_n N_SUM_c_1325_n 0.0153277f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_739 SUM N_VGND_c_1348_n 0.0279732f $X=7.07 $Y=0.425 $X2=0 $Y2=0
cc_740 N_SUM_M1016_d N_VGND_c_1349_n 0.00387172f $X=6.79 $Y=0.235 $X2=0 $Y2=0
cc_741 SUM N_VGND_c_1349_n 0.0153137f $X=7.07 $Y=0.425 $X2=0 $Y2=0
cc_742 N_VGND_c_1349_n A_208_47# 0.00266434f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_743 N_VGND_c_1349_n N_A_382_47#_M1023_d 0.00227466f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_744 N_VGND_c_1349_n N_A_382_47#_M1000_d 0.00204709f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_745 N_VGND_c_1345_n N_A_382_47#_c_1492_n 0.0111986f $X=2.3 $Y=0 $X2=0 $Y2=0
cc_746 N_VGND_c_1349_n N_A_382_47#_c_1492_n 0.00304042f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_747 N_VGND_M1001_d N_A_382_47#_c_1467_n 0.00158918f $X=2.33 $Y=0.235 $X2=0
+ $Y2=0
cc_748 N_VGND_c_1338_n N_A_382_47#_c_1467_n 0.0147553f $X=2.465 $Y=0.36 $X2=0
+ $Y2=0
cc_749 N_VGND_c_1345_n N_A_382_47#_c_1467_n 0.00255672f $X=2.3 $Y=0 $X2=0 $Y2=0
cc_750 N_VGND_c_1346_n N_A_382_47#_c_1467_n 0.00255672f $X=3.24 $Y=0 $X2=0 $Y2=0
cc_751 N_VGND_c_1349_n N_A_382_47#_c_1467_n 0.00461038f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_752 N_VGND_c_1339_n N_A_382_47#_c_1484_n 0.0131643f $X=3.405 $Y=0.405 $X2=0
+ $Y2=0
cc_753 N_VGND_c_1346_n N_A_382_47#_c_1484_n 0.0114f $X=3.24 $Y=0 $X2=0 $Y2=0
cc_754 N_VGND_c_1349_n N_A_382_47#_c_1484_n 0.00304042f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_755 N_VGND_c_1349_n N_A_738_47#_M1026_d 0.00227466f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_756 N_VGND_c_1349_n N_A_738_47#_M1019_d 0.00263427f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_757 N_VGND_c_1347_n N_A_738_47#_c_1524_n 0.0111986f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_758 N_VGND_c_1349_n N_A_738_47#_c_1524_n 0.00304042f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_759 N_VGND_M1014_d N_A_738_47#_c_1502_n 0.00158918f $X=4.11 $Y=0.235 $X2=0
+ $Y2=0
cc_760 N_VGND_c_1340_n N_A_738_47#_c_1502_n 0.0147553f $X=4.245 $Y=0.36 $X2=0
+ $Y2=0
cc_761 N_VGND_c_1342_n N_A_738_47#_c_1502_n 0.00255672f $X=6.265 $Y=0 $X2=0
+ $Y2=0
cc_762 N_VGND_c_1347_n N_A_738_47#_c_1502_n 0.00255672f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_763 N_VGND_c_1349_n N_A_738_47#_c_1502_n 0.00461038f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_764 N_VGND_c_1342_n N_A_738_47#_c_1521_n 0.0114f $X=6.265 $Y=0 $X2=0 $Y2=0
cc_765 N_VGND_c_1349_n N_A_738_47#_c_1521_n 0.00304042f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_766 N_VGND_c_1349_n A_1091_47# 0.00167819f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_767 N_VGND_c_1349_n A_1163_47# 0.002802f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__lpflow_bleeder_1.spice.pex
* Created: Thu Aug 27 14:23:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%SHORT 1 3 4 6 7 9 10 12 13 15 16 27
+ 28
r26 26 28 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.74 $Y=1.16 $X2=2.1
+ $Y2=1.16
r27 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.74
+ $Y=1.16 $X2=1.74 $Y2=1.16
r28 24 26 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.74 $Y2=1.16
r29 23 24 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.38 $Y2=1.16
r30 22 27 17.6812 $w=6.88e-07 $l=1.02e-06 $layer=LI1_cond $X=0.72 $Y=1.385
+ $X2=1.74 $Y2=1.385
r31 21 23 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=0.72 $Y=1.16 $X2=1.02
+ $Y2=1.16
r32 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.72
+ $Y=1.16 $X2=0.72 $Y2=1.16
r33 18 21 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.66 $Y=1.16 $X2=0.72
+ $Y2=1.16
r34 16 22 3.46689 $w=6.88e-07 $l=2e-07 $layer=LI1_cond $X=0.52 $Y=1.385 $X2=0.72
+ $Y2=1.385
r35 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=0.995
+ $X2=2.1 $Y2=1.16
r36 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.1 $Y=0.995 $X2=2.1
+ $Y2=0.705
r37 10 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=0.995
+ $X2=1.74 $Y2=1.16
r38 10 12 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.74 $Y=0.995
+ $X2=1.74 $Y2=0.705
r39 7 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=0.995
+ $X2=1.38 $Y2=1.16
r40 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.38 $Y=0.995 $X2=1.38
+ $Y2=0.705
r41 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=0.995
+ $X2=1.02 $Y2=1.16
r42 4 6 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.02 $Y=0.995 $X2=1.02
+ $Y2=0.705
r43 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.66 $Y=0.995
+ $X2=0.66 $Y2=1.16
r44 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.66 $Y=0.995 $X2=0.66
+ $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%VGND 1 6 9 10 11 20 21
r20 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r21 18 21 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r22 17 20 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r23 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r24 11 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r25 11 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r26 9 14 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.23
+ $Y2=0
r27 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.45
+ $Y2=0
r28 8 17 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.69
+ $Y2=0
r29 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.45
+ $Y2=0
r30 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=0.085 $X2=0.45
+ $Y2=0
r31 4 6 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=0.45 $Y=0.085 $X2=0.45
+ $Y2=0.705
r32 1 6 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.525 $X2=0.45 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%VPWR 1 6 8 9 10 11 22
r13 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r14 19 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r15 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r16 14 18 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r17 11 19 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r18 11 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r19 9 18 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=2.07 $Y2=2.72
r20 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=2.31 $Y2=2.72
r21 8 21 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=2.475 $Y=2.72 $X2=2.53
+ $Y2=2.72
r22 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=2.72
+ $X2=2.31 $Y2=2.72
r23 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=2.635 $X2=2.31
+ $Y2=2.72
r24 4 6 67.4005 $w=3.28e-07 $l=1.93e-06 $layer=LI1_cond $X=2.31 $Y=2.635
+ $X2=2.31 $Y2=0.705
r25 1 6 182 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_NDIFF $count=1 $X=2.175
+ $Y=0.525 $X2=2.31 $Y2=0.705
.ends


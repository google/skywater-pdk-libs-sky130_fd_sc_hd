* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4.pex.spice
* Created: Thu Aug 27 14:26:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VGND 1 2 3 4 5 6 7
+ 8 9 40 54 58 62 66 70 74 78 82 86 97 100 103 106 109 112 114 115 140 147 163
+ 179
c165 78 0 7.6696e-20 $X=5 $Y=0.42
r166 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=5.44
+ $X2=7.13 $Y2=5.44
r167 175 176 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=5.44
+ $X2=4.83 $Y2=5.44
r168 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r169 169 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=5.44
+ $X2=0.23 $Y2=5.44
r170 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r171 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r172 160 163 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r173 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r174 157 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r175 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r176 154 179 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=5.44
+ $X2=7.13 $Y2=5.44
r177 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=5.44
+ $X2=6.67 $Y2=5.44
r178 151 154 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=5.44
+ $X2=6.67 $Y2=5.44
r179 151 176 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=5.44
+ $X2=4.83 $Y2=5.44
r180 150 153 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=5.44
+ $X2=6.67 $Y2=5.44
r181 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=5.44
+ $X2=5.29 $Y2=5.44
r182 148 175 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.955 $Y=5.44
+ $X2=4.7 $Y2=5.44
r183 148 150 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.955 $Y=5.44
+ $X2=5.29 $Y2=5.44
r184 147 178 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=6.985 $Y=5.44
+ $X2=7.172 $Y2=5.44
r185 147 153 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.985 $Y=5.44
+ $X2=6.67 $Y2=5.44
r186 146 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r187 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r188 143 176 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=5.44
+ $X2=4.83 $Y2=5.44
r189 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=5.44
+ $X2=4.37 $Y2=5.44
r190 140 175 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.445 $Y=5.44
+ $X2=4.7 $Y2=5.44
r191 140 142 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.445 $Y=5.44
+ $X2=4.37 $Y2=5.44
r192 139 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r193 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r194 136 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=5.44
+ $X2=4.37 $Y2=5.44
r195 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=5.44
+ $X2=3.45 $Y2=5.44
r196 133 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r197 133 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r198 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r199 130 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0
+ $X2=2.185 $Y2=0
r200 130 132 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.99
+ $Y2=0
r201 129 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=5.44
+ $X2=3.45 $Y2=5.44
r202 128 129 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=5.44
+ $X2=2.53 $Y2=5.44
r203 126 129 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=5.44
+ $X2=2.53 $Y2=5.44
r204 125 128 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=5.44
+ $X2=2.53 $Y2=5.44
r205 125 126 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=5.44
+ $X2=0.69 $Y2=5.44
r206 123 169 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=5.44
+ $X2=0.187 $Y2=5.44
r207 123 125 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=5.44
+ $X2=0.69 $Y2=5.44
r208 122 173 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r209 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r210 119 166 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r211 119 121 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.69 $Y2=0
r212 118 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=0
+ $X2=2.185 $Y2=0
r213 118 121 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=2.02 $Y=0
+ $X2=0.69 $Y2=0
r214 115 122 0.0554856 $w=4.8e-07 $l=1.95e-07 $layer=MET1_cond $X=0.495 $Y=0
+ $X2=0.69 $Y2=0
r215 115 167 0.0754035 $w=4.8e-07 $l=2.65e-07 $layer=MET1_cond $X=0.495 $Y=0
+ $X2=0.23 $Y2=0
r216 114 126 0.0825171 $w=4.8e-07 $l=2.9e-07 $layer=MET1_cond $X=0.4 $Y=5.44
+ $X2=0.69 $Y2=5.44
r217 114 170 0.0483721 $w=4.8e-07 $l=1.7e-07 $layer=MET1_cond $X=0.4 $Y=5.44
+ $X2=0.23 $Y2=5.44
r218 112 159 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.67 $Y2=0
r219 112 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.88 $Y2=0
r220 111 162 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.13 $Y2=0
r221 111 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=6.88 $Y2=0
r222 109 156 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.75 $Y2=0
r223 109 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.99 $Y2=0
r224 108 159 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=6.67 $Y2=0
r225 108 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=5.99 $Y2=0
r226 106 145 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.83 $Y2=0
r227 106 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r228 105 156 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.75 $Y2=0
r229 105 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r230 103 138 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=0
+ $X2=3.91 $Y2=0
r231 103 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0
+ $X2=4.14 $Y2=0
r232 102 145 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.83 $Y2=0
r233 102 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.14 $Y2=0
r234 100 135 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=5.44
+ $X2=3.45 $Y2=5.44
r235 100 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.575 $Y=5.44
+ $X2=3.67 $Y2=5.44
r236 99 142 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.765 $Y=5.44
+ $X2=4.37 $Y2=5.44
r237 99 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.765 $Y=5.44
+ $X2=3.67 $Y2=5.44
r238 97 132 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=0
+ $X2=2.99 $Y2=0
r239 97 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.28
+ $Y2=0
r240 96 138 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.91 $Y2=0
r241 96 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.28
+ $Y2=0
r242 94 128 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.645 $Y=5.44
+ $X2=2.53 $Y2=5.44
r243 94 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.645 $Y=5.44
+ $X2=2.775 $Y2=5.44
r244 93 135 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.905 $Y=5.44
+ $X2=3.45 $Y2=5.44
r245 93 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.905 $Y=5.44
+ $X2=2.775 $Y2=5.44
r246 88 178 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.13 $Y=5.355
+ $X2=7.172 $Y2=5.44
r247 84 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.88 $Y=0.085
+ $X2=6.88 $Y2=0
r248 84 86 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.88 $Y=0.085
+ $X2=6.88 $Y2=0.42
r249 80 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0
r250 80 82 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0.42
r251 76 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r252 76 78 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.42
r253 72 175 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=5.355
+ $X2=4.7 $Y2=5.44
r254 72 74 14.5406 $w=5.08e-07 $l=6.2e-07 $layer=LI1_cond $X=4.7 $Y=5.355
+ $X2=4.7 $Y2=4.735
r255 68 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r256 68 70 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.42
r257 64 101 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=5.355
+ $X2=3.67 $Y2=5.44
r258 64 66 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=3.67 $Y=5.355
+ $X2=3.67 $Y2=4.735
r259 60 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0
r260 60 62 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0.42
r261 56 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=5.355
+ $X2=2.775 $Y2=5.44
r262 56 58 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=2.775 $Y=5.355
+ $X2=2.775 $Y2=4.7
r263 52 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0
r264 52 54 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0.62
r265 47 169 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=5.355
+ $X2=0.187 $Y2=5.44
r266 42 166 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.187 $Y2=0
r267 40 88 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=7.13 $Y=4.8
+ $X2=7.13 $Y2=5.355
r268 40 47 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=0.23 $Y=4.8
+ $X2=0.23 $Y2=5.355
r269 40 42 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=0.23 $Y=0.64
+ $X2=0.23 $Y2=0.085
r270 9 86 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.71
+ $Y=0.235 $X2=6.85 $Y2=0.42
r271 8 82 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.85
+ $Y=0.235 $X2=5.99 $Y2=0.42
r272 7 78 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=0.235 $X2=5 $Y2=0.42
r273 6 74 45.5 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=4 $X=4.39
+ $Y=4.555 $X2=4.87 $Y2=4.735
r274 5 70 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.235 $X2=4.14 $Y2=0.42
r275 4 66 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.53 $Y=4.555
+ $X2=3.67 $Y2=4.735
r276 3 62 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.135
+ $Y=0.235 $X2=3.28 $Y2=0.42
r277 2 58 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.685
+ $Y=4.555 $X2=2.81 $Y2=4.7
r278 1 54 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.41 $X2=2.245 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPB 7 8 11 15 19 22
+ 27 33
r89 19 33 0.00371286 $w=1.4e-07 $l=3e-09 $layer=MET1_cond $X=0.557 $Y=3.57
+ $X2=0.56 $Y2=3.57
r90 18 27 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=7.13 $Y=3.57 $X2=7.13
+ $Y2=3.29
r91 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.075 $Y=3.57
+ $X2=7.075 $Y2=3.57
r92 15 33 7.88365 $w=1.4e-07 $l=6.37e-06 $layer=MET1_cond $X=6.93 $Y=3.57
+ $X2=0.56 $Y2=3.57
r93 15 17 0.0999252 $w=2.12e-07 $l=1.45e-07 $layer=MET1_cond $X=6.93 $Y=3.57
+ $X2=7.075 $Y2=3.57
r94 14 22 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=0.23 $Y=3.57 $X2=0.23
+ $Y2=3.29
r95 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.225 $Y=3.57
+ $X2=0.225 $Y2=3.57
r96 11 19 0.231435 $w=1.4e-07 $l=1.87e-07 $layer=MET1_cond $X=0.37 $Y=3.57
+ $X2=0.557 $Y2=3.57
r97 11 13 0.0980892 $w=2.27e-07 $l=1.45e-07 $layer=MET1_cond $X=0.37 $Y=3.57
+ $X2=0.225 $Y2=3.57
r98 8 27 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=7.045 $Y=3.04 $X2=7.13 $Y2=3.29
r99 7 22 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=0.145 $Y=3.04 $X2=0.23 $Y2=3.29
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPWRIN 1 7 11 16 17
+ 20 25 26 30 32 34
c64 25 0 2.86228e-19 $X=2.225 $Y=2.2
r65 30 32 1.10767 $w=1.4e-07 $l=8.95e-07 $layer=MET1_cond $X=1.36 $Y=2.21
+ $X2=0.465 $Y2=2.21
r66 26 34 2.07418 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.2
+ $X2=2.06 $Y2=2.2
r67 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.225 $Y=2.2
+ $X2=2.225 $Y2=2.2
r68 23 34 23.6891 $w=2.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.505 $Y=2.2
+ $X2=2.06 $Y2=2.2
r69 22 25 0.461955 $w=2.3e-07 $l=7.2e-07 $layer=MET1_cond $X=1.505 $Y=2.2
+ $X2=2.225 $Y2=2.2
r70 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.505 $Y=2.2
+ $X2=1.505 $Y2=2.2
r71 20 30 0.0864037 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=1.475 $Y=2.2
+ $X2=1.36 $Y2=2.2
r72 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=1.475 $Y=2.2
+ $X2=1.505 $Y2=2.2
r73 16 17 17.048 $w=7.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.435 $Y=3.49
+ $X2=2.435 $Y2=2.66
r74 13 26 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.225 $Y=2.335
+ $X2=2.225 $Y2=2.2
r75 13 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.225 $Y=2.335
+ $X2=2.225 $Y2=2.66
r76 9 26 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=2.2
r77 9 11 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=1.79
r78 7 16 91 $w=1.7e-07 $l=6.45697e-07 $layer=licon1_NTAP_notbjt $count=2 $X=2.1
+ $Y=3.27 $X2=2.645 $Y2=3.49
r79 1 11 300 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_PDIFF $count=2 $X=2.1
+ $Y=1.485 $X2=2.225 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_505_297# 1 2 7 9
+ 10 12 13 14 15 17 18 20 22 28 31 35 36 39 40
c84 40 0 1.64106e-19 $X=3.225 $Y=3.84
c85 39 0 1.09489e-19 $X=3.225 $Y=3.84
r86 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=3.84 $X2=3.225 $Y2=3.84
r87 37 39 51.3361 $w=3.28e-07 $l=1.47e-06 $layer=LI1_cond $X=3.225 $Y=2.37
+ $X2=3.225 $Y2=3.84
r88 35 37 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=3.06 $Y=2.25
+ $X2=3.225 $Y2=2.37
r89 35 36 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.06 $Y=2.25 $X2=2.8
+ $Y2=2.25
r90 31 34 56.1816 $w=2.38e-07 $l=1.17e-06 $layer=LI1_cond $X=2.68 $Y=0.62
+ $X2=2.68 $Y2=1.79
r91 29 36 6.81649 $w=2.4e-07 $l=1.69706e-07 $layer=LI1_cond $X=2.68 $Y=2.13
+ $X2=2.8 $Y2=2.25
r92 29 34 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.68 $Y=2.13
+ $X2=2.68 $Y2=1.79
r93 26 40 80.7859 $w=3.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.235 $Y=4.33
+ $X2=3.235 $Y2=3.84
r94 26 27 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.235 $Y=4.405
+ $X2=3.455 $Y2=4.405
r95 23 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.025 $Y=4.405
+ $X2=3.235 $Y2=4.405
r96 20 22 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.315 $Y=4.48
+ $X2=4.315 $Y2=4.88
r97 19 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.96 $Y=4.405
+ $X2=3.885 $Y2=4.405
r98 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.24 $Y=4.405
+ $X2=4.315 $Y2=4.48
r99 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.24 $Y=4.405
+ $X2=3.96 $Y2=4.405
r100 15 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.885 $Y=4.48
+ $X2=3.885 $Y2=4.405
r101 15 17 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.885 $Y=4.48
+ $X2=3.885 $Y2=4.88
r102 14 27 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.53 $Y=4.405
+ $X2=3.455 $Y2=4.405
r103 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.81 $Y=4.405
+ $X2=3.885 $Y2=4.405
r104 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.81 $Y=4.405
+ $X2=3.53 $Y2=4.405
r105 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.455 $Y=4.48
+ $X2=3.455 $Y2=4.405
r106 10 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.455 $Y=4.48
+ $X2=3.455 $Y2=4.88
r107 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.025 $Y=4.48
+ $X2=3.025 $Y2=4.405
r108 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.025 $Y=4.48 $X2=3.025
+ $Y2=4.88
r109 2 34 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=2.525
+ $Y=1.485 $X2=2.675 $Y2=1.79
r110 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.41 $X2=2.675 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_714_47# 1 2 3 10
+ 11 14 19 22 23 24 28 29 30 31 34 38 45
c103 28 0 1.64375e-19 $X=4.105 $Y=2.07
c104 14 0 7.6696e-20 $X=4.78 $Y=1.955
c105 11 0 1.09489e-19 $X=4.27 $Y=2.58
c106 10 0 1.90316e-19 $X=4.705 $Y=2.58
r107 43 45 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.765 $Y=2.49
+ $X2=4.105 $Y2=2.49
r108 40 42 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=3.71 $Y=0.855
+ $X2=4.105 $Y2=0.855
r109 36 38 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=4.57 $Y=0.73
+ $X2=4.57 $Y2=0.42
r110 32 34 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.555 $Y=3.47
+ $X2=4.555 $Y2=3.235
r111 31 42 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.855
+ $X2=4.105 $Y2=0.855
r112 30 36 6.98266 $w=2.5e-07 $l=1.65831e-07 $layer=LI1_cond $X=4.475 $Y=0.855
+ $X2=4.57 $Y2=0.73
r113 30 31 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.475 $Y=0.855
+ $X2=4.19 $Y2=0.855
r114 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.105
+ $Y=2.07 $X2=4.105 $Y2=2.07
r115 26 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.405
+ $X2=4.105 $Y2=2.49
r116 26 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.105 $Y=2.405
+ $X2=4.105 $Y2=2.07
r117 25 42 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.105 $Y=0.98
+ $X2=4.105 $Y2=0.855
r118 25 28 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.105 $Y=0.98
+ $X2=4.105 $Y2=2.07
r119 23 32 9.70995 $w=1.99e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.39 $Y=3.555
+ $X2=4.555 $Y2=3.47
r120 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.39 $Y=3.555
+ $X2=3.85 $Y2=3.555
r121 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=3.47
+ $X2=3.85 $Y2=3.555
r122 21 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=2.575
+ $X2=3.765 $Y2=2.49
r123 21 22 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.765 $Y=2.575
+ $X2=3.765 $Y2=3.47
r124 17 40 2.34666 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.71 $Y=0.73
+ $X2=3.71 $Y2=0.855
r125 17 19 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=3.71 $Y=0.73
+ $X2=3.71 $Y2=0.42
r126 16 29 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=4.105 $Y=2.505
+ $X2=4.105 $Y2=2.07
r127 12 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.78 $Y=2.505
+ $X2=4.78 $Y2=1.955
r128 11 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.27 $Y=2.58
+ $X2=4.105 $Y2=2.505
r129 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.705 $Y=2.58
+ $X2=4.78 $Y2=2.505
r130 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=2.58
+ $X2=4.27 $Y2=2.58
r131 3 34 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=3.09 $X2=4.555 $Y2=3.235
r132 2 38 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.43
+ $Y=0.235 $X2=4.57 $Y2=0.42
r133 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A 3 5 7 8 12 14 15
+ 18 20 24 26 30 32 33 34 35 39
c71 15 0 1.64375e-19 $X=3.63 $Y=1.145
r72 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.25 $X2=3.125 $Y2=1.25
r73 35 39 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=3.13 $Y=1.425
+ $X2=3.13 $Y2=1.25
r74 28 30 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.785 $Y=1.07
+ $X2=4.785 $Y2=0.56
r75 27 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.43 $Y=1.145
+ $X2=4.355 $Y2=1.145
r76 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.71 $Y=1.145
+ $X2=4.785 $Y2=1.07
r77 26 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.71 $Y=1.145
+ $X2=4.43 $Y2=1.145
r78 22 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.355 $Y=1.07
+ $X2=4.355 $Y2=1.145
r79 22 24 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.355 $Y=1.07
+ $X2=4.355 $Y2=0.56
r80 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4 $Y=1.145 $X2=3.925
+ $Y2=1.145
r81 20 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.28 $Y=1.145
+ $X2=4.355 $Y2=1.145
r82 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.28 $Y=1.145 $X2=4
+ $Y2=1.145
r83 16 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=1.07
+ $X2=3.925 $Y2=1.145
r84 16 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.925 $Y=1.07
+ $X2=3.925 $Y2=0.56
r85 14 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.85 $Y=1.145
+ $X2=3.925 $Y2=1.145
r86 14 15 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.85 $Y=1.145
+ $X2=3.63 $Y2=1.145
r87 10 15 33.8325 $w=2.41e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.63 $Y2=1.145
r88 10 38 74 $w=2.41e-07 $l=4.75857e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.125 $Y2=1.312
r89 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.495 $Y2=0.56
r90 9 32 4.83878 $w=1.55e-07 $l=9.38083e-08 $layer=POLY_cond $X=2.535 $Y=1.147
+ $X2=2.455 $Y2=1.117
r91 8 38 39.1212 $w=2.41e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.96 $Y=1.147
+ $X2=3.125 $Y2=1.312
r92 8 9 203.325 $w=1.55e-07 $l=4.25e-07 $layer=POLY_cond $X=2.96 $Y=1.147
+ $X2=2.535 $Y2=1.147
r93 5 32 20.9729 $w=1.5e-07 $l=1.09471e-07 $layer=POLY_cond $X=2.46 $Y=1.01
+ $X2=2.455 $Y2=1.117
r94 5 7 125.32 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.46 $Y=1.01 $X2=2.46
+ $Y2=0.62
r95 1 32 20.9729 $w=1.5e-07 $l=1.10472e-07 $layer=POLY_cond $X=2.45 $Y=1.225
+ $X2=2.455 $Y2=1.117
r96 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.45 $Y=1.225 $X2=2.45
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_620_911# 1 2 3 10
+ 11 12 17 18 20 24 29 31 32 34 38 40 41 44 48 49 53 56 57 60 62 63
c127 60 0 1.02426e-19 $X=4.555 $Y=1.79
c128 44 0 7.14482e-20 $X=4.1 $Y=4.735
c129 38 0 9.26578e-20 $X=3.24 $Y=4.735
c130 31 0 8.23968e-20 $X=4.78 $Y=2.94
c131 24 0 9.10198e-20 $X=5.085 $Y=4.88
c132 18 0 1.25592e-19 $X=5.16 $Y=2.94
c133 11 0 1.76914e-21 $X=4.27 $Y=2.94
c134 10 0 7.64702e-20 $X=4.705 $Y=2.94
r135 58 60 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.555 $Y=2.745
+ $X2=4.555 $Y2=1.79
r136 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.47 $Y=2.83
+ $X2=4.555 $Y2=2.745
r137 56 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.47 $Y=2.83
+ $X2=4.19 $Y2=2.83
r138 54 63 10.0555 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.105 $Y=4.045
+ $X2=4.105 $Y2=3.97
r139 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=3.975 $X2=4.105 $Y2=3.975
r140 51 62 3.70735 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.105 $Y=4.155
+ $X2=3.935 $Y2=4.155
r141 51 53 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.105 $Y=4.155
+ $X2=4.105 $Y2=3.975
r142 49 63 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=4.105 $Y=3.135
+ $X2=4.105 $Y2=3.97
r143 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=3.135 $X2=4.105 $Y2=3.135
r144 46 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.915
+ $X2=4.19 $Y2=2.83
r145 46 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.105 $Y=2.915
+ $X2=4.105 $Y2=3.135
r146 42 62 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=4.1 $Y=4.325
+ $X2=3.935 $Y2=4.155
r147 42 44 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.1 $Y=4.325
+ $X2=4.1 $Y2=4.735
r148 40 62 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=4.24
+ $X2=3.935 $Y2=4.155
r149 40 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.935 $Y=4.24
+ $X2=3.405 $Y2=4.24
r150 36 41 17.4739 $w=1.11e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.24 $Y=4.325
+ $X2=3.405 $Y2=4.24
r151 36 38 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.24 $Y=4.325
+ $X2=3.24 $Y2=4.735
r152 33 34 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.085 $Y=4.045
+ $X2=5.235 $Y2=4.045
r153 30 49 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.105 $Y=3.015
+ $X2=4.105 $Y2=3.135
r154 27 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.235 $Y=3.97
+ $X2=5.235 $Y2=4.045
r155 27 29 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.235 $Y=3.97
+ $X2=5.235 $Y2=3.485
r156 26 29 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.235 $Y=3.015
+ $X2=5.235 $Y2=3.485
r157 22 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.085 $Y=4.12
+ $X2=5.085 $Y2=4.045
r158 22 24 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.085 $Y=4.12
+ $X2=5.085 $Y2=4.88
r159 21 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=4.045
+ $X2=4.78 $Y2=4.045
r160 20 33 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.01 $Y=4.045
+ $X2=5.085 $Y2=4.045
r161 20 21 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.01 $Y=4.045
+ $X2=4.855 $Y2=4.045
r162 19 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=2.94
+ $X2=4.78 $Y2=2.94
r163 18 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.16 $Y=2.94
+ $X2=5.235 $Y2=3.015
r164 18 19 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=5.16 $Y=2.94
+ $X2=4.855 $Y2=2.94
r165 15 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=3.97
+ $X2=4.78 $Y2=4.045
r166 15 17 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.78 $Y=3.97
+ $X2=4.78 $Y2=3.485
r167 14 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=3.015
+ $X2=4.78 $Y2=2.94
r168 14 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.78 $Y=3.015 $X2=4.78
+ $Y2=3.485
r169 13 54 22.122 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=4.045
+ $X2=4.105 $Y2=4.045
r170 12 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=4.045
+ $X2=4.78 $Y2=4.045
r171 12 13 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=4.045
+ $X2=4.27 $Y2=4.045
r172 11 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.27 $Y=2.94
+ $X2=4.105 $Y2=3.015
r173 10 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=2.94
+ $X2=4.78 $Y2=2.94
r174 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=2.94
+ $X2=4.27 $Y2=2.94
r175 3 60 300 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.56 $X2=4.555 $Y2=1.79
r176 2 44 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.96 $Y=4.555
+ $X2=4.1 $Y2=4.735
r177 1 38 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.1 $Y=4.555
+ $X2=3.24 $Y2=4.735
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_1032_911# 1 2 9
+ 11 13 14 18 23 25 26 30 35 36 38 40 45 46 51 52 55 59 62 65
c102 55 0 9.10198e-20 $X=5.455 $Y=3.235
c103 11 0 1.02426e-19 $X=5.255 $Y=1.41
r104 62 64 12.4159 $w=4.52e-07 $l=4.6e-07 $layer=LI1_cond $X=5.45 $Y=4.24
+ $X2=5.45 $Y2=4.7
r105 60 65 19.468 $w=3.59e-07 $l=1.45e-07 $layer=POLY_cond $X=5.92 $Y=4.195
+ $X2=5.775 $Y2=4.195
r106 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.92
+ $Y=4.21 $X2=5.92 $Y2=4.21
r107 57 62 4.69682 $w=2.3e-07 $l=3.15e-07 $layer=LI1_cond $X=5.765 $Y=4.24
+ $X2=5.45 $Y2=4.24
r108 57 59 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.765 $Y=4.24
+ $X2=5.92 $Y2=4.24
r109 53 62 7.30083 $w=4.52e-07 $l=1.17473e-07 $layer=LI1_cond $X=5.455 $Y=4.125
+ $X2=5.45 $Y2=4.24
r110 53 55 51.9522 $w=1.88e-07 $l=8.9e-07 $layer=LI1_cond $X=5.455 $Y=4.125
+ $X2=5.455 $Y2=3.235
r111 43 45 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=6.635 $Y=2.99
+ $X2=6.635 $Y2=1.985
r112 42 45 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.635 $Y=1.41
+ $X2=6.635 $Y2=1.985
r113 38 42 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=6.635 $Y=1.247
+ $X2=6.635 $Y2=1.41
r114 38 40 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.635 $Y=1.085
+ $X2=6.635 $Y2=0.56
r115 37 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.28 $Y=3.065
+ $X2=6.205 $Y2=3.065
r116 36 43 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.56 $Y=3.065
+ $X2=6.635 $Y2=2.99
r117 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.56 $Y=3.065
+ $X2=6.28 $Y2=3.065
r118 33 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.205 $Y=2.99
+ $X2=6.205 $Y2=3.065
r119 33 35 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=6.205 $Y=2.99
+ $X2=6.205 $Y2=1.985
r120 32 35 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.985
r121 28 38 76.3471 $w=3.25e-07 $l=4.3e-07 $layer=POLY_cond $X=6.205 $Y=1.247
+ $X2=6.635 $Y2=1.247
r122 28 32 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=6.205 $Y=1.247
+ $X2=6.205 $Y2=1.41
r123 28 30 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.205 $Y=1.085
+ $X2=6.205 $Y2=0.56
r124 27 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.85 $Y=3.065
+ $X2=5.775 $Y2=3.065
r125 26 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.13 $Y=3.065
+ $X2=6.205 $Y2=3.065
r126 26 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.13 $Y=3.065
+ $X2=5.85 $Y2=3.065
r127 25 65 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.775 $Y=4.015
+ $X2=5.775 $Y2=4.195
r128 24 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.775 $Y=3.14
+ $X2=5.775 $Y2=3.065
r129 24 25 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=5.775 $Y=3.14
+ $X2=5.775 $Y2=4.015
r130 21 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.775 $Y=2.99
+ $X2=5.775 $Y2=3.065
r131 21 23 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=5.775 $Y=2.99
+ $X2=5.775 $Y2=1.985
r132 20 23 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.775 $Y=1.41
+ $X2=5.775 $Y2=1.985
r133 16 28 76.3471 $w=3.25e-07 $l=4.3e-07 $layer=POLY_cond $X=5.775 $Y=1.247
+ $X2=6.205 $Y2=1.247
r134 16 20 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=5.775 $Y=1.247
+ $X2=5.775 $Y2=1.41
r135 16 18 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.775 $Y=1.085
+ $X2=5.775 $Y2=0.56
r136 15 46 4.85217 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.247
+ $X2=5.255 $Y2=1.247
r137 14 16 13.3164 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=5.7 $Y=1.247
+ $X2=5.775 $Y2=1.247
r138 14 15 65.694 $w=3.25e-07 $l=3.7e-07 $layer=POLY_cond $X=5.7 $Y=1.247
+ $X2=5.33 $Y2=1.247
r139 11 46 36.6911 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=5.255 $Y=1.41
+ $X2=5.255 $Y2=1.247
r140 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.255 $Y=1.41
+ $X2=5.255 $Y2=1.985
r141 7 46 36.6911 $w=1.5e-07 $l=1.62e-07 $layer=POLY_cond $X=5.255 $Y=1.085
+ $X2=5.255 $Y2=1.247
r142 7 9 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.255 $Y=1.085
+ $X2=5.255 $Y2=0.56
r143 2 55 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.31
+ $Y=3.09 $X2=5.455 $Y2=3.235
r144 1 64 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.16
+ $Y=4.555 $X2=5.3 $Y2=4.7
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPWR 1 2 3 4 15 19
+ 23 27 30 32 33 35 36 37 44 54 55 62
c108 30 0 1.90316e-19 $X=5.005 $Y=2.72
r109 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r110 52 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r111 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r112 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r113 49 62 0.611765 $w=4.8e-07 $l=2.15e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.6 $Y2=2.72
r114 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 41 45 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r117 40 44 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r118 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r119 37 62 0.13658 $w=4.8e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=2.72
+ $X2=3.6 $Y2=2.72
r120 37 45 0.429658 $w=4.8e-07 $l=1.51e-06 $layer=MET1_cond $X=3.12 $Y=2.72
+ $X2=1.61 $Y2=2.72
r121 35 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=2.72
+ $X2=6.67 $Y2=2.72
r122 35 36 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.755 $Y=2.72
+ $X2=6.845 $Y2=2.72
r123 34 54 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.935 $Y=2.72
+ $X2=7.13 $Y2=2.72
r124 34 36 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.935 $Y=2.72
+ $X2=6.845 $Y2=2.72
r125 32 48 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.75 $Y2=2.72
r126 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.99 $Y2=2.72
r127 31 51 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=6.67 $Y2=2.72
r128 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=5.99 $Y2=2.72
r129 29 48 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.75 $Y2=2.72
r130 29 30 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.005 $Y2=2.72
r131 25 36 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=2.635
+ $X2=6.845 $Y2=2.72
r132 25 27 52.0657 $w=1.78e-07 $l=8.45e-07 $layer=LI1_cond $X=6.845 $Y=2.635
+ $X2=6.845 $Y2=1.79
r133 21 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=2.635
+ $X2=5.99 $Y2=2.72
r134 21 23 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.99 $Y=2.635
+ $X2=5.99 $Y2=1.79
r135 17 30 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.805
+ $X2=5.005 $Y2=2.72
r136 17 19 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.005 $Y=2.805
+ $X2=5.005 $Y2=3.235
r137 13 30 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.635
+ $X2=5.005 $Y2=2.72
r138 13 15 42.3398 $w=2.28e-07 $l=8.45e-07 $layer=LI1_cond $X=5.005 $Y=2.635
+ $X2=5.005 $Y2=1.79
r139 4 27 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=6.71
+ $Y=1.485 $X2=6.85 $Y2=1.79
r140 3 23 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=5.85
+ $Y=1.485 $X2=5.99 $Y2=1.79
r141 2 15 300 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.56 $X2=5.005 $Y2=1.79
r142 1 19 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=3.09 $X2=5.005 $Y2=3.235
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%X 1 2 3 4 15 17 21
+ 25 27 28 29 33 35
r43 33 35 0.628605 $w=2.73e-07 $l=1.5e-08 $layer=LI1_cond $X=5.497 $Y=1.41
+ $X2=5.497 $Y2=1.425
r44 29 33 1.51957 $w=2.81e-07 $l=4.05586e-08 $layer=LI1_cond $X=5.485 $Y=1.375
+ $X2=5.497 $Y2=1.41
r45 29 38 13.8293 $w=2.73e-07 $l=3.3e-07 $layer=LI1_cond $X=5.497 $Y=1.46
+ $X2=5.497 $Y2=1.79
r46 29 35 1.46675 $w=2.73e-07 $l=3.5e-08 $layer=LI1_cond $X=5.497 $Y=1.46
+ $X2=5.497 $Y2=1.425
r47 23 27 6.43939 $w=2.47e-07 $l=1.75442e-07 $layer=LI1_cond $X=6.445 $Y=1.085
+ $X2=6.417 $Y2=1.247
r48 23 25 34.8352 $w=2.18e-07 $l=6.65e-07 $layer=LI1_cond $X=6.445 $Y=1.085
+ $X2=6.445 $Y2=0.42
r49 19 27 6.43939 $w=2.47e-07 $l=1.63e-07 $layer=LI1_cond $X=6.417 $Y=1.41
+ $X2=6.417 $Y2=1.247
r50 19 21 15.9247 $w=2.73e-07 $l=3.8e-07 $layer=LI1_cond $X=6.417 $Y=1.41
+ $X2=6.417 $Y2=1.79
r51 18 29 5.5573 $w=2.81e-07 $l=1.28e-07 $layer=LI1_cond $X=5.485 $Y=1.247
+ $X2=5.485 $Y2=1.375
r52 18 28 8.33594 $w=2.81e-07 $l=1.92e-07 $layer=LI1_cond $X=5.485 $Y=1.247
+ $X2=5.485 $Y2=1.055
r53 17 27 0.38261 $w=3.25e-07 $l=1.37e-07 $layer=LI1_cond $X=6.28 $Y=1.247
+ $X2=6.417 $Y2=1.247
r54 17 18 22.8716 $w=3.23e-07 $l=6.45e-07 $layer=LI1_cond $X=6.28 $Y=1.247
+ $X2=5.635 $Y2=1.247
r55 13 28 9.21519 $w=3e-07 $l=2.25e-07 $layer=LI1_cond $X=5.485 $Y=0.83
+ $X2=5.485 $Y2=1.055
r56 13 15 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=5.485 $Y=0.83
+ $X2=5.485 $Y2=0.42
r57 4 21 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=6.28
+ $Y=1.485 $X2=6.42 $Y2=1.79
r58 3 38 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=5.33
+ $Y=1.485 $X2=5.47 $Y2=1.79
r59 2 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.235 $X2=6.42 $Y2=0.42
r60 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.33
+ $Y=0.235 $X2=5.47 $Y2=0.42
.ends


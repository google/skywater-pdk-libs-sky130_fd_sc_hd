* File: sky130_fd_sc_hd__nand2_2.pxi.spice
* Created: Thu Aug 27 14:28:43 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2_2%B N_B_c_41_n N_B_M1002_g N_B_M1001_g N_B_c_42_n
+ N_B_M1007_g N_B_M1005_g B B N_B_c_44_n PM_SKY130_FD_SC_HD__NAND2_2%B
x_PM_SKY130_FD_SC_HD__NAND2_2%A N_A_c_86_n N_A_M1003_g N_A_M1000_g N_A_c_87_n
+ N_A_M1004_g N_A_M1006_g A A N_A_c_89_n PM_SKY130_FD_SC_HD__NAND2_2%A
x_PM_SKY130_FD_SC_HD__NAND2_2%VPWR N_VPWR_M1001_d N_VPWR_M1005_d N_VPWR_M1006_s
+ N_VPWR_c_132_n N_VPWR_c_133_n N_VPWR_c_134_n N_VPWR_c_135_n N_VPWR_c_136_n
+ N_VPWR_c_137_n N_VPWR_c_138_n VPWR N_VPWR_c_139_n N_VPWR_c_131_n
+ PM_SKY130_FD_SC_HD__NAND2_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND2_2%Y N_Y_M1003_s N_Y_M1001_s N_Y_M1000_d N_Y_c_171_n
+ N_Y_c_175_n N_Y_c_177_n N_Y_c_166_n N_Y_c_178_n N_Y_c_188_n N_Y_c_190_n Y Y Y
+ N_Y_c_168_n N_Y_c_170_n PM_SKY130_FD_SC_HD__NAND2_2%Y
x_PM_SKY130_FD_SC_HD__NAND2_2%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1007_d
+ N_A_27_47#_M1004_d N_A_27_47#_c_219_n N_A_27_47#_c_225_n N_A_27_47#_c_220_n
+ N_A_27_47#_c_231_n N_A_27_47#_c_221_n N_A_27_47#_c_222_n N_A_27_47#_c_236_n
+ PM_SKY130_FD_SC_HD__NAND2_2%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND2_2%VGND N_VGND_M1002_s N_VGND_c_261_n VGND
+ N_VGND_c_262_n N_VGND_c_263_n N_VGND_c_264_n N_VGND_c_265_n
+ PM_SKY130_FD_SC_HD__NAND2_2%VGND
cc_1 VNB N_B_c_41_n 0.0219013f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B_c_42_n 0.0161962f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB B 0.0134006f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_B_c_44_n 0.0377472f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_A_c_86_n 0.0161344f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_A_c_87_n 0.0191995f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_7 VNB A 0.00404378f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_A_c_89_n 0.0331412f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_9 VNB N_VPWR_c_131_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_166_n 0.00400135f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_11 VNB Y 0.0213355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_Y_c_168_n 0.0134647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_219_n 0.0183571f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_14 VNB N_A_27_47#_c_220_n 0.00969418f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_27_47#_c_221_n 0.00152046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_222_n 0.010213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_261_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_18 VNB N_VGND_c_262_n 0.0171188f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_19 VNB N_VGND_c_263_n 0.0385148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_264_n 0.143525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_265_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_22 VPB N_B_M1001_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_23 VPB N_B_M1005_g 0.0188371f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_24 VPB B 0.00508358f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_25 VPB N_B_c_44_n 0.00429053f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_26 VPB N_A_M1000_g 0.0188333f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_27 VPB N_A_M1006_g 0.0219695f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_28 VPB A 0.00214965f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_29 VPB N_A_c_89_n 0.00412921f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_30 VPB N_VPWR_c_132_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_31 VPB N_VPWR_c_133_n 0.0426387f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_32 VPB N_VPWR_c_134_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_135_n 0.0131373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_136_n 0.0294647f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_35 VPB N_VPWR_c_137_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_138_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_37 VPB N_VPWR_c_139_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_131_n 0.0464077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB Y 0.0101999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_Y_c_170_n 0.0125556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 N_B_c_42_n N_A_c_86_n 0.0195944f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_42 N_B_M1005_g N_A_M1000_g 0.0195944f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_43 B A 0.0221072f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_44 N_B_c_44_n A 0.00235002f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_45 N_B_c_44_n N_A_c_89_n 0.0195944f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_46 N_B_M1001_g N_VPWR_c_133_n 0.00321781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_47 B N_VPWR_c_133_n 0.0217397f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_48 N_B_M1005_g N_VPWR_c_134_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_49 N_B_M1001_g N_VPWR_c_137_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_50 N_B_M1005_g N_VPWR_c_137_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_51 N_B_M1001_g N_VPWR_c_131_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_52 N_B_M1005_g N_VPWR_c_131_n 0.00952874f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_53 N_B_M1001_g N_Y_c_171_n 0.00229676f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_54 N_B_M1005_g N_Y_c_171_n 8.84614e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_55 B N_Y_c_171_n 0.0213676f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_56 N_B_c_44_n N_Y_c_171_n 0.00209661f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_57 N_B_M1001_g N_Y_c_175_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_58 N_B_M1005_g N_Y_c_175_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_59 N_B_M1005_g N_Y_c_177_n 0.012321f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_60 N_B_M1005_g N_Y_c_178_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_61 N_B_c_41_n N_A_27_47#_c_219_n 0.00620543f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_62 N_B_c_42_n N_A_27_47#_c_219_n 5.19117e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_63 N_B_c_41_n N_A_27_47#_c_225_n 0.00849378f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_64 N_B_c_42_n N_A_27_47#_c_225_n 0.00969737f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_65 B N_A_27_47#_c_225_n 0.0236508f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B_c_44_n N_A_27_47#_c_225_n 0.00218981f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_c_41_n N_A_27_47#_c_220_n 8.92977e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_68 B N_A_27_47#_c_220_n 0.0240047f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_69 N_B_c_42_n N_A_27_47#_c_231_n 0.00244813f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B_c_41_n N_A_27_47#_c_221_n 4.58193e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_71 N_B_c_42_n N_A_27_47#_c_221_n 0.00507693f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B_c_41_n N_VGND_c_261_n 0.00268723f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_73 N_B_c_42_n N_VGND_c_261_n 0.00268723f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B_c_41_n N_VGND_c_262_n 0.00422241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_75 N_B_c_42_n N_VGND_c_263_n 0.00420723f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_76 N_B_c_41_n N_VGND_c_264_n 0.00665076f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_77 N_B_c_42_n N_VGND_c_264_n 0.00573284f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_VPWR_c_134_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_VPWR_c_136_n 0.00321527f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_VPWR_c_139_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_M1006_g N_VPWR_c_139_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_M1000_g N_VPWR_c_131_n 0.00952874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_VPWR_c_131_n 0.0105388f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1000_g N_Y_c_175_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1000_g N_Y_c_177_n 0.0106747f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_86 A N_Y_c_177_n 0.0227961f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_c_86_n N_Y_c_166_n 0.00382511f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_c_87_n N_Y_c_166_n 0.0137866f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_89 A N_Y_c_166_n 0.0305541f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_89_n N_Y_c_166_n 0.00223984f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_M1000_g N_Y_c_178_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_Y_c_178_n 0.0145598f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_Y_c_188_n 0.0129153f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_94 A N_Y_c_188_n 0.00555408f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_M1000_g N_Y_c_190_n 8.84614e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_M1006_g N_Y_c_190_n 8.84614e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_97 A N_Y_c_190_n 0.0213676f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_98 N_A_c_89_n N_Y_c_190_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_c_87_n Y 0.0200131f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_100 A Y 0.0205554f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_101 A N_A_27_47#_c_221_n 0.0126702f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A_c_87_n N_A_27_47#_c_222_n 0.00157861f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_c_86_n N_A_27_47#_c_236_n 0.0103559f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_87_n N_A_27_47#_c_236_n 0.00750429f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_105 A N_A_27_47#_c_236_n 0.00376413f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A_c_86_n N_VGND_c_263_n 0.00357877f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_87_n N_VGND_c_263_n 0.00357877f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_86_n N_VGND_c_264_n 0.00525237f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_c_87_n N_VGND_c_264_n 0.00626241f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_110 N_VPWR_c_131_n N_Y_M1001_s 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_111 N_VPWR_c_131_n N_Y_M1000_d 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_112 N_VPWR_c_137_n N_Y_c_175_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_113 N_VPWR_c_131_n N_Y_c_175_n 0.0122217f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_114 N_VPWR_M1005_d N_Y_c_177_n 0.00332066f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_115 N_VPWR_c_134_n N_Y_c_177_n 0.0126919f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_116 N_VPWR_c_139_n N_Y_c_178_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_117 N_VPWR_c_131_n N_Y_c_178_n 0.0122217f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_118 N_VPWR_M1006_s N_Y_c_188_n 0.00209819f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_119 N_VPWR_c_136_n N_Y_c_188_n 0.0059027f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_120 N_VPWR_M1006_s N_Y_c_170_n 0.00218031f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_121 N_VPWR_c_136_n N_Y_c_170_n 0.0157986f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_122 N_Y_c_166_n N_A_27_47#_M1004_d 7.4958e-19 $X=1.935 $Y=0.78 $X2=0 $Y2=0
cc_123 N_Y_c_168_n N_A_27_47#_M1004_d 0.00241065f $X=2.075 $Y=0.905 $X2=0 $Y2=0
cc_124 N_Y_c_177_n N_A_27_47#_c_225_n 0.00209359f $X=1.355 $Y=1.58 $X2=0 $Y2=0
cc_125 N_Y_c_177_n N_A_27_47#_c_221_n 7.71103e-19 $X=1.355 $Y=1.58 $X2=0 $Y2=0
cc_126 N_Y_c_166_n N_A_27_47#_c_222_n 0.00728545f $X=1.935 $Y=0.78 $X2=0 $Y2=0
cc_127 N_Y_c_168_n N_A_27_47#_c_222_n 0.0135188f $X=2.075 $Y=0.905 $X2=0 $Y2=0
cc_128 N_Y_M1003_s N_A_27_47#_c_236_n 0.00312175f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_129 N_Y_c_166_n N_A_27_47#_c_236_n 0.0192847f $X=1.935 $Y=0.78 $X2=0 $Y2=0
cc_130 N_Y_c_168_n N_VGND_c_263_n 0.00214403f $X=2.075 $Y=0.905 $X2=0 $Y2=0
cc_131 N_Y_M1003_s N_VGND_c_264_n 0.00216833f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_132 N_Y_c_168_n N_VGND_c_264_n 0.00368014f $X=2.075 $Y=0.905 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_225_n N_VGND_M1002_s 0.00312505f $X=0.935 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_27_47#_c_225_n N_VGND_c_261_n 0.012179f $X=0.935 $Y=0.8 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_219_n N_VGND_c_262_n 0.0216446f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_225_n N_VGND_c_262_n 0.0020257f $X=0.935 $Y=0.8 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_225_n N_VGND_c_263_n 0.0020257f $X=0.935 $Y=0.8 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_231_n N_VGND_c_263_n 0.0151813f $X=1.06 $Y=0.465 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_236_n N_VGND_c_263_n 0.0522346f $X=1.775 $Y=0.37 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1002_d N_VGND_c_264_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_M1007_d N_VGND_c_264_n 0.00215206f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_M1004_d N_VGND_c_264_n 0.00209344f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_c_219_n N_VGND_c_264_n 0.012786f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_225_n N_VGND_c_264_n 0.00841425f $X=0.935 $Y=0.8 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_231_n N_VGND_c_264_n 0.0093992f $X=1.06 $Y=0.465 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_236_n N_VGND_c_264_n 0.0329318f $X=1.775 $Y=0.37 $X2=0 $Y2=0

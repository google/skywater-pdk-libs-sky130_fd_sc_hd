* File: sky130_fd_sc_hd__o211ai_4.pex.spice
* Created: Thu Aug 27 14:35:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O211AI_4%A1 1 3 6 8 10 13 15 17 20 24 28 29 34 38 39
+ 41 48 49 52
c118 52 0 1.81301e-19 $X=3.505 $Y=0.995
c119 48 0 1.10361e-19 $X=1.245 $Y=1.16
c120 39 0 2.62618e-20 $X=3.505 $Y=1.16
c121 38 0 1.15388e-19 $X=3.505 $Y=1.16
c122 24 0 6.54703e-20 $X=3.485 $Y=1.985
r123 47 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.245 $Y=1.16
+ $X2=1.335 $Y2=1.16
r124 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.245
+ $Y=1.16 $X2=1.245 $Y2=1.16
r125 41 59 1.81283 $w=4.43e-07 $l=7e-08 $layer=LI1_cond $X=1.187 $Y=1.53
+ $X2=1.187 $Y2=1.6
r126 39 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.16
+ $X2=3.505 $Y2=1.325
r127 39 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.16
+ $X2=3.505 $Y2=0.995
r128 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.505
+ $Y=1.16 $X2=3.505 $Y2=1.16
r129 36 38 14.6113 $w=2.78e-07 $l=3.55e-07 $layer=LI1_cond $X=3.49 $Y=1.515
+ $X2=3.49 $Y2=1.16
r130 35 59 6.43131 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=1.41 $Y=1.6
+ $X2=1.187 $Y2=1.6
r131 34 36 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.35 $Y=1.6
+ $X2=3.49 $Y2=1.515
r132 34 35 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=3.35 $Y=1.6
+ $X2=1.41 $Y2=1.6
r133 32 47 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.905 $Y=1.16
+ $X2=1.245 $Y2=1.16
r134 32 43 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=1.16
+ $X2=0.475 $Y2=1.16
r135 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.905
+ $Y=1.16 $X2=0.905 $Y2=1.16
r136 29 41 8.49441 $w=4.43e-07 $l=3.28e-07 $layer=LI1_cond $X=1.187 $Y=1.202
+ $X2=1.187 $Y2=1.53
r137 29 48 1.0877 $w=4.43e-07 $l=4.2e-08 $layer=LI1_cond $X=1.187 $Y=1.202
+ $X2=1.187 $Y2=1.16
r138 29 31 2.71163 $w=2.53e-07 $l=6e-08 $layer=LI1_cond $X=0.965 $Y=1.202
+ $X2=0.905 $Y2=1.202
r139 28 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.495 $Y=0.56
+ $X2=3.495 $Y2=0.995
r140 24 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.985
+ $X2=3.485 $Y2=1.325
r141 18 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.16
r142 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.985
r143 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=1.16
r144 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=0.56
r145 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r146 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r147 8 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r148 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r149 4 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.16
r150 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.985
r151 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r152 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 36 37
c77 36 0 6.54703e-20 $X=2.89 $Y=1.16
c78 7 0 1.71138e-19 $X=2.195 $Y=0.995
c79 4 0 1.10361e-19 $X=1.765 $Y=1.375
r80 35 37 24.1488 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=1.185
+ $X2=3.055 $Y2=1.185
r81 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.89
+ $Y=1.16 $X2=2.89 $Y2=1.16
r82 33 35 38.7844 $w=3.8e-07 $l=2.65e-07 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.89 $Y2=1.185
r83 32 33 62.9332 $w=3.8e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.625 $Y2=1.185
r84 30 32 47.5658 $w=3.8e-07 $l=3.25e-07 $layer=POLY_cond $X=1.87 $Y=1.185
+ $X2=2.195 $Y2=1.185
r85 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.87
+ $Y=1.16 $X2=1.87 $Y2=1.16
r86 27 30 15.3674 $w=3.8e-07 $l=1.05e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.87 $Y2=1.185
r87 25 36 34.7867 $w=2.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.075 $Y=1.21
+ $X2=2.89 $Y2=1.21
r88 25 31 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.075 $Y=1.21
+ $X2=1.87 $Y2=1.21
r89 22 37 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.055 $Y=1.375
+ $X2=3.055 $Y2=1.185
r90 22 24 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.055 $Y=1.375
+ $X2=3.055 $Y2=1.985
r91 19 37 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.055 $Y=0.995
+ $X2=3.055 $Y2=1.185
r92 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.055 $Y=0.995
+ $X2=3.055 $Y2=0.56
r93 16 33 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.625 $Y=1.375
+ $X2=2.625 $Y2=1.185
r94 16 18 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.625 $Y=1.375
+ $X2=2.625 $Y2=1.985
r95 13 33 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.625 $Y=0.995
+ $X2=2.625 $Y2=1.185
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.625 $Y=0.995
+ $X2=2.625 $Y2=0.56
r97 10 32 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.195 $Y=1.375
+ $X2=2.195 $Y2=1.185
r98 10 12 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.195 $Y=1.375
+ $X2=2.195 $Y2=1.985
r99 7 32 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.195 $Y=0.995
+ $X2=2.195 $Y2=1.185
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.195 $Y=0.995
+ $X2=2.195 $Y2=0.56
r101 4 27 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.765 $Y=1.375
+ $X2=1.765 $Y2=1.185
r102 4 6 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.765 $Y=1.375
+ $X2=1.765 $Y2=1.985
r103 1 27 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.765 $Y=0.995
+ $X2=1.765 $Y2=1.185
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.765 $Y=0.995
+ $X2=1.765 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%B1 1 3 6 8 10 13 15 17 20 24 28 34 38 39 41
+ 50 53 55 58
c116 24 0 1.88107e-20 $X=6.915 $Y=1.985
c117 15 0 1.91217e-19 $X=4.815 $Y=0.995
r118 49 55 9.94584 $w=6.88e-07 $l=4.65e-07 $layer=LI1_cond $X=4.725 $Y=1.34
+ $X2=4.26 $Y2=1.34
r119 48 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.725 $Y=1.16
+ $X2=4.815 $Y2=1.16
r120 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.725
+ $Y=1.16 $X2=4.725 $Y2=1.16
r121 46 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.385 $Y=1.16
+ $X2=4.725 $Y2=1.16
r122 41 58 10.3075 $w=6.88e-07 $l=1.4e-07 $layer=LI1_cond $X=4.835 $Y=1.34
+ $X2=4.975 $Y2=1.34
r123 41 49 1.90679 $w=6.88e-07 $l=1.1e-07 $layer=LI1_cond $X=4.835 $Y=1.34
+ $X2=4.725 $Y2=1.34
r124 39 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.915 $Y=1.16
+ $X2=6.915 $Y2=0.995
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.915
+ $Y=1.16 $X2=6.915 $Y2=1.16
r126 36 38 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.915 $Y=1.515
+ $X2=6.915 $Y2=1.16
r127 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=1.6
+ $X2=6.915 $Y2=1.515
r128 34 58 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=6.83 $Y=1.6
+ $X2=4.975 $Y2=1.6
r129 32 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=4.385 $Y2=1.16
r130 32 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=3.955 $Y2=1.16
r131 31 55 5.97049 $w=4.13e-07 $l=2.15e-07 $layer=LI1_cond $X=4.045 $Y=1.202
+ $X2=4.26 $Y2=1.202
r132 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.045
+ $Y=1.16 $X2=4.045 $Y2=1.16
r133 28 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.965 $Y=0.56
+ $X2=6.965 $Y2=0.995
r134 22 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.915 $Y=1.325
+ $X2=6.915 $Y2=1.16
r135 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.915 $Y=1.325
+ $X2=6.915 $Y2=1.985
r136 18 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.325
+ $X2=4.815 $Y2=1.16
r137 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.815 $Y=1.325
+ $X2=4.815 $Y2=1.985
r138 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=1.16
r139 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=0.56
r140 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=1.325
+ $X2=4.385 $Y2=1.16
r141 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.385 $Y=1.325
+ $X2=4.385 $Y2=1.985
r142 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=1.16
r143 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=0.56
r144 4 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=1.325
+ $X2=3.955 $Y2=1.16
r145 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.955 $Y=1.325
+ $X2=3.955 $Y2=1.985
r146 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=0.995
+ $X2=3.955 $Y2=1.16
r147 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.955 $Y=0.995
+ $X2=3.955 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 44
c79 29 0 1.88107e-20 $X=6.215 $Y=1.19
c80 22 0 1.73478e-19 $X=6.495 $Y=0.995
r81 42 44 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.275 $Y=1.16
+ $X2=6.495 $Y2=1.16
r82 40 42 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=6.075 $Y=1.16
+ $X2=6.275 $Y2=1.16
r83 38 40 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.935 $Y=1.16
+ $X2=6.075 $Y2=1.16
r84 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.935
+ $Y=1.16 $X2=5.935 $Y2=1.16
r85 36 38 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.655 $Y=1.16
+ $X2=5.935 $Y2=1.16
r86 35 39 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.595 $Y=1.21
+ $X2=5.935 $Y2=1.21
r87 34 36 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.595 $Y=1.16
+ $X2=5.655 $Y2=1.16
r88 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.595
+ $Y=1.16 $X2=5.595 $Y2=1.16
r89 31 34 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=5.235 $Y=1.16
+ $X2=5.595 $Y2=1.16
r90 29 39 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.215 $Y=1.21
+ $X2=5.935 $Y2=1.21
r91 29 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.275
+ $Y=1.16 $X2=6.275 $Y2=1.16
r92 25 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.495 $Y=1.325
+ $X2=6.495 $Y2=1.16
r93 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.495 $Y=1.325
+ $X2=6.495 $Y2=1.985
r94 22 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.495 $Y=0.995
+ $X2=6.495 $Y2=1.16
r95 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.495 $Y=0.995
+ $X2=6.495 $Y2=0.56
r96 18 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.075 $Y=1.325
+ $X2=6.075 $Y2=1.16
r97 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.075 $Y=1.325
+ $X2=6.075 $Y2=1.985
r98 15 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.075 $Y=0.995
+ $X2=6.075 $Y2=1.16
r99 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.075 $Y=0.995
+ $X2=6.075 $Y2=0.56
r100 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.325
+ $X2=5.655 $Y2=1.16
r101 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.655 $Y=1.325
+ $X2=5.655 $Y2=1.985
r102 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=0.995
+ $X2=5.655 $Y2=1.16
r103 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.655 $Y=0.995
+ $X2=5.655 $Y2=0.56
r104 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=1.325
+ $X2=5.235 $Y2=1.16
r105 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.235 $Y=1.325
+ $X2=5.235 $Y2=1.985
r106 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=1.16
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 38 42 46
+ 48 50 53 54 55 56 57 59 74 79 88 91 94 98
r123 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r124 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r126 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 83 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r128 83 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.21 $Y2=2.72
r129 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 80 94 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.455 $Y=2.72
+ $X2=6.287 $Y2=2.72
r131 80 82 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.455 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 79 97 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=7.355 $Y=2.72
+ $X2=7.587 $Y2=2.72
r133 79 82 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.355 $Y=2.72
+ $X2=7.13 $Y2=2.72
r134 78 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r135 78 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r136 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 75 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=2.72
+ $X2=5.445 $Y2=2.72
r138 75 77 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.61 $Y=2.72
+ $X2=5.75 $Y2=2.72
r139 74 94 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=6.12 $Y=2.72
+ $X2=6.287 $Y2=2.72
r140 74 77 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.12 $Y=2.72
+ $X2=5.75 $Y2=2.72
r141 73 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r142 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r143 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r144 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r145 67 70 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r146 67 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r147 66 69 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r148 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 64 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.12 $Y2=2.72
r150 64 66 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 63 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r152 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r153 60 85 4.46799 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r154 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 59 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.12 $Y2=2.72
r156 59 62 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.69 $Y2=2.72
r157 57 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r158 57 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r159 55 72 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.37 $Y2=2.72
r160 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.6 $Y2=2.72
r161 53 69 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.45 $Y2=2.72
r162 53 54 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.75 $Y2=2.72
r163 52 72 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.37 $Y2=2.72
r164 52 54 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.75 $Y2=2.72
r165 48 97 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=7.52 $Y=2.635
+ $X2=7.587 $Y2=2.72
r166 48 50 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.52 $Y=2.635
+ $X2=7.52 $Y2=2.36
r167 44 94 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.287 $Y=2.635
+ $X2=6.287 $Y2=2.72
r168 44 46 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=6.287 $Y=2.635
+ $X2=6.287 $Y2=2.36
r169 40 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=2.635
+ $X2=5.445 $Y2=2.72
r170 40 42 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.445 $Y=2.635
+ $X2=5.445 $Y2=2.36
r171 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=2.72
+ $X2=4.6 $Y2=2.72
r172 38 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.28 $Y=2.72
+ $X2=5.445 $Y2=2.72
r173 38 39 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.28 $Y=2.72
+ $X2=4.765 $Y2=2.72
r174 34 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=2.635 $X2=4.6
+ $Y2=2.72
r175 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.6 $Y=2.635
+ $X2=4.6 $Y2=2.36
r176 30 54 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=2.635
+ $X2=3.75 $Y2=2.72
r177 30 32 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.75 $Y=2.635
+ $X2=3.75 $Y2=2.36
r178 26 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r179 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.36
r180 22 85 3.00953 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.192 $Y2=2.72
r181 22 24 31.448 $w=2.93e-07 $l=8.05e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.237 $Y2=1.83
r182 7 50 600 $w=1.7e-07 $l=1.10877e-06 $layer=licon1_PDIFF $count=1 $X=6.99
+ $Y=1.485 $X2=7.52 $Y2=2.36
r183 6 46 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=6.15
+ $Y=1.485 $X2=6.285 $Y2=2.36
r184 5 42 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=5.31
+ $Y=1.485 $X2=5.445 $Y2=2.36
r185 4 36 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.485 $X2=4.6 $Y2=2.36
r186 3 32 600 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.72 $Y2=2.36
r187 2 28 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=2.36
r188 1 24 300 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%A_110_297# 1 2 3 4 13 19 23 27
c38 4 0 1.10358e-19 $X=3.13 $Y=1.485
r39 21 23 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=2.41 $Y=2.37 $X2=3.27
+ $Y2=2.37
r40 19 21 45.2392 $w=1.88e-07 $l=7.75e-07 $layer=LI1_cond $X=1.635 $Y=2.37
+ $X2=2.41 $Y2=2.37
r41 16 19 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.545 $Y=2.275
+ $X2=1.635 $Y2=2.37
r42 16 18 7.08586 $w=1.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.545 $Y=2.275
+ $X2=1.545 $Y2=2.16
r43 15 18 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.545 $Y=2.105
+ $X2=1.545 $Y2=2.16
r44 14 27 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.775 $Y=2.02
+ $X2=0.665 $Y2=2.02
r45 13 15 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.455 $Y=2.02
+ $X2=1.545 $Y2=2.105
r46 13 14 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.455 $Y=2.02
+ $X2=0.775 $Y2=2.02
r47 4 23 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.485 $X2=3.27 $Y2=2.36
r48 3 21 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.485 $X2=2.41 $Y2=2.36
r49 2 18 600 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=2.16
r50 1 27 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2.025
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%Y 1 2 3 4 5 6 7 8 25 33 40 41 42 45 46 47
+ 48 55
c108 45 0 1.10358e-19 $X=3.47 $Y=1.98
c109 33 0 1.91217e-19 $X=6.565 $Y=0.36
c110 25 0 2.62618e-20 $X=3.345 $Y=1.98
r111 59 61 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=5.865 $Y=1.98
+ $X2=6.705 $Y2=1.98
r112 57 59 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=5.025 $Y=1.98
+ $X2=5.865 $Y2=1.98
r113 54 57 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=4.17 $Y=1.98
+ $X2=5.025 $Y2=1.98
r114 54 55 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.17 $Y=1.98
+ $X2=4.045 $Y2=1.98
r115 51 61 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=7.425 $Y=1.98
+ $X2=6.705 $Y2=1.98
r116 48 51 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=7.595 $Y=1.98
+ $X2=7.425 $Y2=1.98
r117 48 51 0.820838 $w=5.08e-07 $l=3.5e-08 $layer=LI1_cond $X=7.425 $Y=1.82
+ $X2=7.425 $Y2=1.855
r118 46 48 5.27682 $w=5.08e-07 $l=2.25e-07 $layer=LI1_cond $X=7.425 $Y=1.595
+ $X2=7.425 $Y2=1.82
r119 46 47 11.2893 $w=5.08e-07 $l=2.55e-07 $layer=LI1_cond $X=7.425 $Y=1.595
+ $X2=7.425 $Y2=1.34
r120 45 55 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.47 $Y=1.94
+ $X2=4.045 $Y2=1.94
r121 43 47 31.7323 $w=1.78e-07 $l=5.15e-07 $layer=LI1_cond $X=7.26 $Y=0.825
+ $X2=7.26 $Y2=1.34
r122 41 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.17 $Y=0.74
+ $X2=7.26 $Y2=0.825
r123 41 42 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.17 $Y=0.74
+ $X2=6.735 $Y2=0.74
r124 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.65 $Y=0.655
+ $X2=6.735 $Y2=0.74
r125 39 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.65 $Y=0.45
+ $X2=6.65 $Y2=0.655
r126 35 38 51.7576 $w=1.78e-07 $l=8.4e-07 $layer=LI1_cond $X=5.445 $Y=0.36
+ $X2=6.285 $Y2=0.36
r127 33 39 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.565 $Y=0.36
+ $X2=6.65 $Y2=0.45
r128 33 38 17.2525 $w=1.78e-07 $l=2.8e-07 $layer=LI1_cond $X=6.565 $Y=0.36
+ $X2=6.285 $Y2=0.36
r129 27 30 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=1.98 $Y=1.98
+ $X2=2.84 $Y2=1.98
r130 25 45 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=1.98
+ $X2=3.47 $Y2=1.98
r131 25 30 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=3.345 $Y=1.98
+ $X2=2.84 $Y2=1.98
r132 8 61 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=1.485 $X2=6.705 $Y2=1.94
r133 7 59 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=5.73
+ $Y=1.485 $X2=5.865 $Y2=1.94
r134 6 57 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.485 $X2=5.025 $Y2=1.94
r135 5 54 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.485 $X2=4.17 $Y2=1.94
r136 4 30 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.84 $Y2=1.94
r137 3 27 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.485 $X2=1.98 $Y2=1.94
r138 2 38 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=6.15
+ $Y=0.235 $X2=6.285 $Y2=0.365
r139 1 35 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=5.31
+ $Y=0.235 $X2=5.445 $Y2=0.365
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%noxref_10 1 2 3 4 5 6 7 22 26 32 38 40 42
+ 49 50 51 52 53 54 57 60 70
c140 53 0 1.15388e-19 $X=7.45 $Y=0.51
c141 51 0 1.71138e-19 $X=1.795 $Y=0.765
c142 42 0 1.73478e-19 $X=7.51 $Y=0.395
r143 61 70 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.595 $Y=0.51
+ $X2=7.595 $Y2=0.395
r144 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=0.51
+ $X2=7.595 $Y2=0.51
r145 57 66 10.7204 $w=2.13e-07 $l=2e-07 $layer=LI1_cond $X=1.132 $Y=0.51
+ $X2=1.132 $Y2=0.71
r146 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=0.51
+ $X2=1.155 $Y2=0.51
r147 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=0.51
+ $X2=1.155 $Y2=0.51
r148 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=0.51
+ $X2=7.595 $Y2=0.51
r149 53 54 7.61137 $w=1.4e-07 $l=6.15e-06 $layer=MET1_cond $X=7.45 $Y=0.51
+ $X2=1.3 $Y2=0.51
r150 50 51 1.17044 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=1.775 $Y=0.765
+ $X2=1.795 $Y2=0.765
r151 47 49 3.66807 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.26 $Y=0.72
+ $X2=0.355 $Y2=0.72
r152 42 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=0.395
+ $X2=7.595 $Y2=0.395
r153 42 44 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.51 $Y=0.395
+ $X2=7.18 $Y2=0.395
r154 38 40 42.4227 $w=1.98e-07 $l=7.65e-07 $layer=LI1_cond $X=3.835 $Y=0.355
+ $X2=4.6 $Y2=0.355
r155 35 37 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.72 $Y=0.625
+ $X2=3.72 $Y2=0.495
r156 34 38 6.85974 $w=2e-07 $l=1.57242e-07 $layer=LI1_cond $X=3.72 $Y=0.455
+ $X2=3.835 $Y2=0.355
r157 34 37 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=3.72 $Y=0.455
+ $X2=3.72 $Y2=0.495
r158 32 35 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.605 $Y=0.71
+ $X2=3.72 $Y2=0.625
r159 32 52 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=0.71
+ $X2=3.13 $Y2=0.71
r160 29 31 41.2959 $w=2.38e-07 $l=8.6e-07 $layer=LI1_cond $X=1.98 $Y=0.745
+ $X2=2.84 $Y2=0.745
r161 29 51 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=1.98 $Y=0.745
+ $X2=1.795 $Y2=0.745
r162 26 52 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.01 $Y=0.745
+ $X2=3.13 $Y2=0.745
r163 26 31 8.16314 $w=2.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.01 $Y=0.745
+ $X2=2.84 $Y2=0.745
r164 25 68 0.859579 $w=2.1e-07 $l=1.08e-07 $layer=LI1_cond $X=1.24 $Y=0.8
+ $X2=1.132 $Y2=0.8
r165 25 50 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=1.24 $Y=0.8
+ $X2=1.775 $Y2=0.8
r166 22 68 1.87607 $w=2.13e-07 $l=3.5e-08 $layer=LI1_cond $X=1.132 $Y=0.765
+ $X2=1.132 $Y2=0.8
r167 22 66 2.94811 $w=2.13e-07 $l=5.5e-08 $layer=LI1_cond $X=1.132 $Y=0.765
+ $X2=1.132 $Y2=0.71
r168 22 49 27.5763 $w=2.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=0.765
+ $X2=0.355 $Y2=0.765
r169 7 44 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.04
+ $Y=0.235 $X2=7.18 $Y2=0.395
r170 6 40 182 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.235 $X2=4.6 $Y2=0.365
r171 5 37 182 $w=1.7e-07 $l=3.26497e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.72 $Y2=0.495
r172 4 31 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.71
r173 3 29 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.71
r174 2 66 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.71
r175 1 47 182 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
r124 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r125 59 60 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r126 57 60 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=7.59
+ $Y2=0
r127 56 59 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=7.59
+ $Y2=0
r128 56 57 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r129 54 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r130 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r131 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r132 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r133 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r134 48 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r135 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r136 45 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r137 45 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.15
+ $Y2=0
r138 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r139 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r140 38 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r141 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r142 36 53 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.105 $Y=0
+ $X2=2.99 $Y2=0
r143 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.27
+ $Y2=0
r144 35 56 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.45
+ $Y2=0
r145 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.27
+ $Y2=0
r146 33 50 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.07 $Y2=0
r147 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.41
+ $Y2=0
r148 32 53 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.575 $Y=0
+ $X2=2.99 $Y2=0
r149 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.41
+ $Y2=0
r150 30 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.15 $Y2=0
r151 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.55
+ $Y2=0
r152 29 50 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.635 $Y=0
+ $X2=2.07 $Y2=0
r153 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.55
+ $Y2=0
r154 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0
r155 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0.36
r156 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0
r157 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0.36
r158 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r159 17 19 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.36
r160 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r161 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.36
r162 4 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.36
r163 3 23 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.36
r164 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.36
r165 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_4%noxref_12 1 2 11
c23 11 0 1.81301e-19 $X=5.865 $Y=0.725
r24 8 11 104.439 $w=1.78e-07 $l=1.695e-06 $layer=LI1_cond $X=4.17 $Y=0.725
+ $X2=5.865 $Y2=0.725
r25 2 11 182 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_NDIFF $count=1 $X=5.73
+ $Y=0.235 $X2=5.865 $Y2=0.725
r26 1 8 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.235 $X2=4.17 $Y2=0.73
.ends


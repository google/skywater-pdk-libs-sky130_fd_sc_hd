* File: sky130_fd_sc_hd__einvp_1.spice
* Created: Thu Aug 27 14:20:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__einvp_1.pex.spice"
.subckt sky130_fd_sc_hd__einvp_1  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_TE_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 A_204_47# N_TE_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.235625 AS=0.11785 PD=1.375 PS=1.18458 NRD=56.76 NRS=9.228 M=1 R=4.33333
+ SA=75000.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1000 N_Z_M1000_d N_A_M1000_g A_204_47# VNB NSHORT L=0.15 W=0.65 AD=0.1755
+ AS=0.235625 PD=1.84 PS=1.375 NRD=0 NRS=56.76 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_TE_M1003_g N_A_27_47#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.189739 AS=0.1092 PD=0.996761 PS=1.36 NRD=2.3443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 A_276_297# N_A_27_47#_M1002_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1825 AS=0.451761 PD=1.365 PS=2.37324 NRD=25.0978 NRS=11.8003 M=1
+ R=6.66667 SA=75000.7 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g A_276_297# VPB PHIGHVT L=0.15 W=1 AD=0.27
+ AS=0.1825 PD=2.54 PS=1.365 NRD=0.9653 NRS=25.0978 M=1 R=6.66667 SA=75001.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__einvp_1.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__and3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.470000 1.245000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 2.125000 1.370000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.305000 1.295000 0.750000 ;
        RECT 1.065000 0.750000 1.475000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 1.795000 2.245000 2.465000 ;
        RECT 1.980000 0.255000 2.230000 0.715000 ;
        RECT 2.060000 0.715000 2.230000 0.925000 ;
        RECT 2.060000 0.925000 2.675000 1.445000 ;
        RECT 2.075000 1.445000 2.245000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.760000 0.085000 ;
        RECT 1.475000  0.085000 1.805000 0.580000 ;
        RECT 2.400000  0.085000 2.675000 0.745000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.760000 2.805000 ;
        RECT 0.085000 2.130000 0.715000 2.635000 ;
        RECT 0.525000 1.765000 0.855000 1.955000 ;
        RECT 0.525000 1.955000 0.715000 2.130000 ;
        RECT 1.555000 1.790000 1.770000 2.635000 ;
        RECT 2.415000 1.625000 2.675000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.100000 1.425000 1.890000 1.595000 ;
      RECT 0.100000 1.595000 0.355000 1.960000 ;
      RECT 0.105000 0.305000 0.895000 0.570000 ;
      RECT 0.640000 0.570000 0.895000 1.425000 ;
      RECT 1.080000 1.595000 1.330000 1.890000 ;
      RECT 1.660000 0.995000 1.890000 1.425000 ;
  END
END sky130_fd_sc_hd__and3_2
END LIBRARY

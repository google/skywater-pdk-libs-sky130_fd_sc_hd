* File: sky130_fd_sc_hd__dfsbp_2.spice
* Created: Thu Aug 27 14:15:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dfsbp_2.pex.spice"
.subckt sky130_fd_sc_hd__dfsbp_2  VNB VPB CLK D SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1034 N_VGND_M1034_d N_CLK_M1034_g N_A_27_47#_M1034_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_A_193_47#_M1023_d N_A_27_47#_M1023_g N_VGND_M1034_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_381_47#_M1008_d N_D_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.64
+ AD=0.11968 AS=0.1664 PD=1.2352 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1033 N_A_476_47#_M1033_d N_A_27_47#_M1033_g N_A_381_47#_M1008_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.072 AS=0.06732 PD=0.76 PS=0.6948 NRD=23.328 NRS=16.656 M=1
+ R=2.4 SA=75000.7 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1021 A_586_47# N_A_193_47#_M1021_g N_A_476_47#_M1033_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0618923 AS=0.072 PD=0.692308 PS=0.76 NRD=38.964 NRS=16.656 M=1
+ R=2.4 SA=75001.2 SB=75001.6 A=0.054 P=1.02 MULT=1
MM1026 N_VGND_M1026_d N_A_652_21#_M1026_g A_586_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0722077 PD=0.84 PS=0.807692 NRD=41.424 NRS=33.396 M=1 R=2.8
+ SA=75001.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_796_47# N_SET_B_M1003_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1005 N_A_652_21#_M1005_d N_A_476_47#_M1005_g A_796_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75002.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 A_1056_47# N_A_476_47#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 N_A_1028_413#_M1010_d N_A_193_47#_M1010_g A_1056_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0693 AS=0.0441 PD=0.75 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1013 A_1224_47# N_A_27_47#_M1013_g N_A_1028_413#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0693 PD=0.63 PS=0.75 NRD=14.28 NRS=7.14 M=1 R=2.8
+ SA=75001 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1015 A_1296_47# N_A_1178_261#_M1015_g A_1224_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_1296_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0994875 AS=0.0441 PD=0.88375 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8
+ SA=75001.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1018 N_A_1178_261#_M1018_d N_A_1028_413#_M1018_g N_VGND_M1022_d VNB NSHORT
+ L=0.15 W=0.54 AD=0.1404 AS=0.127912 PD=1.6 PS=1.13625 NRD=0 NRS=21.108 M=1
+ R=3.6 SA=75001.9 SB=75000.2 A=0.081 P=1.38 MULT=1
MM1006 N_Q_N_M1006_d N_A_1028_413#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_Q_N_M1006_d N_A_1028_413#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1036 N_VGND_M1036_d N_A_1028_413#_M1036_g N_A_1870_47#_M1036_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 N_Q_M1002_d N_A_1870_47#_M1002_g N_VGND_M1036_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1027 N_Q_M1002_d N_A_1870_47#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1019 N_VPWR_M1019_d N_CLK_M1019_g N_A_27_47#_M1019_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_381_47#_M1029_d N_D_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1666 AS=0.2184 PD=1.56667 PS=2.2 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1009 N_A_476_47#_M1009_d N_A_193_47#_M1009_g N_A_381_47#_M1029_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.0833 PD=0.69 PS=0.783333 NRD=0 NRS=28.1316 M=1
+ R=2.8 SA=75000.7 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1037 A_562_413# N_A_27_47#_M1037_g N_A_476_47#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0945 AS=0.0567 PD=0.87 PS=0.69 NRD=79.7259 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_652_21#_M1007_g A_562_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0945 PD=0.8 PS=0.87 NRD=21.0987 NRS=79.7259 M=1 R=2.8
+ SA=75001.7 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1031 N_A_652_21#_M1031_d N_SET_B_M1031_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0798 PD=0.69 PS=0.8 NRD=0 NRS=25.7873 M=1 R=2.8
+ SA=75002.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_476_47#_M1024_g N_A_652_21#_M1031_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1016 A_956_413# N_A_476_47#_M1016_g N_VPWR_M1024_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.8 SA=75003.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_A_1028_413#_M1004_d N_A_27_47#_M1004_g A_956_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75003.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1030 A_1136_413# N_A_193_47#_M1030_g N_A_1028_413#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=53.9386 M=1 R=2.8
+ SA=75004 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_1178_261#_M1014_g A_1136_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75004.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_SET_B_M1001_g N_A_1028_413#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.1092 PD=0.78 PS=1.36 NRD=25.7873 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1028 N_A_1178_261#_M1028_d N_A_1028_413#_M1028_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2184 AS=0.1638 PD=2.2 PS=1.56 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_A_1028_413#_M1012_g N_Q_N_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1020_d N_A_1028_413#_M1020_g N_Q_N_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1035 N_VPWR_M1035_d N_A_1028_413#_M1035_g N_A_1870_47#_M1035_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1017 N_Q_M1017_d N_A_1870_47#_M1017_g N_VPWR_M1035_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1032 N_Q_M1017_d N_A_1870_47#_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX38_noxref VNB VPB NWDIODE A=18.3291 P=26.05
c_237 VPB 0 9.39049e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dfsbp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__clkdlybuf4s25_2.pex.spice
* Created: Tue Sep  1 19:00:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A 3 7 9 10 14 15
c33 3 0 9.12156e-20 $X=0.475 $Y=0.445
r34 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.385 $Y2=1.325
r35 14 16 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.385 $Y2=0.97
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.355
+ $Y=1.16 $X2=0.355 $Y2=1.16
r37 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=0.29 $Y=1.19 $X2=0.29
+ $Y2=1.53
r38 9 15 0.843251 $w=4.08e-07 $l=3e-08 $layer=LI1_cond $X=0.29 $Y=1.19 $X2=0.29
+ $Y2=1.16
r39 7 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r40 3 16 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_27_47# 1 2 9 12 16 20 21 22 27 29
+ 31 32 33 37
c69 32 0 5.69314e-20 $X=0.95 $Y=1.16
c70 31 0 1.19159e-19 $X=0.95 $Y=1.16
r71 32 38 33.0434 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.16
+ $X2=0.97 $Y2=1.325
r72 32 37 33.0434 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.16
+ $X2=0.97 $Y2=0.995
r73 31 34 5.23542 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=1.16
+ $X2=0.85 $Y2=1.325
r74 31 33 8.35844 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=1.16
+ $X2=0.85 $Y2=0.995
r75 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r76 27 35 11.3402 $w=3.4e-07 $l=2.9e-07 $layer=LI1_cond $X=0.835 $Y=1.58
+ $X2=0.835 $Y2=1.87
r77 27 34 8.64332 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=0.835 $Y=1.58
+ $X2=0.835 $Y2=1.325
r78 24 33 11.7247 $w=1.73e-07 $l=1.85e-07 $layer=LI1_cond $X=0.752 $Y=0.81
+ $X2=0.752 $Y2=0.995
r79 23 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.22 $Y2=1.87
r80 22 35 2.92482 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.665 $Y=1.87
+ $X2=0.835 $Y2=1.87
r81 22 23 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=1.87
+ $X2=0.345 $Y2=1.87
r82 20 24 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.665 $Y=0.725
+ $X2=0.752 $Y2=0.81
r83 20 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=0.725
+ $X2=0.345 $Y2=0.725
r84 14 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=0.64
+ $X2=0.345 $Y2=0.725
r85 14 16 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.22 $Y=0.64
+ $X2=0.22 $Y2=0.47
r86 12 38 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1 $Y=2.075 $X2=1
+ $Y2=1.325
r87 9 37 83.868 $w=2.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1 $Y=0.56 $X2=1
+ $Y2=0.995
r88 2 29 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
r89 1 16 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_225_47# 1 2 9 11 14 18 20 22 25 28
+ 29 31
c61 31 0 9.12156e-20 $X=1.26 $Y=0.78
c62 28 0 1.18904e-19 $X=2.03 $Y=1.16
r63 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=1.16 $X2=2.03 $Y2=1.16
r64 26 28 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.44 $Y=1.16
+ $X2=2.03 $Y2=1.16
r65 25 26 8.4433 $w=2.42e-07 $l=1.68953e-07 $layer=LI1_cond $X=1.315 $Y=0.995
+ $X2=1.307 $Y2=1.16
r66 25 31 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=1.315 $Y=0.995
+ $X2=1.315 $Y2=0.78
r67 20 26 18.3921 $w=2.65e-07 $l=3.97e-07 $layer=LI1_cond $X=1.307 $Y=1.557
+ $X2=1.307 $Y2=1.16
r68 20 22 11.0026 $w=2.63e-07 $l=2.53e-07 $layer=LI1_cond $X=1.307 $Y=1.557
+ $X2=1.307 $Y2=1.81
r69 16 31 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=0.615
+ $X2=1.26 $Y2=0.78
r70 16 18 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.26 $Y=0.615 $X2=1.26
+ $Y2=0.515
r71 12 29 25.545 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.325
+ $X2=2.04 $Y2=1.16
r72 12 14 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.04 $Y=1.325
+ $X2=2.04 $Y2=2.075
r73 9 29 25.545 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.04 $Y2=1.16
r74 9 11 83.868 $w=2.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.04 $Y2=0.56
r75 2 22 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.125
+ $Y=1.665 $X2=1.26 $Y2=1.81
r76 1 18 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.26 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_331_47# 1 2 9 13 17 21 25 29 31 32
+ 33 34 38 42
c89 42 0 1.42295e-19 $X=3.065 $Y=1.162
c90 38 0 1.70937e-19 $X=2.51 $Y=1.16
r91 41 42 68.661 $w=3.51e-07 $l=5e-07 $layer=POLY_cond $X=2.565 $Y=1.162
+ $X2=3.065 $Y2=1.162
r92 39 41 7.55271 $w=3.51e-07 $l=5.5e-08 $layer=POLY_cond $X=2.51 $Y=1.162
+ $X2=2.565 $Y2=1.162
r93 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.16 $X2=2.51 $Y2=1.16
r94 36 38 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.465 $Y=1.5
+ $X2=2.465 $Y2=1.16
r95 35 38 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=2.465 $Y=0.805
+ $X2=2.465 $Y2=1.16
r96 33 36 6.82432 $w=2.45e-07 $l=1.80997e-07 $layer=LI1_cond $X=2.335 $Y=1.622
+ $X2=2.465 $Y2=1.5
r97 33 34 18.345 $w=2.43e-07 $l=3.9e-07 $layer=LI1_cond $X=2.335 $Y=1.622
+ $X2=1.945 $Y2=1.622
r98 31 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.335 $Y=0.72
+ $X2=2.465 $Y2=0.805
r99 31 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.335 $Y=0.72
+ $X2=1.945 $Y2=0.72
r100 27 34 6.8174 $w=2.45e-07 $l=1.76068e-07 $layer=LI1_cond $X=1.82 $Y=1.745
+ $X2=1.945 $Y2=1.622
r101 27 29 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=1.82 $Y=1.745
+ $X2=1.82 $Y2=1.81
r102 23 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.78 $Y=0.635
+ $X2=1.945 $Y2=0.72
r103 23 25 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.78 $Y=0.635
+ $X2=1.78 $Y2=0.41
r104 19 42 22.6971 $w=1.5e-07 $l=1.78e-07 $layer=POLY_cond $X=3.065 $Y=1.34
+ $X2=3.065 $Y2=1.162
r105 19 21 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.065 $Y=1.34
+ $X2=3.065 $Y2=1.985
r106 15 42 22.6971 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=3.065 $Y=0.985
+ $X2=3.065 $Y2=1.162
r107 15 17 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.065 $Y=0.985
+ $X2=3.065 $Y2=0.445
r108 11 41 22.6971 $w=1.5e-07 $l=1.78e-07 $layer=POLY_cond $X=2.565 $Y=1.34
+ $X2=2.565 $Y2=1.162
r109 11 13 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.565 $Y=1.34
+ $X2=2.565 $Y2=1.985
r110 7 41 22.6971 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=2.565 $Y=0.985
+ $X2=2.565 $Y2=1.162
r111 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.565 $Y=0.985
+ $X2=2.565 $Y2=0.445
r112 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.655
+ $Y=1.665 $X2=1.78 $Y2=1.81
r113 1 25 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.78 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%VPWR 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c50 2 0 1.70937e-19 $X=2.165 $Y=1.665
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 39 47 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.472 $Y2=2.72
r56 39 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=0.74 $Y2=2.72
r64 32 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.74 $Y2=2.72
r66 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 23 37 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.07 $Y2=2.72
r70 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.3 $Y2=2.72
r71 22 41 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.3 $Y2=2.72
r73 18 47 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.472 $Y2=2.72
r74 18 20 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.43 $Y2=1.855
r75 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.635 $X2=2.3
+ $Y2=2.72
r76 14 16 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.3 $Y=2.635
+ $X2=2.3 $Y2=2
r77 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=2.635
+ $X2=0.74 $Y2=2.72
r78 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=2.635
+ $X2=0.74 $Y2=2.34
r79 3 20 300 $w=1.7e-07 $l=4.63249e-07 $layer=licon1_PDIFF $count=2 $X=3.14
+ $Y=1.485 $X2=3.35 $Y2=1.855
r80 2 16 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=2.165
+ $Y=1.665 $X2=2.3 $Y2=2
r81 1 12 600 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.74 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%X 1 2 7 8 10 11 12 26 28 40 55
c35 8 0 1.42295e-19 $X=3.01 $Y=1.19
r36 26 28 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=2.932 $Y=1.79
+ $X2=2.932 $Y2=1.87
r37 24 26 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=2.932 $Y=1.787
+ $X2=2.932 $Y2=1.79
r38 10 24 0.0354598 $w=3.23e-07 $l=1e-09 $layer=LI1_cond $X=2.932 $Y=1.786
+ $X2=2.932 $Y2=1.787
r39 10 55 6.70896 $w=3.23e-07 $l=1.61e-07 $layer=LI1_cond $X=2.932 $Y=1.786
+ $X2=2.932 $Y2=1.625
r40 10 11 12.0209 $w=3.23e-07 $l=3.39e-07 $layer=LI1_cond $X=2.932 $Y=1.871
+ $X2=2.932 $Y2=2.21
r41 10 28 0.0354598 $w=3.23e-07 $l=1e-09 $layer=LI1_cond $X=2.932 $Y=1.871
+ $X2=2.932 $Y2=1.87
r42 8 12 10.7882 $w=5.08e-07 $l=4.6e-07 $layer=LI1_cond $X=3.01 $Y=1.02 $X2=3.47
+ $Y2=1.02
r43 8 45 0.703576 $w=5.08e-07 $l=3e-08 $layer=LI1_cond $X=3.01 $Y=1.02 $X2=2.98
+ $Y2=1.02
r44 8 45 5.41923 $w=2.3e-07 $l=2.55e-07 $layer=LI1_cond $X=2.98 $Y=1.275
+ $X2=2.98 $Y2=1.02
r45 8 45 5.41923 $w=2.3e-07 $l=2.55e-07 $layer=LI1_cond $X=2.98 $Y=0.765
+ $X2=2.98 $Y2=1.02
r46 8 55 11.3371 $w=3.98e-07 $l=3.5e-07 $layer=LI1_cond $X=2.98 $Y=1.275
+ $X2=2.98 $Y2=1.625
r47 8 44 5.57489 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.98 $Y=0.765
+ $X2=2.98 $Y2=0.615
r48 7 44 4.72321 $w=3.23e-07 $l=1.05e-07 $layer=LI1_cond $X=2.932 $Y=0.51
+ $X2=2.932 $Y2=0.615
r49 7 40 2.12759 $w=3.23e-07 $l=6e-08 $layer=LI1_cond $X=2.932 $Y=0.51 $X2=2.932
+ $Y2=0.45
r50 2 26 300 $w=1.7e-07 $l=3.98246e-07 $layer=licon1_PDIFF $count=2 $X=2.64
+ $Y=1.485 $X2=2.855 $Y2=1.79
r51 1 40 182 $w=1.7e-07 $l=3.04056e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.235 $X2=2.855 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%VGND 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c55 12 0 5.69314e-20 $X=0.74 $Y=0.385
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r58 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r59 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r60 39 47 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.472
+ $Y2=0
r61 39 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=2.99
+ $Y2=0
r62 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r63 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r64 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r65 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r66 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r67 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r68 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r69 32 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.15
+ $Y2=0
r70 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r71 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.23
+ $Y2=0
r72 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r73 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r74 23 37 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.07
+ $Y2=0
r75 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.3
+ $Y2=0
r76 22 41 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.99
+ $Y2=0
r77 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.3
+ $Y2=0
r78 18 47 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.472 $Y2=0
r79 18 20 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.43 $Y=0.085 $X2=3.43
+ $Y2=0.385
r80 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.085 $X2=2.3
+ $Y2=0
r81 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.3 $Y=0.085
+ $X2=2.3 $Y2=0.38
r82 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r83 10 12 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0.385
r84 3 20 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=3.14
+ $Y=0.235 $X2=3.35 $Y2=0.385
r85 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.235 $X2=2.3 $Y2=0.38
r86 1 12 182 $w=1.7e-07 $l=2.54165e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.74 $Y2=0.385
.ends


* File: sky130_fd_sc_hd__o21bai_2.spice
* Created: Thu Aug 27 14:36:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21bai_2.pex.spice"
.subckt sky130_fd_sc_hd__o21bai_2  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_A_28_297#_M1005_d N_B1_N_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A_28_297#_M1007_g N_A_229_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1007_d N_A_28_297#_M1009_g N_A_229_47#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1012 N_A_229_47#_M1009_s N_A2_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1013 N_A_229_47#_M1013_d N_A2_M1013_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1001 N_A_229_47#_M1013_d N_A1_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_229_47#_M1002_d N_A1_M1002_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_B1_N_M1006_g N_A_28_297#_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=70.4866 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1006_d N_A_28_297#_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.205282 AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_28_297#_M1011_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_397_297#_M1003_d N_A2_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_A_397_297#_M1004_d N_A2_M1004_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_397_297#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1000_d N_A1_M1010_g N_A_397_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__o21bai_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__or3_1.pxi.spice
* Created: Thu Aug 27 14:43:17 2020
* 
x_PM_SKY130_FD_SC_HD__OR3_1%C N_C_M1004_g N_C_M1003_g C N_C_c_58_n
+ PM_SKY130_FD_SC_HD__OR3_1%C
x_PM_SKY130_FD_SC_HD__OR3_1%B N_B_M1001_g N_B_M1000_g N_B_c_83_n N_B_c_84_n B B
+ N_B_c_86_n N_B_c_87_n PM_SKY130_FD_SC_HD__OR3_1%B
x_PM_SKY130_FD_SC_HD__OR3_1%A N_A_M1005_g N_A_M1007_g A A A N_A_c_124_n
+ N_A_c_125_n N_A_c_126_n PM_SKY130_FD_SC_HD__OR3_1%A
x_PM_SKY130_FD_SC_HD__OR3_1%A_29_53# N_A_29_53#_M1004_s N_A_29_53#_M1000_d
+ N_A_29_53#_M1003_s N_A_29_53#_M1006_g N_A_29_53#_M1002_g N_A_29_53#_c_175_n
+ N_A_29_53#_c_176_n N_A_29_53#_c_177_n N_A_29_53#_c_185_n N_A_29_53#_c_259_p
+ N_A_29_53#_c_178_n N_A_29_53#_c_217_n N_A_29_53#_c_186_n N_A_29_53#_c_187_n
+ N_A_29_53#_c_179_n N_A_29_53#_c_188_n N_A_29_53#_c_180_n N_A_29_53#_c_181_n
+ N_A_29_53#_c_182_n N_A_29_53#_c_183_n PM_SKY130_FD_SC_HD__OR3_1%A_29_53#
x_PM_SKY130_FD_SC_HD__OR3_1%VPWR N_VPWR_M1007_d N_VPWR_c_273_n VPWR
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_272_n N_VPWR_c_277_n VPWR
+ PM_SKY130_FD_SC_HD__OR3_1%VPWR
x_PM_SKY130_FD_SC_HD__OR3_1%X N_X_M1006_d N_X_M1002_d N_X_c_298_n N_X_c_300_n
+ N_X_c_299_n X PM_SKY130_FD_SC_HD__OR3_1%X
x_PM_SKY130_FD_SC_HD__OR3_1%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_c_316_n
+ N_VGND_c_317_n VGND N_VGND_c_318_n N_VGND_c_319_n N_VGND_c_320_n
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n VGND
+ PM_SKY130_FD_SC_HD__OR3_1%VGND
cc_1 VNB N_C_M1004_g 0.0346235f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.475
cc_2 VNB C 0.0123316f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_C_c_58_n 0.0351857f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_4 VNB N_B_M1001_g 0.0163624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_B_c_83_n 0.013575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_B_c_84_n 0.0110772f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_7 VNB N_A_M1005_g 0.0266374f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.475
cc_8 VNB N_A_c_124_n 0.0206834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_c_125_n 0.00216296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_126_n 0.00335991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_29_53#_c_175_n 0.0135183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_29_53#_c_176_n 0.00380326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_29_53#_c_177_n 0.00918699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_29_53#_c_178_n 0.00106516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_29_53#_c_179_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_29_53#_c_180_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_29_53#_c_181_n 0.0234012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_29_53#_c_182_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_29_53#_c_183_n 0.0197196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_272_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_298_n 0.013635f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_22 VNB N_X_c_299_n 0.0241196f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_23 VNB N_VGND_c_316_n 0.00101984f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_24 VNB N_VGND_c_317_n 6.33941e-19 $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_25 VNB N_VGND_c_318_n 0.0151077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_319_n 0.0115649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_320_n 0.0167832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_321_n 0.147339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_322_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_323_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_C_M1003_g 0.025409f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.695
cc_32 VPB C 0.00162495f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_33 VPB N_C_c_58_n 0.00868279f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_34 VPB N_B_M1001_g 0.0242366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_B_c_86_n 0.0370191f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_36 VPB N_B_c_87_n 0.0353191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_M1007_g 0.0214042f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.695
cc_38 VPB A 0.00145597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_c_124_n 0.00403484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_c_125_n 0.00327409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_29_53#_M1002_g 0.0244726f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_42 VPB N_A_29_53#_c_185_n 0.00300673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_29_53#_c_186_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_29_53#_c_187_n 0.0208029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_29_53#_c_188_n 0.00130908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_29_53#_c_181_n 0.00544454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_273_n 0.0125577f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.695
cc_48 VPB N_VPWR_c_274_n 0.0379933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_275_n 0.0178726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_272_n 0.0573406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_277_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_300_n 0.00521594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_X_c_299_n 0.00880306f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_54 VPB X 0.0319967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 C N_B_M1001_g 2.51577e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_56 N_C_c_58_n N_B_M1001_g 0.0395923f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_57 N_C_M1004_g N_B_c_83_n 0.0136742f $X=0.48 $Y=0.475 $X2=0 $Y2=0
cc_58 N_C_M1004_g N_B_c_84_n 0.0395923f $X=0.48 $Y=0.475 $X2=0 $Y2=0
cc_59 N_C_M1003_g N_B_c_87_n 0.00441056f $X=0.48 $Y=1.695 $X2=0 $Y2=0
cc_60 N_C_M1003_g A 0.00420104f $X=0.48 $Y=1.695 $X2=0 $Y2=0
cc_61 C N_A_c_126_n 0.0278765f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_62 N_C_c_58_n N_A_c_126_n 0.00274214f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_63 N_C_M1004_g N_A_29_53#_c_176_n 0.0163464f $X=0.48 $Y=0.475 $X2=0 $Y2=0
cc_64 C N_A_29_53#_c_176_n 0.00550551f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_65 N_C_c_58_n N_A_29_53#_c_176_n 0.00111883f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_66 C N_A_29_53#_c_177_n 0.0211211f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_67 N_C_c_58_n N_A_29_53#_c_177_n 0.00542346f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_68 N_C_M1003_g N_A_29_53#_c_185_n 0.0104454f $X=0.48 $Y=1.695 $X2=0 $Y2=0
cc_69 N_C_M1003_g N_A_29_53#_c_187_n 0.0073535f $X=0.48 $Y=1.695 $X2=0 $Y2=0
cc_70 C N_A_29_53#_c_187_n 0.0234604f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_71 N_C_c_58_n N_A_29_53#_c_187_n 0.00639808f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C_M1004_g N_VGND_c_316_n 0.00953333f $X=0.48 $Y=0.475 $X2=0 $Y2=0
cc_73 N_C_M1004_g N_VGND_c_318_n 0.00322006f $X=0.48 $Y=0.475 $X2=0 $Y2=0
cc_74 N_C_M1004_g N_VGND_c_321_n 0.00465668f $X=0.48 $Y=0.475 $X2=0 $Y2=0
cc_75 N_B_M1001_g N_A_M1005_g 0.0033853f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_76 N_B_c_83_n N_A_M1005_g 0.0187947f $X=0.87 $Y=0.76 $X2=0 $Y2=0
cc_77 N_B_M1001_g N_A_M1007_g 0.0246912f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_78 N_B_c_87_n N_A_M1007_g 8.96507e-19 $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_79 N_B_M1001_g A 0.00692006f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_80 N_B_M1001_g N_A_c_124_n 0.0167622f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_A_c_125_n 0.0117813f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_82 N_B_c_84_n N_A_c_125_n 0.00177283f $X=0.87 $Y=0.91 $X2=0 $Y2=0
cc_83 N_B_M1001_g N_A_c_126_n 0.00332338f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_84 N_B_c_83_n N_A_29_53#_c_176_n 0.00683722f $X=0.87 $Y=0.76 $X2=0 $Y2=0
cc_85 N_B_c_84_n N_A_29_53#_c_176_n 0.0060465f $X=0.87 $Y=0.91 $X2=0 $Y2=0
cc_86 N_B_M1001_g N_A_29_53#_c_185_n 0.0107454f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_87 N_B_c_86_n N_A_29_53#_c_185_n 0.00120401f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_88 N_B_c_87_n N_A_29_53#_c_185_n 0.0497523f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_89 N_B_M1001_g N_A_29_53#_c_187_n 6.82547e-19 $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_90 N_B_c_87_n N_A_29_53#_c_187_n 0.0264475f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_91 N_B_M1001_g N_A_29_53#_c_188_n 0.00287525f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_92 N_B_c_87_n N_A_29_53#_c_188_n 0.0136891f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_93 N_B_M1001_g N_VPWR_c_273_n 0.00249809f $X=0.84 $Y=1.695 $X2=0 $Y2=0
cc_94 N_B_c_86_n N_VPWR_c_273_n 7.14013e-19 $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_95 N_B_c_87_n N_VPWR_c_273_n 0.0251801f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_96 N_B_c_86_n N_VPWR_c_274_n 0.00736312f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_97 N_B_c_87_n N_VPWR_c_274_n 0.0596585f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_98 N_B_c_86_n N_VPWR_c_272_n 0.0106165f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_99 N_B_c_87_n N_VPWR_c_272_n 0.0433365f $X=0.9 $Y=2.28 $X2=0 $Y2=0
cc_100 N_B_c_83_n N_VGND_c_316_n 0.00679416f $X=0.87 $Y=0.76 $X2=0 $Y2=0
cc_101 N_B_c_84_n N_VGND_c_316_n 2.19529e-19 $X=0.87 $Y=0.91 $X2=0 $Y2=0
cc_102 N_B_c_83_n N_VGND_c_317_n 5.25642e-19 $X=0.87 $Y=0.76 $X2=0 $Y2=0
cc_103 N_B_c_83_n N_VGND_c_319_n 0.00322006f $X=0.87 $Y=0.76 $X2=0 $Y2=0
cc_104 N_B_c_83_n N_VGND_c_321_n 0.00390029f $X=0.87 $Y=0.76 $X2=0 $Y2=0
cc_105 N_A_M1007_g N_A_29_53#_M1002_g 0.0189405f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_106 N_A_c_125_n N_A_29_53#_c_176_n 0.0169885f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_c_126_n N_A_29_53#_c_176_n 0.0160986f $X=0.697 $Y=1.325 $X2=0 $Y2=0
cc_108 N_A_M1007_g N_A_29_53#_c_185_n 2.22963e-19 $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_109 A N_A_29_53#_c_185_n 0.00994382f $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_110 N_A_c_125_n N_A_29_53#_c_185_n 0.0100971f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_M1005_g N_A_29_53#_c_178_n 0.0116406f $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_112 N_A_c_124_n N_A_29_53#_c_178_n 0.00220162f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_c_125_n N_A_29_53#_c_178_n 0.0166868f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_M1007_g N_A_29_53#_c_217_n 0.011218f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_115 N_A_c_125_n N_A_29_53#_c_217_n 0.00969518f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_M1007_g N_A_29_53#_c_186_n 0.0034529f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_117 N_A_c_124_n N_A_29_53#_c_179_n 5.77159e-19 $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_c_125_n N_A_29_53#_c_179_n 0.0146254f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_M1007_g N_A_29_53#_c_188_n 0.0100989f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_120 A N_A_29_53#_c_188_n 0.00536946f $X=0.6 $Y=1.445 $X2=0 $Y2=0
cc_121 N_A_c_124_n N_A_29_53#_c_188_n 0.00156816f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_125_n N_A_29_53#_c_188_n 0.0112207f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_124_n N_A_29_53#_c_180_n 0.00186332f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_125_n N_A_29_53#_c_180_n 0.0271506f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_124_n N_A_29_53#_c_181_n 0.0202671f $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_125_n N_A_29_53#_c_181_n 3.55971e-19 $X=1.305 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_M1005_g N_A_29_53#_c_182_n 0.0034529f $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_A_29_53#_c_183_n 0.0172443f $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_129 A A_111_297# 0.00106198f $X=0.6 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_130 N_A_M1007_g N_VPWR_c_273_n 0.00293484f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_131 N_A_M1007_g N_VPWR_c_274_n 0.00264561f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_132 N_A_M1007_g N_VPWR_c_272_n 0.00333991f $X=1.32 $Y=1.695 $X2=0 $Y2=0
cc_133 N_A_M1005_g N_VGND_c_316_n 5.2354e-19 $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_134 N_A_M1005_g N_VGND_c_317_n 0.00709299f $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_135 N_A_M1005_g N_VGND_c_319_n 0.00322006f $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_136 N_A_M1005_g N_VGND_c_321_n 0.00390029f $X=1.32 $Y=0.475 $X2=0 $Y2=0
cc_137 N_A_29_53#_c_185_n A_111_297# 0.0010205f $X=1.105 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_29_53#_c_185_n A_183_297# 0.00258288f $X=1.105 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_139 N_A_29_53#_c_188_n A_183_297# 0.00486567f $X=1.19 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_29_53#_c_217_n N_VPWR_M1007_d 0.00526233f $X=1.595 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_29_53#_M1002_g N_VPWR_c_273_n 0.00485906f $X=1.81 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_29_53#_c_217_n N_VPWR_c_273_n 0.0190361f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A_29_53#_c_188_n N_VPWR_c_273_n 0.00605542f $X=1.19 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A_29_53#_c_181_n N_VPWR_c_273_n 2.11345e-19 $X=1.785 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_29_53#_M1002_g N_VPWR_c_275_n 0.00585385f $X=1.81 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_29_53#_M1002_g N_VPWR_c_272_n 0.012849f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_29_53#_M1002_g N_X_c_299_n 0.00349311f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_29_53#_c_178_n N_X_c_299_n 0.0035218f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_29_53#_c_186_n N_X_c_299_n 0.00841221f $X=1.68 $Y=1.495 $X2=0 $Y2=0
cc_150 N_A_29_53#_c_180_n N_X_c_299_n 0.024459f $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_29_53#_c_181_n N_X_c_299_n 0.00753248f $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_29_53#_c_182_n N_X_c_299_n 0.00836618f $X=1.732 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_29_53#_c_183_n N_X_c_299_n 0.00441003f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_29_53#_c_176_n N_VGND_M1004_d 0.00160115f $X=1.025 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_29_53#_c_178_n N_VGND_M1005_d 0.00482895f $X=1.595 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_29_53#_c_182_n N_VGND_M1005_d 6.98847e-19 $X=1.732 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_29_53#_c_176_n N_VGND_c_316_n 0.0160613f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_29_53#_c_178_n N_VGND_c_317_n 0.020701f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_29_53#_c_181_n N_VGND_c_317_n 2.33671e-19 $X=1.785 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A_29_53#_c_183_n N_VGND_c_317_n 0.0132447f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A_29_53#_c_175_n N_VGND_c_318_n 0.0131002f $X=0.27 $Y=0.47 $X2=0 $Y2=0
cc_162 N_A_29_53#_c_176_n N_VGND_c_318_n 0.00232396f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_163 N_A_29_53#_c_176_n N_VGND_c_319_n 0.00232396f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_164 N_A_29_53#_c_259_p N_VGND_c_319_n 0.00846569f $X=1.11 $Y=0.47 $X2=0 $Y2=0
cc_165 N_A_29_53#_c_178_n N_VGND_c_319_n 0.00232396f $X=1.595 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_29_53#_c_178_n N_VGND_c_320_n 3.34073e-19 $X=1.595 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_29_53#_c_183_n N_VGND_c_320_n 0.00524631f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_29_53#_c_175_n N_VGND_c_321_n 0.00942308f $X=0.27 $Y=0.47 $X2=0 $Y2=0
cc_169 N_A_29_53#_c_176_n N_VGND_c_321_n 0.00970544f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_29_53#_c_259_p N_VGND_c_321_n 0.00625722f $X=1.11 $Y=0.47 $X2=0 $Y2=0
cc_171 N_A_29_53#_c_178_n N_VGND_c_321_n 0.00637905f $X=1.595 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_29_53#_c_183_n N_VGND_c_321_n 0.00952212f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_272_n N_X_M1002_d 0.00403568f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_174 N_VPWR_c_275_n X 0.019049f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_175 N_VPWR_c_272_n X 0.0105137f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_176 N_X_c_298_n N_VGND_c_320_n 0.00892181f $X=2.125 $Y=0.587 $X2=0 $Y2=0
cc_177 N_X_M1006_d N_VGND_c_321_n 0.00420587f $X=1.885 $Y=0.235 $X2=0 $Y2=0
cc_178 N_X_c_298_n N_VGND_c_321_n 0.00941771f $X=2.125 $Y=0.587 $X2=0 $Y2=0

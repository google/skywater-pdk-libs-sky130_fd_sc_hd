* File: sky130_fd_sc_hd__a31oi_2.spice.pex
* Created: Thu Aug 27 14:05:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A31OI_2%A3 1 3 6 8 10 13 15 17 28
r40 26 28 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=0.605 $Y=1.16
+ $X2=0.89 $Y2=1.16
r41 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.16 $X2=0.605 $Y2=1.16
r42 23 26 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.605 $Y2=1.16
r43 17 27 1.73624 $w=6.18e-07 $l=9e-08 $layer=LI1_cond $X=0.695 $Y=1.305
+ $X2=0.605 $Y2=1.305
r44 15 27 7.13789 $w=6.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.305
+ $X2=0.605 $Y2=1.305
r45 11 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r47 8 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r49 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r51 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%A2 1 3 6 8 10 13 15 17 27 28
c46 28 0 2.97772e-20 $X=1.73 $Y=1.16
r47 26 28 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.67 $Y=1.16 $X2=1.73
+ $Y2=1.16
r48 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r49 23 26 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.67 $Y2=1.16
r50 17 27 1.06104 $w=6.18e-07 $l=5.5e-08 $layer=LI1_cond $X=1.615 $Y=1.305
+ $X2=1.67 $Y2=1.305
r51 15 17 8.87413 $w=6.18e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.305
+ $X2=1.615 $Y2=1.305
r52 11 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r54 8 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r56 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r58 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%A1 3 5 7 8 10 13 15 18 21 23 29 32 35
c64 15 0 2.97772e-20 $X=2.225 $Y=1.16
r65 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.58
+ $Y=1.16 $X2=2.58 $Y2=1.16
r66 29 33 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.67 $Y2=1.16
r67 29 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.58 $Y2=1.16
r68 23 32 0.48229 $w=6.18e-07 $l=2.5e-08 $layer=LI1_cond $X=2.555 $Y=1.305
+ $X2=2.58 $Y2=1.305
r69 21 23 9.25996 $w=6.18e-07 $l=4.8e-07 $layer=LI1_cond $X=2.075 $Y=1.305
+ $X2=2.555 $Y2=1.305
r70 18 35 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.99 $Y=1.16 $X2=3.12
+ $Y2=1.16
r71 18 33 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=2.67 $Y2=1.16
r72 15 31 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.58 $Y2=1.16
r73 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.325
+ $X2=3.12 $Y2=1.16
r74 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=1.325
+ $X2=3.12 $Y2=1.985
r75 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=1.16
r76 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=0.56
r77 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=1.16
r78 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995 $X2=2.67
+ $Y2=0.56
r79 1 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.225 $Y2=1.16
r80 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%B1 1 3 6 8 10 12 15 17 18 19 20 27 30
c55 30 0 1.70053e-19 $X=4.265 $Y=1.175
r56 25 27 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.13 $Y=1.16
+ $X2=4.325 $Y2=1.16
r57 19 30 3.6174 $w=2e-07 $l=1.12e-07 $layer=LI1_cond $X=4.377 $Y=1.175
+ $X2=4.265 $Y2=1.175
r58 19 20 9.55671 $w=3.93e-07 $l=2.55e-07 $layer=LI1_cond $X=4.377 $Y=1.275
+ $X2=4.377 $Y2=1.53
r59 19 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.325
+ $Y=1.16 $X2=4.325 $Y2=1.16
r60 18 30 19.9636 $w=1.98e-07 $l=3.6e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=4.265 $Y2=1.175
r61 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.325
+ $X2=4.13 $Y2=1.16
r62 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.13 $Y=1.325
+ $X2=4.13 $Y2=1.985
r63 10 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=0.995
+ $X2=4.13 $Y2=1.16
r64 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.995
+ $X2=4.13 $Y2=0.56
r65 9 17 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.705 $Y=1.16
+ $X2=3.63 $Y2=1.16
r66 8 25 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.055 $Y=1.16
+ $X2=4.13 $Y2=1.16
r67 8 9 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=4.055 $Y=1.16
+ $X2=3.705 $Y2=1.16
r68 4 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.325
+ $X2=3.63 $Y2=1.16
r69 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.63 $Y=1.325 $X2=3.63
+ $Y2=1.985
r70 1 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=0.995
+ $X2=3.63 $Y2=1.16
r71 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.63 $Y=0.995 $X2=3.63
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%A_27_297# 1 2 3 4 5 18 22 26 28 29 30 31 34
+ 37 39 41
c59 41 0 2.97772e-20 $X=1.94 $Y=1.95
c60 39 0 2.97772e-20 $X=1.1 $Y=1.95
c61 34 0 1.70053e-19 $X=4.34 $Y=1.96
r62 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.34 $Y=2.295
+ $X2=4.34 $Y2=1.96
r63 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.255 $Y=2.38
+ $X2=4.34 $Y2=2.295
r64 30 31 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.255 $Y=2.38
+ $X2=3.505 $Y2=2.38
r65 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=2.295
+ $X2=3.505 $Y2=2.38
r66 28 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.955
+ $X2=3.42 $Y2=1.87
r67 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.42 $Y=1.955
+ $X2=3.42 $Y2=2.295
r68 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.87
+ $X2=1.94 $Y2=1.87
r69 26 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.87
+ $X2=3.42 $Y2=1.87
r70 26 27 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.335 $Y=1.87
+ $X2=2.025 $Y2=1.87
r71 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.87 $X2=1.1
+ $Y2=1.87
r72 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=1.87
+ $X2=1.94 $Y2=1.87
r73 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=1.87
+ $X2=1.185 $Y2=1.87
r74 19 37 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.26 $Y2=1.87
r75 18 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=1.87 $X2=1.1
+ $Y2=1.87
r76 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=1.87
+ $X2=0.345 $Y2=1.87
r77 5 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=1.96
r78 4 43 300 $w=1.7e-07 $l=5.66436e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=1.485 $X2=3.42 $Y2=1.95
r79 3 41 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.95
r80 2 39 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.95
r81 1 37 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%VPWR 1 2 3 12 16 19 20 21 23 32 41 42 45 48
r66 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r67 48 51 9.10448 $w=6.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.645 $Y=2.21
+ $X2=2.645 $Y2=2.72
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r70 39 42 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r71 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 38 41 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 36 51 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=2.645 $Y2=2.72
r75 36 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.98 $Y=2.72 $X2=2.99
+ $Y2=2.72
r76 35 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r78 32 51 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.645 $Y2=2.72
r79 32 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 31 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r81 31 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 28 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r84 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 23 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r86 23 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 21 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 21 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 19 30 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.15 $Y2=2.72
r90 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.52 $Y2=2.72
r91 18 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=2.07 $Y2=2.72
r92 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.52 $Y2=2.72
r93 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r94 14 16 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.21
r95 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r96 10 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.21
r97 3 48 300 $w=1.7e-07 $l=9.76409e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.815 $Y2=2.21
r98 2 16 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.21
r99 1 12 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%Y 1 2 3 4 13 19 21 23 27 31 33 34 35 44
r70 41 44 0.914637 $w=3.13e-07 $l=2.5e-08 $layer=LI1_cond $X=3.412 $Y=0.825
+ $X2=3.412 $Y2=0.85
r71 34 35 7.75597 $w=4.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.412 $Y=1.19
+ $X2=3.412 $Y2=1.445
r72 33 41 2.04209 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.412 $Y=0.74
+ $X2=3.412 $Y2=0.825
r73 33 34 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=3.412 $Y=0.88
+ $X2=3.412 $Y2=1.19
r74 33 44 1.09756 $w=3.13e-07 $l=3e-08 $layer=LI1_cond $X=3.412 $Y=0.88
+ $X2=3.412 $Y2=0.85
r75 29 31 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.34 $Y=0.655
+ $X2=4.34 $Y2=0.38
r76 25 27 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.92 $Y=1.615
+ $X2=3.92 $Y2=1.63
r77 24 35 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.57 $Y=1.53
+ $X2=3.412 $Y2=1.53
r78 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.755 $Y=1.53
+ $X2=3.92 $Y2=1.615
r79 23 24 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.755 $Y=1.53
+ $X2=3.57 $Y2=1.53
r80 22 33 4.19666 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.57 $Y=0.74
+ $X2=3.412 $Y2=0.74
r81 21 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.175 $Y=0.74
+ $X2=4.34 $Y2=0.655
r82 21 22 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.175 $Y=0.74
+ $X2=3.57 $Y2=0.74
r83 17 33 2.04209 $w=1.7e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.34 $Y=0.655
+ $X2=3.412 $Y2=0.74
r84 17 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.34 $Y=0.655
+ $X2=3.34 $Y2=0.42
r85 13 33 4.19666 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=3.255 $Y=0.74
+ $X2=3.412 $Y2=0.74
r86 13 15 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.255 $Y=0.74
+ $X2=2.46 $Y2=0.74
r87 4 27 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=3.705
+ $Y=1.485 $X2=3.92 $Y2=1.63
r88 3 31 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=0.235 $X2=4.34 $Y2=0.38
r89 2 33 182 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.34 $Y2=0.76
r90 2 19 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.34 $Y2=0.42
r91 1 15 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%A_27_47# 1 2 3 16
r23 14 16 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=0.74 $X2=1.94
+ $Y2=0.74
r24 11 14 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.26 $Y=0.74 $X2=1.1
+ $Y2=0.74
r25 3 16 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.74
r26 2 14 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.74
r27 1 11 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r60 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r62 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r63 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r64 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=3.84
+ $Y2=0
r65 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.37
+ $Y2=0
r66 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r67 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r68 26 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r69 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r70 25 28 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r71 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r72 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r73 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r74 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.84
+ $Y2=0
r75 22 28 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.45
+ $Y2=0
r76 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r77 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r78 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r79 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r80 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0
r81 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0.38
r82 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r83 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r84 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.235 $X2=3.84 $Y2=0.38
r85 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_2%A_277_47# 1 2 11
r20 8 11 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.52 $Y=0.38
+ $X2=2.91 $Y2=0.38
r21 2 11 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.91 $Y2=0.38
r22 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
.ends


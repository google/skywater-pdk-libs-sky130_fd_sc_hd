* File: sky130_fd_sc_hd__a21bo_4.spice
* Created: Thu Aug 27 14:00:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21bo_4.pex.spice"
.subckt sky130_fd_sc_hd__a21bo_4  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_B1_N_M1021_g N_A_42_47#_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.25025 PD=0.93 PS=2.07 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75000.3
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1021_d N_A_205_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_205_21#_M1007_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1007_d N_A_205_21#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A_205_21#_M1019_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.26325 AS=0.091 PD=1.46 PS=0.93 NRD=20.304 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_205_21#_M1014_d N_A_42_47#_M1014_g N_VGND_M1019_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.26325 PD=0.92 PS=1.46 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75003 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1020 N_A_205_21#_M1014_d N_A_42_47#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.10075 PD=0.92 PS=0.96 NRD=0 NRS=6.456 M=1 R=4.33333
+ SA=75003.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1020_s N_A2_M1004_g A_861_47# VNB NSHORT L=0.15 W=0.65 AD=0.10075
+ AS=0.07475 PD=0.96 PS=0.88 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75003.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 A_861_47# N_A1_M1002_g N_A_205_21#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.07475 AS=0.08775 PD=0.88 PS=0.92 NRD=11.076 NRS=0 M=1 R=4.33333
+ SA=75004.2 SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 A_1021_47# N_A1_M1012_g N_A_205_21#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75004.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A2_M1013_g A_1021_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75005.1 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1017 N_VPWR_M1017_d N_B1_N_M1017_g N_A_42_47#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_X_M1006_d N_A_205_21#_M1006_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1006_d N_A_205_21#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1010 N_X_M1010_d N_A_205_21#_M1010_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1018 N_X_M1010_d N_A_205_21#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_603_297#_M1000_d N_A_42_47#_M1000_g N_A_205_21#_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1003 N_A_603_297#_M1003_d N_A_42_47#_M1003_g N_A_205_21#_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 N_A_603_297#_M1003_d N_A2_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1015_s N_A1_M1001_g N_A_603_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g N_A_603_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_603_297#_M1016_d N_A2_M1016_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_46 VNB 0 9.49649e-20 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__a21bo_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__clkdlybuf4s15_2.pex.spice
* Created: Thu Aug 27 14:11:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A 3 7 9 10 14 15
r34 14 17 41.0874 $w=3.35e-07 $l=1.35e-07 $layer=POLY_cond $X=0.387 $Y=1.16
+ $X2=0.387 $Y2=1.295
r35 14 16 41.0874 $w=3.35e-07 $l=1.35e-07 $layer=POLY_cond $X=0.387 $Y=1.16
+ $X2=0.387 $Y2=1.025
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.16 $X2=0.385 $Y2=1.16
r37 9 10 8.65248 $w=4.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.32 $Y=1.19 $X2=0.32
+ $Y2=1.53
r38 9 15 0.763454 $w=4.68e-07 $l=3e-08 $layer=LI1_cond $X=0.32 $Y=1.19 $X2=0.32
+ $Y2=1.16
r39 7 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.48 $Y=1.985
+ $X2=0.48 $Y2=1.295
r40 3 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.48 $Y=0.445
+ $X2=0.48 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_27_47# 1 2 9 13 17 21 22 23 26 28
+ 30 34 35
c77 34 0 1.45867e-19 $X=1.155 $Y=1.16
c78 28 0 3.38757e-20 $X=0.975 $Y=1.795
r79 35 39 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.155 $Y=1.16
+ $X2=1.155 $Y2=1.295
r80 35 38 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.155 $Y=1.16
+ $X2=1.155 $Y2=1.025
r81 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.16 $X2=1.155 $Y2=1.16
r82 31 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.975 $Y=1.16
+ $X2=1.155 $Y2=1.16
r83 27 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=1.245
+ $X2=0.975 $Y2=1.16
r84 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=1.245
+ $X2=0.975 $Y2=1.795
r85 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=1.075
+ $X2=0.975 $Y2=1.16
r86 25 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.975 $Y=0.89
+ $X2=0.975 $Y2=1.075
r87 24 30 5.29321 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.43 $Y=1.88
+ $X2=0.257 $Y2=1.88
r88 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.89 $Y=1.88
+ $X2=0.975 $Y2=1.795
r89 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.89 $Y=1.88
+ $X2=0.43 $Y2=1.88
r90 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.89 $Y=0.805
+ $X2=0.975 $Y2=0.89
r91 21 22 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.89 $Y=0.805
+ $X2=0.415 $Y2=0.805
r92 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.25 $Y=0.72
+ $X2=0.415 $Y2=0.805
r93 15 17 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.25 $Y=0.72 $X2=0.25
+ $Y2=0.42
r94 13 39 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.065 $Y=2.075
+ $X2=1.065 $Y2=1.295
r95 9 38 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.065 $Y=0.56
+ $X2=1.065 $Y2=1.025
r96 2 30 300 $w=1.7e-07 $l=5.36074e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=1.96
r97 1 17 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_228_47# 1 2 9 13 19 22 30 31 34 35
+ 36 37 38
c74 38 0 1.79743e-19 $X=2.075 $Y=1.16
c75 31 0 1.84487e-19 $X=2.25 $Y=1.16
r76 38 41 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=1.16
+ $X2=2.15 $Y2=1.16
r77 34 35 9.0529 $w=4.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.445 $Y=1.96
+ $X2=1.445 $Y2=1.785
r78 31 41 22.2174 $w=2.7e-07 $l=1e-07 $layer=POLY_cond $X=2.25 $Y=1.16 $X2=2.15
+ $Y2=1.16
r79 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r80 28 38 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.16
+ $X2=2.075 $Y2=1.16
r81 27 30 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.91 $Y=1.28
+ $X2=2.25 $Y2=1.28
r82 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.16 $X2=1.91 $Y2=1.16
r83 25 37 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=1.28
+ $X2=1.575 $Y2=1.28
r84 25 27 7.02709 $w=4.08e-07 $l=2.5e-07 $layer=LI1_cond $X=1.66 $Y=1.28
+ $X2=1.91 $Y2=1.28
r85 23 37 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.575 $Y=1.485
+ $X2=1.575 $Y2=1.28
r86 23 35 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.575 $Y=1.485
+ $X2=1.575 $Y2=1.785
r87 22 37 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.575 $Y=1.075
+ $X2=1.575 $Y2=1.28
r88 22 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.575 $Y=1.075
+ $X2=1.575 $Y2=0.905
r89 17 36 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=1.47 $Y=0.715
+ $X2=1.47 $Y2=0.905
r90 17 19 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.47 $Y=0.715
+ $X2=1.47 $Y2=0.42
r91 11 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r92 11 13 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=2.075
r93 7 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r94 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r95 2 34 300 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.665 $X2=1.395 $Y2=1.96
r96 1 19 182 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.235 $X2=1.42 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_362_333# 1 2 9 13 15 19 23 25 28
+ 32 33 34 37 39 42 43 46 47
c91 43 0 9.88072e-20 $X=3.02 $Y=1.16
c92 39 0 1.84487e-19 $X=2.815 $Y=1.79
c93 9 0 1.39978e-20 $X=3.01 $Y=0.445
r94 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.16 $X2=3.02 $Y2=1.16
r95 40 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=1.16 $X2=2.815
+ $Y2=1.16
r96 40 42 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.9 $Y=1.16 $X2=3.02
+ $Y2=1.16
r97 38 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=1.245
+ $X2=2.815 $Y2=1.16
r98 38 39 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.815 $Y=1.245
+ $X2=2.815 $Y2=1.79
r99 37 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=1.075
+ $X2=2.815 $Y2=1.16
r100 36 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.815 $Y=0.905
+ $X2=2.815 $Y2=1.075
r101 35 46 4.376 $w=1.75e-07 $l=1.35e-07 $layer=LI1_cond $X=2.1 $Y=1.877
+ $X2=1.965 $Y2=1.877
r102 34 39 6.81835 $w=1.75e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.73 $Y=1.877
+ $X2=2.815 $Y2=1.79
r103 34 35 39.9273 $w=1.73e-07 $l=6.3e-07 $layer=LI1_cond $X=2.73 $Y=1.877
+ $X2=2.1 $Y2=1.877
r104 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.73 $Y=0.82
+ $X2=2.815 $Y2=0.905
r105 32 33 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.73 $Y=0.82
+ $X2=2.1 $Y2=0.82
r106 26 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.965 $Y=0.735
+ $X2=2.1 $Y2=0.82
r107 26 28 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.965 $Y=0.735
+ $X2=1.965 $Y2=0.42
r108 21 25 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.44 $Y=1.295
+ $X2=3.44 $Y2=1.16
r109 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.44 $Y=1.295
+ $X2=3.44 $Y2=1.985
r110 17 25 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.44 $Y=1.025
+ $X2=3.44 $Y2=1.16
r111 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.44 $Y=1.025
+ $X2=3.44 $Y2=0.445
r112 16 43 2.60871 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=3.085 $Y=1.16
+ $X2=2.97 $Y2=1.16
r113 15 25 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.16
+ $X2=3.44 $Y2=1.16
r114 15 16 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=3.365 $Y=1.16
+ $X2=3.085 $Y2=1.16
r115 11 43 32.2453 $w=1.5e-07 $l=1.53704e-07 $layer=POLY_cond $X=3.01 $Y=1.295
+ $X2=2.97 $Y2=1.16
r116 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.01 $Y=1.295
+ $X2=3.01 $Y2=1.985
r117 7 43 32.2453 $w=1.5e-07 $l=1.53704e-07 $layer=POLY_cond $X=3.01 $Y=1.025
+ $X2=2.97 $Y2=1.16
r118 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.01 $Y=1.025
+ $X2=3.01 $Y2=0.445
r119 2 46 300 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=1.665 $X2=1.935 $Y2=1.96
r120 1 28 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.235 $X2=1.94 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%VPWR 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 39 47 4.85147 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.72 $Y=2.72 $X2=3.93
+ $Y2=2.72
r56 39 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.72 $Y=2.72 $X2=3.45
+ $Y2=2.72
r57 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.765 $Y2=2.72
r64 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.765 $Y2=2.72
r66 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r67 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 23 37 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.55 $Y=2.72 $X2=2.53
+ $Y2=2.72
r70 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=2.72
+ $X2=2.715 $Y2=2.72
r71 22 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.88 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=2.72
+ $X2=2.715 $Y2=2.72
r73 18 47 2.95709 $w=3.35e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.887 $Y=2.635
+ $X2=3.93 $Y2=2.72
r74 18 20 26.833 $w=3.33e-07 $l=7.8e-07 $layer=LI1_cond $X=3.887 $Y=2.635
+ $X2=3.887 $Y2=1.855
r75 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=2.635
+ $X2=2.715 $Y2=2.72
r76 14 16 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.715 $Y=2.635
+ $X2=2.715 $Y2=2.3
r77 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.72
r78 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.3
r79 3 20 300 $w=1.7e-07 $l=5.21488e-07 $layer=licon1_PDIFF $count=2 $X=3.515
+ $Y=1.485 $X2=3.88 $Y2=1.855
r80 2 16 600 $w=1.7e-07 $l=8.45207e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.665 $X2=2.715 $Y2=2.3
r81 1 12 600 $w=1.7e-07 $l=9.13989e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.485 $X2=0.765 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%X 1 2 7 8 9 10 11 12 29 40 43
r29 43 44 5.46507 $w=4.78e-07 $l=4.5e-08 $layer=LI1_cond $X=3.31 $Y=1.53
+ $X2=3.31 $Y2=1.485
r30 27 29 3.23938 $w=4.78e-07 $l=1.3e-07 $layer=LI1_cond $X=3.31 $Y=1.725
+ $X2=3.31 $Y2=1.855
r31 20 40 4.74025 $w=1.95e-07 $l=1.93e-07 $layer=LI1_cond $X=3.452 $Y=0.64
+ $X2=3.452 $Y2=0.447
r32 11 12 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.31 $Y=1.87
+ $X2=3.31 $Y2=2.21
r33 11 29 0.373774 $w=4.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.31 $Y=1.87
+ $X2=3.31 $Y2=1.855
r34 10 27 4.3607 $w=4.78e-07 $l=1.75e-07 $layer=LI1_cond $X=3.31 $Y=1.55
+ $X2=3.31 $Y2=1.725
r35 10 43 0.498366 $w=4.78e-07 $l=2e-08 $layer=LI1_cond $X=3.31 $Y=1.55 $X2=3.31
+ $Y2=1.53
r36 10 44 1.13753 $w=1.93e-07 $l=2e-08 $layer=LI1_cond $X=3.452 $Y=1.465
+ $X2=3.452 $Y2=1.485
r37 9 10 15.641 $w=1.93e-07 $l=2.75e-07 $layer=LI1_cond $X=3.452 $Y=1.19
+ $X2=3.452 $Y2=1.465
r38 8 9 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=3.452 $Y=0.85 $X2=3.452
+ $Y2=1.19
r39 8 20 11.9441 $w=1.93e-07 $l=2.1e-07 $layer=LI1_cond $X=3.452 $Y=0.85
+ $X2=3.452 $Y2=0.64
r40 7 40 0.0598672 $w=3.83e-07 $l=2e-09 $layer=LI1_cond $X=3.45 $Y=0.447
+ $X2=3.452 $Y2=0.447
r41 7 36 6.73506 $w=3.83e-07 $l=2.25e-07 $layer=LI1_cond $X=3.45 $Y=0.447
+ $X2=3.225 $Y2=0.447
r42 2 29 300 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=2 $X=3.085
+ $Y=1.485 $X2=3.225 $Y2=1.855
r43 1 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.225 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%VGND 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c49 20 0 1.39978e-20 $X=3.88 $Y=0.42
c50 16 0 9.88072e-20 $X=2.715 $Y=0.4
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r55 39 47 4.85147 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.93
+ $Y2=0
r56 39 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.45
+ $Y2=0
r57 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r58 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r59 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r60 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r61 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r62 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r64 32 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.15
+ $Y2=0
r65 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r66 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.23
+ $Y2=0
r67 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r68 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 23 37 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.53
+ $Y2=0
r70 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.715
+ $Y2=0
r71 22 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.45
+ $Y2=0
r72 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.715
+ $Y2=0
r73 18 47 2.95709 $w=3.35e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.887 $Y=0.085
+ $X2=3.93 $Y2=0
r74 18 20 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=3.887 $Y=0.085
+ $X2=3.887 $Y2=0.42
r75 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0
r76 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0.4
r77 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r78 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.42
r79 3 20 182 $w=1.7e-07 $l=4.48051e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.88 $Y2=0.42
r80 2 16 182 $w=1.7e-07 $l=5.66524e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.715 $Y2=0.4
r81 1 12 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.75 $Y2=0.42
.ends


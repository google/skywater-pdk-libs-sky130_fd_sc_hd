* File: sky130_fd_sc_hd__mux2_4.spice
* Created: Tue Sep  1 19:14:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2_4.pex.spice"
.subckt sky130_fd_sc_hd__mux2_4  VNB VPB S A0 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_S_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.169 PD=0.985 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1005 A_206_47# N_A_27_47#_M1005_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.65
+ AD=0.26 AS=0.108875 PD=1.45 PS=0.985 NRD=63.684 NRS=11.076 M=1 R=4.33333
+ SA=75000.7 SB=75004.3 A=0.0975 P=1.6 MULT=1
MM1007 N_A_396_47#_M1007_d N_A0_M1007_g A_206_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.26 PD=0.97 PS=1.45 NRD=3.684 NRS=63.684 M=1 R=4.33333 SA=75001.6
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1002 A_490_47# N_A1_M1002_g N_A_396_47#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.274625 AS=0.104 PD=1.495 PS=0.97 NRD=67.836 NRS=3.684 M=1 R=4.33333
+ SA=75002.1 SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_S_M1011_g A_490_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.274625 PD=0.92 PS=1.495 NRD=0 NRS=67.836 M=1 R=4.33333 SA=75003.1
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_396_47#_M1008_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1008_d N_A_396_47#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.9
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 N_X_M1012_d N_A_396_47#_M1012_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.3
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1014 N_X_M1012_d N_A_396_47#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 N_VPWR_M1015_d N_S_M1015_g N_A_27_47#_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1625 AS=0.26 PD=1.325 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1000 N_A_204_297#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=1 AD=0.28 AS=0.1625 PD=2.56 PS=1.325 NRD=0.9653 NRS=9.8303 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_396_47#_M1004_d N_A0_M1004_g N_A_314_297#_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.16 AS=0.26 PD=1.32 PS=2.52 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_A_204_297#_M1001_d N_A1_M1001_g N_A_396_47#_M1004_d VPB PHIGHVT L=0.15
+ W=1 AD=0.3 AS=0.16 PD=2.6 PS=1.32 NRD=2.9353 NRS=2.9353 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_S_M1016_g N_A_314_297#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_396_47#_M1003_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1006 N_X_M1003_d N_A_396_47#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1010 N_X_M1010_d N_A_396_47#_M1010_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1010_d N_A_396_47#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_707 A_490_47# 0 1.83477e-19 $X=2.45 $Y=0.235
*
.include "sky130_fd_sc_hd__mux2_4.pxi.spice"
*
.ends
*
*

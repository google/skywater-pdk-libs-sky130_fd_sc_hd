* File: sky130_fd_sc_hd__nor4_4.pex.spice
* Created: Tue Sep  1 19:19:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r74 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.6 $Y=1.16 $X2=1.75
+ $Y2=1.16
r75 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.6 $Y=1.16
+ $X2=1.6 $Y2=1.16
r76 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.33 $Y=1.16 $X2=1.6
+ $Y2=1.16
r77 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r78 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.58 $Y=1.16
+ $X2=0.91 $Y2=1.16
r79 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r80 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.58
+ $Y2=1.16
r81 29 40 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=1.6 $Y2=1.18
r82 29 35 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=0.58 $Y2=1.18
r83 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r85 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r87 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r89 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r91 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r93 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r95 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r97 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 45
r78 43 45 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.28 $Y=1.16
+ $X2=3.43 $Y2=1.16
r79 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.28
+ $Y=1.16 $X2=3.28 $Y2=1.16
r80 41 43 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.28 $Y2=1.16
r81 40 41 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=3.01 $Y2=1.16
r82 38 40 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.59 $Y2=1.16
r83 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r84 35 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.17 $Y=1.16 $X2=2.26
+ $Y2=1.16
r85 30 31 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=3.455 $Y=1.18
+ $X2=3.915 $Y2=1.18
r86 30 44 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=3.455 $Y=1.18
+ $X2=3.28 $Y2=1.18
r87 29 44 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.995 $Y=1.18
+ $X2=3.28 $Y2=1.18
r88 29 39 38.8182 $w=2.08e-07 $l=7.35e-07 $layer=LI1_cond $X=2.995 $Y=1.18
+ $X2=2.26 $Y2=1.18
r89 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r90 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.985
r91 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r93 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r94 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.985
r95 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.16
r96 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r97 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.16
r98 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.985
r99 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r100 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r101 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r102 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r103 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r77 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.48 $Y=1.16
+ $X2=5.63 $Y2=1.16
r78 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.48
+ $Y=1.16 $X2=5.48 $Y2=1.16
r79 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.21 $Y=1.16
+ $X2=5.48 $Y2=1.16
r80 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=5.21 $Y2=1.16
r81 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.79 $Y2=1.16
r82 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r83 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.37 $Y=1.16 $X2=4.46
+ $Y2=1.16
r84 29 40 34.0649 $w=2.08e-07 $l=6.45e-07 $layer=LI1_cond $X=4.835 $Y=1.18
+ $X2=5.48 $Y2=1.18
r85 29 35 19.8052 $w=2.08e-07 $l=3.75e-07 $layer=LI1_cond $X=4.835 $Y=1.18
+ $X2=4.46 $Y2=1.18
r86 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.16
r87 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.985
r88 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=1.16
r89 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=0.56
r90 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.16
r91 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.985
r92 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=1.16
r93 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=0.56
r94 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.16
r95 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.985
r96 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=1.16
r97 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=0.56
r98 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.16
r99 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.37 $Y=1.325 $X2=4.37
+ $Y2=1.985
r100 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=1.16
r101 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%D 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r78 39 41 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.13 $Y=1.16 $X2=7.31
+ $Y2=1.16
r79 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.13
+ $Y=1.16 $X2=7.13 $Y2=1.16
r80 37 39 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=6.89 $Y=1.16
+ $X2=7.13 $Y2=1.16
r81 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.47 $Y=1.16
+ $X2=6.89 $Y2=1.16
r82 34 36 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=6.11 $Y=1.16
+ $X2=6.47 $Y2=1.16
r83 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.11
+ $Y=1.16 $X2=6.11 $Y2=1.16
r84 31 34 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.05 $Y=1.16 $X2=6.11
+ $Y2=1.16
r85 29 40 24.0303 $w=2.08e-07 $l=4.55e-07 $layer=LI1_cond $X=6.675 $Y=1.18
+ $X2=7.13 $Y2=1.18
r86 29 35 29.8398 $w=2.08e-07 $l=5.65e-07 $layer=LI1_cond $X=6.675 $Y=1.18
+ $X2=6.11 $Y2=1.18
r87 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=1.325
+ $X2=7.31 $Y2=1.16
r88 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.31 $Y=1.325
+ $X2=7.31 $Y2=1.985
r89 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=0.995
+ $X2=7.31 $Y2=1.16
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.31 $Y=0.995
+ $X2=7.31 $Y2=0.56
r91 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.16
r92 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.985
r93 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=1.16
r94 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=0.56
r95 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=1.325
+ $X2=6.47 $Y2=1.16
r96 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.47 $Y=1.325
+ $X2=6.47 $Y2=1.985
r97 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=0.995
+ $X2=6.47 $Y2=1.16
r98 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.47 $Y=0.995
+ $X2=6.47 $Y2=0.56
r99 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=1.325
+ $X2=6.05 $Y2=1.16
r100 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.05 $Y=1.325
+ $X2=6.05 $Y2=1.985
r101 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=0.995
+ $X2=6.05 $Y2=1.16
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.05 $Y=0.995
+ $X2=6.05 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 36 40 45 50
r62 38 40 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=3.667 $Y=2.295
+ $X2=3.667 $Y2=1.96
r63 37 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.925 $Y=2.38
+ $X2=2.8 $Y2=2.38
r64 36 38 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=3.515 $Y=2.38
+ $X2=3.667 $Y2=2.295
r65 36 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.515 $Y=2.38
+ $X2=2.925 $Y2=2.38
r66 32 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=2.295
+ $X2=2.8 $Y2=2.38
r67 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.8 $Y=2.295
+ $X2=2.8 $Y2=1.96
r68 31 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=2.38
+ $X2=1.96 $Y2=2.38
r69 30 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.675 $Y=2.38
+ $X2=2.8 $Y2=2.38
r70 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.675 $Y=2.38
+ $X2=2.085 $Y2=2.38
r71 29 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.295
+ $X2=1.96 $Y2=2.38
r72 28 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=1.625
+ $X2=1.96 $Y2=1.54
r73 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.96 $Y=1.625
+ $X2=1.96 $Y2=2.295
r74 27 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.54
+ $X2=1.12 $Y2=1.54
r75 26 47 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.96 $Y2=1.54
r76 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.245 $Y2=1.54
r77 22 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=1.54
r78 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=2.3
r79 21 43 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.247 $Y2=1.54
r80 20 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=1.12 $Y2=1.54
r81 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=0.405 $Y2=1.54
r82 16 43 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=1.54
r83 16 18 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=2.3
r84 5 40 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=1.96
r85 4 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=1.96
r86 3 49 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.3
r87 3 47 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r88 2 45 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r89 2 24 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r90 1 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r91 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%VPWR 1 2 9 13 15 17 22 29 30 33 36
r93 36 37 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 30 37 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=1.61 $Y2=2.72
r96 29 30 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r97 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.54 $Y2=2.72
r98 27 29 386.551 $w=1.68e-07 $l=5.925e-06 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=7.59 $Y2=2.72
r99 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r100 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r101 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r103 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r104 22 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.54 $Y2=2.72
r105 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r107 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r108 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r109 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r110 11 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.72
r111 11 13 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=1.96
r112 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r113 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r114 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
r115 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%A_449_297# 1 2 3 4 15 19 23 28 30 32 34
r58 24 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.705 $Y=1.54
+ $X2=4.58 $Y2=1.54
r59 23 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=1.54
+ $X2=5.42 $Y2=1.54
r60 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.295 $Y=1.54
+ $X2=4.705 $Y2=1.54
r61 20 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=1.54
+ $X2=3.22 $Y2=1.54
r62 19 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.455 $Y=1.54
+ $X2=4.58 $Y2=1.54
r63 19 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.455 $Y=1.54
+ $X2=3.345 $Y2=1.54
r64 16 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=1.54
+ $X2=2.38 $Y2=1.54
r65 15 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=1.54
+ $X2=3.22 $Y2=1.54
r66 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.095 $Y=1.54
+ $X2=2.505 $Y2=1.54
r67 4 34 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.485 $X2=5.42 $Y2=1.62
r68 3 32 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=1.485 $X2=4.58 $Y2=1.62
r69 2 30 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.62
r70 1 28 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%A_807_297# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 45 46
r57 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.52 $Y=2.295
+ $X2=7.52 $Y2=1.96
r58 39 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.805 $Y=2.38
+ $X2=6.68 $Y2=2.38
r59 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.395 $Y=2.38
+ $X2=7.52 $Y2=2.295
r60 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.395 $Y=2.38
+ $X2=6.805 $Y2=2.38
r61 34 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.68 $Y=2.295
+ $X2=6.68 $Y2=2.38
r62 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.68 $Y=2.295
+ $X2=6.68 $Y2=1.96
r63 33 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.965 $Y=2.38
+ $X2=5.84 $Y2=2.38
r64 32 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.555 $Y=2.38
+ $X2=6.68 $Y2=2.38
r65 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.555 $Y=2.38
+ $X2=5.965 $Y2=2.38
r66 28 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.84 $Y=2.295
+ $X2=5.84 $Y2=2.38
r67 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.84 $Y=2.295
+ $X2=5.84 $Y2=1.96
r68 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.125 $Y=2.38 $X2=5
+ $Y2=2.38
r69 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.715 $Y=2.38
+ $X2=5.84 $Y2=2.38
r70 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.715 $Y=2.38
+ $X2=5.125 $Y2=2.38
r71 22 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=2.295 $X2=5
+ $Y2=2.38
r72 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5 $Y=2.295 $X2=5
+ $Y2=1.96
r73 20 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.875 $Y=2.38 $X2=5
+ $Y2=2.38
r74 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.875 $Y=2.38
+ $X2=4.285 $Y2=2.38
r75 16 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.145 $Y=2.295
+ $X2=4.285 $Y2=2.38
r76 16 18 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.145 $Y=2.295
+ $X2=4.145 $Y2=1.96
r77 5 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.385
+ $Y=1.485 $X2=7.52 $Y2=1.96
r78 4 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.545
+ $Y=1.485 $X2=6.68 $Y2=1.96
r79 3 30 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.705
+ $Y=1.485 $X2=5.84 $Y2=1.96
r80 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5 $Y2=1.96
r81 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=1.485 $X2=4.16 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 41 45 47
+ 51 53 57 59 63 65 69 73 75 79 83 85 87 88 89 90 91 92 94 95 97 99 102
r211 99 102 2.87089 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=7.6 $Y=0.815 $X2=7.6
+ $Y2=0.905
r212 99 102 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.6 $Y=0.92
+ $X2=7.6 $Y2=0.905
r213 98 99 22.8354 $w=2.68e-07 $l=5.35e-07 $layer=LI1_cond $X=7.6 $Y=1.455
+ $X2=7.6 $Y2=0.92
r214 86 95 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=0.815
+ $X2=7.1 $Y2=0.815
r215 85 99 4.30634 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=7.465 $Y=0.815
+ $X2=7.6 $Y2=0.815
r216 85 86 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=7.465 $Y=0.815
+ $X2=7.265 $Y2=0.815
r217 84 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.225 $Y=1.54
+ $X2=7.1 $Y2=1.54
r218 83 98 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.465 $Y=1.54
+ $X2=7.6 $Y2=1.455
r219 83 84 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.465 $Y=1.54
+ $X2=7.225 $Y2=1.54
r220 77 95 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.1 $Y=0.725 $X2=7.1
+ $Y2=0.815
r221 77 79 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.1 $Y=0.725
+ $X2=7.1 $Y2=0.39
r222 76 92 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=0.815
+ $X2=6.26 $Y2=0.815
r223 75 95 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.935 $Y=0.815
+ $X2=7.1 $Y2=0.815
r224 75 76 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.935 $Y=0.815
+ $X2=6.425 $Y2=0.815
r225 74 94 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.385 $Y=1.54
+ $X2=6.26 $Y2=1.54
r226 73 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.975 $Y=1.54
+ $X2=7.1 $Y2=1.54
r227 73 74 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.975 $Y=1.54
+ $X2=6.385 $Y2=1.54
r228 67 92 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.26 $Y=0.725
+ $X2=6.26 $Y2=0.815
r229 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.26 $Y=0.725
+ $X2=6.26 $Y2=0.39
r230 66 91 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=0.815
+ $X2=5.42 $Y2=0.815
r231 65 92 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=0.815
+ $X2=6.26 $Y2=0.815
r232 65 66 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.095 $Y=0.815
+ $X2=5.585 $Y2=0.815
r233 61 91 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.42 $Y=0.725
+ $X2=5.42 $Y2=0.815
r234 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.42 $Y=0.725
+ $X2=5.42 $Y2=0.39
r235 60 90 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=0.815
+ $X2=4.58 $Y2=0.815
r236 59 91 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=0.815
+ $X2=5.42 $Y2=0.815
r237 59 60 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.255 $Y=0.815
+ $X2=4.745 $Y2=0.815
r238 55 90 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.58 $Y=0.725
+ $X2=4.58 $Y2=0.815
r239 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.58 $Y=0.725
+ $X2=4.58 $Y2=0.39
r240 54 89 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.815
+ $X2=3.22 $Y2=0.815
r241 53 90 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=0.815
+ $X2=4.58 $Y2=0.815
r242 53 54 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=4.415 $Y=0.815
+ $X2=3.385 $Y2=0.815
r243 49 89 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.815
r244 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.39
r245 48 88 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0.815
+ $X2=2.38 $Y2=0.815
r246 47 89 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=3.22 $Y2=0.815
r247 47 48 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=2.545 $Y2=0.815
r248 43 88 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.815
r249 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.39
r250 42 87 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r251 41 88 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=2.38 $Y2=0.815
r252 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=1.705 $Y2=0.815
r253 37 87 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r254 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r255 35 87 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r256 35 36 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r257 31 36 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r258 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r259 10 97 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=1.62
r260 9 94 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.125
+ $Y=1.485 $X2=6.26 $Y2=1.62
r261 8 79 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.965
+ $Y=0.235 $X2=7.1 $Y2=0.39
r262 7 69 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.125
+ $Y=0.235 $X2=6.26 $Y2=0.39
r263 6 63 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.235 $X2=5.42 $Y2=0.39
r264 5 57 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.39
r265 4 51 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.39
r266 3 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.39
r267 2 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r268 1 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_4%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 52 56 58 60 63 64 66 67 69 70 72 73 74 75 76 99 110 113 115 119
r144 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r145 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r146 112 113 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=0.235
+ $X2=4.245 $Y2=0.235
r147 108 112 4.67218 $w=6.38e-07 $l=2.5e-07 $layer=LI1_cond $X=3.91 $Y=0.235
+ $X2=4.16 $Y2=0.235
r148 108 110 13.9677 $w=6.38e-07 $l=3.55e-07 $layer=LI1_cond $X=3.91 $Y=0.235
+ $X2=3.555 $Y2=0.235
r149 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r150 103 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r151 103 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.67 $Y2=0
r152 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r153 100 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=6.68 $Y2=0
r154 100 102 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=7.13 $Y2=0
r155 99 118 3.40825 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=7.435 $Y=0
+ $X2=7.627 $Y2=0
r156 99 102 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.435 $Y=0
+ $X2=7.13 $Y2=0
r157 98 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r158 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r159 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r160 95 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=3.91 $Y2=0
r161 94 113 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=4.245 $Y2=0
r162 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r163 91 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r164 90 110 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=3.555 $Y2=0
r165 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r166 87 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r167 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r168 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r169 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r170 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r171 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r172 78 105 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r173 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.69 $Y2=0
r174 76 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r175 76 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r176 74 97 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.75
+ $Y2=0
r177 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.84
+ $Y2=0
r178 72 94 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0 $X2=4.83
+ $Y2=0
r179 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0 $X2=5
+ $Y2=0
r180 71 97 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.085 $Y=0 $X2=5.75
+ $Y2=0
r181 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=0 $X2=5
+ $Y2=0
r182 69 86 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=2.53 $Y2=0
r183 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.8
+ $Y2=0
r184 68 90 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r185 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.8
+ $Y2=0
r186 66 83 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r187 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r188 65 86 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.53 $Y2=0
r189 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r190 63 80 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r191 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r192 62 83 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r193 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r194 58 118 3.40825 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=7.52 $Y=0.085
+ $X2=7.627 $Y2=0
r195 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.52 $Y=0.085
+ $X2=7.52 $Y2=0.39
r196 54 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.68 $Y=0.085
+ $X2=6.68 $Y2=0
r197 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.68 $Y=0.085
+ $X2=6.68 $Y2=0.39
r198 53 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=0 $X2=5.84
+ $Y2=0
r199 52 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.68
+ $Y2=0
r200 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.595 $Y=0
+ $X2=5.925 $Y2=0
r201 48 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.84 $Y=0.085
+ $X2=5.84 $Y2=0
r202 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.84 $Y=0.085
+ $X2=5.84 $Y2=0.39
r203 44 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r204 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.39
r205 40 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r206 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.39
r207 36 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r208 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r209 32 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r210 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r211 28 105 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r212 28 30 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r213 9 60 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.385
+ $Y=0.235 $X2=7.52 $Y2=0.39
r214 8 56 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.545
+ $Y=0.235 $X2=6.68 $Y2=0.39
r215 7 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.84 $Y2=0.39
r216 6 46 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.39
r217 5 112 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.235 $X2=4.16 $Y2=0.39
r218 4 42 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.39
r219 3 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r220 2 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r221 1 30 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


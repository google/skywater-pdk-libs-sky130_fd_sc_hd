* File: sky130_fd_sc_hd__o211a_4.pxi.spice
* Created: Thu Aug 27 14:34:41 2020
* 
x_PM_SKY130_FD_SC_HD__O211A_4%A_79_21# N_A_79_21#_M1017_d N_A_79_21#_M1006_d
+ N_A_79_21#_M1007_d N_A_79_21#_M1019_s N_A_79_21#_c_101_n N_A_79_21#_M1010_g
+ N_A_79_21#_M1004_g N_A_79_21#_c_102_n N_A_79_21#_M1013_g N_A_79_21#_M1008_g
+ N_A_79_21#_c_103_n N_A_79_21#_M1016_g N_A_79_21#_M1018_g N_A_79_21#_c_104_n
+ N_A_79_21#_M1021_g N_A_79_21#_M1020_g N_A_79_21#_c_212_p N_A_79_21#_c_105_n
+ N_A_79_21#_c_106_n N_A_79_21#_c_107_n N_A_79_21#_c_122_p N_A_79_21#_c_118_p
+ N_A_79_21#_c_168_p N_A_79_21#_c_149_p N_A_79_21#_c_145_p N_A_79_21#_c_184_p
+ N_A_79_21#_c_119_p N_A_79_21#_c_108_n N_A_79_21#_c_129_p N_A_79_21#_c_138_p
+ N_A_79_21#_c_156_p N_A_79_21#_c_109_n PM_SKY130_FD_SC_HD__O211A_4%A_79_21#
x_PM_SKY130_FD_SC_HD__O211A_4%B1 N_B1_M1006_g N_B1_M1000_g N_B1_M1022_g
+ N_B1_M1009_g N_B1_c_262_n N_B1_c_263_n N_B1_c_290_n B1 N_B1_c_264_n
+ N_B1_c_265_n N_B1_c_273_n N_B1_c_266_n N_B1_c_274_n B1
+ PM_SKY130_FD_SC_HD__O211A_4%B1
x_PM_SKY130_FD_SC_HD__O211A_4%C1 N_C1_c_356_n N_C1_M1017_g N_C1_M1003_g
+ N_C1_c_357_n N_C1_M1011_g N_C1_M1007_g C1 N_C1_c_358_n N_C1_c_359_n
+ PM_SKY130_FD_SC_HD__O211A_4%C1
x_PM_SKY130_FD_SC_HD__O211A_4%A1 N_A1_M1014_g N_A1_M1005_g N_A1_M1015_g
+ N_A1_M1012_g N_A1_c_402_n N_A1_c_403_n N_A1_c_417_n N_A1_c_420_n A1
+ N_A1_c_404_n N_A1_c_405_n N_A1_c_412_n N_A1_c_406_n N_A1_c_451_p
+ PM_SKY130_FD_SC_HD__O211A_4%A1
x_PM_SKY130_FD_SC_HD__O211A_4%A2 N_A2_c_484_n N_A2_M1001_g N_A2_M1019_g
+ N_A2_c_485_n N_A2_M1002_g N_A2_M1023_g A2 N_A2_c_486_n N_A2_c_487_n
+ PM_SKY130_FD_SC_HD__O211A_4%A2
x_PM_SKY130_FD_SC_HD__O211A_4%VPWR N_VPWR_M1004_s N_VPWR_M1008_s N_VPWR_M1020_s
+ N_VPWR_M1003_s N_VPWR_M1009_s N_VPWR_M1012_d N_VPWR_c_537_n N_VPWR_c_538_n
+ N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n
+ N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n
+ VPWR N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_536_n PM_SKY130_FD_SC_HD__O211A_4%VPWR
x_PM_SKY130_FD_SC_HD__O211A_4%X N_X_M1010_s N_X_M1016_s N_X_M1004_d N_X_M1018_d
+ N_X_c_652_n N_X_c_647_n N_X_c_648_n N_X_c_692_p N_X_c_657_n N_X_c_678_n
+ N_X_c_649_n N_X_c_695_p N_X_c_682_n N_X_c_667_n N_X_c_650_n X N_X_c_645_n X
+ PM_SKY130_FD_SC_HD__O211A_4%X
x_PM_SKY130_FD_SC_HD__O211A_4%VGND N_VGND_M1010_d N_VGND_M1013_d N_VGND_M1021_d
+ N_VGND_M1014_d N_VGND_M1002_s N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n
+ N_VGND_c_713_n N_VGND_c_714_n N_VGND_c_715_n VGND N_VGND_c_716_n
+ N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n
+ N_VGND_c_722_n N_VGND_c_723_n N_VGND_c_724_n N_VGND_c_725_n
+ PM_SKY130_FD_SC_HD__O211A_4%VGND
x_PM_SKY130_FD_SC_HD__O211A_4%A_474_47# N_A_474_47#_M1000_s N_A_474_47#_M1022_s
+ N_A_474_47#_M1001_d N_A_474_47#_M1015_s N_A_474_47#_c_812_n
+ N_A_474_47#_c_830_n N_A_474_47#_c_819_n N_A_474_47#_c_832_n
+ N_A_474_47#_c_820_n N_A_474_47#_c_838_n N_A_474_47#_c_813_n
+ N_A_474_47#_c_814_n N_A_474_47#_c_854_n PM_SKY130_FD_SC_HD__O211A_4%A_474_47#
cc_1 VNB N_A_79_21#_c_101_n 0.0182637f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_102_n 0.0157727f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_103_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_104_n 0.0188049f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_105_n 0.00434115f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.065
cc_6 VNB N_A_79_21#_c_106_n 2.29655e-19 $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.855
cc_7 VNB N_A_79_21#_c_107_n 0.00522718f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.725
cc_8 VNB N_A_79_21#_c_108_n 0.00120371f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.165
cc_9 VNB N_A_79_21#_c_109_n 0.0936275f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.16
cc_10 VNB N_B1_c_262_n 0.0036285f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.985
cc_11 VNB N_B1_c_263_n 0.0226435f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.985
cc_12 VNB N_B1_c_264_n 0.0190789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B1_c_265_n 0.0261696f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_14 VNB N_B1_c_266_n 0.0170444f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=1.985
cc_15 VNB N_C1_c_356_n 0.0171751f $X=-0.19 $Y=-0.24 $X2=3.145 $Y2=0.235
cc_16 VNB N_C1_c_357_n 0.0178707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C1_c_358_n 0.00159247f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_18 VNB N_C1_c_359_n 0.0401802f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.325
cc_19 VNB N_A1_c_402_n 0.00191336f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.985
cc_20 VNB N_A1_c_403_n 0.0238912f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.985
cc_21 VNB N_A1_c_404_n 0.0179853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_405_n 0.0403853f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_23 VNB N_A1_c_406_n 0.0223198f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=1.985
cc_24 VNB N_A2_c_484_n 0.0173848f $X=-0.19 $Y=-0.24 $X2=3.145 $Y2=0.235
cc_25 VNB N_A2_c_485_n 0.0164438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A2_c_486_n 0.0322691f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_27 VNB N_A2_c_487_n 0.00366561f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_28 VNB N_VPWR_c_536_n 0.269736f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.16
cc_29 VNB N_X_c_645_n 0.0076991f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.16
cc_30 VNB X 0.0253091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_710_n 0.0102584f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.325
cc_32 VNB N_VGND_c_711_n 0.0118704f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.985
cc_33 VNB N_VGND_c_712_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_34 VNB N_VGND_c_713_n 0.00556717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_714_n 0.00491058f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=1.325
cc_36 VNB N_VGND_c_715_n 0.00422004f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_37 VNB N_VGND_c_716_n 0.0109337f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_38 VNB N_VGND_c_717_n 0.0116974f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=1.16
cc_39 VNB N_VGND_c_718_n 0.0581773f $X=-0.19 $Y=-0.24 $X2=2.06 $Y2=1.16
cc_40 VNB N_VGND_c_719_n 0.0165909f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.725
cc_41 VNB N_VGND_c_720_n 0.0171884f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=2.3
cc_42 VNB N_VGND_c_721_n 0.317934f $X=-0.19 $Y=-0.24 $X2=2.895 $Y2=2.3
cc_43 VNB N_VGND_c_722_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=2.3
cc_44 VNB N_VGND_c_723_n 0.00574413f $X=-0.19 $Y=-0.24 $X2=4.12 $Y2=1.94
cc_45 VNB N_VGND_c_724_n 0.00602253f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.165
cc_46 VNB N_VGND_c_725_n 0.00361995f $X=-0.19 $Y=-0.24 $X2=5.32 $Y2=1.94
cc_47 VNB N_A_474_47#_c_812_n 0.00255878f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_48 VNB N_A_474_47#_c_813_n 0.00872789f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.985
cc_49 VNB N_A_474_47#_c_814_n 0.0172776f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_50 VPB N_A_79_21#_M1004_g 0.0217968f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.985
cc_51 VPB N_A_79_21#_M1008_g 0.0180969f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.985
cc_52 VPB N_A_79_21#_M1018_g 0.0180889f $X=-0.19 $Y=1.305 $X2=1.72 $Y2=1.985
cc_53 VPB N_A_79_21#_M1020_g 0.0178732f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_54 VPB N_A_79_21#_c_106_n 0.00106471f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=1.855
cc_55 VPB N_A_79_21#_c_109_n 0.0215037f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.16
cc_56 VPB N_B1_M1006_g 0.0201829f $X=-0.19 $Y=1.305 $X2=3.74 $Y2=1.485
cc_57 VPB N_B1_M1009_g 0.0197154f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_58 VPB N_B1_c_262_n 0.00159694f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.985
cc_59 VPB N_B1_c_263_n 0.0053819f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.985
cc_60 VPB B1 2.77229e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_61 VPB N_B1_c_265_n 0.00647903f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_62 VPB N_B1_c_273_n 0.00127557f $X=-0.19 $Y=1.305 $X2=1.72 $Y2=1.325
cc_63 VPB N_B1_c_274_n 0.0136495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_C1_M1003_g 0.0204388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_C1_M1007_g 0.0194958f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_66 VPB N_C1_c_359_n 0.00882602f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.325
cc_67 VPB N_A1_M1005_g 0.0179515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A1_M1012_g 0.0225654f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_69 VPB N_A1_c_402_n 0.00287769f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.985
cc_70 VPB N_A1_c_403_n 0.00633775f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.985
cc_71 VPB N_A1_c_405_n 0.00932547f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_72 VPB N_A1_c_412_n 0.00610505f $X=-0.19 $Y=1.305 $X2=1.72 $Y2=1.325
cc_73 VPB N_A2_M1019_g 0.0190317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A2_M1023_g 0.0190427f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_75 VPB N_A2_c_486_n 0.0058739f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_76 VPB N_A2_c_487_n 4.7433e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_77 VPB N_VPWR_c_537_n 0.026733f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_78 VPB N_VPWR_c_538_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.985
cc_79 VPB N_VPWR_c_539_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_80 VPB N_VPWR_c_540_n 4.21859e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_541_n 0.0158785f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_82 VPB N_VPWR_c_542_n 0.00473001f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_83 VPB N_VPWR_c_543_n 0.0103398f $X=-0.19 $Y=1.305 $X2=2.2 $Y2=1.165
cc_84 VPB N_VPWR_c_544_n 0.0263776f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=1.16
cc_85 VPB N_VPWR_c_545_n 0.0130339f $X=-0.19 $Y=1.305 $X2=2.06 $Y2=1.165
cc_86 VPB N_VPWR_c_546_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.06 $Y2=1.16
cc_87 VPB N_VPWR_c_547_n 0.0129398f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=0.815
cc_88 VPB N_VPWR_c_548_n 0.00436475f $X=-0.19 $Y=1.305 $X2=2.285 $Y2=1.065
cc_89 VPB N_VPWR_c_549_n 0.0174178f $X=-0.19 $Y=1.305 $X2=2.37 $Y2=0.725
cc_90 VPB N_VPWR_c_550_n 0.0169255f $X=-0.19 $Y=1.305 $X2=3.952 $Y2=2.025
cc_91 VPB N_VPWR_c_551_n 0.0396606f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=1.94
cc_92 VPB N_VPWR_c_552_n 0.00510842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_93 VPB N_VPWR_c_553_n 0.00436502f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.16
cc_94 VPB N_VPWR_c_554_n 0.00506838f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_95 VPB N_VPWR_c_536_n 0.0596437f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.16
cc_96 VPB N_X_c_647_n 0.00960895f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_97 VPB N_X_c_648_n 0.0248561f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.325
cc_98 VPB N_X_c_649_n 0.00496901f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_99 VPB N_X_c_650_n 0.00135109f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_100 VPB X 0.00756881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 N_A_79_21#_M1020_g N_B1_M1006_g 0.0390217f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_106_n N_B1_M1006_g 0.00578089f $X=2.285 $Y=1.855 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_118_p N_B1_M1006_g 0.0138053f $X=2.7 $Y=1.94 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_119_p N_B1_M1009_g 0.0127781f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_105_n N_B1_c_262_n 0.00517151f $X=2.285 $Y=1.065 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_106_n N_B1_c_262_n 0.0132839f $X=2.285 $Y=1.855 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_122_p N_B1_c_262_n 0.0180373f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_108_n N_B1_c_262_n 0.0167177f $X=2.285 $Y=1.165 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_109_n N_B1_c_262_n 4.16906e-19 $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_105_n N_B1_c_263_n 4.54171e-19 $X=2.285 $Y=1.065 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_106_n N_B1_c_263_n 3.88943e-19 $X=2.285 $Y=1.855 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_122_p N_B1_c_263_n 0.00256568f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_108_n N_B1_c_263_n 0.00149504f $X=2.285 $Y=1.165 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_129_p N_B1_c_263_n 2.90672e-19 $X=2.88 $Y=1.94 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_109_n N_B1_c_263_n 0.0151048f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_79_21#_M1006_d N_B1_c_290_n 0.00129533f $X=2.655 $Y=1.485 $X2=0 $Y2=0
cc_117 N_A_79_21#_M1020_g N_B1_c_290_n 2.27197e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_106_n N_B1_c_290_n 0.0189163f $X=2.285 $Y=1.855 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_118_p N_B1_c_290_n 0.00872871f $X=2.7 $Y=1.94 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_129_p N_B1_c_290_n 0.0105655f $X=2.88 $Y=1.94 $X2=0 $Y2=0
cc_121 N_A_79_21#_M1007_d B1 0.00134822f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_119_p B1 0.0113072f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_138_p B1 0.0109646f $X=3.952 $Y=1.94 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_105_n N_B1_c_264_n 0.00553512f $X=2.285 $Y=1.065 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_122_p N_B1_c_264_n 0.0121531f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_138_p N_B1_c_265_n 5.45953e-19 $X=3.952 $Y=1.94 $X2=0 $Y2=0
cc_127 N_A_79_21#_M1006_d N_B1_c_274_n 0.00437665f $X=2.655 $Y=1.485 $X2=0 $Y2=0
cc_128 N_A_79_21#_M1007_d N_B1_c_274_n 0.00192038f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_122_p N_B1_c_274_n 0.00556051f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_145_p N_B1_c_274_n 0.036434f $X=3.785 $Y=1.94 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_129_p N_B1_c_274_n 0.0189546f $X=2.88 $Y=1.94 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_138_p N_B1_c_274_n 0.0125956f $X=3.952 $Y=1.94 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_122_p N_C1_c_356_n 0.0117025f $X=3.355 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_79_21#_c_149_p N_C1_M1003_g 0.0075892f $X=2.895 $Y=2.3 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_145_p N_C1_M1003_g 0.0127965f $X=3.785 $Y=1.94 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_122_p N_C1_c_357_n 0.00315994f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_145_p N_C1_M1007_g 0.0123549f $X=3.785 $Y=1.94 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_122_p N_C1_c_358_n 0.0256515f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_122_p N_C1_c_359_n 0.00667699f $X=3.355 $Y=0.73 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_119_p N_A1_M1005_g 0.0122497f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_156_p N_A1_M1005_g 0.00164393f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_156_p N_A1_M1012_g 0.00190709f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_119_p N_A1_c_403_n 4.56052e-19 $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_144 N_A_79_21#_M1019_s N_A1_c_417_n 0.00331619f $X=5.18 $Y=1.485 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_119_p N_A1_c_417_n 0.0178501f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_156_p N_A1_c_417_n 0.0172104f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_119_p N_A1_c_420_n 0.0186703f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_119_p N_A2_M1019_g 0.00866486f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_156_p N_A2_M1019_g 0.00900867f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_156_p N_A2_M1023_g 0.0112998f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_106_n N_VPWR_M1020_s 0.00357053f $X=2.285 $Y=1.855 $X2=0
+ $Y2=0
cc_152 N_A_79_21#_c_118_p N_VPWR_M1020_s 0.00374269f $X=2.7 $Y=1.94 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_168_p N_VPWR_M1020_s 9.4656e-19 $X=2.37 $Y=1.94 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_145_p N_VPWR_M1003_s 0.0033738f $X=3.785 $Y=1.94 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_119_p N_VPWR_M1009_s 0.00846156f $X=5.155 $Y=1.94 $X2=0
+ $Y2=0
cc_156 N_A_79_21#_M1004_g N_VPWR_c_537_n 0.0114143f $X=0.86 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_79_21#_M1008_g N_VPWR_c_537_n 6.1315e-19 $X=1.29 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_79_21#_M1004_g N_VPWR_c_538_n 6.22378e-19 $X=0.86 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_79_21#_M1008_g N_VPWR_c_538_n 0.0104876f $X=1.29 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_79_21#_M1018_g N_VPWR_c_538_n 0.0103509f $X=1.72 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_79_21#_M1020_g N_VPWR_c_538_n 6.1315e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_79_21#_M1018_g N_VPWR_c_539_n 5.1979e-19 $X=1.72 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_79_21#_M1020_g N_VPWR_c_539_n 0.00698285f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_79_21#_c_118_p N_VPWR_c_539_n 0.00753139f $X=2.7 $Y=1.94 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_168_p N_VPWR_c_539_n 0.00915804f $X=2.37 $Y=1.94 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_149_p N_VPWR_c_540_n 0.0170139f $X=2.895 $Y=2.3 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_145_p N_VPWR_c_540_n 0.0162971f $X=3.785 $Y=1.94 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_145_p N_VPWR_c_541_n 0.00215462f $X=3.785 $Y=1.94 $X2=0
+ $Y2=0
cc_169 N_A_79_21#_c_184_p N_VPWR_c_541_n 0.0212772f $X=3.95 $Y=2.3 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_119_p N_VPWR_c_541_n 0.00229661f $X=5.155 $Y=1.94 $X2=0
+ $Y2=0
cc_171 N_A_79_21#_c_119_p N_VPWR_c_542_n 0.0159967f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_172 N_A_79_21#_c_156_p N_VPWR_c_544_n 0.0164451f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_173 N_A_79_21#_M1004_g N_VPWR_c_545_n 0.00486043f $X=0.86 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_79_21#_M1008_g N_VPWR_c_545_n 0.00486043f $X=1.29 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_79_21#_M1018_g N_VPWR_c_547_n 0.00486043f $X=1.72 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_79_21#_M1020_g N_VPWR_c_547_n 0.00486043f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_79_21#_c_118_p N_VPWR_c_550_n 0.00215462f $X=2.7 $Y=1.94 $X2=0 $Y2=0
cc_178 N_A_79_21#_c_149_p N_VPWR_c_550_n 0.0245983f $X=2.895 $Y=2.3 $X2=0 $Y2=0
cc_179 N_A_79_21#_c_145_p N_VPWR_c_550_n 0.00291008f $X=3.785 $Y=1.94 $X2=0
+ $Y2=0
cc_180 N_A_79_21#_c_119_p N_VPWR_c_551_n 0.00780235f $X=5.155 $Y=1.94 $X2=0
+ $Y2=0
cc_181 N_A_79_21#_c_156_p N_VPWR_c_551_n 0.0188082f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_182 N_A_79_21#_M1006_d N_VPWR_c_536_n 0.00471965f $X=2.655 $Y=1.485 $X2=0
+ $Y2=0
cc_183 N_A_79_21#_M1007_d N_VPWR_c_536_n 0.00335196f $X=3.74 $Y=1.485 $X2=0
+ $Y2=0
cc_184 N_A_79_21#_M1019_s N_VPWR_c_536_n 0.00223231f $X=5.18 $Y=1.485 $X2=0
+ $Y2=0
cc_185 N_A_79_21#_M1004_g N_VPWR_c_536_n 0.00822531f $X=0.86 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_79_21#_M1008_g N_VPWR_c_536_n 0.00822531f $X=1.29 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_79_21#_M1018_g N_VPWR_c_536_n 0.00822531f $X=1.72 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_79_21#_M1020_g N_VPWR_c_536_n 0.00822531f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_79_21#_c_118_p N_VPWR_c_536_n 0.00463328f $X=2.7 $Y=1.94 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_168_p N_VPWR_c_536_n 7.65976e-19 $X=2.37 $Y=1.94 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_149_p N_VPWR_c_536_n 0.0137481f $X=2.895 $Y=2.3 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_145_p N_VPWR_c_536_n 0.0107826f $X=3.785 $Y=1.94 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_184_p N_VPWR_c_536_n 0.012788f $X=3.95 $Y=2.3 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_119_p N_VPWR_c_536_n 0.0196162f $X=5.155 $Y=1.94 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_156_p N_VPWR_c_536_n 0.0122321f $X=5.32 $Y=2.02 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_101_n N_X_c_652_n 0.014584f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_79_21#_c_212_p N_X_c_652_n 0.00172614f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_198 N_A_79_21#_M1004_g N_X_c_647_n 0.0207716f $X=0.86 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_79_21#_c_212_p N_X_c_647_n 0.0327402f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_200 N_A_79_21#_c_109_n N_X_c_647_n 0.0115443f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_79_21#_c_102_n N_X_c_657_n 0.0125611f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_79_21#_c_103_n N_X_c_657_n 0.0121263f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_212_p N_X_c_657_n 0.0373312f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_204 N_A_79_21#_c_109_n N_X_c_657_n 0.00433322f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_79_21#_M1008_g N_X_c_649_n 0.0175819f $X=1.29 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_79_21#_M1018_g N_X_c_649_n 0.0170821f $X=1.72 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_79_21#_M1020_g N_X_c_649_n 0.00111897f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_212_p N_X_c_649_n 0.0652299f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_209 N_A_79_21#_c_106_n N_X_c_649_n 0.0113079f $X=2.285 $Y=1.855 $X2=0 $Y2=0
cc_210 N_A_79_21#_c_109_n N_X_c_649_n 0.00502261f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_79_21#_c_212_p N_X_c_667_n 0.00917312f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_212 N_A_79_21#_c_109_n N_X_c_667_n 0.00214922f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_79_21#_c_212_p N_X_c_650_n 0.0146791f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_214 N_A_79_21#_c_109_n N_X_c_650_n 0.00263158f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_79_21#_c_101_n X 0.0191249f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_79_21#_M1004_g X 0.00304213f $X=0.86 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_79_21#_c_212_p X 0.0164096f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_218 N_A_79_21#_c_119_p A_950_297# 0.00483504f $X=5.155 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_79_21#_c_101_n N_VGND_c_711_n 0.00774571f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_79_21#_c_102_n N_VGND_c_711_n 5.08801e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_79_21#_c_101_n N_VGND_c_712_n 5.02907e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_79_21#_c_102_n N_VGND_c_712_n 0.00643498f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_79_21#_c_103_n N_VGND_c_712_n 0.00643498f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_79_21#_c_104_n N_VGND_c_712_n 5.02907e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_c_103_n N_VGND_c_713_n 5.1088e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_79_21#_c_104_n N_VGND_c_713_n 0.00821699f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_79_21#_c_212_p N_VGND_c_713_n 0.00960079f $X=2.2 $Y=1.165 $X2=0 $Y2=0
cc_228 N_A_79_21#_c_109_n N_VGND_c_713_n 0.00655194f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_79_21#_c_101_n N_VGND_c_716_n 0.00339367f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A_79_21#_c_102_n N_VGND_c_716_n 0.00337001f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_c_103_n N_VGND_c_717_n 0.00337001f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_c_104_n N_VGND_c_717_n 0.0046653f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_79_21#_c_107_n N_VGND_c_718_n 0.00263957f $X=2.37 $Y=0.725 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_M1017_d N_VGND_c_721_n 0.00358802f $X=3.145 $Y=0.235 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_c_101_n N_VGND_c_721_n 0.00394406f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_102_n N_VGND_c_721_n 0.00390568f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_103_n N_VGND_c_721_n 0.00390568f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_79_21#_c_104_n N_VGND_c_721_n 0.00789179f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_79_21#_c_107_n N_VGND_c_721_n 0.00401338f $X=2.37 $Y=0.725 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_c_122_p N_A_474_47#_M1000_s 0.00844235f $X=3.355 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_241 N_A_79_21#_M1017_d N_A_474_47#_c_812_n 0.0074793f $X=3.145 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_79_21#_c_107_n N_A_474_47#_c_812_n 0.00323932f $X=2.37 $Y=0.725 $X2=0
+ $Y2=0
cc_243 N_A_79_21#_c_122_p N_A_474_47#_c_812_n 0.0634213f $X=3.355 $Y=0.73 $X2=0
+ $Y2=0
cc_244 N_A_79_21#_c_122_p N_A_474_47#_c_819_n 0.00188177f $X=3.355 $Y=0.73 $X2=0
+ $Y2=0
cc_245 N_A_79_21#_c_122_p N_A_474_47#_c_820_n 0.00408942f $X=3.355 $Y=0.73 $X2=0
+ $Y2=0
cc_246 N_A_79_21#_c_122_p A_748_47# 0.00295109f $X=3.355 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_247 N_B1_c_264_n N_C1_c_356_n 0.0399566f $X=2.637 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_248 N_B1_M1006_g N_C1_M1003_g 0.0248212f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B1_c_262_n N_C1_M1003_g 0.00246052f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B1_c_274_n N_C1_M1003_g 0.014578f $X=3.95 $Y=1.565 $X2=0 $Y2=0
cc_251 N_B1_c_266_n N_C1_c_357_n 0.0411449f $X=4.115 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_M1009_g N_C1_M1007_g 0.0315817f $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_253 N_B1_c_273_n N_C1_M1007_g 0.0027946f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_c_274_n N_C1_M1007_g 0.0139524f $X=3.95 $Y=1.565 $X2=0 $Y2=0
cc_255 N_B1_c_262_n N_C1_c_358_n 0.0160184f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_263_n N_C1_c_358_n 2.49806e-19 $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B1_c_265_n N_C1_c_358_n 8.27404e-19 $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_273_n N_C1_c_358_n 0.0160381f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B1_c_274_n N_C1_c_358_n 0.0504691f $X=3.95 $Y=1.565 $X2=0 $Y2=0
cc_260 N_B1_c_262_n N_C1_c_359_n 0.00380744f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B1_c_263_n N_C1_c_359_n 0.0399566f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_262 N_B1_c_265_n N_C1_c_359_n 0.0219138f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_c_273_n N_C1_c_359_n 6.8991e-19 $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_c_274_n N_C1_c_359_n 0.00736789f $X=3.95 $Y=1.565 $X2=0 $Y2=0
cc_265 N_B1_M1009_g N_A1_M1005_g 0.038511f $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_266 B1 N_A1_M1005_g 2.61793e-19 $X=3.82 $Y=1.445 $X2=0 $Y2=0
cc_267 N_B1_M1009_g N_A1_c_402_n 9.53614e-19 $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_268 B1 N_A1_c_402_n 0.00354633f $X=3.82 $Y=1.445 $X2=0 $Y2=0
cc_269 N_B1_c_265_n N_A1_c_402_n 0.0010097f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B1_c_273_n N_A1_c_402_n 0.0265747f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B1_c_265_n N_A1_c_403_n 0.020645f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_273_n N_A1_c_403_n 0.00101004f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B1_M1009_g N_A1_c_420_n 8.26999e-19 $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_274 B1 N_A1_c_420_n 0.0140905f $X=3.82 $Y=1.445 $X2=0 $Y2=0
cc_275 N_B1_c_266_n N_A1_c_404_n 0.0105489f $X=4.115 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B1_c_274_n N_VPWR_M1003_s 0.00178782f $X=3.95 $Y=1.565 $X2=0 $Y2=0
cc_277 N_B1_M1006_g N_VPWR_c_539_n 0.00826871f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1006_g N_VPWR_c_540_n 8.85136e-19 $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_M1009_g N_VPWR_c_540_n 4.91952e-19 $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B1_M1009_g N_VPWR_c_541_n 0.00433717f $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B1_M1009_g N_VPWR_c_542_n 0.00177885f $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B1_M1006_g N_VPWR_c_550_n 0.00360664f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_283 N_B1_M1006_g N_VPWR_c_536_n 0.00477256f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B1_M1009_g N_VPWR_c_536_n 0.00615213f $X=4.205 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B1_c_264_n N_VGND_c_713_n 0.002364f $X=2.637 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B1_c_264_n N_VGND_c_718_n 0.00357877f $X=2.637 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B1_c_266_n N_VGND_c_718_n 0.00357877f $X=4.115 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B1_c_264_n N_VGND_c_721_n 0.00641668f $X=2.637 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B1_c_266_n N_VGND_c_721_n 0.00542429f $X=4.115 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B1_c_264_n N_A_474_47#_c_812_n 0.00812316f $X=2.637 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_B1_c_265_n N_A_474_47#_c_812_n 0.00102667f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_273_n N_A_474_47#_c_812_n 0.00548502f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_293 N_B1_c_266_n N_A_474_47#_c_812_n 0.0106221f $X=4.115 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B1_c_265_n N_A_474_47#_c_820_n 0.00296796f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_295 N_B1_c_273_n N_A_474_47#_c_820_n 0.00688852f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_296 N_C1_M1003_g N_VPWR_c_539_n 8.71023e-19 $X=3.235 $Y=1.985 $X2=0 $Y2=0
cc_297 N_C1_M1003_g N_VPWR_c_540_n 0.00871505f $X=3.235 $Y=1.985 $X2=0 $Y2=0
cc_298 N_C1_M1007_g N_VPWR_c_540_n 0.00743575f $X=3.665 $Y=1.985 $X2=0 $Y2=0
cc_299 N_C1_M1007_g N_VPWR_c_541_n 0.00360664f $X=3.665 $Y=1.985 $X2=0 $Y2=0
cc_300 N_C1_M1003_g N_VPWR_c_550_n 0.00360664f $X=3.235 $Y=1.985 $X2=0 $Y2=0
cc_301 N_C1_M1003_g N_VPWR_c_536_n 0.00477256f $X=3.235 $Y=1.985 $X2=0 $Y2=0
cc_302 N_C1_M1007_g N_VPWR_c_536_n 0.00455826f $X=3.665 $Y=1.985 $X2=0 $Y2=0
cc_303 N_C1_c_356_n N_VGND_c_718_n 0.00357877f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_304 N_C1_c_357_n N_VGND_c_718_n 0.00357877f $X=3.665 $Y=0.995 $X2=0 $Y2=0
cc_305 N_C1_c_356_n N_VGND_c_721_n 0.00554055f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_306 N_C1_c_357_n N_VGND_c_721_n 0.0057288f $X=3.665 $Y=0.995 $X2=0 $Y2=0
cc_307 N_C1_c_356_n N_A_474_47#_c_812_n 0.0116665f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_308 N_C1_c_357_n N_A_474_47#_c_812_n 0.0141822f $X=3.665 $Y=0.995 $X2=0 $Y2=0
cc_309 N_C1_c_358_n N_A_474_47#_c_812_n 0.00504034f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A1_c_404_n N_A2_c_484_n 0.0216207f $X=4.655 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_311 N_A1_M1005_g N_A2_M1019_g 0.0580745f $X=4.675 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A1_c_417_n N_A2_M1019_g 0.0112197f $X=5.89 $Y=1.59 $X2=0 $Y2=0
cc_313 N_A1_c_406_n N_A2_c_485_n 0.0264199f $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A1_M1012_g N_A2_M1023_g 0.0571498f $X=5.965 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A1_c_417_n N_A2_M1023_g 0.0151007f $X=5.89 $Y=1.59 $X2=0 $Y2=0
cc_316 N_A1_c_412_n N_A2_M1023_g 0.00105271f $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A1_c_402_n N_A2_c_486_n 0.00496582f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A1_c_403_n N_A2_c_486_n 0.0220248f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A1_c_417_n N_A2_c_486_n 0.00369289f $X=5.89 $Y=1.59 $X2=0 $Y2=0
cc_320 N_A1_c_405_n N_A2_c_486_n 0.0217001f $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A1_c_412_n N_A2_c_486_n 3.39822e-19 $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A1_c_402_n N_A2_c_487_n 0.022781f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A1_c_403_n N_A2_c_487_n 3.42061e-19 $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A1_c_417_n N_A2_c_487_n 0.0428079f $X=5.89 $Y=1.59 $X2=0 $Y2=0
cc_325 N_A1_c_405_n N_A2_c_487_n 0.0018092f $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A1_c_412_n N_A2_c_487_n 0.0230799f $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A1_c_420_n N_VPWR_M1009_s 0.00239683f $X=4.845 $Y=1.59 $X2=0 $Y2=0
cc_328 N_A1_c_412_n N_VPWR_M1012_d 3.80768e-19 $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A1_c_451_p N_VPWR_M1012_d 0.0116956f $X=6.09 $Y=1.495 $X2=0 $Y2=0
cc_330 N_A1_M1005_g N_VPWR_c_542_n 0.00291543f $X=4.675 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A1_M1012_g N_VPWR_c_544_n 0.0162084f $X=5.965 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A1_c_405_n N_VPWR_c_544_n 8.5021e-19 $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A1_c_451_p N_VPWR_c_544_n 0.0153578f $X=6.09 $Y=1.495 $X2=0 $Y2=0
cc_334 N_A1_M1005_g N_VPWR_c_551_n 0.00433717f $X=4.675 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A1_M1012_g N_VPWR_c_551_n 0.00486043f $X=5.965 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A1_M1005_g N_VPWR_c_536_n 0.00604372f $X=4.675 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A1_M1012_g N_VPWR_c_536_n 0.0083285f $X=5.965 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A1_c_417_n A_950_297# 0.00396291f $X=5.89 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_339 N_A1_c_420_n A_950_297# 4.09894e-19 $X=4.845 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_340 N_A1_c_417_n A_1122_297# 0.00942166f $X=5.89 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_341 N_A1_c_404_n N_VGND_c_714_n 0.00315768f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A1_c_406_n N_VGND_c_715_n 0.00275982f $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A1_c_404_n N_VGND_c_718_n 0.00428647f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A1_c_406_n N_VGND_c_720_n 0.0042256f $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A1_c_404_n N_VGND_c_721_n 0.00615671f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A1_c_406_n N_VGND_c_721_n 0.00668068f $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_347 N_A1_c_404_n N_A_474_47#_c_830_n 0.00202761f $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_348 N_A1_c_404_n N_A_474_47#_c_819_n 0.00374965f $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A1_c_402_n N_A_474_47#_c_832_n 0.0245945f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A1_c_403_n N_A_474_47#_c_832_n 0.00454565f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A1_c_417_n N_A_474_47#_c_832_n 0.00349677f $X=5.89 $Y=1.59 $X2=0 $Y2=0
cc_352 N_A1_c_404_n N_A_474_47#_c_832_n 0.0100368f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_353 N_A1_c_402_n N_A_474_47#_c_820_n 7.53006e-19 $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A1_c_404_n N_A_474_47#_c_820_n 2.73532e-19 $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A1_c_404_n N_A_474_47#_c_838_n 5.15871e-19 $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A1_c_406_n N_A_474_47#_c_838_n 5.11235e-19 $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A1_c_417_n N_A_474_47#_c_813_n 0.0035106f $X=5.89 $Y=1.59 $X2=0 $Y2=0
cc_358 N_A1_c_405_n N_A_474_47#_c_813_n 0.00591814f $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A1_c_412_n N_A_474_47#_c_813_n 0.0304103f $X=6.085 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A1_c_406_n N_A_474_47#_c_813_n 0.00936114f $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A1_c_406_n N_A_474_47#_c_814_n 0.00587404f $X=6.09 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A2_M1023_g N_VPWR_c_544_n 0.00273322f $X=5.535 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A2_M1019_g N_VPWR_c_551_n 0.0042256f $X=5.105 $Y=1.985 $X2=0 $Y2=0
cc_364 N_A2_M1023_g N_VPWR_c_551_n 0.0054895f $X=5.535 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A2_M1019_g N_VPWR_c_536_n 0.00592932f $X=5.105 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A2_M1023_g N_VPWR_c_536_n 0.00996518f $X=5.535 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A2_c_484_n N_VGND_c_714_n 0.00339147f $X=5.105 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A2_c_485_n N_VGND_c_715_n 0.00151324f $X=5.535 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A2_c_484_n N_VGND_c_719_n 0.0042256f $X=5.105 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A2_c_485_n N_VGND_c_719_n 0.0042256f $X=5.535 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A2_c_484_n N_VGND_c_721_n 0.00604526f $X=5.105 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A2_c_485_n N_VGND_c_721_n 0.00574807f $X=5.535 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A2_c_484_n N_A_474_47#_c_819_n 5.28584e-19 $X=5.105 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A2_c_484_n N_A_474_47#_c_832_n 0.00923148f $X=5.105 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A2_c_487_n N_A_474_47#_c_832_n 0.00880077f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_376 N_A2_c_484_n N_A_474_47#_c_838_n 0.00634828f $X=5.105 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A2_c_485_n N_A_474_47#_c_838_n 0.00587404f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A2_c_485_n N_A_474_47#_c_813_n 0.00866486f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A2_c_486_n N_A_474_47#_c_813_n 0.00150953f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_380 N_A2_c_487_n N_A_474_47#_c_813_n 0.0137766f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_381 N_A2_c_485_n N_A_474_47#_c_814_n 5.11235e-19 $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A2_c_484_n N_A_474_47#_c_854_n 7.16038e-19 $X=5.105 $Y=0.995 $X2=0
+ $Y2=0
cc_383 N_A2_c_485_n N_A_474_47#_c_854_n 7.16038e-19 $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_384 N_A2_c_486_n N_A_474_47#_c_854_n 0.00243264f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A2_c_487_n N_A_474_47#_c_854_n 0.0215186f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_386 N_VPWR_c_536_n N_X_M1004_d 0.00570388f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_536_n N_X_M1018_d 0.00535672f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_M1004_s N_X_c_647_n 0.00324835f $X=0.52 $Y=1.485 $X2=0 $Y2=0
cc_389 N_VPWR_c_537_n N_X_c_647_n 0.0226846f $X=0.645 $Y=1.955 $X2=0 $Y2=0
cc_390 N_VPWR_c_545_n N_X_c_678_n 0.012099f $X=1.34 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_536_n N_X_c_678_n 0.00684987f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_M1008_s N_X_c_649_n 0.00178891f $X=1.365 $Y=1.485 $X2=0 $Y2=0
cc_393 N_VPWR_c_538_n N_X_c_649_n 0.0176092f $X=1.505 $Y=1.955 $X2=0 $Y2=0
cc_394 N_VPWR_c_547_n N_X_c_682_n 0.0124538f $X=2.2 $Y=2.72 $X2=0 $Y2=0
cc_395 N_VPWR_c_536_n N_X_c_682_n 0.00724021f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_c_536_n A_950_297# 0.00351559f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_397 N_VPWR_c_536_n A_1122_297# 0.0119688f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_398 N_X_c_645_n N_VGND_M1010_d 0.00291379f $X=0.225 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_399 X N_VGND_M1010_d 3.49814e-19 $X=0.23 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_400 N_X_c_657_n N_VGND_M1013_d 0.00335113f $X=1.435 $Y=0.71 $X2=0 $Y2=0
cc_401 N_X_c_645_n N_VGND_c_710_n 2.03606e-19 $X=0.225 $Y=0.805 $X2=0 $Y2=0
cc_402 N_X_c_652_n N_VGND_c_711_n 0.0020301f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_403 N_X_c_645_n N_VGND_c_711_n 0.0205224f $X=0.225 $Y=0.805 $X2=0 $Y2=0
cc_404 N_X_c_657_n N_VGND_c_712_n 0.0159757f $X=1.435 $Y=0.71 $X2=0 $Y2=0
cc_405 N_X_c_652_n N_VGND_c_716_n 0.00244309f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_406 N_X_c_692_p N_VGND_c_716_n 0.0112274f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_407 N_X_c_657_n N_VGND_c_716_n 0.00257772f $X=1.435 $Y=0.71 $X2=0 $Y2=0
cc_408 N_X_c_657_n N_VGND_c_717_n 0.00257772f $X=1.435 $Y=0.71 $X2=0 $Y2=0
cc_409 N_X_c_695_p N_VGND_c_717_n 0.0112274f $X=1.52 $Y=0.42 $X2=0 $Y2=0
cc_410 N_X_M1010_s N_VGND_c_721_n 0.00247944f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_411 N_X_M1016_s N_VGND_c_721_n 0.0040445f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_412 N_X_c_652_n N_VGND_c_721_n 0.00445306f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_413 N_X_c_692_p N_VGND_c_721_n 0.00643448f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_414 N_X_c_657_n N_VGND_c_721_n 0.0101011f $X=1.435 $Y=0.71 $X2=0 $Y2=0
cc_415 N_X_c_695_p N_VGND_c_721_n 0.00643448f $X=1.52 $Y=0.42 $X2=0 $Y2=0
cc_416 N_X_c_645_n N_VGND_c_721_n 0.00170408f $X=0.225 $Y=0.805 $X2=0 $Y2=0
cc_417 N_VGND_c_721_n N_A_474_47#_M1000_s 0.00213443f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_418 N_VGND_c_721_n N_A_474_47#_M1022_s 0.0025535f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_c_721_n N_A_474_47#_M1001_d 0.00223231f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_721_n N_A_474_47#_M1015_s 0.00213418f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_713_n N_A_474_47#_c_812_n 0.0171306f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_422 N_VGND_c_718_n N_A_474_47#_c_812_n 0.105565f $X=4.67 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_721_n N_A_474_47#_c_812_n 0.0660081f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_718_n N_A_474_47#_c_830_n 0.0190605f $X=4.67 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_721_n N_A_474_47#_c_830_n 0.0125165f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_M1014_d N_A_474_47#_c_832_n 0.00699963f $X=4.64 $Y=0.235 $X2=0
+ $Y2=0
cc_427 N_VGND_c_714_n N_A_474_47#_c_832_n 0.0214325f $X=4.82 $Y=0.36 $X2=0 $Y2=0
cc_428 N_VGND_c_718_n N_A_474_47#_c_832_n 0.00223745f $X=4.67 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_719_n N_A_474_47#_c_832_n 0.0021487f $X=5.655 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_721_n N_A_474_47#_c_832_n 0.0090689f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_719_n N_A_474_47#_c_838_n 0.0188082f $X=5.655 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_721_n N_A_474_47#_c_838_n 0.0122321f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_M1002_s N_A_474_47#_c_813_n 0.0047036f $X=5.61 $Y=0.235 $X2=0
+ $Y2=0
cc_434 N_VGND_c_715_n N_A_474_47#_c_813_n 0.0128906f $X=5.75 $Y=0.36 $X2=0 $Y2=0
cc_435 N_VGND_c_719_n N_A_474_47#_c_813_n 0.0021487f $X=5.655 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_720_n N_A_474_47#_c_813_n 0.0021487f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_721_n N_A_474_47#_c_813_n 0.00860478f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_720_n N_A_474_47#_c_814_n 0.0208978f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_721_n N_A_474_47#_c_814_n 0.0124141f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_721_n A_748_47# 0.00168648f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_441 N_VGND_c_721_n A_557_47# 0.00224864f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_442 N_A_474_47#_c_812_n A_748_47# 0.00193721f $X=4.17 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_443 N_A_474_47#_c_812_n A_557_47# 0.00775585f $X=4.17 $Y=0.36 $X2=-0.19
+ $Y2=-0.24

* File: sky130_fd_sc_hd__a21bo_1.spice
* Created: Thu Aug 27 14:00:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21bo_1.pex.spice"
.subckt sky130_fd_sc_hd__a21bo_1  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B1_N_M1005_g N_A_27_413#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.106688 AS=0.1113 PD=0.863551 PS=1.37 NRD=22.14 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_215_297#_M1009_d N_A_27_413#_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.165112 PD=0.92 PS=1.33645 NRD=0 NRS=17.532 M=1
+ R=4.33333 SA=75000.6 SB=75002 A=0.0975 P=1.6 MULT=1
MM1008 A_382_47# N_A1_M1008_g N_A_215_297#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.08775 PD=0.93 PS=0.92 NRD=15.684 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_382_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.258375 AS=0.091 PD=1.445 PS=0.93 NRD=14.76 NRS=15.684 M=1 R=4.33333
+ SA=75001.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_215_297#_M1007_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.258375 PD=1.82 PS=1.445 NRD=0 NRS=15.684 M=1 R=4.33333
+ SA=75002.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_B1_N_M1002_g N_A_27_413#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_298_297#_M1000_d N_A_27_413#_M1000_g N_A_215_297#_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.265 PD=1.27 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_298_297#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_298_297#_M1003_d N_A2_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_215_297#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_65 VPB 0 1.83237e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a21bo_1.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__or2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__or2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.765000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.500000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.180000 0.825000 ;
        RECT 1.645000 1.845000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.300000 0.085000 ;
        RECT 0.250000  0.085000 0.490000 0.595000 ;
        RECT 1.180000  0.085000 1.395000 0.595000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.300000 2.805000 ;
        RECT 1.145000 1.835000 1.475000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.270000 1.495000 1.695000 1.665000 ;
      RECT 0.270000 1.665000 0.660000 1.840000 ;
      RECT 0.670000 0.265000 0.950000 0.595000 ;
      RECT 0.670000 0.595000 0.840000 1.495000 ;
      RECT 1.525000 0.995000 1.695000 1.495000 ;
  END
END sky130_fd_sc_hd__or2_1

* File: sky130_fd_sc_hd__sdfxbp_2.pex.spice
* Created: Tue Sep  1 19:31:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%CLK 1 2 3 5 6 8 11 13
c42 1 0 2.71124e-20 $X=0.31 $Y=1.325
r43 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.475 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=2.135
r47 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r50 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_27_47# 1 2 9 13 17 19 20 25 29 31 35 39
+ 43 44 45 49 50 52 55 56 57 58 59 60 69 75 78 79 80 82 86
c247 86 0 1.77381e-19 $X=6.69 $Y=1.41
c248 52 0 8.70797e-20 $X=0.76 $Y=1.235
c249 50 0 1.81794e-19 $X=0.73 $Y=1.795
c250 45 0 3.29888e-20 $X=0.615 $Y=1.88
c251 29 0 4.21632e-20 $X=6.695 $Y=2.275
c252 19 0 1.57835e-19 $X=5.005 $Y=1.32
r253 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.41
+ $X2=6.69 $Y2=1.575
r254 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.69
+ $Y=1.41 $X2=6.69 $Y2=1.41
r255 82 85 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.69 $Y=1.32 $X2=6.69
+ $Y2=1.41
r256 78 81 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.74
+ $X2=5.14 $Y2=1.905
r257 78 80 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.74
+ $X2=5.14 $Y2=1.575
r258 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.74 $X2=5.14 $Y2=1.74
r259 74 75 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=0.89 $Y=1.235
+ $X2=0.895 $Y2=1.235
r260 70 86 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.7 $Y=1.87 $X2=6.7
+ $Y2=1.41
r261 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=1.87
+ $X2=6.71 $Y2=1.87
r262 66 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r263 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.87
r264 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r265 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.565 $Y=1.87
+ $X2=6.71 $Y2=1.87
r266 59 60 1.39851 $w=1.4e-07 $l=1.13e-06 $layer=MET1_cond $X=6.565 $Y=1.87
+ $X2=5.435 $Y2=1.87
r267 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=1.87
+ $X2=0.73 $Y2=1.87
r268 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r269 57 58 5.28464 $w=1.4e-07 $l=4.27e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=0.875 $Y2=1.87
r270 53 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r271 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r272 50 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r273 50 52 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r274 49 56 6.0623 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=0.97
r275 49 52 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=1.235
r276 47 56 9.38461 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=0.805
+ $X2=0.712 $Y2=0.97
r277 46 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r278 45 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r279 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.35 $Y2=1.88
r280 43 47 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.712 $Y2=0.805
r281 43 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r282 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r283 37 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r284 33 35 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.34 $Y=1.245
+ $X2=7.34 $Y2=0.415
r285 32 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.825 $Y=1.32
+ $X2=6.69 $Y2=1.32
r286 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.265 $Y=1.32
+ $X2=7.34 $Y2=1.245
r287 31 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.265 $Y=1.32
+ $X2=6.825 $Y2=1.32
r288 29 87 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.695 $Y=2.275
+ $X2=6.695 $Y2=1.575
r289 25 81 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.08 $Y=2.275
+ $X2=5.08 $Y2=1.905
r290 21 80 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.08 $Y=1.395
+ $X2=5.08 $Y2=1.575
r291 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.005 $Y=1.32
+ $X2=5.08 $Y2=1.395
r292 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=5.005 $Y=1.32
+ $X2=4.695 $Y2=1.32
r293 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.62 $Y=1.245
+ $X2=4.695 $Y2=1.32
r294 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.62 $Y=1.245
+ $X2=4.62 $Y2=0.415
r295 11 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=1.235
r296 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=2.135
r297 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r298 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r299 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r300 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%SCE 3 7 11 15 19 20 22 23 24 28 29 32 33
c110 24 0 1.66251e-19 $X=3.085 $Y=0.7
c111 22 0 1.76484e-19 $X=2.475 $Y=0.7
r112 35 36 3.41038 $w=2.12e-07 $l=1.5e-08 $layer=POLY_cond $X=1.835 $Y=1.52
+ $X2=1.85 $Y2=1.52
r113 31 33 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.51
r114 31 32 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.7
r115 29 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=0.95
+ $X2=3.17 $Y2=0.785
r116 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=0.95 $X2=3.17 $Y2=0.95
r117 26 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0.785
+ $X2=3.17 $Y2=0.95
r118 25 32 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.65 $Y=0.7
+ $X2=2.562 $Y2=0.7
r119 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=0.7
+ $X2=3.17 $Y2=0.785
r120 24 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.085 $Y=0.7
+ $X2=2.65 $Y2=0.7
r121 22 32 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=2.562 $Y2=0.7
r122 22 23 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=1.95 $Y2=0.7
r123 20 38 88.6698 $w=2.12e-07 $l=3.9e-07 $layer=POLY_cond $X=1.865 $Y=1.52
+ $X2=2.255 $Y2=1.52
r124 20 36 3.41038 $w=2.12e-07 $l=1.5e-08 $layer=POLY_cond $X=1.865 $Y=1.52
+ $X2=1.85 $Y2=1.52
r125 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=1.52 $X2=1.865 $Y2=1.52
r126 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=0.785
+ $X2=1.95 $Y2=0.7
r127 17 19 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.865 $Y=0.785
+ $X2=1.865 $Y2=1.52
r128 15 40 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.23 $Y=0.445
+ $X2=3.23 $Y2=0.785
r129 9 38 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.255 $Y=1.655
+ $X2=2.255 $Y2=1.52
r130 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.255 $Y=1.655
+ $X2=2.255 $Y2=2.165
r131 5 36 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.85 $Y=1.385
+ $X2=1.85 $Y2=1.52
r132 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.85 $Y=1.385 $X2=1.85
+ $Y2=0.445
r133 1 35 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.835 $Y=1.655
+ $X2=1.835 $Y2=1.52
r134 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.835 $Y=1.655
+ $X2=1.835 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_299_47# 1 2 9 13 16 19 21 24 25 28 32 34
+ 38 39 41 43 44
c126 43 0 1.84493e-19 $X=3.19 $Y=1.52
c127 39 0 1.12087e-19 $X=2.3 $Y=1.04
c128 24 0 1.60762e-19 $X=2.205 $Y=1.86
c129 9 0 1.20015e-19 $X=2.36 $Y=0.445
r130 44 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.52
+ $X2=3.19 $Y2=1.685
r131 43 46 9.59627 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.177 $Y=1.52
+ $X2=3.177 $Y2=1.685
r132 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.52 $X2=3.19 $Y2=1.52
r133 39 48 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.3 $Y=1.04
+ $X2=2.3 $Y2=0.905
r134 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.04 $X2=2.3 $Y2=1.04
r135 35 38 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.205 $Y=1.04
+ $X2=2.3 $Y2=1.04
r136 29 32 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.52 $Y=0.36
+ $X2=1.64 $Y2=0.36
r137 28 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.165 $Y=1.86
+ $X2=3.165 $Y2=1.685
r138 26 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=1.967
+ $X2=2.205 $Y2=1.967
r139 25 28 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.08 $Y=1.967
+ $X2=3.165 $Y2=1.86
r140 25 26 42.3456 $w=2.13e-07 $l=7.9e-07 $layer=LI1_cond $X=3.08 $Y=1.967
+ $X2=2.29 $Y2=1.967
r141 24 41 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.205 $Y=1.86
+ $X2=2.205 $Y2=1.967
r142 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=1.125
+ $X2=2.205 $Y2=1.04
r143 23 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.205 $Y=1.125
+ $X2=2.205 $Y2=1.86
r144 22 34 1.46632 $w=2.15e-07 $l=1.38e-07 $layer=LI1_cond $X=1.71 $Y=1.967
+ $X2=1.572 $Y2=1.967
r145 21 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=1.967
+ $X2=2.205 $Y2=1.967
r146 21 22 21.9768 $w=2.13e-07 $l=4.1e-07 $layer=LI1_cond $X=2.12 $Y=1.967
+ $X2=1.71 $Y2=1.967
r147 17 34 5.02022 $w=2.22e-07 $l=1.08e-07 $layer=LI1_cond $X=1.572 $Y=2.075
+ $X2=1.572 $Y2=1.967
r148 17 19 4.1907 $w=2.73e-07 $l=1e-07 $layer=LI1_cond $X=1.572 $Y=2.075
+ $X2=1.572 $Y2=2.175
r149 16 34 5.02022 $w=2.22e-07 $l=1.30434e-07 $layer=LI1_cond $X=1.52 $Y=1.86
+ $X2=1.572 $Y2=1.967
r150 15 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.445
+ $X2=1.52 $Y2=0.36
r151 15 16 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.52 $Y=0.445
+ $X2=1.52 $Y2=1.86
r152 13 52 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.145 $Y=2.165
+ $X2=3.145 $Y2=1.685
r153 9 48 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.36 $Y=0.445
+ $X2=2.36 $Y2=0.905
r154 2 19 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.845 $X2=1.625 $Y2=2.175
r155 1 32 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.64 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%D 3 7 9 12 13
c49 13 0 2.8857e-19 $X=2.71 $Y=1.52
r50 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.52
+ $X2=2.71 $Y2=1.685
r51 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.52
+ $X2=2.71 $Y2=1.355
r52 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.52 $X2=2.71 $Y2=1.52
r53 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.56 $Y=1.52 $X2=2.71
+ $Y2=1.52
r54 7 14 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.75 $Y=0.445
+ $X2=2.75 $Y2=1.355
r55 3 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.725 $Y=2.165
+ $X2=2.725 $Y2=1.685
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%SCD 3 7 9 12
c48 7 0 1.84493e-19 $X=3.61 $Y=2.165
c49 3 0 1.66251e-19 $X=3.61 $Y=0.445
r50 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.355
+ $X2=3.67 $Y2=1.52
r51 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.355
+ $X2=3.67 $Y2=1.19
r52 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.67
+ $Y=1.355 $X2=3.67 $Y2=1.355
r53 9 13 5.20873 $w=6.18e-07 $l=2.7e-07 $layer=LI1_cond $X=3.94 $Y=1.345
+ $X2=3.67 $Y2=1.345
r54 7 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.61 $Y=2.165
+ $X2=3.61 $Y2=1.52
r55 3 14 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.61 $Y=0.445
+ $X2=3.61 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_193_47# 1 2 9 13 14 16 19 23 24 27 30 33
+ 37 38 40 41 42 43 46 52 59 60 61 66
c215 66 0 1.77381e-19 $X=6.92 $Y=0.87
c216 42 0 1.57835e-19 $X=6.58 $Y=0.85
r217 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.92
+ $Y=0.87 $X2=6.92 $Y2=0.87
r218 63 66 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.825 $Y=0.87
+ $X2=6.92 $Y2=0.87
r219 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.04 $Y=0.87
+ $X2=5.04 $Y2=0.705
r220 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=0.87 $X2=5.04 $Y2=0.87
r221 53 67 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.725 $Y=0.87
+ $X2=6.92 $Y2=0.87
r222 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.725 $Y=0.85
+ $X2=6.725 $Y2=0.85
r223 50 60 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=0.87
+ $X2=5.04 $Y2=0.87
r224 50 80 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0.87
+ $X2=4.665 $Y2=0.87
r225 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0.85
+ $X2=4.83 $Y2=0.85
r226 46 75 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.132 $Y=0.85
+ $X2=1.132 $Y2=1.96
r227 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.135 $Y=0.85
+ $X2=1.135 $Y2=0.85
r228 43 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=0.85
+ $X2=4.83 $Y2=0.85
r229 42 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.58 $Y=0.85
+ $X2=6.725 $Y2=0.85
r230 42 43 1.98638 $w=1.4e-07 $l=1.605e-06 $layer=MET1_cond $X=6.58 $Y=0.85
+ $X2=4.975 $Y2=0.85
r231 41 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.28 $Y=0.85
+ $X2=1.135 $Y2=0.85
r232 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=4.83 $Y2=0.85
r233 40 41 4.2141 $w=1.4e-07 $l=3.405e-06 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=1.28 $Y2=0.85
r234 38 69 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=7.2 $Y=1.74
+ $X2=7.115 $Y2=1.74
r235 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.2
+ $Y=1.74 $X2=7.2 $Y2=1.74
r236 34 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.06 $Y=1.74
+ $X2=7.2 $Y2=1.74
r237 33 67 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.965 $Y=0.87
+ $X2=6.92 $Y2=0.87
r238 32 46 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=1.132 $Y=0.715
+ $X2=1.132 $Y2=0.85
r239 30 32 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.13 $Y=0.51
+ $X2=1.13 $Y2=0.715
r240 27 34 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.06 $Y=1.575
+ $X2=7.06 $Y2=1.74
r241 26 33 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.06 $Y=1.035
+ $X2=6.965 $Y2=0.87
r242 26 27 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.06 $Y=1.035
+ $X2=7.06 $Y2=1.575
r243 24 57 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.63 $Y=1.74
+ $X2=4.63 $Y2=1.875
r244 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.63
+ $Y=1.74 $X2=4.63 $Y2=1.74
r245 21 80 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=1.035
+ $X2=4.665 $Y2=0.87
r246 21 23 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.665 $Y=1.035
+ $X2=4.665 $Y2=1.74
r247 17 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.115 $Y=1.875
+ $X2=7.115 $Y2=1.74
r248 17 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.115 $Y=1.875
+ $X2=7.115 $Y2=2.275
r249 14 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.705
+ $X2=6.825 $Y2=0.87
r250 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.825 $Y=0.705
+ $X2=6.825 $Y2=0.415
r251 13 61 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.1 $Y=0.415
+ $X2=5.1 $Y2=0.705
r252 9 57 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.615 $Y=2.275
+ $X2=4.615 $Y2=1.875
r253 2 75 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.815 $X2=1.105 $Y2=1.96
r254 1 30 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_1097_183# 1 2 9 13 15 18 21 23 29 30 32
+ 33 36
r95 35 36 5.54023 $w=2.61e-07 $l=3e-08 $layer=POLY_cond $X=5.56 $Y=0.93 $X2=5.59
+ $Y2=0.93
r96 32 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.39 $Y=2.3
+ $X2=6.39 $Y2=2.135
r97 27 36 24.0077 $w=2.61e-07 $l=1.3e-07 $layer=POLY_cond $X=5.72 $Y=0.93
+ $X2=5.59 $Y2=0.93
r98 26 29 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=0.93
+ $X2=5.805 $Y2=0.93
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.72
+ $Y=0.93 $X2=5.72 $Y2=0.93
r100 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.435 $Y=0.45
+ $X2=6.56 $Y2=0.45
r101 19 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.35 $Y=1.065
+ $X2=6.35 $Y2=0.915
r102 19 33 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.35 $Y=1.065
+ $X2=6.35 $Y2=2.135
r103 18 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.35 $Y=0.765
+ $X2=6.35 $Y2=0.915
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.35 $Y=0.535
+ $X2=6.435 $Y2=0.45
r105 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.35 $Y=0.535
+ $X2=6.35 $Y2=0.765
r106 15 30 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.265 $Y=0.915
+ $X2=6.35 $Y2=0.915
r107 15 29 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.265 $Y=0.915
+ $X2=5.805 $Y2=0.915
r108 11 36 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.59 $Y=0.795
+ $X2=5.59 $Y2=0.93
r109 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.59 $Y=0.795
+ $X2=5.59 $Y2=0.445
r110 7 35 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.56 $Y=1.065
+ $X2=5.56 $Y2=0.93
r111 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.56 $Y=1.065
+ $X2=5.56 $Y2=2.275
r112 2 32 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.735 $X2=6.43 $Y2=2.3
r113 1 23 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.395
+ $Y=0.235 $X2=6.56 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_938_413# 1 2 8 11 13 15 18 20 21 22 26 31
+ 33 35
c108 31 0 1.42307e-19 $X=5.38 $Y=1.315
r109 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.01
+ $Y=1.41 $X2=6.01 $Y2=1.41
r110 35 37 17.1405 $w=2.42e-07 $l=3.4e-07 $layer=LI1_cond $X=5.67 $Y=1.41
+ $X2=6.01 $Y2=1.41
r111 32 35 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=1.575
+ $X2=5.67 $Y2=1.41
r112 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.67 $Y=1.575
+ $X2=5.67 $Y2=2.19
r113 31 35 14.6198 $w=2.42e-07 $l=2.9e-07 $layer=LI1_cond $X=5.38 $Y=1.41
+ $X2=5.67 $Y2=1.41
r114 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.38 $Y=0.535
+ $X2=5.38 $Y2=1.315
r115 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.295 $Y=0.45
+ $X2=5.38 $Y2=0.535
r116 26 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.295 $Y=0.45
+ $X2=4.89 $Y2=0.45
r117 22 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.585 $Y=2.275
+ $X2=5.67 $Y2=2.19
r118 22 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.585 $Y=2.275
+ $X2=4.85 $Y2=2.275
r119 20 38 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.145 $Y=1.41
+ $X2=6.01 $Y2=1.41
r120 20 21 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.145 $Y=1.41
+ $X2=6.22 $Y2=1.41
r121 16 18 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.22 $Y=1.025
+ $X2=6.32 $Y2=1.025
r122 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.32 $Y=0.95
+ $X2=6.32 $Y2=1.025
r123 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.32 $Y=0.95
+ $X2=6.32 $Y2=0.555
r124 9 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.22 $Y=1.545
+ $X2=6.22 $Y2=1.41
r125 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.22 $Y=1.545
+ $X2=6.22 $Y2=2.11
r126 8 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.22 $Y=1.275
+ $X2=6.22 $Y2=1.41
r127 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.22 $Y=1.1 $X2=6.22
+ $Y2=1.025
r128 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.22 $Y=1.1 $X2=6.22
+ $Y2=1.275
r129 2 24 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=2.065 $X2=4.85 $Y2=2.275
r130 1 28 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.235 $X2=4.89 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_1525_315# 1 2 9 13 15 17 20 22 24 27 29
+ 30 31 33 35 38 41 42 43 46 50 53 55 58 62 66 67
c136 41 0 1.53472e-19 $X=10.552 $Y=1.515
c137 31 0 1.26281e-19 $X=10.525 $Y=1.325
c138 30 0 1.02967e-19 $X=9.705 $Y=1.16
r139 75 76 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=9.21 $Y=1.16
+ $X2=9.63 $Y2=1.16
r140 68 70 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.7 $Y=1.74
+ $X2=7.815 $Y2=1.74
r141 62 64 16.6896 $w=3.63e-07 $l=4.4e-07 $layer=LI1_cond $X=8.542 $Y=0.385
+ $X2=8.542 $Y2=0.825
r142 59 75 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=9.19 $Y=1.16 $X2=9.21
+ $Y2=1.16
r143 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.19
+ $Y=1.16 $X2=9.19 $Y2=1.16
r144 56 67 0.63164 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=8.725 $Y=1.16
+ $X2=8.632 $Y2=1.16
r145 56 58 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.725 $Y=1.16
+ $X2=9.19 $Y2=1.16
r146 55 66 6.31733 $w=2.57e-07 $l=1.9775e-07 $layer=LI1_cond $X=8.632 $Y=1.575
+ $X2=8.56 $Y2=1.74
r147 54 67 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=8.632 $Y=1.325
+ $X2=8.632 $Y2=1.16
r148 54 55 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=8.632 $Y=1.325
+ $X2=8.632 $Y2=1.575
r149 53 67 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=8.632 $Y=0.995
+ $X2=8.632 $Y2=1.16
r150 53 64 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=8.632 $Y=0.995
+ $X2=8.632 $Y2=0.825
r151 48 66 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=8.56 $Y=1.905
+ $X2=8.56 $Y2=1.74
r152 48 50 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=8.56 $Y=1.905
+ $X2=8.56 $Y2=2.34
r153 46 70 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.88 $Y=1.74
+ $X2=7.815 $Y2=1.74
r154 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.88
+ $Y=1.74 $X2=7.88 $Y2=1.74
r155 43 66 0.466467 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.395 $Y=1.74
+ $X2=8.56 $Y2=1.74
r156 43 45 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=8.395 $Y=1.74
+ $X2=7.88 $Y2=1.74
r157 41 42 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=10.552 $Y=1.515
+ $X2=10.552 $Y2=1.665
r158 38 42 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=10.58 $Y=2.165
+ $X2=10.58 $Y2=1.665
r159 33 35 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.58 $Y=0.73
+ $X2=10.58 $Y2=0.445
r160 31 41 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.525 $Y=1.325
+ $X2=10.525 $Y2=1.515
r161 30 76 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.705 $Y=1.16
+ $X2=9.63 $Y2=1.16
r162 29 31 49.1818 $w=1.63e-07 $l=1.77989e-07 $layer=POLY_cond $X=10.552 $Y=1.16
+ $X2=10.525 $Y2=1.325
r163 29 33 127.544 $w=1.63e-07 $l=4.43779e-07 $layer=POLY_cond $X=10.552 $Y=1.16
+ $X2=10.58 $Y2=0.73
r164 29 30 130.272 $w=3.3e-07 $l=7.45e-07 $layer=POLY_cond $X=10.45 $Y=1.16
+ $X2=9.705 $Y2=1.16
r165 25 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=1.325
+ $X2=9.63 $Y2=1.16
r166 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.63 $Y=1.325
+ $X2=9.63 $Y2=1.985
r167 22 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=0.995
+ $X2=9.63 $Y2=1.16
r168 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.63 $Y=0.995
+ $X2=9.63 $Y2=0.56
r169 18 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=1.325
+ $X2=9.21 $Y2=1.16
r170 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.21 $Y=1.325
+ $X2=9.21 $Y2=1.985
r171 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=0.995
+ $X2=9.21 $Y2=1.16
r172 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.21 $Y=0.995
+ $X2=9.21 $Y2=0.56
r173 11 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=1.575
+ $X2=7.815 $Y2=1.74
r174 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.815 $Y=1.575
+ $X2=7.815 $Y2=0.445
r175 7 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.7 $Y=1.905
+ $X2=7.7 $Y2=1.74
r176 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.7 $Y=1.905 $X2=7.7
+ $Y2=2.275
r177 2 66 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.435
+ $Y=1.485 $X2=8.56 $Y2=1.66
r178 2 50 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=8.435
+ $Y=1.485 $X2=8.56 $Y2=2.34
r179 1 62 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=8.435
+ $Y=0.235 $X2=8.56 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_1354_413# 1 2 7 9 12 14 15 16 20 27 30 33
+ 34
c87 30 0 1.02967e-19 $X=8.285 $Y=1.16
c88 27 0 4.21632e-20 $X=7.54 $Y=2.165
c89 15 0 1.26247e-19 $X=8.77 $Y=1.16
c90 12 0 1.04554e-19 $X=8.77 $Y=1.985
c91 7 0 1.04554e-19 $X=8.77 $Y=0.995
r92 33 35 11.5578 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=7.475 $Y=1.16
+ $X2=7.475 $Y2=1.405
r93 33 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=1.16
+ $X2=7.475 $Y2=0.995
r94 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.285
+ $Y=1.16 $X2=8.285 $Y2=1.16
r95 28 33 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.625 $Y=1.16
+ $X2=7.475 $Y2=1.16
r96 28 30 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=7.625 $Y=1.16
+ $X2=8.285 $Y2=1.16
r97 27 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.54 $Y=2.165
+ $X2=7.54 $Y2=1.405
r98 24 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.41 $Y=0.535
+ $X2=7.41 $Y2=0.995
r99 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.325 $Y=0.45
+ $X2=7.41 $Y2=0.535
r100 20 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.325 $Y=0.45
+ $X2=7.12 $Y2=0.45
r101 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.455 $Y=2.25
+ $X2=7.54 $Y2=2.165
r102 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.455 $Y=2.25
+ $X2=6.905 $Y2=2.25
r103 14 31 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=8.695 $Y=1.16
+ $X2=8.285 $Y2=1.16
r104 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.695 $Y=1.16
+ $X2=8.77 $Y2=1.16
r105 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.77 $Y=1.325
+ $X2=8.77 $Y2=1.16
r106 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.77 $Y=1.325
+ $X2=8.77 $Y2=1.985
r107 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.77 $Y=0.995
+ $X2=8.77 $Y2=1.16
r108 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.77 $Y=0.995
+ $X2=8.77 $Y2=0.56
r109 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=2.065 $X2=6.905 $Y2=2.25
r110 1 22 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.235 $X2=7.12 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_2049_47# 1 2 7 9 12 14 16 19 23 27 31 34
+ 38
c69 38 0 3.00828e-19 $X=11.485 $Y=1.16
r70 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.065 $Y=1.16
+ $X2=11.485 $Y2=1.16
r71 32 37 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=10.98 $Y=1.16
+ $X2=11.065 $Y2=1.16
r72 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.98
+ $Y=1.16 $X2=10.98 $Y2=1.16
r73 29 34 0.881669 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.535 $Y=1.16
+ $X2=10.37 $Y2=1.16
r74 29 31 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=10.535 $Y=1.16
+ $X2=10.98 $Y2=1.16
r75 25 34 5.74456 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=10.37 $Y=1.325
+ $X2=10.37 $Y2=1.16
r76 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.37 $Y=1.325
+ $X2=10.37 $Y2=2
r77 21 34 5.74456 $w=2.9e-07 $l=1.83916e-07 $layer=LI1_cond $X=10.33 $Y=0.995
+ $X2=10.37 $Y2=1.16
r78 21 23 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=10.33 $Y=0.995
+ $X2=10.33 $Y2=0.51
r79 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.485 $Y=1.325
+ $X2=11.485 $Y2=1.16
r80 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.485 $Y=1.325
+ $X2=11.485 $Y2=1.985
r81 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.485 $Y=0.995
+ $X2=11.485 $Y2=1.16
r82 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.485 $Y=0.995
+ $X2=11.485 $Y2=0.56
r83 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.065 $Y=1.325
+ $X2=11.065 $Y2=1.16
r84 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.065 $Y=1.325
+ $X2=11.065 $Y2=1.985
r85 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.065 $Y=0.995
+ $X2=11.065 $Y2=1.16
r86 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.065 $Y=0.995
+ $X2=11.065 $Y2=0.56
r87 2 27 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=10.245
+ $Y=1.845 $X2=10.37 $Y2=2
r88 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=10.245
+ $Y=0.235 $X2=10.37 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 48 52
+ 56 60 64 66 71 72 74 75 76 78 83 88 100 111 115 121 124 127 130 133 136 140
c191 140 0 1.81794e-19 $X=11.73 $Y=2.72
c192 60 0 1.53472e-19 $X=10.855 $Y=1.66
c193 2 0 1.60762e-19 $X=1.91 $Y=1.845
c194 1 0 3.29888e-20 $X=0.55 $Y=1.815
r195 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r196 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r197 133 134 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r198 131 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r199 130 131 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r200 127 128 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r201 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r202 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r203 119 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r204 119 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=10.81 $Y2=2.72
r205 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r206 116 136 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=11.02 $Y=2.72
+ $X2=10.867 $Y2=2.72
r207 116 118 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=11.02 $Y=2.72
+ $X2=11.27 $Y2=2.72
r208 115 139 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=11.61 $Y=2.72
+ $X2=11.785 $Y2=2.72
r209 115 118 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.61 $Y=2.72
+ $X2=11.27 $Y2=2.72
r210 114 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r211 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r212 111 136 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=10.715 $Y=2.72
+ $X2=10.867 $Y2=2.72
r213 111 113 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=10.715 $Y=2.72
+ $X2=10.35 $Y2=2.72
r214 110 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r215 110 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r216 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r217 107 133 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.075 $Y=2.72
+ $X2=8.985 $Y2=2.72
r218 107 109 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.075 $Y=2.72
+ $X2=9.43 $Y2=2.72
r219 106 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r220 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r221 103 106 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r222 102 105 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r223 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r224 100 130 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.805 $Y=2.72
+ $X2=7.957 $Y2=2.72
r225 100 105 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.805 $Y=2.72
+ $X2=7.59 $Y2=2.72
r226 99 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r227 99 128 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r228 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r229 96 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=2.72
+ $X2=3.845 $Y2=2.72
r230 96 98 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=3.93 $Y=2.72
+ $X2=5.75 $Y2=2.72
r231 95 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r232 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r233 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r234 92 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r235 91 94 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r236 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r237 89 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.045 $Y2=2.72
r238 89 91 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.53 $Y2=2.72
r239 88 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=2.72
+ $X2=3.845 $Y2=2.72
r240 88 94 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=2.72
+ $X2=3.45 $Y2=2.72
r241 87 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r242 87 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r243 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r244 84 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=0.685 $Y2=2.72
r245 84 86 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r246 83 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=2.045 $Y2=2.72
r247 83 86 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=1.61 $Y2=2.72
r248 78 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.685 $Y2=2.72
r249 78 80 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r250 76 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r251 76 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r252 74 109 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.765 $Y=2.72
+ $X2=9.43 $Y2=2.72
r253 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.765 $Y=2.72
+ $X2=9.85 $Y2=2.72
r254 73 113 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.935 $Y=2.72
+ $X2=10.35 $Y2=2.72
r255 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.935 $Y=2.72
+ $X2=9.85 $Y2=2.72
r256 71 98 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r257 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=2.72
+ $X2=6.01 $Y2=2.72
r258 70 102 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.21 $Y2=2.72
r259 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.01 $Y2=2.72
r260 66 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.695 $Y=1.66
+ $X2=11.695 $Y2=2.34
r261 64 139 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=11.695 $Y=2.635
+ $X2=11.785 $Y2=2.72
r262 64 69 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.695 $Y=2.635
+ $X2=11.695 $Y2=2.34
r263 60 63 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=10.867 $Y=1.66
+ $X2=10.867 $Y2=2
r264 58 136 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=10.867 $Y=2.635
+ $X2=10.867 $Y2=2.72
r265 58 63 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=10.867 $Y=2.635
+ $X2=10.867 $Y2=2
r266 54 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.85 $Y=2.635
+ $X2=9.85 $Y2=2.72
r267 54 56 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=9.85 $Y=2.635
+ $X2=9.85 $Y2=1.78
r268 50 133 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.985 $Y=2.635
+ $X2=8.985 $Y2=2.72
r269 50 52 52.0657 $w=1.78e-07 $l=8.45e-07 $layer=LI1_cond $X=8.985 $Y=2.635
+ $X2=8.985 $Y2=1.79
r270 49 130 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.11 $Y=2.72
+ $X2=7.957 $Y2=2.72
r271 48 133 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.895 $Y=2.72
+ $X2=8.985 $Y2=2.72
r272 48 49 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.895 $Y=2.72
+ $X2=8.11 $Y2=2.72
r273 44 130 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.957 $Y=2.635
+ $X2=7.957 $Y2=2.72
r274 44 46 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=7.957 $Y=2.635
+ $X2=7.957 $Y2=2.3
r275 40 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=2.635
+ $X2=6.01 $Y2=2.72
r276 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.01 $Y=2.635
+ $X2=6.01 $Y2=2
r277 36 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.72
r278 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.33
r279 32 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.72
r280 32 34 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.33
r281 28 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.72
r282 28 30 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.22
r283 9 69 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=11.56
+ $Y=1.485 $X2=11.695 $Y2=2.34
r284 9 66 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=11.56
+ $Y=1.485 $X2=11.695 $Y2=1.66
r285 8 63 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=10.655
+ $Y=1.845 $X2=10.855 $Y2=2
r286 8 60 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=1.845 $X2=10.855 $Y2=1.66
r287 7 56 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=9.705
+ $Y=1.485 $X2=9.85 $Y2=1.78
r288 6 52 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=8.845
+ $Y=1.485 $X2=8.99 $Y2=1.79
r289 5 46 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=2.065 $X2=8.02 $Y2=2.3
r290 4 42 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=5.635
+ $Y=2.065 $X2=6.01 $Y2=2
r291 3 38 600 $w=1.7e-07 $l=5.59308e-07 $layer=licon1_PDIFF $count=1 $X=3.685
+ $Y=1.845 $X2=3.845 $Y2=2.33
r292 2 34 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.845 $X2=2.045 $Y2=2.33
r293 1 30 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.815 $X2=0.685 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%A_560_369# 1 2 3 4 13 17 22 24 25 26 27 28
+ 30 32 36 38 39
c111 17 0 1.20015e-19 $X=3.425 $Y=0.36
r112 39 41 18.789 $w=2.37e-07 $l=3.65e-07 $layer=LI1_cond $X=4.345 $Y=1.91
+ $X2=4.345 $Y2=2.275
r113 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.29 $Y=0.45 $X2=4.39
+ $Y2=0.45
r114 32 39 5.36951 $w=2.37e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.29 $Y=1.825
+ $X2=4.345 $Y2=1.91
r115 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0.865
+ $X2=4.29 $Y2=0.78
r116 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.29 $Y=0.865
+ $X2=4.29 $Y2=1.825
r117 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0.695
+ $X2=4.29 $Y2=0.78
r118 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0.535
+ $X2=4.29 $Y2=0.45
r119 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.29 $Y=0.535
+ $X2=4.29 $Y2=0.695
r120 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=0.78
+ $X2=4.29 $Y2=0.78
r121 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.205 $Y=0.78
+ $X2=3.595 $Y2=0.78
r122 25 39 2.684 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.205 $Y=1.91
+ $X2=4.345 $Y2=1.91
r123 25 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.205 $Y=1.91
+ $X2=3.59 $Y2=1.91
r124 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.51 $Y=0.695
+ $X2=3.595 $Y2=0.78
r125 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.51 $Y=0.445
+ $X2=3.51 $Y2=0.695
r126 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=1.995
+ $X2=3.59 $Y2=1.91
r127 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.505 $Y=1.995
+ $X2=3.505 $Y2=2.245
r128 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=0.36
+ $X2=3.51 $Y2=0.445
r129 17 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.425 $Y=0.36
+ $X2=3.015 $Y2=0.36
r130 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=2.33
+ $X2=3.505 $Y2=2.245
r131 13 15 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.42 $Y=2.33
+ $X2=2.935 $Y2=2.33
r132 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=2.065 $X2=4.4 $Y2=2.275
r133 3 15 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.845 $X2=2.935 $Y2=2.33
r134 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.235 $X2=4.39 $Y2=0.45
r135 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=3.015 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%Q 1 2 9 14 15 16 19
c39 15 0 1.04554e-19 $X=9.42 $Y=0.79
c40 14 0 2.30802e-19 $X=9.53 $Y=1.43
r41 16 19 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=9.42 $Y=0.51
+ $X2=9.42 $Y2=0.36
r42 15 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=9.42 $Y=0.79 $X2=9.42
+ $Y2=0.51
r43 13 15 4.71042 $w=2.59e-07 $l=1.51987e-07 $layer=LI1_cond $X=9.53 $Y=0.89
+ $X2=9.42 $Y2=0.79
r44 13 14 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=9.53 $Y=0.89
+ $X2=9.53 $Y2=1.43
r45 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.42 $Y=1.63 $X2=9.42
+ $Y2=2.31
r46 7 14 4.71042 $w=2.59e-07 $l=1.51987e-07 $layer=LI1_cond $X=9.42 $Y=1.53
+ $X2=9.53 $Y2=1.43
r47 7 9 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=9.42 $Y=1.53 $X2=9.42
+ $Y2=1.63
r48 2 11 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.285
+ $Y=1.485 $X2=9.42 $Y2=2.31
r49 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.285
+ $Y=1.485 $X2=9.42 $Y2=1.63
r50 1 19 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=9.285
+ $Y=0.235 $X2=9.42 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%Q_N 1 2 7 11 12 26
c20 12 0 2.86308e-19 $X=11.235 $Y=1.445
c21 11 0 1.408e-19 $X=11.315 $Y=0.795
r22 16 26 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=11.315 $Y=1.57
+ $X2=11.315 $Y2=1.53
r23 12 26 1.06025 $w=2.48e-07 $l=2.3e-08 $layer=LI1_cond $X=11.315 $Y=1.507
+ $X2=11.315 $Y2=1.53
r24 12 19 10.5103 $w=2.48e-07 $l=2.28e-07 $layer=LI1_cond $X=11.315 $Y=1.592
+ $X2=11.315 $Y2=1.82
r25 12 16 1.01415 $w=2.48e-07 $l=2.2e-08 $layer=LI1_cond $X=11.315 $Y=1.592
+ $X2=11.315 $Y2=1.57
r26 11 12 21.282 $w=3.73e-07 $l=6.5e-07 $layer=LI1_cond $X=11.337 $Y=0.795
+ $X2=11.337 $Y2=1.445
r27 7 11 6.16968 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.315 $Y=0.67
+ $X2=11.315 $Y2=0.795
r28 7 9 1.952 $w=2.5e-07 $l=4e-08 $layer=LI1_cond $X=11.315 $Y=0.67 $X2=11.315
+ $Y2=0.63
r29 2 19 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=11.14
+ $Y=1.485 $X2=11.275 $Y2=1.82
r30 1 9 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=11.14
+ $Y=0.235 $X2=11.275 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 40 44 48 50
+ 54 58 62 64 66 68 70 75 80 88 96 101 106 112 115 118 121 124 127 130 133 137
c193 137 0 2.71124e-20 $X=11.73 $Y=0
r194 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r195 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r196 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r197 127 128 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r198 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r199 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r200 121 122 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r201 119 122 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r202 118 119 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r203 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r204 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r205 110 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r206 110 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=10.81 $Y2=0
r207 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r208 107 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.02 $Y=0
+ $X2=10.855 $Y2=0
r209 107 109 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=11.02 $Y=0
+ $X2=11.27 $Y2=0
r210 106 136 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=11.61 $Y=0
+ $X2=11.785 $Y2=0
r211 106 109 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.61 $Y=0
+ $X2=11.27 $Y2=0
r212 105 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r213 105 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.89 $Y2=0
r214 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r215 102 130 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=9.87 $Y2=0
r216 102 104 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=10.35 $Y2=0
r217 101 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.69 $Y=0
+ $X2=10.855 $Y2=0
r218 101 104 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.69 $Y=0
+ $X2=10.35 $Y2=0
r219 100 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r220 100 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r221 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r222 97 127 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.085 $Y=0 $X2=8.99
+ $Y2=0
r223 97 99 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.085 $Y=0 $X2=9.43
+ $Y2=0
r224 96 130 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.755 $Y=0
+ $X2=9.87 $Y2=0
r225 96 99 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.755 $Y=0
+ $X2=9.43 $Y2=0
r226 95 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r227 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r228 92 95 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r229 92 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r230 91 94 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=7.59
+ $Y2=0
r231 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r232 89 121 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=5.9
+ $Y2=0
r233 89 91 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=6.21 $Y2=0
r234 88 124 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.74 $Y=0
+ $X2=7.925 $Y2=0
r235 88 94 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.59
+ $Y2=0
r236 87 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r237 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r238 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r239 84 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r240 83 86 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r241 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r242 81 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.14 $Y2=0
r243 81 83 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r244 80 118 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.865
+ $Y2=0
r245 80 86 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.765 $Y=0
+ $X2=3.45 $Y2=0
r246 79 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r247 79 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r248 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r249 76 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r250 76 78 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r251 75 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=2.14 $Y2=0
r252 75 78 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r253 70 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r254 70 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r255 68 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r256 68 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r257 64 136 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=11.695 $Y=0.085
+ $X2=11.785 $Y2=0
r258 64 66 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.695 $Y=0.085
+ $X2=11.695 $Y2=0.38
r259 60 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.855 $Y=0.085
+ $X2=10.855 $Y2=0
r260 60 62 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.855 $Y=0.085
+ $X2=10.855 $Y2=0.38
r261 56 130 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.87 $Y=0.085
+ $X2=9.87 $Y2=0
r262 56 58 22.0467 $w=2.28e-07 $l=4.4e-07 $layer=LI1_cond $X=9.87 $Y=0.085
+ $X2=9.87 $Y2=0.525
r263 52 127 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=0.085
+ $X2=8.99 $Y2=0
r264 52 54 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=8.99 $Y=0.085
+ $X2=8.99 $Y2=0.53
r265 51 124 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.11 $Y=0
+ $X2=7.925 $Y2=0
r266 50 127 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.895 $Y=0 $X2=8.99
+ $Y2=0
r267 50 51 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.895 $Y=0
+ $X2=8.11 $Y2=0
r268 46 124 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.925 $Y=0.085
+ $X2=7.925 $Y2=0
r269 46 48 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.925 $Y=0.085
+ $X2=7.925 $Y2=0.45
r270 42 121 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0
r271 42 44 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0.42
r272 41 118 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.865
+ $Y2=0
r273 40 121 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.9
+ $Y2=0
r274 40 41 114.171 $w=1.68e-07 $l=1.75e-06 $layer=LI1_cond $X=5.715 $Y=0
+ $X2=3.965 $Y2=0
r275 36 118 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0
r276 36 38 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0.36
r277 32 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r278 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.36
r279 28 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r280 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r281 9 66 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=11.56
+ $Y=0.235 $X2=11.695 $Y2=0.38
r282 8 62 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=10.655
+ $Y=0.235 $X2=10.855 $Y2=0.38
r283 7 58 182 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_NDIFF $count=1 $X=9.705
+ $Y=0.235 $X2=9.85 $Y2=0.525
r284 6 54 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=8.845
+ $Y=0.235 $X2=8.99 $Y2=0.53
r285 5 48 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=7.89
+ $Y=0.235 $X2=8.025 $Y2=0.45
r286 4 44 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=5.665
+ $Y=0.235 $X2=5.97 $Y2=0.42
r287 3 38 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.235 $X2=3.85 $Y2=0.36
r288 2 34 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.14 $Y2=0.36
r289 1 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


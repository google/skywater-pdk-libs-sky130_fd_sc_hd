* File: sky130_fd_sc_hd__o41a_4.spice
* Created: Thu Aug 27 14:41:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o41a_4.spice.pex"
.subckt sky130_fd_sc_hd__o41a_4  VNB VPB B1 A4 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_79_21#_M1013_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A_79_21#_M1018_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1018_d N_A_79_21#_M1019_g N_X_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_A_79_21#_M1025_g N_X_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_467_47#_M1014_d N_B1_M1014_g N_A_79_21#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1015 N_A_467_47#_M1015_d N_B1_M1015_g N_A_79_21#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1002 N_A_467_47#_M1015_d N_A4_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1026 N_A_467_47#_M1026_d N_A4_M1026_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1007 N_A_467_47#_M1026_d N_A3_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1009 N_A_467_47#_M1009_d N_A3_M1009_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_A2_M1022_g N_A_467_47#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.09425 PD=1.26 PS=0.94 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75002.7
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1022_d N_A2_M1027_g N_A_467_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.15275 PD=1.26 PS=1.12 NRD=0 NRS=22.152 M=1 R=4.33333
+ SA=75003.5 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1000 N_A_467_47#_M1027_s N_A1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15275 AS=0.08775 PD=1.12 PS=0.92 NRD=12.912 NRS=0 M=1 R=4.33333
+ SA=75004.1 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1012 N_A_467_47#_M1012_d N_A1_M1012_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.3185 AS=0.08775 PD=2.28 PS=0.92 NRD=34.152 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_79_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1001_d N_A_79_21#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1020 N_X_M1020_d N_A_79_21#_M1020_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1023 N_X_M1020_d N_A_79_21#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1023_s N_B1_M1004_g N_A_79_21#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_B1_M1021_g N_A_79_21#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.145 PD=2.52 PS=1.29 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_639_297#_M1006_d N_A4_M1006_g N_A_79_21#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1010 N_A_639_297#_M1010_d N_A4_M1010_g N_A_79_21#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1003 N_A_889_297#_M1003_d N_A3_M1003_g N_A_639_297#_M1010_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1024 N_A_889_297#_M1003_d N_A3_M1024_g N_A_639_297#_M1024_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_A_1083_297#_M1011_d N_A2_M1011_g N_A_889_297#_M1011_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1016 N_A_1083_297#_M1016_d N_A2_M1016_g N_A_889_297#_M1011_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_1083_297#_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1008_d N_A1_M1017_g N_A_1083_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.49 PD=1.27 PS=2.98 NRD=0 NRS=36.445 M=1 R=6.66667 SA=75001.5
+ SB=75000.4 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__o41a_4.spice.SKY130_FD_SC_HD__O41A_4.pxi"
*
.ends
*
*

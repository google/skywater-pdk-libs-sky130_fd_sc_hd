* File: sky130_fd_sc_hd__or2_2.spice
* Created: Thu Aug 27 14:42:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or2_2.spice.pex"
.subckt sky130_fd_sc_hd__or2_2  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1007 N_A_39_297#_M1007_d N_B_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_39_297#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0838037 AS=0.0567 PD=0.788972 PS=0.69 NRD=21.42 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_39_297#_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.129696 PD=0.92 PS=1.22103 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1000_d N_A_39_297#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 A_121_297# N_B_M1004_g N_A_39_297#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_121_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0921338 AS=0.0441 PD=0.801549 PS=0.63 NRD=77.0861 NRS=23.443 M=1 R=2.8
+ SA=75000.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1001_d N_A_39_297#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.219366 AS=0.135 PD=1.90845 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_39_297#_M1005_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_174 A_121_297# 0 1.02064e-19 $X=0.605 $Y=1.485
*
.include "sky130_fd_sc_hd__or2_2.spice.SKY130_FD_SC_HD__OR2_2.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__dlrbn_2.spice.SKY130_FD_SC_HD__DLRBN_2.pxi
* Created: Thu Aug 27 14:16:47 2020
* 
x_PM_SKY130_FD_SC_HD__DLRBN_2%GATE_N N_GATE_N_c_180_n N_GATE_N_c_175_n
+ N_GATE_N_M1024_g N_GATE_N_c_181_n N_GATE_N_M1014_g N_GATE_N_c_176_n
+ N_GATE_N_c_182_n GATE_N GATE_N N_GATE_N_c_178_n N_GATE_N_c_179_n
+ PM_SKY130_FD_SC_HD__DLRBN_2%GATE_N
x_PM_SKY130_FD_SC_HD__DLRBN_2%A_27_47# N_A_27_47#_M1024_s N_A_27_47#_M1014_s
+ N_A_27_47#_M1015_g N_A_27_47#_M1000_g N_A_27_47#_M1019_g N_A_27_47#_M1005_g
+ N_A_27_47#_c_219_n N_A_27_47#_c_220_n N_A_27_47#_c_221_n N_A_27_47#_c_231_n
+ N_A_27_47#_c_232_n N_A_27_47#_c_233_n N_A_27_47#_c_222_n N_A_27_47#_c_223_n
+ N_A_27_47#_c_224_n N_A_27_47#_c_225_n N_A_27_47#_c_235_n N_A_27_47#_c_236_n
+ N_A_27_47#_c_237_n N_A_27_47#_c_238_n N_A_27_47#_c_239_n N_A_27_47#_c_226_n
+ N_A_27_47#_c_227_n N_A_27_47#_c_241_n N_A_27_47#_c_228_n
+ PM_SKY130_FD_SC_HD__DLRBN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRBN_2%D N_D_M1006_g N_D_M1022_g D N_D_c_388_n
+ N_D_c_389_n PM_SKY130_FD_SC_HD__DLRBN_2%D
x_PM_SKY130_FD_SC_HD__DLRBN_2%A_299_47# N_A_299_47#_M1006_s N_A_299_47#_M1022_s
+ N_A_299_47#_M1013_g N_A_299_47#_M1017_g N_A_299_47#_c_434_n
+ N_A_299_47#_c_427_n N_A_299_47#_c_435_n N_A_299_47#_c_436_n
+ N_A_299_47#_c_428_n N_A_299_47#_c_429_n N_A_299_47#_c_430_n
+ N_A_299_47#_c_431_n N_A_299_47#_c_432_n PM_SKY130_FD_SC_HD__DLRBN_2%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRBN_2%A_193_47# N_A_193_47#_M1015_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1001_g N_A_193_47#_c_509_n N_A_193_47#_c_510_n
+ N_A_193_47#_M1011_g N_A_193_47#_c_516_n N_A_193_47#_c_512_n
+ N_A_193_47#_c_518_n N_A_193_47#_c_519_n N_A_193_47#_c_520_n
+ N_A_193_47#_c_521_n N_A_193_47#_c_522_n N_A_193_47#_c_523_n
+ N_A_193_47#_c_524_n PM_SKY130_FD_SC_HD__DLRBN_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRBN_2%A_724_21# N_A_724_21#_M1012_s N_A_724_21#_M1004_d
+ N_A_724_21#_M1020_g N_A_724_21#_M1009_g N_A_724_21#_c_622_n
+ N_A_724_21#_M1018_g N_A_724_21#_M1007_g N_A_724_21#_c_623_n
+ N_A_724_21#_M1025_g N_A_724_21#_M1026_g N_A_724_21#_c_624_n
+ N_A_724_21#_c_625_n N_A_724_21#_c_626_n N_A_724_21#_c_637_n
+ N_A_724_21#_c_627_n N_A_724_21#_M1021_g N_A_724_21#_c_638_n
+ N_A_724_21#_M1010_g N_A_724_21#_c_639_n N_A_724_21#_c_640_n
+ N_A_724_21#_c_641_n N_A_724_21#_c_649_p N_A_724_21#_c_709_p
+ N_A_724_21#_c_671_p N_A_724_21#_c_642_n N_A_724_21#_c_655_p
+ N_A_724_21#_c_676_p N_A_724_21#_c_628_n N_A_724_21#_c_629_n
+ PM_SKY130_FD_SC_HD__DLRBN_2%A_724_21#
x_PM_SKY130_FD_SC_HD__DLRBN_2%A_561_413# N_A_561_413#_M1019_d
+ N_A_561_413#_M1001_d N_A_561_413#_c_768_n N_A_561_413#_M1012_g
+ N_A_561_413#_M1004_g N_A_561_413#_c_769_n N_A_561_413#_c_770_n
+ N_A_561_413#_c_779_n N_A_561_413#_c_782_n N_A_561_413#_c_771_n
+ N_A_561_413#_c_772_n N_A_561_413#_c_777_n N_A_561_413#_c_773_n
+ PM_SKY130_FD_SC_HD__DLRBN_2%A_561_413#
x_PM_SKY130_FD_SC_HD__DLRBN_2%RESET_B N_RESET_B_c_849_n N_RESET_B_M1008_g
+ N_RESET_B_M1016_g RESET_B N_RESET_B_c_850_n N_RESET_B_c_851_n
+ PM_SKY130_FD_SC_HD__DLRBN_2%RESET_B
x_PM_SKY130_FD_SC_HD__DLRBN_2%A_1313_47# N_A_1313_47#_M1021_s
+ N_A_1313_47#_M1010_s N_A_1313_47#_c_886_n N_A_1313_47#_M1003_g
+ N_A_1313_47#_M1002_g N_A_1313_47#_c_887_n N_A_1313_47#_c_888_n
+ N_A_1313_47#_M1027_g N_A_1313_47#_M1023_g N_A_1313_47#_c_891_n
+ N_A_1313_47#_c_892_n N_A_1313_47#_c_897_n N_A_1313_47#_c_893_n
+ N_A_1313_47#_c_913_n PM_SKY130_FD_SC_HD__DLRBN_2%A_1313_47#
x_PM_SKY130_FD_SC_HD__DLRBN_2%VPWR N_VPWR_M1014_d N_VPWR_M1022_d N_VPWR_M1009_d
+ N_VPWR_M1004_s N_VPWR_M1016_d N_VPWR_M1026_s N_VPWR_M1010_d N_VPWR_M1023_s
+ N_VPWR_c_964_n N_VPWR_c_965_n N_VPWR_c_966_n N_VPWR_c_967_n N_VPWR_c_968_n
+ N_VPWR_c_969_n N_VPWR_c_970_n N_VPWR_c_971_n N_VPWR_c_972_n VPWR
+ N_VPWR_c_973_n N_VPWR_c_974_n N_VPWR_c_975_n N_VPWR_c_976_n N_VPWR_c_977_n
+ N_VPWR_c_978_n N_VPWR_c_979_n N_VPWR_c_980_n N_VPWR_c_981_n N_VPWR_c_982_n
+ N_VPWR_c_983_n N_VPWR_c_963_n PM_SKY130_FD_SC_HD__DLRBN_2%VPWR
x_PM_SKY130_FD_SC_HD__DLRBN_2%Q N_Q_M1018_s N_Q_M1007_d N_Q_c_1096_n
+ N_Q_c_1098_n N_Q_c_1110_n Q Q Q N_Q_c_1114_n PM_SKY130_FD_SC_HD__DLRBN_2%Q
x_PM_SKY130_FD_SC_HD__DLRBN_2%Q_N N_Q_N_M1003_d N_Q_N_M1002_d N_Q_N_c_1130_n
+ N_Q_N_c_1139_n N_Q_N_c_1132_n Q_N Q_N Q_N Q_N Q_N
+ PM_SKY130_FD_SC_HD__DLRBN_2%Q_N
x_PM_SKY130_FD_SC_HD__DLRBN_2%VGND N_VGND_M1024_d N_VGND_M1006_d N_VGND_M1020_d
+ N_VGND_M1008_d N_VGND_M1025_d N_VGND_M1021_d N_VGND_M1027_s N_VGND_c_1159_n
+ N_VGND_c_1160_n N_VGND_c_1161_n N_VGND_c_1162_n N_VGND_c_1163_n
+ N_VGND_c_1164_n N_VGND_c_1165_n N_VGND_c_1166_n VGND N_VGND_c_1167_n
+ N_VGND_c_1168_n N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n
+ N_VGND_c_1176_n N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n
+ N_VGND_c_1180_n PM_SKY130_FD_SC_HD__DLRBN_2%VGND
cc_1 VNB N_GATE_N_c_175_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_176_n 0.0231103f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0128731f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_178_n 0.0212735f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_179_n 0.0148043f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1015_g 0.0397896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_219_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_8 VNB N_A_27_47#_c_220_n 0.00222599f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_9 VNB N_A_27_47#_c_221_n 0.00793517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_222_n 7.842e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_223_n 0.00418741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_224_n 0.0271287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_225_n 0.00378508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_226_n 0.0230814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_227_n 0.0176114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_228_n 0.00469707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1006_g 0.025905f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_18 VNB N_D_M1022_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_19 VNB N_D_c_388_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_20 VNB N_D_c_389_n 0.0421785f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_21 VNB N_A_299_47#_M1017_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_427_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_428_n 0.00496114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_299_47#_c_429_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_25 VNB N_A_299_47#_c_430_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_26 VNB N_A_299_47#_c_431_n 0.0274388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_299_47#_c_432_n 0.01709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_509_n 0.0133385f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_29 VNB N_A_193_47#_c_510_n 0.00520223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_M1011_g 0.0464035f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_31 VNB N_A_193_47#_c_512_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_724_21#_M1020_g 0.0506249f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_33 VNB N_A_724_21#_c_622_n 0.0155418f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_34 VNB N_A_724_21#_c_623_n 0.019441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_724_21#_c_624_n 0.0397733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_724_21#_c_625_n 0.0274505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_724_21#_c_626_n 0.0342609f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_38 VNB N_A_724_21#_c_627_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_724_21#_c_628_n 0.00183535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_724_21#_c_629_n 0.00105339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_561_413#_c_768_n 0.0222234f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_42 VNB N_A_561_413#_c_769_n 0.0434828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_561_413#_c_770_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_44 VNB N_A_561_413#_c_771_n 0.00691811f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_45 VNB N_A_561_413#_c_772_n 0.0118438f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_46 VNB N_A_561_413#_c_773_n 0.00194757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_849_n 0.0161955f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_48 VNB N_RESET_B_c_850_n 0.0200304f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_49 VNB N_RESET_B_c_851_n 0.0019514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1313_47#_c_886_n 0.0169457f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_51 VNB N_A_1313_47#_c_887_n 0.01318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1313_47#_c_888_n 0.0191396f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_53 VNB N_A_1313_47#_M1027_g 0.0238416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1313_47#_M1023_g 5.18715e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1313_47#_c_891_n 0.0128325f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_56 VNB N_A_1313_47#_c_892_n 0.00901723f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_57 VNB N_A_1313_47#_c_893_n 0.00489864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_963_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_Q_c_1096_n 0.0023168f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_60 VNB N_Q_N_c_1130_n 0.00121852f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_61 VNB Q_N 0.0157064f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_62 VNB N_VGND_c_1159_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_63 VNB N_VGND_c_1160_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_64 VNB N_VGND_c_1161_n 0.012582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1162_n 4.11979e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1163_n 0.00765821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1164_n 0.00201517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1165_n 0.0101024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1166_n 0.0320347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1167_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1168_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1169_n 0.0412073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1170_n 0.0278531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1171_n 0.0160822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1172_n 0.0180452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1173_n 0.0153174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1174_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1175_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1176_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1177_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1178_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1179_n 0.00459225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1180_n 0.417662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VPB N_GATE_N_c_180_n 0.0128858f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_85 VPB N_GATE_N_c_181_n 0.0186097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_86 VPB N_GATE_N_c_182_n 0.023868f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_87 VPB GATE_N 0.0128465f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_88 VPB N_GATE_N_c_178_n 0.01087f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_89 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_90 VPB N_A_27_47#_M1005_g 0.0212472f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_91 VPB N_A_27_47#_c_231_n 0.00124413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_47#_c_232_n 0.00556025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_27_47#_c_233_n 0.0300266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_47#_c_222_n 5.99662e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_c_235_n 0.0280095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_27_47#_c_236_n 0.00366942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_47#_c_237_n 0.00546122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_27_47#_c_238_n 0.0035222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_47#_c_239_n 0.0037442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_c_226_n 0.0115924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_47#_c_241_n 0.0330434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_c_228_n 2.971e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_D_M1022_g 0.0462846f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_104 VPB N_D_c_388_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_105 VPB N_A_299_47#_M1017_g 0.0366887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_299_47#_c_434_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_299_47#_c_435_n 0.00415091f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_108 VPB N_A_299_47#_c_436_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_299_47#_c_429_n 0.00361895f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_110 VPB N_A_193_47#_M1001_g 0.0316829f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_111 VPB N_A_193_47#_c_509_n 0.0172364f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_112 VPB N_A_193_47#_c_510_n 0.00687211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_193_47#_c_516_n 0.0117991f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_114 VPB N_A_193_47#_c_512_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_193_47#_c_518_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_116 VPB N_A_193_47#_c_519_n 0.00515533f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_117 VPB N_A_193_47#_c_520_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_118 VPB N_A_193_47#_c_521_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_193_47#_c_522_n 0.00114133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_193_47#_c_523_n 0.0104341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_193_47#_c_524_n 0.0126899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_724_21#_M1020_g 0.0180275f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_123 VPB N_A_724_21#_M1009_g 0.0275278f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_124 VPB N_A_724_21#_M1007_g 0.0184875f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_125 VPB N_A_724_21#_M1026_g 0.0231478f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_126 VPB N_A_724_21#_c_624_n 0.019214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_724_21#_c_625_n 0.0053174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_724_21#_c_626_n 6.08077e-19 $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_129 VPB N_A_724_21#_c_637_n 0.0171146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_724_21#_c_638_n 0.0183859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_724_21#_c_639_n 0.0185209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_724_21#_c_640_n 0.00725325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_724_21#_c_641_n 0.0414048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_724_21#_c_642_n 0.00153659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_561_413#_M1004_g 0.0254462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_561_413#_c_769_n 0.0148072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_561_413#_c_770_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_138 VPB N_A_561_413#_c_777_n 0.00517422f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_139 VPB N_A_561_413#_c_773_n 0.00161757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_M1016_g 0.018858f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_141 VPB N_RESET_B_c_850_n 0.00399554f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_142 VPB N_RESET_B_c_851_n 0.00194848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_1313_47#_M1002_g 0.0198362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_1313_47#_c_888_n 0.00570712f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_145 VPB N_A_1313_47#_M1023_g 0.0265634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_1313_47#_c_897_n 0.0150366f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_147 VPB N_A_1313_47#_c_893_n 0.0054092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_964_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_149 VPB N_VPWR_c_965_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_150 VPB N_VPWR_c_966_n 0.00226627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_967_n 0.0121273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_968_n 0.00281522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_969_n 0.0100765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_970_n 0.0432338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_971_n 0.0125756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_972_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_973_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_974_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_975_n 0.0207222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_976_n 0.0183604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_977_n 0.0153174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_978_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_979_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_980_n 0.0406078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_981_n 0.0250891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_982_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_983_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_963_n 0.0597682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_Q_c_1096_n 0.00354692f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_170 VPB N_Q_c_1098_n 0.00121379f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_171 VPB N_Q_N_c_1132_n 0.00222192f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_172 VPB Q_N 0.00519938f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_173 N_GATE_N_c_175_n N_A_27_47#_M1015_g 0.018782f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_174 N_GATE_N_c_179_n N_A_27_47#_M1015_g 0.00419152f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_175 N_GATE_N_c_182_n N_A_27_47#_M1000_g 0.0260324f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_176 N_GATE_N_c_178_n N_A_27_47#_M1000_g 0.0052657f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_177 N_GATE_N_c_175_n N_A_27_47#_c_220_n 0.00674622f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_178 N_GATE_N_c_176_n N_A_27_47#_c_220_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_179 N_GATE_N_c_176_n N_A_27_47#_c_221_n 0.00672951f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_180 GATE_N N_A_27_47#_c_221_n 0.0202563f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_181 N_GATE_N_c_178_n N_A_27_47#_c_221_n 7.62625e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_182 N_GATE_N_c_181_n N_A_27_47#_c_231_n 0.0135762f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_183 N_GATE_N_c_182_n N_A_27_47#_c_231_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_184 N_GATE_N_c_181_n N_A_27_47#_c_233_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_185 N_GATE_N_c_182_n N_A_27_47#_c_233_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_186 GATE_N N_A_27_47#_c_233_n 0.0221922f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_187 N_GATE_N_c_178_n N_A_27_47#_c_233_n 5.90345e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_188 N_GATE_N_c_178_n N_A_27_47#_c_222_n 0.0032236f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_189 N_GATE_N_c_176_n N_A_27_47#_c_223_n 0.00181464f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_190 GATE_N N_A_27_47#_c_223_n 0.0293747f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_191 N_GATE_N_c_179_n N_A_27_47#_c_223_n 0.0015333f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_192 N_GATE_N_c_180_n N_A_27_47#_c_236_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_193 N_GATE_N_c_182_n N_A_27_47#_c_236_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_194 GATE_N N_A_27_47#_c_236_n 0.0065266f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_195 N_GATE_N_c_180_n N_A_27_47#_c_237_n 7.65064e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_182_n N_A_27_47#_c_237_n 0.00432523f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_197 GATE_N N_A_27_47#_c_226_n 9.03754e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_198 N_GATE_N_c_178_n N_A_27_47#_c_226_n 0.0165848f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_199 N_GATE_N_c_181_n N_VPWR_c_964_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_200 N_GATE_N_c_181_n N_VPWR_c_973_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_201 N_GATE_N_c_181_n N_VPWR_c_963_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_202 N_GATE_N_c_175_n N_VGND_c_1159_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_203 N_GATE_N_c_175_n N_VGND_c_1167_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_204 N_GATE_N_c_176_n N_VGND_c_1167_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_205 N_GATE_N_c_175_n N_VGND_c_1180_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_235_n N_D_M1022_g 0.00583826f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_235_n N_D_c_388_n 0.0087134f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1015_g N_D_c_389_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_235_n N_A_299_47#_M1017_g 0.00493352f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_228_n N_A_299_47#_M1017_g 0.00369716f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_211 N_A_27_47#_c_235_n N_A_299_47#_c_435_n 0.0116478f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_235_n N_A_299_47#_c_436_n 0.0115067f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_224_n N_A_299_47#_c_428_n 9.56555e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_225_n N_A_299_47#_c_428_n 0.0129081f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_235_n N_A_299_47#_c_428_n 0.00675641f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_228_n N_A_299_47#_c_428_n 0.00178567f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_217 N_A_27_47#_c_235_n N_A_299_47#_c_429_n 0.0108506f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_224_n N_A_299_47#_c_431_n 0.0117556f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_225_n N_A_299_47#_c_431_n 9.50608e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_235_n N_A_299_47#_c_431_n 0.00107604f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_228_n N_A_299_47#_c_431_n 9.9633e-19 $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_224_n N_A_299_47#_c_432_n 0.00200147f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_225_n N_A_299_47#_c_432_n 2.04855e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_227_n N_A_299_47#_c_432_n 0.0197936f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_M1005_g N_A_193_47#_M1001_g 0.014011f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_232_n N_A_193_47#_M1001_g 0.00220245f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_225_n N_A_193_47#_c_509_n 7.03475e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_235_n N_A_193_47#_c_509_n 0.00144279f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_238_n N_A_193_47#_c_509_n 0.00140497f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_239_n N_A_193_47#_c_509_n 0.0049391f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_241_n N_A_193_47#_c_509_n 0.0184089f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_228_n N_A_193_47#_c_509_n 0.01293f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_224_n N_A_193_47#_c_510_n 0.0186665f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_225_n N_A_193_47#_c_510_n 0.00136525f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_224_n N_A_193_47#_M1011_g 0.0192792f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_225_n N_A_193_47#_M1011_g 0.00256371f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_227_n N_A_193_47#_M1011_g 0.0126141f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_228_n N_A_193_47#_M1011_g 0.0049729f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_235_n N_A_193_47#_c_516_n 0.00274258f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_238_n N_A_193_47#_c_516_n 7.88621e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_239_n N_A_193_47#_c_516_n 0.00220245f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_241_n N_A_193_47#_c_516_n 0.0160512f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_M1015_g N_A_193_47#_c_512_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_220_n N_A_193_47#_c_512_n 0.0100297f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_222_n N_A_193_47#_c_512_n 0.0235786f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_223_n N_A_193_47#_c_512_n 0.0158689f $X=0.722 $Y=1.07 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_235_n N_A_193_47#_c_512_n 0.0184539f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_236_n N_A_193_47#_c_512_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_237_n N_A_193_47#_c_512_n 0.0208435f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_231_n N_A_193_47#_c_518_n 0.00294892f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_235_n N_A_193_47#_c_518_n 0.00195186f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_226_n N_A_193_47#_c_518_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_235_n N_A_193_47#_c_519_n 0.0871075f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1000_g N_A_193_47#_c_520_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_231_n N_A_193_47#_c_520_n 0.00551586f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_235_n N_A_193_47#_c_520_n 0.0259095f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_237_n N_A_193_47#_c_520_n 0.00110596f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1000_g N_A_193_47#_c_521_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_232_n N_A_193_47#_c_522_n 0.00155445f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_235_n N_A_193_47#_c_522_n 0.0255946f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_235_n N_A_193_47#_c_523_n 0.00169866f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_238_n N_A_193_47#_c_523_n 0.00124306f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_228_n N_A_193_47#_c_523_n 0.00220245f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_264 N_A_27_47#_c_224_n N_A_193_47#_c_524_n 4.0812e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_225_n N_A_193_47#_c_524_n 0.00161882f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_235_n N_A_193_47#_c_524_n 0.0240266f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_238_n N_A_193_47#_c_524_n 0.00272314f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_241_n N_A_193_47#_c_524_n 2.5966e-19 $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_228_n N_A_193_47#_c_524_n 0.0454941f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_239_n N_A_724_21#_M1020_g 4.9921e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_228_n N_A_724_21#_M1020_g 2.17095e-19 $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_272 N_A_27_47#_M1005_g N_A_724_21#_M1009_g 0.0313444f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_232_n N_A_724_21#_c_641_n 8.09252e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_241_n N_A_724_21#_c_641_n 0.0313444f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_224_n N_A_561_413#_c_779_n 0.00144439f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_225_n N_A_561_413#_c_779_n 0.0162478f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_227_n N_A_561_413#_c_779_n 0.00412044f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1005_g N_A_561_413#_c_782_n 0.0116262f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_279 N_A_27_47#_c_232_n N_A_561_413#_c_782_n 0.016081f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_238_n N_A_561_413#_c_782_n 0.00173361f $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_241_n N_A_561_413#_c_782_n 0.00111122f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_282 N_A_27_47#_c_225_n N_A_561_413#_c_771_n 0.0184898f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_225_n N_A_561_413#_c_772_n 0.0027819f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_241_n N_A_561_413#_c_772_n 0.00291146f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_285 N_A_27_47#_c_228_n N_A_561_413#_c_772_n 0.016104f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_238_n N_A_561_413#_c_777_n 0.00130345f $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_239_n N_A_561_413#_c_777_n 0.0359174f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_241_n N_A_561_413#_c_777_n 0.00856317f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_228_n N_A_561_413#_c_777_n 0.00353544f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_231_n N_VPWR_M1014_d 0.00191359f $X=0.605 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_291 N_A_27_47#_M1000_g N_VPWR_c_964_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_231_n N_VPWR_c_964_n 0.0150624f $X=0.605 $Y=1.88 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_233_n N_VPWR_c_964_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_236_n N_VPWR_c_964_n 0.00311191f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_235_n N_VPWR_c_965_n 0.0019389f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_231_n N_VPWR_c_973_n 0.0018545f $X=0.605 $Y=1.88 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_233_n N_VPWR_c_973_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_298 N_A_27_47#_M1000_g N_VPWR_c_974_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1005_g N_VPWR_c_980_n 0.00366111f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1000_g N_VPWR_c_963_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1005_g N_VPWR_c_963_n 0.00549379f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_231_n N_VPWR_c_963_n 0.00483604f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_233_n N_VPWR_c_963_n 0.00993215f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_220_n N_VGND_M1024_d 0.00164702f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_305 N_A_27_47#_M1015_g N_VGND_c_1159_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_220_n N_VGND_c_1159_n 0.0150545f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_222_n N_VGND_c_1159_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_226_n N_VGND_c_1159_n 5.88506e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_227_n N_VGND_c_1160_n 0.00174223f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_219_n N_VGND_c_1167_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_220_n N_VGND_c_1167_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_M1015_g N_VGND_c_1168_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_224_n N_VGND_c_1169_n 9.43262e-19 $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_314 N_A_27_47#_c_225_n N_VGND_c_1169_n 0.00182549f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_227_n N_VGND_c_1169_n 0.00425892f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_M1024_s N_VGND_c_1180_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_M1015_g N_VGND_c_1180_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_219_n N_VGND_c_1180_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_220_n N_VGND_c_1180_n 0.00549621f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_224_n N_VGND_c_1180_n 0.00121904f $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_321 N_A_27_47#_c_225_n N_VGND_c_1180_n 0.00328555f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_227_n N_VGND_c_1180_n 0.00628992f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_323 N_D_c_389_n N_A_299_47#_M1017_g 0.0382098f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_324 N_D_M1022_g N_A_299_47#_c_434_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_325 N_D_M1006_g N_A_299_47#_c_427_n 0.0144498f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_326 N_D_c_388_n N_A_299_47#_c_427_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_327 N_D_c_389_n N_A_299_47#_c_427_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_328 N_D_M1022_g N_A_299_47#_c_435_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_329 N_D_M1022_g N_A_299_47#_c_436_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_330 N_D_c_388_n N_A_299_47#_c_436_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_331 N_D_c_389_n N_A_299_47#_c_436_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_332 N_D_M1006_g N_A_299_47#_c_428_n 0.00563568f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_333 N_D_c_388_n N_A_299_47#_c_428_n 0.0107593f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_334 N_D_c_388_n N_A_299_47#_c_429_n 0.0164827f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_335 N_D_c_389_n N_A_299_47#_c_429_n 0.00552652f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_336 N_D_M1006_g N_A_299_47#_c_430_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_337 N_D_c_388_n N_A_299_47#_c_430_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_338 N_D_c_389_n N_A_299_47#_c_430_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_339 N_D_M1006_g N_A_299_47#_c_431_n 0.0197208f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_340 N_D_M1006_g N_A_299_47#_c_432_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_341 N_D_M1006_g N_A_193_47#_c_512_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_342 N_D_M1022_g N_A_193_47#_c_512_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_343 N_D_c_388_n N_A_193_47#_c_512_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_344 N_D_c_389_n N_A_193_47#_c_512_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_345 N_D_M1022_g N_A_193_47#_c_518_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_346 N_D_M1022_g N_A_193_47#_c_519_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_347 N_D_M1022_g N_VPWR_c_965_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_348 N_D_M1022_g N_VPWR_c_974_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_349 N_D_M1022_g N_VPWR_c_963_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_350 N_D_M1006_g N_VGND_c_1160_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_351 N_D_M1006_g N_VGND_c_1168_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_352 N_D_M1006_g N_VGND_c_1180_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_353 N_D_c_389_n N_VGND_c_1180_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_354 N_A_299_47#_M1017_g N_A_193_47#_M1001_g 0.0342299f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_355 N_A_299_47#_M1017_g N_A_193_47#_c_510_n 0.0248238f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_356 N_A_299_47#_c_434_n N_A_193_47#_c_512_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_357 N_A_299_47#_c_436_n N_A_193_47#_c_512_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_358 N_A_299_47#_c_430_n N_A_193_47#_c_512_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_359 N_A_299_47#_c_434_n N_A_193_47#_c_518_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_360 N_A_299_47#_M1017_g N_A_193_47#_c_519_n 0.00365242f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_361 N_A_299_47#_c_434_n N_A_193_47#_c_519_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_362 N_A_299_47#_c_435_n N_A_193_47#_c_519_n 0.00551435f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_363 N_A_299_47#_c_434_n N_A_193_47#_c_520_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_364 N_A_299_47#_M1017_g N_A_193_47#_c_522_n 0.00149195f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_365 N_A_299_47#_M1017_g N_A_193_47#_c_524_n 0.00673436f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_366 N_A_299_47#_c_435_n N_A_193_47#_c_524_n 0.00754519f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_367 N_A_299_47#_c_429_n N_A_193_47#_c_524_n 0.00645446f $X=2.055 $Y=1.495
+ $X2=0 $Y2=0
cc_368 N_A_299_47#_c_432_n N_A_561_413#_c_779_n 6.54613e-19 $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_369 N_A_299_47#_M1017_g N_VPWR_c_965_n 0.0223997f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_370 N_A_299_47#_c_434_n N_VPWR_c_965_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_371 N_A_299_47#_c_435_n N_VPWR_c_965_n 0.013562f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_372 N_A_299_47#_c_434_n N_VPWR_c_974_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_373 N_A_299_47#_M1017_g N_VPWR_c_980_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_374 N_A_299_47#_M1022_s N_VPWR_c_963_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_375 N_A_299_47#_M1017_g N_VPWR_c_963_n 0.00262666f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_376 N_A_299_47#_c_434_n N_VPWR_c_963_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_377 N_A_299_47#_c_428_n N_VGND_M1006_d 0.00156939f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_378 N_A_299_47#_c_427_n N_VGND_c_1160_n 0.00259081f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_379 N_A_299_47#_c_428_n N_VGND_c_1160_n 0.0141976f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_380 N_A_299_47#_c_432_n N_VGND_c_1160_n 0.00964732f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_381 N_A_299_47#_c_427_n N_VGND_c_1168_n 0.00255672f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_382 N_A_299_47#_c_430_n N_VGND_c_1168_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_383 N_A_299_47#_c_431_n N_VGND_c_1169_n 9.84895e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_384 N_A_299_47#_c_432_n N_VGND_c_1169_n 0.0046653f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_385 N_A_299_47#_M1006_s N_VGND_c_1180_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_386 N_A_299_47#_c_427_n N_VGND_c_1180_n 0.00473142f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_387 N_A_299_47#_c_428_n N_VGND_c_1180_n 0.00552372f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_388 N_A_299_47#_c_430_n N_VGND_c_1180_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_389 N_A_299_47#_c_431_n N_VGND_c_1180_n 0.00117722f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_390 N_A_299_47#_c_432_n N_VGND_c_1180_n 0.00454932f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_391 N_A_193_47#_M1011_g N_A_724_21#_M1020_g 0.0429763f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_392 N_A_193_47#_M1011_g N_A_561_413#_c_779_n 0.0125662f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_393 N_A_193_47#_M1001_g N_A_561_413#_c_782_n 0.00281839f $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_394 N_A_193_47#_M1011_g N_A_561_413#_c_771_n 0.00562201f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_395 N_A_193_47#_M1011_g N_A_561_413#_c_772_n 0.00348305f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_396 N_A_193_47#_M1001_g N_A_561_413#_c_777_n 8.05921e-19 $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_397 N_A_193_47#_c_509_n N_A_561_413#_c_777_n 6.71539e-19 $X=3.145 $Y=1.32
+ $X2=0 $Y2=0
cc_398 N_A_193_47#_c_519_n N_VPWR_M1022_d 6.81311e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_399 N_A_193_47#_c_521_n N_VPWR_c_964_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_400 N_A_193_47#_M1001_g N_VPWR_c_965_n 0.00357414f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_401 N_A_193_47#_c_519_n N_VPWR_c_965_n 0.0171797f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_402 N_A_193_47#_c_522_n N_VPWR_c_965_n 0.0013481f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_403 N_A_193_47#_c_524_n N_VPWR_c_965_n 0.00972665f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_404 N_A_193_47#_c_521_n N_VPWR_c_974_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_405 N_A_193_47#_M1001_g N_VPWR_c_980_n 0.00487021f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_406 N_A_193_47#_c_524_n N_VPWR_c_980_n 0.00456724f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_407 N_A_193_47#_M1001_g N_VPWR_c_963_n 0.00815857f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_408 N_A_193_47#_c_519_n N_VPWR_c_963_n 0.0516753f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_409 N_A_193_47#_c_520_n N_VPWR_c_963_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_410 N_A_193_47#_c_521_n N_VPWR_c_963_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_411 N_A_193_47#_c_522_n N_VPWR_c_963_n 0.0151013f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_412 N_A_193_47#_c_524_n N_VPWR_c_963_n 0.00403974f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_413 N_A_193_47#_c_519_n A_465_369# 0.00119229f $X=2.41 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_414 N_A_193_47#_c_522_n A_465_369# 0.00120144f $X=2.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_415 N_A_193_47#_c_524_n A_465_369# 0.0030615f $X=2.67 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_416 N_A_193_47#_M1011_g N_VGND_c_1161_n 0.0018373f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_417 N_A_193_47#_c_512_n N_VGND_c_1168_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_418 N_A_193_47#_M1011_g N_VGND_c_1169_n 0.0037981f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_419 N_A_193_47#_M1015_d N_VGND_c_1180_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_A_193_47#_M1011_g N_VGND_c_1180_n 0.00555936f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_421 N_A_193_47#_c_512_n N_VGND_c_1180_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_422 N_A_724_21#_c_649_p N_A_561_413#_c_768_n 0.00981052f $X=5.31 $Y=0.74
+ $X2=0 $Y2=0
cc_423 N_A_724_21#_c_640_n N_A_561_413#_M1004_g 0.0184636f $X=4.76 $Y=1.68 $X2=0
+ $Y2=0
cc_424 N_A_724_21#_c_641_n N_A_561_413#_M1004_g 0.00639026f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_425 N_A_724_21#_M1020_g N_A_561_413#_c_769_n 0.0214321f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_426 N_A_724_21#_c_640_n N_A_561_413#_c_769_n 0.0145535f $X=4.76 $Y=1.68 $X2=0
+ $Y2=0
cc_427 N_A_724_21#_c_641_n N_A_561_413#_c_769_n 0.00500108f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_428 N_A_724_21#_c_655_p N_A_561_413#_c_769_n 0.00514482f $X=4.425 $Y=0.58
+ $X2=0 $Y2=0
cc_429 N_A_724_21#_M1020_g N_A_561_413#_c_779_n 0.00148607f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_430 N_A_724_21#_M1009_g N_A_561_413#_c_782_n 0.00369339f $X=3.695 $Y=2.275
+ $X2=0 $Y2=0
cc_431 N_A_724_21#_M1020_g N_A_561_413#_c_771_n 0.00598699f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_432 N_A_724_21#_M1020_g N_A_561_413#_c_772_n 0.00570022f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_433 N_A_724_21#_M1020_g N_A_561_413#_c_777_n 0.0103141f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_434 N_A_724_21#_M1009_g N_A_561_413#_c_777_n 0.0144032f $X=3.695 $Y=2.275
+ $X2=0 $Y2=0
cc_435 N_A_724_21#_c_640_n N_A_561_413#_c_777_n 0.0257766f $X=4.76 $Y=1.68 $X2=0
+ $Y2=0
cc_436 N_A_724_21#_c_641_n N_A_561_413#_c_777_n 0.00825753f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_437 N_A_724_21#_M1020_g N_A_561_413#_c_773_n 0.0170014f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_438 N_A_724_21#_c_640_n N_A_561_413#_c_773_n 0.0293281f $X=4.76 $Y=1.68 $X2=0
+ $Y2=0
cc_439 N_A_724_21#_c_641_n N_A_561_413#_c_773_n 0.00373366f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_440 N_A_724_21#_c_622_n N_RESET_B_c_849_n 0.0262014f $X=5.475 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_441 N_A_724_21#_c_649_p N_RESET_B_c_849_n 0.0114332f $X=5.31 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_442 N_A_724_21#_c_629_n N_RESET_B_c_849_n 0.00341753f $X=5.465 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_443 N_A_724_21#_M1007_g N_RESET_B_M1016_g 0.0287414f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_724_21#_c_671_p N_RESET_B_M1016_g 0.012767f $X=5.31 $Y=1.58 $X2=0
+ $Y2=0
cc_445 N_A_724_21#_c_642_n N_RESET_B_M1016_g 0.00341753f $X=5.395 $Y=1.495 $X2=0
+ $Y2=0
cc_446 N_A_724_21#_c_625_n N_RESET_B_c_850_n 0.0202849f $X=6.025 $Y=1.16 $X2=0
+ $Y2=0
cc_447 N_A_724_21#_c_649_p N_RESET_B_c_850_n 0.00245514f $X=5.31 $Y=0.74 $X2=0
+ $Y2=0
cc_448 N_A_724_21#_c_671_p N_RESET_B_c_850_n 0.00123496f $X=5.31 $Y=1.58 $X2=0
+ $Y2=0
cc_449 N_A_724_21#_c_676_p N_RESET_B_c_850_n 2.11627e-19 $X=4.845 $Y=1.755 $X2=0
+ $Y2=0
cc_450 N_A_724_21#_c_628_n N_RESET_B_c_850_n 0.00202421f $X=5.535 $Y=1.16 $X2=0
+ $Y2=0
cc_451 N_A_724_21#_c_625_n N_RESET_B_c_851_n 3.10361e-19 $X=6.025 $Y=1.16 $X2=0
+ $Y2=0
cc_452 N_A_724_21#_c_640_n N_RESET_B_c_851_n 0.0243889f $X=4.76 $Y=1.68 $X2=0
+ $Y2=0
cc_453 N_A_724_21#_c_649_p N_RESET_B_c_851_n 0.0384591f $X=5.31 $Y=0.74 $X2=0
+ $Y2=0
cc_454 N_A_724_21#_c_671_p N_RESET_B_c_851_n 0.0129632f $X=5.31 $Y=1.58 $X2=0
+ $Y2=0
cc_455 N_A_724_21#_c_655_p N_RESET_B_c_851_n 0.0110762f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_456 N_A_724_21#_c_676_p N_RESET_B_c_851_n 0.014068f $X=4.845 $Y=1.755 $X2=0
+ $Y2=0
cc_457 N_A_724_21#_c_628_n N_RESET_B_c_851_n 0.0273934f $X=5.535 $Y=1.16 $X2=0
+ $Y2=0
cc_458 N_A_724_21#_c_626_n N_A_1313_47#_c_886_n 0.00249753f $X=6.77 $Y=1.325
+ $X2=0 $Y2=0
cc_459 N_A_724_21#_c_627_n N_A_1313_47#_c_886_n 0.0159717f $X=6.9 $Y=0.73 $X2=0
+ $Y2=0
cc_460 N_A_724_21#_c_637_n N_A_1313_47#_M1002_g 0.00638756f $X=6.77 $Y=1.62
+ $X2=0 $Y2=0
cc_461 N_A_724_21#_c_639_n N_A_1313_47#_M1002_g 0.0124781f $X=6.9 $Y=1.695 $X2=0
+ $Y2=0
cc_462 N_A_724_21#_c_626_n N_A_1313_47#_c_888_n 0.0132452f $X=6.77 $Y=1.325
+ $X2=0 $Y2=0
cc_463 N_A_724_21#_c_623_n N_A_1313_47#_c_892_n 0.00450382f $X=5.95 $Y=0.995
+ $X2=0 $Y2=0
cc_464 N_A_724_21#_c_626_n N_A_1313_47#_c_892_n 0.0140183f $X=6.77 $Y=1.325
+ $X2=0 $Y2=0
cc_465 N_A_724_21#_c_627_n N_A_1313_47#_c_892_n 0.00963175f $X=6.9 $Y=0.73 $X2=0
+ $Y2=0
cc_466 N_A_724_21#_M1026_g N_A_1313_47#_c_897_n 0.00512189f $X=5.95 $Y=1.985
+ $X2=0 $Y2=0
cc_467 N_A_724_21#_c_637_n N_A_1313_47#_c_897_n 0.0102214f $X=6.77 $Y=1.62 $X2=0
+ $Y2=0
cc_468 N_A_724_21#_c_638_n N_A_1313_47#_c_897_n 0.00975787f $X=6.9 $Y=1.77 $X2=0
+ $Y2=0
cc_469 N_A_724_21#_c_639_n N_A_1313_47#_c_897_n 0.0102619f $X=6.9 $Y=1.695 $X2=0
+ $Y2=0
cc_470 N_A_724_21#_c_626_n N_A_1313_47#_c_893_n 0.00562989f $X=6.77 $Y=1.325
+ $X2=0 $Y2=0
cc_471 N_A_724_21#_c_639_n N_A_1313_47#_c_893_n 0.0046403f $X=6.9 $Y=1.695 $X2=0
+ $Y2=0
cc_472 N_A_724_21#_c_624_n N_A_1313_47#_c_913_n 0.0139585f $X=6.695 $Y=1.16
+ $X2=0 $Y2=0
cc_473 N_A_724_21#_c_626_n N_A_1313_47#_c_913_n 0.00895211f $X=6.77 $Y=1.325
+ $X2=0 $Y2=0
cc_474 N_A_724_21#_c_640_n N_VPWR_M1004_s 0.0064585f $X=4.76 $Y=1.68 $X2=0 $Y2=0
cc_475 N_A_724_21#_c_671_p N_VPWR_M1016_d 0.00411552f $X=5.31 $Y=1.58 $X2=0
+ $Y2=0
cc_476 N_A_724_21#_M1007_g N_VPWR_c_966_n 0.00279634f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_477 N_A_724_21#_c_671_p N_VPWR_c_966_n 0.0138527f $X=5.31 $Y=1.58 $X2=0 $Y2=0
cc_478 N_A_724_21#_M1026_g N_VPWR_c_967_n 0.00675978f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_479 N_A_724_21#_c_624_n N_VPWR_c_967_n 0.001594f $X=6.695 $Y=1.16 $X2=0 $Y2=0
cc_480 N_A_724_21#_c_638_n N_VPWR_c_967_n 0.00331619f $X=6.9 $Y=1.77 $X2=0 $Y2=0
cc_481 N_A_724_21#_c_638_n N_VPWR_c_968_n 0.00537515f $X=6.9 $Y=1.77 $X2=0 $Y2=0
cc_482 N_A_724_21#_c_709_p N_VPWR_c_971_n 0.00955594f $X=4.845 $Y=2.27 $X2=0
+ $Y2=0
cc_483 N_A_724_21#_M1007_g N_VPWR_c_975_n 0.00585385f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_484 N_A_724_21#_M1026_g N_VPWR_c_975_n 0.00526178f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A_724_21#_c_638_n N_VPWR_c_976_n 0.00541359f $X=6.9 $Y=1.77 $X2=0 $Y2=0
cc_486 N_A_724_21#_M1009_g N_VPWR_c_980_n 0.00541489f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_487 N_A_724_21#_M1009_g N_VPWR_c_981_n 0.00483063f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_488 N_A_724_21#_c_640_n N_VPWR_c_981_n 0.0394174f $X=4.76 $Y=1.68 $X2=0 $Y2=0
cc_489 N_A_724_21#_c_641_n N_VPWR_c_981_n 0.00547013f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_490 N_A_724_21#_M1004_d N_VPWR_c_963_n 0.00428563f $X=4.71 $Y=1.485 $X2=0
+ $Y2=0
cc_491 N_A_724_21#_M1009_g N_VPWR_c_963_n 0.0106954f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_492 N_A_724_21#_M1007_g N_VPWR_c_963_n 0.0107033f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_724_21#_M1026_g N_VPWR_c_963_n 0.0106219f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A_724_21#_c_638_n N_VPWR_c_963_n 0.0110094f $X=6.9 $Y=1.77 $X2=0 $Y2=0
cc_495 N_A_724_21#_c_640_n N_VPWR_c_963_n 0.00827674f $X=4.76 $Y=1.68 $X2=0
+ $Y2=0
cc_496 N_A_724_21#_c_641_n N_VPWR_c_963_n 0.00109376f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_497 N_A_724_21#_c_709_p N_VPWR_c_963_n 0.00637538f $X=4.845 $Y=2.27 $X2=0
+ $Y2=0
cc_498 N_A_724_21#_c_622_n N_Q_c_1096_n 0.00568165f $X=5.475 $Y=0.995 $X2=0
+ $Y2=0
cc_499 N_A_724_21#_c_623_n N_Q_c_1096_n 0.0192656f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_500 N_A_724_21#_c_624_n N_Q_c_1096_n 0.0241513f $X=6.695 $Y=1.16 $X2=0 $Y2=0
cc_501 N_A_724_21#_c_625_n N_Q_c_1096_n 0.0183105f $X=6.025 $Y=1.16 $X2=0 $Y2=0
cc_502 N_A_724_21#_c_626_n N_Q_c_1096_n 3.59924e-19 $X=6.77 $Y=1.325 $X2=0 $Y2=0
cc_503 N_A_724_21#_c_649_p N_Q_c_1096_n 0.0140495f $X=5.31 $Y=0.74 $X2=0 $Y2=0
cc_504 N_A_724_21#_c_628_n N_Q_c_1096_n 0.0258372f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_505 N_A_724_21#_c_629_n N_Q_c_1096_n 0.00849233f $X=5.465 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_724_21#_M1007_g N_Q_c_1098_n 0.00112899f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_507 N_A_724_21#_M1026_g N_Q_c_1098_n 0.00533048f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_508 N_A_724_21#_c_642_n N_Q_c_1098_n 0.00772738f $X=5.395 $Y=1.495 $X2=0
+ $Y2=0
cc_509 N_A_724_21#_M1007_g N_Q_c_1110_n 0.00845677f $X=5.475 $Y=1.985 $X2=0
+ $Y2=0
cc_510 N_A_724_21#_M1026_g N_Q_c_1110_n 0.00886344f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_511 N_A_724_21#_c_625_n N_Q_c_1110_n 0.00402417f $X=6.025 $Y=1.16 $X2=0 $Y2=0
cc_512 N_A_724_21#_c_671_p N_Q_c_1110_n 0.013948f $X=5.31 $Y=1.58 $X2=0 $Y2=0
cc_513 N_A_724_21#_M1026_g N_Q_c_1114_n 0.0125087f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_514 N_A_724_21#_c_649_p N_VGND_M1008_d 0.00398929f $X=5.31 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_724_21#_c_629_n N_VGND_M1008_d 6.88945e-19 $X=5.465 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_A_724_21#_M1020_g N_VGND_c_1161_n 0.018542f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_517 N_A_724_21#_c_655_p N_VGND_c_1161_n 0.0233849f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_518 N_A_724_21#_c_622_n N_VGND_c_1162_n 0.0113761f $X=5.475 $Y=0.995 $X2=0
+ $Y2=0
cc_519 N_A_724_21#_c_623_n N_VGND_c_1162_n 0.00103437f $X=5.95 $Y=0.995 $X2=0
+ $Y2=0
cc_520 N_A_724_21#_c_649_p N_VGND_c_1162_n 0.0204969f $X=5.31 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_724_21#_c_655_p N_VGND_c_1162_n 0.0022543f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_522 N_A_724_21#_c_623_n N_VGND_c_1163_n 0.0050871f $X=5.95 $Y=0.995 $X2=0
+ $Y2=0
cc_523 N_A_724_21#_c_624_n N_VGND_c_1163_n 0.00138822f $X=6.695 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_A_724_21#_c_627_n N_VGND_c_1163_n 0.00226455f $X=6.9 $Y=0.73 $X2=0
+ $Y2=0
cc_525 N_A_724_21#_c_627_n N_VGND_c_1164_n 0.0016211f $X=6.9 $Y=0.73 $X2=0 $Y2=0
cc_526 N_A_724_21#_M1020_g N_VGND_c_1169_n 0.0046653f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_527 N_A_724_21#_c_649_p N_VGND_c_1170_n 0.00787618f $X=5.31 $Y=0.74 $X2=0
+ $Y2=0
cc_528 N_A_724_21#_c_655_p N_VGND_c_1170_n 0.00639536f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_529 N_A_724_21#_c_622_n N_VGND_c_1171_n 0.00271402f $X=5.475 $Y=0.995 $X2=0
+ $Y2=0
cc_530 N_A_724_21#_c_623_n N_VGND_c_1171_n 0.00471997f $X=5.95 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_724_21#_c_626_n N_VGND_c_1172_n 2.96334e-19 $X=6.77 $Y=1.325 $X2=0
+ $Y2=0
cc_532 N_A_724_21#_c_627_n N_VGND_c_1172_n 0.00541359f $X=6.9 $Y=0.73 $X2=0
+ $Y2=0
cc_533 N_A_724_21#_M1012_s N_VGND_c_1180_n 0.00370868f $X=4.3 $Y=0.235 $X2=0
+ $Y2=0
cc_534 N_A_724_21#_M1020_g N_VGND_c_1180_n 0.00813035f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_535 N_A_724_21#_c_622_n N_VGND_c_1180_n 0.00511345f $X=5.475 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_A_724_21#_c_623_n N_VGND_c_1180_n 0.00874256f $X=5.95 $Y=0.995 $X2=0
+ $Y2=0
cc_537 N_A_724_21#_c_627_n N_VGND_c_1180_n 0.0110742f $X=6.9 $Y=0.73 $X2=0 $Y2=0
cc_538 N_A_724_21#_c_649_p N_VGND_c_1180_n 0.0154165f $X=5.31 $Y=0.74 $X2=0
+ $Y2=0
cc_539 N_A_724_21#_c_655_p N_VGND_c_1180_n 0.00751733f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_540 N_A_724_21#_c_649_p A_942_47# 0.00441372f $X=5.31 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_541 N_A_561_413#_c_768_n N_RESET_B_c_849_n 0.0427304f $X=4.635 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_542 N_A_561_413#_M1004_g N_RESET_B_M1016_g 0.0236754f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_543 N_A_561_413#_c_770_n N_RESET_B_c_850_n 0.0214963f $X=4.635 $Y=1.16 $X2=0
+ $Y2=0
cc_544 N_A_561_413#_c_769_n N_RESET_B_c_851_n 0.011692f $X=4.56 $Y=1.16 $X2=0
+ $Y2=0
cc_545 N_A_561_413#_c_770_n N_RESET_B_c_851_n 0.0118703f $X=4.635 $Y=1.16 $X2=0
+ $Y2=0
cc_546 N_A_561_413#_c_773_n N_RESET_B_c_851_n 0.0254258f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_547 N_A_561_413#_c_782_n N_VPWR_c_965_n 0.00489615f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_548 N_A_561_413#_M1004_g N_VPWR_c_966_n 6.7327e-19 $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_549 N_A_561_413#_M1004_g N_VPWR_c_971_n 0.0046653f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_550 N_A_561_413#_c_782_n N_VPWR_c_980_n 0.0343719f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_551 N_A_561_413#_M1004_g N_VPWR_c_981_n 0.0101248f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_552 N_A_561_413#_M1001_d N_VPWR_c_963_n 0.00699187f $X=2.805 $Y=2.065 $X2=0
+ $Y2=0
cc_553 N_A_561_413#_M1004_g N_VPWR_c_963_n 0.00443606f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_554 N_A_561_413#_c_782_n N_VPWR_c_963_n 0.0265731f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_555 N_A_561_413#_c_782_n A_682_413# 0.00145479f $X=3.48 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_556 N_A_561_413#_c_777_n A_682_413# 0.00208506f $X=3.565 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_557 N_A_561_413#_c_779_n N_VGND_c_1160_n 0.00209539f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_558 N_A_561_413#_c_768_n N_VGND_c_1161_n 0.00697233f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_559 N_A_561_413#_c_769_n N_VGND_c_1161_n 0.00207331f $X=4.56 $Y=1.16 $X2=0
+ $Y2=0
cc_560 N_A_561_413#_c_779_n N_VGND_c_1161_n 0.01074f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_561 N_A_561_413#_c_771_n N_VGND_c_1161_n 0.0166369f $X=3.415 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_A_561_413#_c_773_n N_VGND_c_1161_n 0.0283975f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_563 N_A_561_413#_c_768_n N_VGND_c_1162_n 0.00214771f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_564 N_A_561_413#_c_779_n N_VGND_c_1169_n 0.0221606f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_565 N_A_561_413#_c_768_n N_VGND_c_1170_n 0.00428022f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_566 N_A_561_413#_M1019_d N_VGND_c_1180_n 0.00237979f $X=2.865 $Y=0.235 $X2=0
+ $Y2=0
cc_567 N_A_561_413#_c_768_n N_VGND_c_1180_n 0.00733083f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_568 N_A_561_413#_c_779_n N_VGND_c_1180_n 0.0222941f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_569 N_A_561_413#_c_779_n A_659_47# 0.00369541f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_570 N_A_561_413#_c_771_n A_659_47# 0.00128174f $X=3.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_571 N_RESET_B_M1016_g N_VPWR_c_966_n 0.0106738f $X=5.055 $Y=1.985 $X2=0 $Y2=0
cc_572 N_RESET_B_M1016_g N_VPWR_c_971_n 0.0046653f $X=5.055 $Y=1.985 $X2=0 $Y2=0
cc_573 N_RESET_B_M1016_g N_VPWR_c_981_n 6.14765e-19 $X=5.055 $Y=1.985 $X2=0
+ $Y2=0
cc_574 N_RESET_B_M1016_g N_VPWR_c_963_n 0.00799591f $X=5.055 $Y=1.985 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_849_n N_VGND_c_1162_n 0.00988605f $X=5.055 $Y=0.995 $X2=0
+ $Y2=0
cc_576 N_RESET_B_c_849_n N_VGND_c_1170_n 0.00341689f $X=5.055 $Y=0.995 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_849_n N_VGND_c_1180_n 0.00405445f $X=5.055 $Y=0.995 $X2=0
+ $Y2=0
cc_578 N_A_1313_47#_c_897_n N_VPWR_c_967_n 0.0520844f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_579 N_A_1313_47#_M1002_g N_VPWR_c_968_n 0.0114729f $X=7.375 $Y=1.985 $X2=0
+ $Y2=0
cc_580 N_A_1313_47#_c_888_n N_VPWR_c_968_n 0.00244466f $X=7.45 $Y=1.16 $X2=0
+ $Y2=0
cc_581 N_A_1313_47#_M1023_g N_VPWR_c_968_n 7.50282e-19 $X=7.8 $Y=1.985 $X2=0
+ $Y2=0
cc_582 N_A_1313_47#_c_897_n N_VPWR_c_968_n 0.0464059f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_583 N_A_1313_47#_c_893_n N_VPWR_c_968_n 0.00959603f $X=7.29 $Y=1.16 $X2=0
+ $Y2=0
cc_584 N_A_1313_47#_M1023_g N_VPWR_c_970_n 0.00313327f $X=7.8 $Y=1.985 $X2=0
+ $Y2=0
cc_585 N_A_1313_47#_c_897_n N_VPWR_c_976_n 0.0210382f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_586 N_A_1313_47#_M1002_g N_VPWR_c_977_n 0.0046653f $X=7.375 $Y=1.985 $X2=0
+ $Y2=0
cc_587 N_A_1313_47#_M1023_g N_VPWR_c_977_n 0.00541359f $X=7.8 $Y=1.985 $X2=0
+ $Y2=0
cc_588 N_A_1313_47#_M1010_s N_VPWR_c_963_n 0.00209319f $X=6.565 $Y=1.845 $X2=0
+ $Y2=0
cc_589 N_A_1313_47#_M1002_g N_VPWR_c_963_n 0.00798142f $X=7.375 $Y=1.985 $X2=0
+ $Y2=0
cc_590 N_A_1313_47#_M1023_g N_VPWR_c_963_n 0.0105179f $X=7.8 $Y=1.985 $X2=0
+ $Y2=0
cc_591 N_A_1313_47#_c_897_n N_VPWR_c_963_n 0.0124268f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_592 N_A_1313_47#_c_892_n N_Q_c_1096_n 0.0202336f $X=6.69 $Y=0.51 $X2=0 $Y2=0
cc_593 N_A_1313_47#_c_913_n N_Q_c_1096_n 0.0275465f $X=6.69 $Y=1.16 $X2=0 $Y2=0
cc_594 N_A_1313_47#_c_897_n N_Q_c_1098_n 0.0107084f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_595 N_A_1313_47#_c_897_n N_Q_c_1114_n 0.00503216f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_596 N_A_1313_47#_c_886_n N_Q_N_c_1130_n 0.00421369f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_597 N_A_1313_47#_c_887_n N_Q_N_c_1130_n 0.00306399f $X=7.725 $Y=1.16 $X2=0
+ $Y2=0
cc_598 N_A_1313_47#_M1027_g N_Q_N_c_1130_n 0.00803505f $X=7.8 $Y=0.56 $X2=0
+ $Y2=0
cc_599 N_A_1313_47#_c_891_n N_Q_N_c_1130_n 0.00120998f $X=7.8 $Y=1.16 $X2=0
+ $Y2=0
cc_600 N_A_1313_47#_c_893_n N_Q_N_c_1130_n 0.00463694f $X=7.29 $Y=1.16 $X2=0
+ $Y2=0
cc_601 N_A_1313_47#_M1027_g N_Q_N_c_1139_n 0.00202845f $X=7.8 $Y=0.56 $X2=0
+ $Y2=0
cc_602 N_A_1313_47#_M1002_g N_Q_N_c_1132_n 9.04394e-19 $X=7.375 $Y=1.985 $X2=0
+ $Y2=0
cc_603 N_A_1313_47#_c_887_n N_Q_N_c_1132_n 0.00976675f $X=7.725 $Y=1.16 $X2=0
+ $Y2=0
cc_604 N_A_1313_47#_c_888_n N_Q_N_c_1132_n 0.00309314f $X=7.45 $Y=1.16 $X2=0
+ $Y2=0
cc_605 N_A_1313_47#_M1023_g N_Q_N_c_1132_n 0.0104283f $X=7.8 $Y=1.985 $X2=0
+ $Y2=0
cc_606 N_A_1313_47#_c_891_n N_Q_N_c_1132_n 6.77984e-19 $X=7.8 $Y=1.16 $X2=0
+ $Y2=0
cc_607 N_A_1313_47#_c_897_n N_Q_N_c_1132_n 0.00268711f $X=6.69 $Y=2 $X2=0 $Y2=0
cc_608 N_A_1313_47#_c_893_n N_Q_N_c_1132_n 0.022823f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_609 N_A_1313_47#_M1027_g Q_N 0.0061015f $X=7.8 $Y=0.56 $X2=0 $Y2=0
cc_610 N_A_1313_47#_M1023_g Q_N 0.0115188f $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_611 N_A_1313_47#_M1023_g Q_N 0.00643843f $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_612 N_A_1313_47#_c_891_n Q_N 0.0131132f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_613 N_A_1313_47#_c_892_n N_VGND_c_1163_n 0.0237866f $X=6.69 $Y=0.51 $X2=0
+ $Y2=0
cc_614 N_A_1313_47#_c_886_n N_VGND_c_1164_n 0.00789409f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_615 N_A_1313_47#_c_888_n N_VGND_c_1164_n 0.00255976f $X=7.45 $Y=1.16 $X2=0
+ $Y2=0
cc_616 N_A_1313_47#_M1027_g N_VGND_c_1164_n 6.51904e-19 $X=7.8 $Y=0.56 $X2=0
+ $Y2=0
cc_617 N_A_1313_47#_c_893_n N_VGND_c_1164_n 0.0107987f $X=7.29 $Y=1.16 $X2=0
+ $Y2=0
cc_618 N_A_1313_47#_M1027_g N_VGND_c_1166_n 0.00313327f $X=7.8 $Y=0.56 $X2=0
+ $Y2=0
cc_619 N_A_1313_47#_c_892_n N_VGND_c_1172_n 0.0210709f $X=6.69 $Y=0.51 $X2=0
+ $Y2=0
cc_620 N_A_1313_47#_c_886_n N_VGND_c_1173_n 0.0046653f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_621 N_A_1313_47#_M1027_g N_VGND_c_1173_n 0.00541359f $X=7.8 $Y=0.56 $X2=0
+ $Y2=0
cc_622 N_A_1313_47#_M1021_s N_VGND_c_1180_n 0.00210122f $X=6.565 $Y=0.235 $X2=0
+ $Y2=0
cc_623 N_A_1313_47#_c_886_n N_VGND_c_1180_n 0.00798142f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_624 N_A_1313_47#_M1027_g N_VGND_c_1180_n 0.0105179f $X=7.8 $Y=0.56 $X2=0
+ $Y2=0
cc_625 N_A_1313_47#_c_892_n N_VGND_c_1180_n 0.0124992f $X=6.69 $Y=0.51 $X2=0
+ $Y2=0
cc_626 N_VPWR_c_963_n A_465_369# 0.00373974f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_627 N_VPWR_c_963_n A_682_413# 0.00170472f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_628 N_VPWR_c_963_n N_Q_M1007_d 0.00606522f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_629 N_VPWR_c_967_n N_Q_c_1096_n 0.00981369f $X=6.17 $Y=2 $X2=0 $Y2=0
cc_630 N_VPWR_c_967_n N_Q_c_1114_n 0.0477523f $X=6.17 $Y=2 $X2=0 $Y2=0
cc_631 N_VPWR_c_975_n N_Q_c_1114_n 0.0163923f $X=6.085 $Y=2.72 $X2=0 $Y2=0
cc_632 N_VPWR_c_963_n N_Q_c_1114_n 0.00987779f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_633 N_VPWR_c_963_n N_Q_N_M1002_d 0.00397872f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_634 N_VPWR_c_977_n Q_N 0.0155342f $X=7.925 $Y=2.72 $X2=0 $Y2=0
cc_635 N_VPWR_c_963_n Q_N 0.00961085f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_636 N_VPWR_c_970_n Q_N 0.0227331f $X=8.01 $Y=1.66 $X2=0 $Y2=0
cc_637 N_Q_c_1096_n N_VGND_M1025_d 0.00578085f $X=5.882 $Y=1.325 $X2=0 $Y2=0
cc_638 N_Q_c_1096_n N_VGND_c_1162_n 0.00542068f $X=5.882 $Y=1.325 $X2=0 $Y2=0
cc_639 N_Q_c_1096_n N_VGND_c_1163_n 0.0237291f $X=5.882 $Y=1.325 $X2=0 $Y2=0
cc_640 N_Q_c_1096_n N_VGND_c_1171_n 0.00887161f $X=5.882 $Y=1.325 $X2=0 $Y2=0
cc_641 N_Q_M1018_s N_VGND_c_1180_n 0.0062991f $X=5.55 $Y=0.235 $X2=0 $Y2=0
cc_642 N_Q_c_1096_n N_VGND_c_1180_n 0.0104396f $X=5.882 $Y=1.325 $X2=0 $Y2=0
cc_643 Q_N N_VGND_c_1166_n 0.0227331f $X=7.985 $Y=1.105 $X2=0 $Y2=0
cc_644 Q_N N_VGND_c_1173_n 0.0155f $X=7.525 $Y=0.425 $X2=0 $Y2=0
cc_645 N_Q_N_M1003_d N_VGND_c_1180_n 0.00397872f $X=7.45 $Y=0.235 $X2=0 $Y2=0
cc_646 Q_N N_VGND_c_1180_n 0.0096031f $X=7.525 $Y=0.425 $X2=0 $Y2=0
cc_647 N_VGND_c_1180_n A_465_47# 0.0139156f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_648 N_VGND_c_1180_n A_659_47# 0.00687059f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_649 N_VGND_c_1180_n A_942_47# 0.00323135f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24

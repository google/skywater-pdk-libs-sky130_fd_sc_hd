* File: sky130_fd_sc_hd__xnor2_1.spice.SKY130_FD_SC_HD__XNOR2_1.pxi
* Created: Thu Aug 27 14:48:57 2020
* 
x_PM_SKY130_FD_SC_HD__XNOR2_1%B N_B_M1008_g N_B_M1005_g N_B_M1004_g N_B_M1006_g
+ N_B_c_58_n N_B_c_59_n N_B_c_60_n N_B_c_61_n N_B_c_70_n B N_B_c_62_n N_B_c_63_n
+ N_B_c_64_n N_B_c_65_n B PM_SKY130_FD_SC_HD__XNOR2_1%B
x_PM_SKY130_FD_SC_HD__XNOR2_1%A N_A_c_149_n N_A_M1007_g N_A_M1003_g N_A_c_150_n
+ N_A_M1001_g N_A_M1002_g A N_A_c_161_n N_A_c_151_n
+ PM_SKY130_FD_SC_HD__XNOR2_1%A
x_PM_SKY130_FD_SC_HD__XNOR2_1%A_47_47# N_A_47_47#_M1005_s N_A_47_47#_M1008_d
+ N_A_47_47#_M1000_g N_A_47_47#_c_198_n N_A_47_47#_M1009_g N_A_47_47#_c_199_n
+ N_A_47_47#_c_219_n N_A_47_47#_c_205_n N_A_47_47#_c_222_n N_A_47_47#_c_223_n
+ N_A_47_47#_c_226_n N_A_47_47#_c_206_n N_A_47_47#_c_207_n N_A_47_47#_c_200_n
+ N_A_47_47#_c_201_n N_A_47_47#_c_202_n N_A_47_47#_c_244_n
+ PM_SKY130_FD_SC_HD__XNOR2_1%A_47_47#
x_PM_SKY130_FD_SC_HD__XNOR2_1%VPWR N_VPWR_M1008_s N_VPWR_M1003_d N_VPWR_M1000_d
+ N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n VPWR
+ N_VPWR_c_308_n N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_303_n
+ PM_SKY130_FD_SC_HD__XNOR2_1%VPWR
x_PM_SKY130_FD_SC_HD__XNOR2_1%Y N_Y_M1009_d N_Y_M1004_d N_Y_c_359_n N_Y_c_356_n
+ N_Y_c_371_n N_Y_c_360_n N_Y_c_357_n Y N_Y_c_379_n
+ PM_SKY130_FD_SC_HD__XNOR2_1%Y
x_PM_SKY130_FD_SC_HD__XNOR2_1%VGND N_VGND_M1007_d N_VGND_M1006_s N_VGND_c_398_n
+ N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n VGND N_VGND_c_402_n
+ N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n PM_SKY130_FD_SC_HD__XNOR2_1%VGND
x_PM_SKY130_FD_SC_HD__XNOR2_1%A_285_47# N_A_285_47#_M1001_d N_A_285_47#_M1006_d
+ N_A_285_47#_c_443_n N_A_285_47#_c_444_n N_A_285_47#_c_445_n
+ N_A_285_47#_c_462_n PM_SKY130_FD_SC_HD__XNOR2_1%A_285_47#
cc_1 VNB N_B_c_58_n 5.704e-19 $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.445
cc_2 VNB N_B_c_59_n 7.48283e-19 $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.16
cc_3 VNB N_B_c_60_n 0.00485988f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=1.16
cc_4 VNB N_B_c_61_n 0.0200129f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=1.16
cc_5 VNB N_B_c_62_n 0.0223964f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_6 VNB N_B_c_63_n 0.00413128f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_7 VNB N_B_c_64_n 0.0190329f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_8 VNB N_B_c_65_n 0.0209219f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=0.995
cc_9 VNB N_A_c_149_n 0.0156421f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.325
cc_10 VNB N_A_c_150_n 0.0215746f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.325
cc_11 VNB N_A_c_151_n 0.0560839f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_12 VNB N_A_47_47#_c_198_n 0.0195351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_47_47#_c_199_n 0.0222048f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.245
cc_14 VNB N_A_47_47#_c_200_n 4.4441e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_15 VNB N_A_47_47#_c_201_n 0.024826f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=1.16
cc_16 VNB N_A_47_47#_c_202_n 0.0253194f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.53
cc_17 VNB N_VPWR_c_303_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_356_n 0.0219408f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.985
cc_19 VNB N_Y_c_357_n 0.0191091f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=1.16
cc_20 VNB N_VGND_c_398_n 0.00576786f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.985
cc_21 VNB N_VGND_c_399_n 0.00534711f $X=-0.19 $Y=-0.24 $X2=2.29 $Y2=0.56
cc_22 VNB N_VGND_c_400_n 0.0315674f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.445
cc_23 VNB N_VGND_c_401_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.16
cc_24 VNB N_VGND_c_402_n 0.0174177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_403_n 0.0266107f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_26 VNB N_VGND_c_404_n 0.183838f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=1.16
cc_27 VNB N_VGND_c_405_n 0.00545658f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.53
cc_28 VNB N_A_285_47#_c_443_n 0.00569684f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.985
cc_29 VNB N_A_285_47#_c_444_n 0.00815854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_285_47#_c_445_n 0.00235789f $X=-0.19 $Y=-0.24 $X2=2.29 $Y2=0.995
cc_31 VPB N_B_M1008_g 0.0223541f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_32 VPB N_B_M1004_g 0.0186332f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_33 VPB N_B_c_58_n 0.00122864f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.445
cc_34 VPB N_B_c_61_n 0.00425883f $X=-0.19 $Y=1.305 $X2=2.23 $Y2=1.16
cc_35 VPB N_B_c_70_n 0.0124667f $X=-0.19 $Y=1.305 $X2=1.795 $Y2=1.53
cc_36 VPB B 3.66229e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_37 VPB N_B_c_62_n 0.00472483f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_38 VPB N_B_c_63_n 0.00251016f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_39 VPB N_A_M1003_g 0.0252636f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=0.56
cc_40 VPB N_A_M1002_g 0.0238287f $X=-0.19 $Y=1.305 $X2=2.29 $Y2=0.56
cc_41 VPB N_A_c_151_n 0.0161566f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_42 VPB N_A_47_47#_M1000_g 0.0235501f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_43 VPB N_A_47_47#_c_199_n 0.0191394f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.245
cc_44 VPB N_A_47_47#_c_205_n 0.00766781f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.16
cc_45 VPB N_A_47_47#_c_206_n 0.00410862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_47_47#_c_207_n 3.56375e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_47 VPB N_A_47_47#_c_200_n 8.17603e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_48 VPB N_A_47_47#_c_201_n 0.00482079f $X=-0.19 $Y=1.305 $X2=2.23 $Y2=1.16
cc_49 VPB N_VPWR_c_304_n 0.0106536f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_50 VPB N_VPWR_c_305_n 0.019142f $X=-0.19 $Y=1.305 $X2=2.29 $Y2=0.995
cc_51 VPB N_VPWR_c_306_n 0.0112167f $X=-0.19 $Y=1.305 $X2=2.29 $Y2=0.56
cc_52 VPB N_VPWR_c_307_n 0.0192743f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.445
cc_53 VPB N_VPWR_c_308_n 0.0333321f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_309_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.53
cc_55 VPB N_VPWR_c_310_n 0.018848f $X=-0.19 $Y=1.305 $X2=0.547 $Y2=1.53
cc_56 VPB N_VPWR_c_303_n 0.0424524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_Y_c_356_n 0.0271223f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_58 N_B_c_64_n N_A_c_149_n 0.037632f $X=0.51 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_59 N_B_M1008_g N_A_M1003_g 0.0272756f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_60 N_B_c_70_n N_A_M1003_g 0.0147159f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_61 N_B_M1004_g N_A_M1002_g 0.0509111f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_62 N_B_c_58_n N_A_M1002_g 0.00582672f $X=1.88 $Y=1.445 $X2=0 $Y2=0
cc_63 N_B_c_70_n N_A_M1002_g 0.0105003f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_64 N_B_c_58_n N_A_c_161_n 0.00217909f $X=1.88 $Y=1.445 $X2=0 $Y2=0
cc_65 N_B_c_59_n N_A_c_161_n 0.0141956f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_66 N_B_c_70_n N_A_c_161_n 0.0500238f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_67 N_B_c_62_n N_A_c_161_n 2.12332e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B_c_63_n N_A_c_161_n 0.0118218f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B_c_58_n N_A_c_151_n 0.00359482f $X=1.88 $Y=1.445 $X2=0 $Y2=0
cc_70 N_B_c_59_n N_A_c_151_n 0.00604726f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B_c_61_n N_A_c_151_n 0.0509111f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B_c_70_n N_A_c_151_n 0.0141615f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_73 N_B_c_62_n N_A_c_151_n 0.037632f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_74 N_B_c_63_n N_A_c_151_n 0.00688395f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B_c_70_n N_A_47_47#_M1008_d 0.00135003f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_76 B N_A_47_47#_M1008_d 2.97948e-19 $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_77 N_B_M1004_g N_A_47_47#_M1000_g 0.0327045f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B_c_65_n N_A_47_47#_c_198_n 0.0235629f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B_M1008_g N_A_47_47#_c_199_n 0.00776159f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_80 B N_A_47_47#_c_199_n 0.00807294f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_81 N_B_c_62_n N_A_47_47#_c_199_n 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B_c_63_n N_A_47_47#_c_199_n 0.0334999f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B_c_64_n N_A_47_47#_c_199_n 0.00442653f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B_M1008_g N_A_47_47#_c_219_n 0.00961786f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_85 B N_A_47_47#_c_219_n 0.00903642f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_86 N_B_c_62_n N_A_47_47#_c_219_n 7.98519e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B_M1008_g N_A_47_47#_c_222_n 0.0113712f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_88 N_B_M1004_g N_A_47_47#_c_223_n 0.00950123f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B_c_60_n N_A_47_47#_c_223_n 0.00434139f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_c_70_n N_A_47_47#_c_223_n 0.0653957f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_A_47_47#_c_226_n 0.00550752f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B_c_70_n N_A_47_47#_c_226_n 0.00233386f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_93 N_B_c_60_n N_A_47_47#_c_206_n 0.00651241f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B_c_61_n N_A_47_47#_c_206_n 0.00173414f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B_M1004_g N_A_47_47#_c_207_n 0.00652275f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_96 N_B_c_58_n N_A_47_47#_c_207_n 0.00235384f $X=1.88 $Y=1.445 $X2=0 $Y2=0
cc_97 N_B_c_60_n N_A_47_47#_c_207_n 0.0129647f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_98 N_B_c_61_n N_A_47_47#_c_207_n 0.00178505f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B_c_70_n N_A_47_47#_c_207_n 0.0122795f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_100 N_B_M1004_g N_A_47_47#_c_200_n 3.22764e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B_c_58_n N_A_47_47#_c_200_n 0.00425475f $X=1.88 $Y=1.445 $X2=0 $Y2=0
cc_102 N_B_c_60_n N_A_47_47#_c_200_n 0.0107022f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_c_61_n N_A_47_47#_c_200_n 0.00101515f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B_c_60_n N_A_47_47#_c_201_n 0.00112113f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B_c_61_n N_A_47_47#_c_201_n 0.0208698f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B_c_62_n N_A_47_47#_c_202_n 0.00255604f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B_c_63_n N_A_47_47#_c_202_n 0.0078258f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B_c_64_n N_A_47_47#_c_202_n 0.0114653f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_M1008_g N_A_47_47#_c_244_n 8.68888e-19 $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B_c_70_n N_A_47_47#_c_244_n 0.0126206f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_111 B N_A_47_47#_c_244_n 0.00498744f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_112 N_B_c_70_n N_VPWR_M1003_d 0.00920603f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_113 N_B_M1008_g N_VPWR_c_305_n 0.00362074f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B_M1004_g N_VPWR_c_308_n 0.00585385f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B_M1008_g N_VPWR_c_309_n 0.00541359f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B_M1008_g N_VPWR_c_303_n 0.00681316f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B_M1004_g N_VPWR_c_303_n 0.00623606f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B_c_70_n A_377_297# 0.00136153f $X=1.795 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_119 N_B_M1004_g N_Y_c_359_n 0.00295401f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B_M1004_g N_Y_c_360_n 7.11336e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B_c_65_n N_VGND_c_399_n 0.00910793f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_64_n N_VGND_c_400_n 0.00505274f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_65_n N_VGND_c_403_n 0.00341574f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_64_n N_VGND_c_404_n 0.00968079f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B_c_65_n N_VGND_c_404_n 0.00405248f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B_c_65_n N_A_285_47#_c_443_n 0.00388209f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_59_n N_A_285_47#_c_444_n 0.0136907f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B_c_60_n N_A_285_47#_c_444_n 0.0286943f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B_c_61_n N_A_285_47#_c_444_n 0.00349202f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_c_70_n N_A_285_47#_c_444_n 0.0020966f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_131 N_B_c_65_n N_A_285_47#_c_444_n 0.0159419f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B_c_70_n N_A_285_47#_c_445_n 0.00373857f $X=1.795 $Y=1.53 $X2=0 $Y2=0
cc_133 N_A_M1003_g N_A_47_47#_c_222_n 0.0113952f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1003_g N_A_47_47#_c_223_n 0.0101664f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1002_g N_A_47_47#_c_223_n 0.013248f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1002_g N_A_47_47#_c_226_n 0.00106399f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_c_149_n N_A_47_47#_c_202_n 0.00162052f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_A_47_47#_c_244_n 8.70118e-19 $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1002_g N_VPWR_c_308_n 0.00585385f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1003_g N_VPWR_c_309_n 0.00541359f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_VPWR_c_310_n 0.00334593f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_VPWR_c_310_n 0.00478724f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1003_g N_VPWR_c_303_n 0.0071463f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1002_g N_VPWR_c_303_n 0.00721936f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_c_149_n N_VGND_c_398_n 0.00314514f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_150_n N_VGND_c_398_n 0.00159991f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_161_n N_VGND_c_398_n 0.0137004f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_c_151_n N_VGND_c_398_n 0.00231083f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_c_150_n N_VGND_c_399_n 0.00150459f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_149_n N_VGND_c_400_n 0.00585385f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_150_n N_VGND_c_402_n 0.00541359f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_149_n N_VGND_c_404_n 0.0104784f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_150_n N_VGND_c_404_n 0.0108276f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_150_n N_A_285_47#_c_443_n 0.0052355f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_151_n N_A_285_47#_c_444_n 0.00493251f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_150_n N_A_285_47#_c_445_n 0.00265987f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_161_n N_A_285_47#_c_445_n 0.018547f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_c_151_n N_A_285_47#_c_445_n 0.00862609f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_47_47#_c_199_n N_VPWR_M1008_s 0.00501491f $X=0.17 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_47_47#_c_219_n N_VPWR_M1008_s 0.00581182f $X=0.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_47_47#_c_205_n N_VPWR_M1008_s 0.00242f $X=0.255 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_47_47#_c_223_n N_VPWR_M1003_d 0.0157189f $X=2.135 $Y=1.87 $X2=0 $Y2=0
cc_163 N_A_47_47#_c_206_n N_VPWR_M1000_d 0.00124088f $X=2.625 $Y=1.5 $X2=0 $Y2=0
cc_164 N_A_47_47#_c_219_n N_VPWR_c_305_n 0.00968766f $X=0.555 $Y=1.87 $X2=0
+ $Y2=0
cc_165 N_A_47_47#_c_205_n N_VPWR_c_305_n 0.0148845f $X=0.255 $Y=1.87 $X2=0 $Y2=0
cc_166 N_A_47_47#_M1000_g N_VPWR_c_307_n 0.0088127f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_47_47#_M1000_g N_VPWR_c_308_n 0.0049461f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_47_47#_c_222_n N_VPWR_c_309_n 0.0189039f $X=0.72 $Y=1.96 $X2=0 $Y2=0
cc_169 N_A_47_47#_c_223_n N_VPWR_c_310_n 0.0484396f $X=2.135 $Y=1.87 $X2=0 $Y2=0
cc_170 N_A_47_47#_M1008_d N_VPWR_c_303_n 0.00215201f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_171 N_A_47_47#_M1000_g N_VPWR_c_303_n 0.00697363f $X=2.65 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_47_47#_c_219_n N_VPWR_c_303_n 0.00576828f $X=0.555 $Y=1.87 $X2=0
+ $Y2=0
cc_173 N_A_47_47#_c_205_n N_VPWR_c_303_n 6.8277e-19 $X=0.255 $Y=1.87 $X2=0 $Y2=0
cc_174 N_A_47_47#_c_222_n N_VPWR_c_303_n 0.0122217f $X=0.72 $Y=1.96 $X2=0 $Y2=0
cc_175 N_A_47_47#_c_223_n N_VPWR_c_303_n 0.0271519f $X=2.135 $Y=1.87 $X2=0 $Y2=0
cc_176 N_A_47_47#_c_223_n A_377_297# 0.00343157f $X=2.135 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_47_47#_c_223_n N_Y_M1004_d 0.00153429f $X=2.135 $Y=1.87 $X2=0 $Y2=0
cc_178 N_A_47_47#_c_226_n N_Y_M1004_d 0.00285214f $X=2.22 $Y=1.785 $X2=0 $Y2=0
cc_179 N_A_47_47#_c_206_n N_Y_M1004_d 0.00363776f $X=2.625 $Y=1.5 $X2=0 $Y2=0
cc_180 N_A_47_47#_M1000_g N_Y_c_359_n 0.00826103f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_47_47#_M1000_g N_Y_c_356_n 0.00526114f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_47_47#_c_198_n N_Y_c_356_n 0.00491405f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_47_47#_c_226_n N_Y_c_356_n 0.00439683f $X=2.22 $Y=1.785 $X2=0 $Y2=0
cc_184 N_A_47_47#_c_206_n N_Y_c_356_n 0.0140129f $X=2.625 $Y=1.5 $X2=0 $Y2=0
cc_185 N_A_47_47#_c_200_n N_Y_c_356_n 0.03034f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_47_47#_c_201_n N_Y_c_356_n 0.00753248f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_47_47#_M1000_g N_Y_c_371_n 0.00360286f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_47_47#_c_223_n N_Y_c_371_n 2.31245e-19 $X=2.135 $Y=1.87 $X2=0 $Y2=0
cc_189 N_A_47_47#_c_206_n N_Y_c_371_n 0.0052308f $X=2.625 $Y=1.5 $X2=0 $Y2=0
cc_190 N_A_47_47#_M1000_g N_Y_c_360_n 0.00371962f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_47_47#_c_223_n N_Y_c_360_n 0.0152933f $X=2.135 $Y=1.87 $X2=0 $Y2=0
cc_192 N_A_47_47#_c_226_n N_Y_c_360_n 0.00239828f $X=2.22 $Y=1.785 $X2=0 $Y2=0
cc_193 N_A_47_47#_c_206_n N_Y_c_360_n 0.00848651f $X=2.625 $Y=1.5 $X2=0 $Y2=0
cc_194 N_A_47_47#_c_201_n N_Y_c_357_n 6.53374e-19 $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_47_47#_M1000_g N_Y_c_379_n 0.00859959f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_47_47#_c_206_n N_Y_c_379_n 0.00711419f $X=2.625 $Y=1.5 $X2=0 $Y2=0
cc_197 N_A_47_47#_c_201_n N_Y_c_379_n 0.00166165f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_47_47#_c_198_n N_VGND_c_399_n 0.00125667f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_47_47#_c_202_n N_VGND_c_400_n 0.0261949f $X=0.36 $Y=0.39 $X2=0 $Y2=0
cc_200 N_A_47_47#_c_198_n N_VGND_c_403_n 0.00571722f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_47_47#_M1005_s N_VGND_c_404_n 0.00210425f $X=0.235 $Y=0.235 $X2=0
+ $Y2=0
cc_202 N_A_47_47#_c_198_n N_VGND_c_404_n 0.0115356f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_47_47#_c_202_n N_VGND_c_404_n 0.0172239f $X=0.36 $Y=0.39 $X2=0 $Y2=0
cc_204 N_A_47_47#_c_198_n N_A_285_47#_c_444_n 0.00290848f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_47_47#_c_206_n N_A_285_47#_c_444_n 0.00613834f $X=2.625 $Y=1.5 $X2=0
+ $Y2=0
cc_206 N_A_47_47#_c_200_n N_A_285_47#_c_444_n 0.00120016f $X=2.71 $Y=1.16 $X2=0
+ $Y2=0
cc_207 N_A_47_47#_c_201_n N_A_285_47#_c_444_n 0.00125943f $X=2.71 $Y=1.16 $X2=0
+ $Y2=0
cc_208 N_A_47_47#_c_198_n N_A_285_47#_c_462_n 0.00761101f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_303_n A_377_297# 0.00285576f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_210 N_VPWR_c_303_n N_Y_M1004_d 0.0030672f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_M1000_d N_Y_c_356_n 0.00780139f $X=2.725 $Y=1.485 $X2=0 $Y2=0
cc_212 N_VPWR_c_306_n N_Y_c_356_n 3.08556e-19 $X=2.965 $Y=2.635 $X2=0 $Y2=0
cc_213 N_VPWR_c_307_n N_Y_c_356_n 0.0130694f $X=2.9 $Y=2.29 $X2=0 $Y2=0
cc_214 N_VPWR_c_303_n N_Y_c_356_n 0.00118299f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_c_307_n N_Y_c_371_n 0.0131484f $X=2.9 $Y=2.29 $X2=0 $Y2=0
cc_216 N_VPWR_c_308_n N_Y_c_371_n 0.0101981f $X=2.815 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_303_n N_Y_c_371_n 0.0122729f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_M1000_d N_Y_c_379_n 0.00833142f $X=2.725 $Y=1.485 $X2=0 $Y2=0
cc_219 N_VPWR_c_307_n N_Y_c_379_n 0.0118674f $X=2.9 $Y=2.29 $X2=0 $Y2=0
cc_220 N_VPWR_c_303_n N_Y_c_379_n 0.00626494f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_221 N_Y_c_357_n N_VGND_c_403_n 0.0134936f $X=2.96 $Y=0.555 $X2=0 $Y2=0
cc_222 N_Y_M1009_d N_VGND_c_404_n 0.00359348f $X=2.785 $Y=0.235 $X2=0 $Y2=0
cc_223 N_Y_c_357_n N_VGND_c_404_n 0.011609f $X=2.96 $Y=0.555 $X2=0 $Y2=0
cc_224 N_Y_c_356_n N_A_285_47#_c_444_n 0.00213471f $X=3.05 $Y=1.755 $X2=0 $Y2=0
cc_225 A_129_47# N_VGND_c_404_n 0.00897657f $X=0.645 $Y=0.235 $X2=2.99 $Y2=0
cc_226 N_VGND_c_404_n N_A_285_47#_M1001_d 0.00209319f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_227 N_VGND_c_404_n N_A_285_47#_M1006_d 0.00235622f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_399_n N_A_285_47#_c_443_n 0.0184009f $X=2.08 $Y=0.39 $X2=0 $Y2=0
cc_229 N_VGND_c_402_n N_A_285_47#_c_443_n 0.0209752f $X=1.895 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_404_n N_A_285_47#_c_443_n 0.0124119f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_M1006_s N_A_285_47#_c_444_n 0.00430809f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_VGND_c_399_n N_A_285_47#_c_444_n 0.0167347f $X=2.08 $Y=0.39 $X2=0 $Y2=0
cc_233 N_VGND_c_402_n N_A_285_47#_c_444_n 0.00252694f $X=1.895 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_403_n N_A_285_47#_c_444_n 0.00235386f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_404_n N_A_285_47#_c_444_n 0.0102478f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_398_n N_A_285_47#_c_445_n 0.00787895f $X=1.14 $Y=0.39 $X2=0
+ $Y2=0
cc_237 N_VGND_c_403_n N_A_285_47#_c_462_n 0.0136708f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_404_n N_A_285_47#_c_462_n 0.00869934f $X=2.99 $Y=0 $X2=0 $Y2=0

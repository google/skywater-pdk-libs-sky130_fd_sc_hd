* File: sky130_fd_sc_hd__o41a_2.spice
* Created: Tue Sep  1 19:26:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o41a_2.pex.spice"
.subckt sky130_fd_sc_hd__o41a_2  VNB VPB B1 A4 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_79_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_79_21#_M1012_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_393_47#_M1002_d N_B1_M1002_g N_A_79_21#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.118625 AS=0.208 PD=1.015 PS=1.94 NRD=8.304 NRS=10.152 M=1
+ R=4.33333 SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A4_M1003_g N_A_393_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.118625 PD=1.005 PS=1.015 NRD=0 NRS=7.38 M=1 R=4.33333
+ SA=75000.8 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1013 N_A_393_47#_M1013_d N_A3_M1013_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.115375 PD=1 PS=1.005 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75001.3
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_393_47#_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.11375 PD=1 PS=1 NRD=2.76 NRS=13.836 M=1 R=4.33333 SA=75001.8
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_393_47#_M1009_d N_A1_M1009_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2665 AS=0.11375 PD=2.12 PS=1 NRD=19.38 NRS=10.152 M=1 R=4.33333
+ SA=75002.3 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_79_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.8 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A_79_21#_M1008_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.305 AS=0.135 PD=1.61 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1005 N_A_79_21#_M1005_d N_B1_M1005_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.3025 AS=0.305 PD=1.605 PS=1.61 NRD=0 NRS=21.3351 M=1 R=6.66667 SA=75001.4
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1006 A_496_297# N_A4_M1006_g N_A_79_21#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1775 AS=0.3025 PD=1.355 PS=1.605 NRD=24.1128 NRS=64.9903 M=1 R=6.66667
+ SA=75002.1 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1007 A_597_297# N_A3_M1007_g A_496_297# VPB PHIGHVT L=0.15 W=1 AD=0.175
+ AS=0.1775 PD=1.35 PS=1.355 NRD=23.6203 NRS=24.1128 M=1 R=6.66667 SA=75002.6
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1011 A_697_297# N_A2_M1011_g A_597_297# VPB PHIGHVT L=0.15 W=1 AD=0.175
+ AS=0.175 PD=1.35 PS=1.35 NRD=23.6203 NRS=23.6203 M=1 R=6.66667 SA=75003.1
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_697_297# VPB PHIGHVT L=0.15 W=1 AD=0.41
+ AS=0.175 PD=2.82 PS=1.35 NRD=20.685 NRS=23.6203 M=1 R=6.66667 SA=75003.6
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__o41a_2.pxi.spice"
*
.ends
*
*

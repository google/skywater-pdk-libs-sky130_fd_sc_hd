* File: sky130_fd_sc_hd__clkinv_16.spice
* Created: Tue Sep  1 19:01:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkinv_16.pex.spice"
.subckt sky130_fd_sc_hd__clkinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75006.8 A=0.063
+ P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75006.4 A=0.063
+ P=1.14 MULT=1
MM1008 N_VGND_M1007_d N_A_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75006 A=0.063
+ P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75005.5 A=0.063
+ P=1.14 MULT=1
MM1016 N_VGND_M1011_d N_A_M1016_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75005.1 A=0.063
+ P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_M1017_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.0588 PD=0.735 PS=0.7 NRD=7.14 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75004.7 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1017_d N_A_M1018_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.09135 PD=0.735 PS=0.855 NRD=2.856 NRS=8.568 M=1 R=2.8
+ SA=75002.8 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_M1021_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.09135 PD=0.7 PS=0.855 NRD=0 NRS=35.712 M=1 R=2.8 SA=75003.4 SB=75003.6
+ A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1021_d N_A_M1023_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.8 SB=75003.2 A=0.063
+ P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_M1024_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.2 SB=75002.8 A=0.063
+ P=1.14 MULT=1
MM1026 N_VGND_M1024_d N_A_M1026_g N_Y_M1026_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.7 SB=75002.3 A=0.063
+ P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_M1032_g N_Y_M1026_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.1 SB=75001.9 A=0.063
+ P=1.14 MULT=1
MM1033 N_VGND_M1032_d N_A_M1033_g N_Y_M1033_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.5 SB=75001.5 A=0.063
+ P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_M1035_g N_Y_M1033_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006 SB=75001.1 A=0.063
+ P=1.14 MULT=1
MM1036 N_VGND_M1035_d N_A_M1036_g N_Y_M1036_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.4 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_M1037_g N_Y_M1036_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.8 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.275
+ AS=0.14 PD=2.55 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75010.3 A=0.15
+ P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75009.8 A=0.15
+ P=2.3 MULT=1
MM1002 N_VPWR_M1001_d N_A_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1 SB=75009.4 A=0.15
+ P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75009 A=0.15
+ P=2.3 MULT=1
MM1005 N_VPWR_M1003_d N_A_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75008.5 A=0.15
+ P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75008.1 A=0.15
+ P=2.3 MULT=1
MM1009 N_VPWR_M1006_d N_A_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8 SB=75007.7 A=0.15
+ P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2 SB=75007.3 A=0.15
+ P=2.3 MULT=1
MM1012 N_VPWR_M1010_d N_A_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6 SB=75006.8 A=0.15
+ P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.1575
+ AS=0.14 PD=1.315 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75006.4
+ A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1013_d N_A_M1014_g N_Y_M1014_s VPB PHIGHVT L=0.15 W=1 AD=0.1575
+ AS=0.2175 PD=1.315 PS=1.435 NRD=2.9353 NRS=25.5903 M=1 R=6.66667 SA=75004.5
+ SB=75005.9 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_Y_M1014_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.2175 PD=1.28 PS=1.435 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75005.1
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1015_d N_A_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75005.5 SB=75004.9
+ A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_Y_M1019_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006 SB=75004.5 A=0.15
+ P=2.3 MULT=1
MM1022 N_VPWR_M1020_d N_A_M1022_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.4 SB=75004.1 A=0.15
+ P=2.3 MULT=1
MM1025 N_VPWR_M1025_d N_A_M1025_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.8 SB=75003.6 A=0.15
+ P=2.3 MULT=1
MM1027 N_VPWR_M1025_d N_A_M1027_g N_Y_M1027_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.3 SB=75003.2 A=0.15
+ P=2.3 MULT=1
MM1028 N_VPWR_M1028_d N_A_M1028_g N_Y_M1027_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.7 SB=75002.8 A=0.15
+ P=2.3 MULT=1
MM1029 N_VPWR_M1028_d N_A_M1029_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.1 SB=75002.3 A=0.15
+ P=2.3 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.6 SB=75001.9 A=0.15
+ P=2.3 MULT=1
MM1031 N_VPWR_M1030_d N_A_M1031_g N_Y_M1031_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75009 SB=75001.5 A=0.15
+ P=2.3 MULT=1
MM1034 N_VPWR_M1034_d N_A_M1034_g N_Y_M1031_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.4 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1038 N_VPWR_M1034_d N_A_M1038_g N_Y_M1038_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.8 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1039 N_VPWR_M1039_d N_A_M1039_g N_Y_M1038_s VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75010.3 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=18.3291 P=26.05
*
.include "sky130_fd_sc_hd__clkinv_16.pxi.spice"
*
.ends
*
*

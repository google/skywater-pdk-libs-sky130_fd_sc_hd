* File: sky130_fd_sc_hd__lpflow_decapkapwr_6.pxi.spice
* Created: Thu Aug 27 14:24:42 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%VGND N_VGND_M1001_s N_VGND_c_18_n VGND
+ N_VGND_c_19_n N_VGND_M1000_g N_VGND_c_20_n N_VGND_c_21_n N_VGND_c_22_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%KAPWR N_KAPWR_M1000_s N_KAPWR_M1001_g
+ KAPWR N_KAPWR_c_40_n N_KAPWR_c_41_n N_KAPWR_c_42_n N_KAPWR_c_44_n
+ N_KAPWR_c_45_n N_KAPWR_c_46_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%VPWR VPWR N_VPWR_c_69_n N_VPWR_c_68_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%VPWR
cc_1 VNB N_VGND_c_18_n 0.0120582f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=0.385
cc_2 VNB N_VGND_c_19_n 0.0332598f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.29
cc_3 VNB N_VGND_c_20_n 0.0745147f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.475
cc_4 VNB N_VGND_c_21_n 0.0439657f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=0.475
cc_5 VNB N_VGND_c_22_n 0.159975f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0
cc_6 VNB N_KAPWR_c_40_n 0.121206f $X=-0.19 $Y=-0.24 $X2=0.647 $Y2=0
cc_7 VNB N_KAPWR_c_41_n 0.0178046f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0
cc_8 VNB N_KAPWR_c_42_n 0.0831515f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0
cc_9 VNB N_VPWR_c_68_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=-0.085
cc_10 VPB N_VGND_c_19_n 0.183789f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.29
cc_11 VPB N_VGND_c_20_n 0.00687586f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.475
cc_12 VPB N_KAPWR_c_41_n 0.0451006f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0
cc_13 VPB N_KAPWR_c_44_n 0.0353425f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=0
cc_14 VPB N_KAPWR_c_45_n 0.0111567f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=0
cc_15 VPB N_KAPWR_c_46_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_16 VPB N_VPWR_c_69_n 0.0671091f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.385
cc_17 VPB N_VPWR_c_68_n 0.0420602f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=-0.085
cc_18 N_VGND_c_18_n N_KAPWR_c_40_n 0.0738934f $X=2.205 $Y=0.385 $X2=0 $Y2=0
cc_19 N_VGND_c_19_n N_KAPWR_c_40_n 0.0673714f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_20 N_VGND_c_20_n N_KAPWR_c_40_n 0.00648994f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_21 N_VGND_c_21_n N_KAPWR_c_40_n 0.0237188f $X=2.5 $Y=0.475 $X2=0 $Y2=0
cc_22 N_VGND_c_18_n N_KAPWR_c_41_n 0.0622608f $X=2.205 $Y=0.385 $X2=0 $Y2=0
cc_23 N_VGND_c_19_n N_KAPWR_c_41_n 0.116191f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_24 N_VGND_c_20_n N_KAPWR_c_41_n 0.0326482f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_25 N_VGND_c_21_n N_KAPWR_c_41_n 0.0424967f $X=2.5 $Y=0.475 $X2=0 $Y2=0
cc_26 N_VGND_c_18_n N_KAPWR_c_42_n 0.0203211f $X=2.205 $Y=0.385 $X2=0 $Y2=0
cc_27 N_VGND_c_19_n N_KAPWR_c_42_n 0.0617911f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_28 N_VGND_c_20_n N_KAPWR_c_42_n 0.105038f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_29 N_VGND_c_19_n N_KAPWR_c_44_n 0.123992f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_30 N_VGND_c_20_n N_KAPWR_c_44_n 0.104838f $X=0.26 $Y=0.475 $X2=0 $Y2=0
cc_31 N_VGND_c_19_n N_VPWR_c_69_n 0.0470038f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_32 N_VGND_c_19_n N_VPWR_c_68_n 0.0437167f $X=1.11 $Y=1.29 $X2=0 $Y2=0
cc_33 N_KAPWR_c_41_n N_VPWR_c_69_n 0.0810717f $X=2.2 $Y=1.11 $X2=0 $Y2=0
cc_34 N_KAPWR_c_44_n N_VPWR_c_69_n 0.0922017f $X=1.465 $Y=2.005 $X2=0 $Y2=0
cc_35 N_KAPWR_c_45_n N_VPWR_c_69_n 9.05775e-19 $X=2.53 $Y=2.21 $X2=0 $Y2=0
cc_36 N_KAPWR_c_46_n N_VPWR_c_69_n 0.00102011f $X=0.215 $Y=2.21 $X2=0 $Y2=0
cc_37 N_KAPWR_M1000_s N_VPWR_c_68_n 0.00214089f $X=0.135 $Y=1.615 $X2=0 $Y2=0
cc_38 N_KAPWR_c_41_n N_VPWR_c_68_n 0.0102288f $X=2.2 $Y=1.11 $X2=0 $Y2=0
cc_39 N_KAPWR_c_44_n N_VPWR_c_68_n 0.0116508f $X=1.465 $Y=2.005 $X2=0 $Y2=0
cc_40 N_KAPWR_c_46_n N_VPWR_c_68_n 0.267826f $X=0.215 $Y=2.21 $X2=0 $Y2=0

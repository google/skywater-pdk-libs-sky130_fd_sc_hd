* File: sky130_fd_sc_hd__dlclkp_1.spice
* Created: Thu Aug 27 14:16:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlclkp_1.spice.pex"
.subckt sky130_fd_sc_hd__dlclkp_1  VNB VPB CLK GATE VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* GATE	GATE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_CLK_M1019_g N_A_27_47#_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_193_47#_M1010_d N_A_27_47#_M1010_g N_VGND_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_396_119# N_GATE_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.117125 AS=0.1281 PD=1.085 PS=1.45 NRD=63.96 NRS=11.424 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_476_413#_M1009_d N_A_27_47#_M1009_g A_396_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.123615 AS=0.117125 PD=1.13037 PS=1.085 NRD=81.42 NRS=63.96 M=1
+ R=2.8 SA=75000.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 A_651_47# N_A_193_47#_M1014_g N_A_476_413#_M1009_d VNB NSHORT L=0.15
+ W=0.39 AD=0.0646389 AS=0.114785 PD=0.717407 PS=1.04963 NRD=34.068 NRS=3.072
+ M=1 R=2.6 SA=75000.9 SB=75001.2 A=0.0585 P=1.08 MULT=1
MM1004 N_VGND_M1004_d N_A_642_307#_M1004_g A_651_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.0696111 PD=0.816449 PS=0.772593 NRD=32.856 NRS=31.632 M=1
+ R=2.8 SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_A_642_307#_M1011_d N_A_476_413#_M1011_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.143516 PD=1.82 PS=1.26355 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 A_1042_47# N_A_642_307#_M1001_g N_A_957_369#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_CLK_M1016_g A_1042_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.0441 PD=0.765421 PS=0.63 NRD=12.852 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_GCLK_M1006_d N_A_957_369#_M1006_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_CLK_M1008_g N_A_27_47#_M1008_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 A_381_369# N_GATE_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.115623 AS=0.1664 PD=1.16528 PS=1.8 NRD=38.6711 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_476_413#_M1005_d N_A_193_47#_M1005_g A_381_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0987 AS=0.0758774 PD=0.89 PS=0.764717 NRD=56.2829 NRS=58.9227 M=1
+ R=2.8 SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 A_600_413# N_A_27_47#_M1002_g N_A_476_413#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0987 PD=0.63 PS=0.89 NRD=23.443 NRS=32.8202 M=1 R=2.8
+ SA=75001.3 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_642_307#_M1003_g A_600_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_476_413#_M1018_g N_A_642_307#_M1018_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.181707 AS=0.27 PD=1.61585 PS=2.54 NRD=1.9503 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1007 N_A_957_369#_M1007_d N_A_642_307#_M1007_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2032 AS=0.116293 PD=1.275 PS=1.03415 NRD=75.4116
+ NRS=10.7562 M=1 R=4.26667 SA=75000.7 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1013 N_VPWR_M1013_d N_CLK_M1013_g N_A_957_369#_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.116293 AS=0.2032 PD=1.03415 PS=1.275 NRD=15.3857 NRS=33.8446 M=1
+ R=4.26667 SA=75001.5 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1012 N_GCLK_M1012_d N_A_957_369#_M1012_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.8648 P=16.95
c_141 VPB 0 4.14077e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dlclkp_1.spice.SKY130_FD_SC_HD__DLCLKP_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__dlxtn_2.spice.pex
* Created: Thu Aug 27 14:18:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLXTN_2%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%A_27_47# 1 2 9 13 17 20 24 28 29 30 38 42 45
+ 47 52 54 56 57 60 63 64 68 71 75 79
c167 20 0 1.41946e-19 $X=3.355 $Y=2.275
c168 13 0 2.6965e-20 $X=0.89 $Y=2.135
c169 9 0 2.6965e-20 $X=0.89 $Y=0.445
r170 64 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.115 $Y=1.53
+ $X2=3.115 $Y2=1.415
r171 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.035 $Y=1.53
+ $X2=3.035 $Y2=1.53
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r173 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.89 $Y=1.53
+ $X2=3.035 $Y2=1.53
r175 56 57 2.53712 $w=1.4e-07 $l=2.05e-06 $layer=MET1_cond $X=2.89 $Y=1.53
+ $X2=0.84 $Y2=1.53
r176 52 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=0.87
+ $X2=2.82 $Y2=0.705
r177 51 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.82 $Y=0.87
+ $X2=3.03 $Y2=0.87
r178 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=0.87 $X2=2.82 $Y2=0.87
r179 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r180 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r181 46 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r182 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r183 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r184 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r185 39 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.2 $Y=1.74
+ $X2=3.355 $Y2=1.74
r186 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.74 $X2=3.2 $Y2=1.74
r187 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.115 $Y=1.585
+ $X2=3.115 $Y2=1.53
r188 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.115 $Y=1.585
+ $X2=3.115 $Y2=1.74
r189 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=1.035
+ $X2=3.03 $Y2=0.87
r190 34 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.03 $Y=1.035
+ $X2=3.03 $Y2=1.415
r191 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r192 31 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r193 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r194 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r195 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r196 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r197 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r198 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r199 18 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.355 $Y=1.875
+ $X2=3.355 $Y2=1.74
r200 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.355 $Y=1.875
+ $X2=3.355 $Y2=2.275
r201 17 71 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.81 $Y=0.415
+ $X2=2.81 $Y2=0.705
r202 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r203 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r204 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r206 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.645 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.645 $Y=1.04
+ $X2=1.85 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.04 $X2=1.645 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.645 $Y=1.19
+ $X2=1.645 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.205
+ $X2=1.85 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.85 $Y=1.205 $X2=1.85
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=0.875
+ $X2=1.85 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.85 $Y=0.875 $X2=1.85
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%A_303_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 32 0 1.12109e-19 $X=2.275 $Y=0.93
c84 18 0 7.13094e-20 $X=1.99 $Y=0.7
r85 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.93
+ $X2=2.275 $Y2=1.095
r86 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.93
+ $X2=2.275 $Y2=0.765
r87 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=0.93 $X2=2.275 $Y2=0.93
r88 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.64 $Y=0.51
+ $X2=1.64 $Y2=0.7
r89 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.075 $Y=1.095
+ $X2=2.175 $Y2=0.93
r90 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.075 $Y=1.095
+ $X2=2.075 $Y2=1.495
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.99 $Y=1.58
+ $X2=2.075 $Y2=1.495
r92 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.99 $Y=1.58
+ $X2=1.805 $Y2=1.58
r93 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.7
+ $X2=1.64 $Y2=0.7
r94 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.99 $Y=0.7
+ $X2=2.175 $Y2=0.93
r95 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.99 $Y=0.7
+ $X2=1.725 $Y2=0.7
r96 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=1.665
+ $X2=1.805 $Y2=1.58
r97 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.64 $Y=1.665
+ $X2=1.64 $Y2=1.99
r98 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.27 $Y=2.165
+ $X2=2.27 $Y2=1.095
r99 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.27 $Y=0.445
+ $X2=2.27 $Y2=0.765
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=1.845 $X2=1.64 $Y2=1.99
r101 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.235 $X2=1.64 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c112 38 0 1.41946e-19 $X=2.69 $Y=1.52
r113 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.52 $X2=2.69 $Y2=1.52
r114 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.632 $Y=1.87
+ $X2=2.632 $Y2=1.52
r115 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.575 $Y=1.87
+ $X2=2.575 $Y2=1.87
r116 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r117 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.43 $Y=1.87
+ $X2=2.575 $Y2=1.87
r119 26 27 1.39851 $w=1.4e-07 $l=1.13e-06 $layer=MET1_cond $X=2.43 $Y=1.87
+ $X2=1.3 $Y2=1.87
r120 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r121 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r122 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r123 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.69 $Y=1.55 $X2=2.69
+ $Y2=1.52
r124 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.69 $Y=1.55
+ $X2=2.69 $Y2=1.685
r125 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.69 $Y=1.395
+ $X2=2.69 $Y2=1.52
r126 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.24 $Y=1.245
+ $X2=3.24 $Y2=0.415
r127 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.825 $Y=1.32
+ $X2=2.69 $Y2=1.395
r128 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.165 $Y=1.32
+ $X2=3.24 $Y2=1.245
r129 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.165 $Y=1.32
+ $X2=2.825 $Y2=1.32
r130 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.75 $Y=2.275
+ $X2=2.75 $Y2=1.685
r131 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r132 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%A_728_21# 1 2 9 13 15 17 20 22 24 27 29 32
+ 36 40 43 45 48 51 53 54 62
r96 61 62 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.51 $Y2=1.16
r97 49 61 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.075 $Y=1.16
+ $X2=5.09 $Y2=1.16
r98 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.075
+ $Y=1.16 $X2=5.075 $Y2=1.16
r99 46 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=1.16
+ $X2=4.495 $Y2=1.16
r100 46 48 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.58 $Y=1.16
+ $X2=5.075 $Y2=1.16
r101 45 53 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.495 $Y=1.535
+ $X2=4.47 $Y2=1.7
r102 44 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=1.325
+ $X2=4.495 $Y2=1.16
r103 44 45 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.495 $Y=1.325
+ $X2=4.495 $Y2=1.535
r104 43 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.995
+ $X2=4.495 $Y2=1.16
r105 43 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.495 $Y=0.995
+ $X2=4.495 $Y2=0.825
r106 38 53 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=1.865
+ $X2=4.47 $Y2=1.7
r107 38 40 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.47 $Y=1.865
+ $X2=4.47 $Y2=2.27
r108 34 51 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=4.47 $Y=0.715
+ $X2=4.47 $Y2=0.825
r109 34 36 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=4.47 $Y=0.715
+ $X2=4.47 $Y2=0.58
r110 32 55 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.945 $Y=1.7
+ $X2=3.715 $Y2=1.7
r111 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.945
+ $Y=1.7 $X2=3.945 $Y2=1.7
r112 29 53 0.463323 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.36 $Y=1.7
+ $X2=4.47 $Y2=1.7
r113 29 31 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.36 $Y=1.7
+ $X2=3.945 $Y2=1.7
r114 25 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=1.325
+ $X2=5.51 $Y2=1.16
r115 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.51 $Y=1.325
+ $X2=5.51 $Y2=1.985
r116 22 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=0.995
+ $X2=5.51 $Y2=1.16
r117 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.51 $Y=0.995
+ $X2=5.51 $Y2=0.56
r118 18 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.325
+ $X2=5.09 $Y2=1.16
r119 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.09 $Y=1.325
+ $X2=5.09 $Y2=1.985
r120 15 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=0.995
+ $X2=5.09 $Y2=1.16
r121 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.09 $Y=0.995
+ $X2=5.09 $Y2=0.56
r122 11 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.715 $Y=1.865
+ $X2=3.715 $Y2=1.7
r123 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.715 $Y=1.865
+ $X2=3.715 $Y2=2.275
r124 7 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.715 $Y=1.535
+ $X2=3.715 $Y2=1.7
r125 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.715 $Y=1.535
+ $X2=3.715 $Y2=0.445
r126 2 53 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.485 $X2=4.445 $Y2=1.755
r127 2 40 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.485 $X2=4.445 $Y2=2.27
r128 1 36 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.235 $X2=4.445 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%A_565_413# 1 2 7 9 12 14 15 16 20 25 26 27
+ 30
c83 26 0 1.57048e-19 $X=3.585 $Y=1.325
c84 15 0 1.24415e-19 $X=4.655 $Y=1.16
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.16 $X2=4.135 $Y2=1.16
r86 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.67 $Y=1.16
+ $X2=4.135 $Y2=1.16
r87 26 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.585 $Y=1.325
+ $X2=3.51 $Y2=1.16
r88 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.585 $Y=1.325
+ $X2=3.585 $Y2=2.255
r89 25 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.435 $Y=0.995
+ $X2=3.51 $Y2=1.16
r90 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.435 $Y=0.535
+ $X2=3.435 $Y2=0.995
r91 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=2.34
+ $X2=3.585 $Y2=2.255
r92 20 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.5 $Y=2.34
+ $X2=3.085 $Y2=2.34
r93 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.35 $Y=0.45
+ $X2=3.435 $Y2=0.535
r94 16 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.35 $Y=0.45
+ $X2=3.025 $Y2=0.45
r95 14 31 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.58 $Y=1.16
+ $X2=4.135 $Y2=1.16
r96 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.58 $Y=1.16
+ $X2=4.655 $Y2=1.16
r97 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.325
+ $X2=4.655 $Y2=1.16
r98 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.655 $Y=1.325
+ $X2=4.655 $Y2=1.985
r99 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=0.995
+ $X2=4.655 $Y2=1.16
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.655 $Y=0.995
+ $X2=4.655 $Y2=0.56
r101 2 22 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=2.065 $X2=3.085 $Y2=2.34
r102 1 18 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.235 $X2=3.025 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%VPWR 1 2 3 4 5 18 22 26 28 32 34 36 38 40 45
+ 50 55 61 64 67 70 74
r94 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r95 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r96 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r97 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r99 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r100 59 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 59 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r103 56 70 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=4.902 $Y2=2.72
r104 56 58 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=5.29 $Y2=2.72
r105 55 73 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.807 $Y2=2.72
r106 55 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.29 $Y2=2.72
r107 54 68 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r108 54 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r110 51 64 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.29 $Y=2.72
+ $X2=2.132 $Y2=2.72
r111 51 53 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.29 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 50 67 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.84 $Y=2.72
+ $X2=3.99 $Y2=2.72
r113 50 53 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.84 $Y=2.72
+ $X2=2.53 $Y2=2.72
r114 49 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r115 49 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r117 46 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r118 46 48 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r119 45 64 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.132 $Y2=2.72
r120 45 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r121 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r122 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r123 38 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r125 34 73 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.765 $Y=2.635
+ $X2=5.807 $Y2=2.72
r126 34 36 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=5.765 $Y=2.635
+ $X2=5.765 $Y2=2
r127 30 70 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.902 $Y=2.635
+ $X2=4.902 $Y2=2.72
r128 30 32 36.3929 $w=2.83e-07 $l=9e-07 $layer=LI1_cond $X=4.902 $Y=2.635
+ $X2=4.902 $Y2=1.735
r129 29 67 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.14 $Y=2.72
+ $X2=3.99 $Y2=2.72
r130 28 70 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.76 $Y=2.72
+ $X2=4.902 $Y2=2.72
r131 28 29 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.76 $Y=2.72
+ $X2=4.14 $Y2=2.72
r132 24 67 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=2.635
+ $X2=3.99 $Y2=2.72
r133 24 26 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.99 $Y=2.635
+ $X2=3.99 $Y2=2.3
r134 20 64 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.132 $Y=2.635
+ $X2=2.132 $Y2=2.72
r135 20 22 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.132 $Y=2.635
+ $X2=2.132 $Y2=2
r136 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r137 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r138 5 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=2
r139 4 32 300 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=2 $X=4.73
+ $Y=1.485 $X2=4.88 $Y2=1.735
r140 3 26 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.79
+ $Y=2.065 $X2=3.925 $Y2=2.3
r141 2 22 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=1.845 $X2=2.06 $Y2=2
r142 1 18 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%Q 1 2 7 8 12 13 14 15 16 17
c25 17 0 1.24415e-19 $X=5.78 $Y=1.19
r26 17 31 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.78 $Y=1.16
+ $X2=5.415 $Y2=1.16
r27 15 16 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=5.34 $Y=1.835
+ $X2=5.34 $Y2=2.21
r28 13 15 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=5.34 $Y=1.64
+ $X2=5.34 $Y2=1.835
r29 12 13 7.87132 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=5.357 $Y=1.495
+ $X2=5.357 $Y2=1.64
r30 9 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=1.325
+ $X2=5.415 $Y2=1.16
r31 9 12 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=1.325
+ $X2=5.415 $Y2=1.495
r32 8 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=0.995
+ $X2=5.415 $Y2=1.16
r33 7 14 16.2055 $w=2.61e-07 $l=3.42775e-07 $layer=LI1_cond $X=5.415 $Y=0.825
+ $X2=5.357 $Y2=0.51
r34 7 8 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=0.825
+ $X2=5.415 $Y2=0.995
r35 2 15 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=1.835
r36 1 14 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.165
+ $Y=0.235 $X2=5.3 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_2%VGND 1 2 3 4 5 18 22 26 28 32 34 36 38 40 45
+ 50 58 64 67 70 73 77
c97 77 0 2.71124e-20 $X=5.75 $Y=0
c98 2 0 7.13094e-20 $X=1.925 $Y=0.235
r99 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r100 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r101 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r102 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r103 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r104 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r105 62 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r106 62 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r107 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r108 59 73 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=4.902 $Y2=0
r109 59 61 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.29
+ $Y2=0
r110 58 76 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.635 $Y=0
+ $X2=5.807 $Y2=0
r111 58 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.635 $Y=0 $X2=5.29
+ $Y2=0
r112 57 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r113 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r114 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r115 54 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r116 53 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r117 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r118 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.06
+ $Y2=0
r119 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.53 $Y2=0
r120 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.925
+ $Y2=0
r121 50 56 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.45
+ $Y2=0
r122 49 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r123 49 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r124 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r125 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r126 46 48 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r127 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.06
+ $Y2=0
r128 45 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.61 $Y2=0
r129 40 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r130 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r131 38 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r132 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r133 34 76 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.765 $Y=0.085
+ $X2=5.807 $Y2=0
r134 34 36 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.765 $Y=0.085
+ $X2=5.765 $Y2=0.38
r135 30 73 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.902 $Y=0.085
+ $X2=4.902 $Y2=0
r136 30 32 18.803 $w=2.83e-07 $l=4.65e-07 $layer=LI1_cond $X=4.902 $Y=0.085
+ $X2=4.902 $Y2=0.55
r137 29 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.925
+ $Y2=0
r138 28 73 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.76 $Y=0 $X2=4.902
+ $Y2=0
r139 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.76 $Y=0 $X2=4.09
+ $Y2=0
r140 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r141 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.445
r142 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0
r143 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0.36
r144 16 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r145 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r146 5 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.38
r147 4 32 182 $w=1.7e-07 $l=3.82721e-07 $layer=licon1_NDIFF $count=1 $X=4.73
+ $Y=0.235 $X2=4.88 $Y2=0.55
r148 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.79
+ $Y=0.235 $X2=3.925 $Y2=0.445
r149 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.06 $Y2=0.36
r150 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.195000 1.445000 ;
        RECT 0.855000 1.445000 1.240000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.500000 0.255000 6.830000 0.445000 ;
        RECT 6.580000 0.445000 6.830000 0.715000 ;
        RECT 6.580000 0.715000 7.220000 0.885000 ;
        RECT 6.580000 1.485000 7.220000 1.655000 ;
        RECT 6.580000 1.655000 6.830000 2.465000 ;
        RECT 7.050000 0.885000 7.220000 1.055000 ;
        RECT 7.050000 1.055000 8.195000 1.315000 ;
        RECT 7.050000 1.315000 7.220000 1.485000 ;
        RECT 7.420000 0.255000 7.720000 1.055000 ;
        RECT 7.420000 1.315000 7.720000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.345000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.725000 0.995000 4.945000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.685000 0.995000 6.065000 1.325000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.710000 1.075000 5.000000 1.120000 ;
        RECT 4.710000 1.120000 5.940000 1.260000 ;
        RECT 4.710000 1.260000 5.000000 1.305000 ;
        RECT 5.650000 1.075000 5.940000 1.120000 ;
        RECT 5.650000 1.260000 5.940000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.445000 ;
        RECT 2.670000  0.085000 3.015000 0.825000 ;
        RECT 4.095000  0.085000 4.425000 0.445000 ;
        RECT 5.605000  0.085000 6.330000 0.445000 ;
        RECT 7.000000  0.085000 7.250000 0.545000 ;
        RECT 7.890000  0.085000 8.195000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 0.085000 1.835000 0.345000 2.635000 ;
        RECT 2.375000 2.075000 3.015000 2.635000 ;
        RECT 3.595000 2.255000 5.515000 2.635000 ;
        RECT 6.055000 2.255000 6.385000 2.635000 ;
        RECT 7.000000 1.825000 7.250000 2.635000 ;
        RECT 7.890000 1.485000 8.195000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.345000 0.615000 ;
      RECT 0.085000 0.615000 1.195000 0.785000 ;
      RECT 0.515000 0.785000 0.685000 2.125000 ;
      RECT 0.515000 2.125000 1.260000 2.465000 ;
      RECT 1.015000 0.255000 1.195000 0.615000 ;
      RECT 1.365000 0.255000 2.500000 0.535000 ;
      RECT 1.365000 0.705000 1.705000 1.205000 ;
      RECT 1.365000 1.205000 1.865000 1.325000 ;
      RECT 1.410000 1.325000 1.865000 1.955000 ;
      RECT 1.430000 2.125000 2.205000 2.465000 ;
      RECT 1.875000 0.705000 2.160000 1.035000 ;
      RECT 2.035000 1.205000 3.015000 1.375000 ;
      RECT 2.035000 1.375000 2.205000 2.125000 ;
      RECT 2.330000 0.535000 2.500000 0.995000 ;
      RECT 2.330000 0.995000 3.015000 1.205000 ;
      RECT 2.375000 1.575000 2.545000 1.635000 ;
      RECT 2.375000 1.635000 3.405000 1.905000 ;
      RECT 3.185000 0.255000 3.405000 1.635000 ;
      RECT 3.185000 1.905000 3.405000 1.915000 ;
      RECT 3.185000 1.915000 5.515000 2.085000 ;
      RECT 3.185000 2.085000 3.405000 2.465000 ;
      RECT 3.595000 0.255000 3.925000 0.765000 ;
      RECT 3.595000 0.765000 4.020000 0.935000 ;
      RECT 3.595000 0.935000 3.765000 1.575000 ;
      RECT 3.595000 1.575000 4.005000 1.745000 ;
      RECT 3.935000 1.105000 4.480000 1.275000 ;
      RECT 4.175000 1.275000 4.480000 1.495000 ;
      RECT 4.175000 1.495000 4.975000 1.745000 ;
      RECT 4.190000 0.615000 4.845000 0.785000 ;
      RECT 4.190000 0.785000 4.480000 1.105000 ;
      RECT 4.595000 0.255000 4.845000 0.615000 ;
      RECT 5.015000 0.255000 5.435000 0.615000 ;
      RECT 5.015000 0.615000 6.410000 0.785000 ;
      RECT 5.165000 0.995000 5.515000 1.915000 ;
      RECT 5.685000 1.495000 6.410000 2.085000 ;
      RECT 5.685000 2.085000 5.855000 2.465000 ;
      RECT 6.240000 0.785000 6.410000 1.055000 ;
      RECT 6.240000 1.055000 6.880000 1.315000 ;
      RECT 6.240000 1.315000 6.410000 1.495000 ;
    LAYER mcon ;
      RECT 1.530000 1.445000 1.700000 1.615000 ;
      RECT 1.990000 0.765000 2.160000 0.935000 ;
      RECT 3.850000 0.765000 4.020000 0.935000 ;
      RECT 4.310000 1.445000 4.480000 1.615000 ;
    LAYER met1 ;
      RECT 1.470000 1.415000 1.760000 1.460000 ;
      RECT 1.470000 1.460000 4.540000 1.600000 ;
      RECT 1.470000 1.600000 1.760000 1.645000 ;
      RECT 1.930000 0.735000 2.220000 0.780000 ;
      RECT 1.930000 0.780000 4.080000 0.920000 ;
      RECT 1.930000 0.920000 2.220000 0.965000 ;
      RECT 3.790000 0.735000 4.080000 0.780000 ;
      RECT 3.790000 0.920000 4.080000 0.965000 ;
      RECT 4.250000 1.415000 4.540000 1.460000 ;
      RECT 4.250000 1.600000 4.540000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_4
END LIBRARY

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.5898e+12p ps=1.527e+07u
M1001 a_725_21# a_562_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1002 VPWR a_725_21# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6.15e+11p ps=5.23e+06u
M1003 a_943_47# a_562_413# a_725_21# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=1.69e+11p ps=1.82e+06u
M1004 a_683_413# a_27_47# a_562_413# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.911e+11p ps=1.75e+06u
M1005 a_466_47# a_300_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.62e+06u as=9.0475e+11p ps=9.77e+06u
M1006 VPWR a_725_21# a_683_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_725_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.9975e+11p ps=3.83e+06u
M1008 a_562_413# a_27_47# a_466_47# VNB nshort w=360000u l=150000u
+  ad=1.008e+11p pd=1.28e+06u as=0p ps=0u
M1009 VGND a_725_21# a_660_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1010 VPWR RESET_B a_725_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR GATE_N a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1012 a_466_369# a_300_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.936e+11p pd=1.94e+06u as=0p ps=0u
M1013 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1014 Q a_725_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_725_21# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR D a_300_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1017 VGND a_725_21# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_725_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_660_47# a_193_47# a_562_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q a_725_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND RESET_B a_943_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND D a_300_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1023 Q a_725_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND GATE_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1025 a_562_413# a_193_47# a_466_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__einvp_1.pex.spice
* Created: Thu Aug 27 14:20:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVP_1%TE 3 7 9 10 11 13 14 15
c38 10 0 1.48222e-19 $X=0.545 $Y=1.035
r39 19 21 30.5162 $w=3.08e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.132
+ $X2=0.47 $Y2=1.132
r40 14 15 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=1.16
+ $X2=0.315 $Y2=1.53
r41 14 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r42 11 13 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.945 $Y=0.96
+ $X2=0.945 $Y2=0.56
r43 10 21 24.4482 $w=3.08e-07 $l=1.29167e-07 $layer=POLY_cond $X=0.545 $Y=1.035
+ $X2=0.47 $Y2=1.132
r44 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.87 $Y=1.035
+ $X2=0.945 $Y2=0.96
r45 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.87 $Y=1.035
+ $X2=0.545 $Y2=1.035
r46 5 21 19.5884 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.132
r47 5 7 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=2.275
r48 1 21 19.5884 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.47 $Y2=1.132
r49 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_1%A_27_47# 1 2 9 13 17 19 20 21 22 26 27
c66 21 0 1.48222e-19 $X=0.715 $Y=1.98
r67 27 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.16
+ $X2=1.365 $Y2=1.325
r68 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.365
+ $Y=1.16 $X2=1.365 $Y2=1.16
r69 24 26 11.9608 $w=7.33e-07 $l=7.35e-07 $layer=LI1_cond $X=1.082 $Y=1.895
+ $X2=1.082 $Y2=1.16
r70 23 26 5.45151 $w=7.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.082 $Y=0.825
+ $X2=1.082 $Y2=1.16
r71 21 24 11.0548 $w=1.7e-07 $l=4.07289e-07 $layer=LI1_cond $X=0.715 $Y=1.98
+ $X2=1.082 $Y2=1.895
r72 21 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=1.98
+ $X2=0.345 $Y2=1.98
r73 19 23 11.0548 $w=1.7e-07 $l=4.07289e-07 $layer=LI1_cond $X=0.715 $Y=0.74
+ $X2=1.082 $Y2=0.825
r74 19 20 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.74
+ $X2=0.345 $Y2=0.74
r75 15 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=2.065
+ $X2=0.345 $Y2=1.98
r76 15 17 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=2.065
+ $X2=0.215 $Y2=2.275
r77 11 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.345 $Y2=0.74
r78 11 13 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r79 9 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.305 $Y=1.985
+ $X2=1.305 $Y2=1.325
r80 2 17 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.275
r81 1 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_1%A 1 3 6 8 9 10 17
r29 14 17 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=2.06 $Y2=1.16
r30 9 10 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.095 $Y=1.53
+ $X2=2.095 $Y2=1.87
r31 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=1.16
+ $X2=2.095 $Y2=1.53
r32 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r33 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.325
+ $X2=1.82 $Y2=1.16
r34 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.82 $Y=1.325 $X2=1.82
+ $Y2=1.985
r35 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.82 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_1%VPWR 1 4 6 8 9 10 22 23
r28 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 20 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r30 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r31 17 19 2.51806 $w=5.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.03 $Y=2.52
+ $X2=1.15 $Y2=2.52
r32 10 20 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 10 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r34 9 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=2.72 $X2=2.07
+ $Y2=2.72
r35 8 19 0.314757 $w=5.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=2.52
+ $X2=1.15 $Y2=2.52
r36 8 9 12.4791 $w=5.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.165 $Y=2.52
+ $X2=1.45 $Y2=2.52
r37 6 13 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r38 4 17 4.82628 $w=5.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.8 $Y=2.52 $X2=1.03
+ $Y2=2.52
r39 4 6 12.4791 $w=5.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.8 $Y=2.52 $X2=0.515
+ $Y2=2.52
r40 1 17 300 $w=1.7e-07 $l=6.13086e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=2.065 $X2=1.03 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_1%Z 1 2 8 9 10 14
r34 19 22 11.2872 $w=3.38e-07 $l=3.33e-07 $layer=LI1_cond $X=1.707 $Y=2.295
+ $X2=2.04 $Y2=2.295
r35 10 22 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=2.075 $Y=2.295
+ $X2=2.04 $Y2=2.295
r36 9 18 12.5286 $w=5.93e-07 $l=2.95e-07 $layer=LI1_cond $X=1.917 $Y=0.51
+ $X2=1.917 $Y2=0.805
r37 9 14 2.61328 $w=5.93e-07 $l=1.3e-07 $layer=LI1_cond $X=1.917 $Y=0.51
+ $X2=1.917 $Y2=0.38
r38 8 19 4.64683 $w=1.75e-07 $l=1.7e-07 $layer=LI1_cond $X=1.707 $Y=2.125
+ $X2=1.707 $Y2=2.295
r39 8 18 83.6571 $w=1.73e-07 $l=1.32e-06 $layer=LI1_cond $X=1.707 $Y=2.125
+ $X2=1.707 $Y2=0.805
r40 2 22 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.04 $Y2=2.3
r41 1 14 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.895
+ $Y=0.235 $X2=2.03 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_1%VGND 1 4 13 14 18 25
r27 23 25 12.7938 $w=5.68e-07 $l=3e-07 $layer=LI1_cond $X=1.15 $Y=0.2 $X2=1.45
+ $Y2=0.2
r28 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r29 21 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r30 20 23 9.65256 $w=5.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.2 $X2=1.15
+ $Y2=0.2
r31 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r32 17 20 0.209838 $w=5.68e-07 $l=1e-08 $layer=LI1_cond $X=0.68 $Y=0.2 $X2=0.69
+ $Y2=0.2
r33 17 18 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.2
+ $X2=0.515 $Y2=0.2
r34 14 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r35 13 25 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.45
+ $Y2=0
r36 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r37 8 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.515
+ $Y2=0
r38 4 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r39 4 8 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r40 1 17 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


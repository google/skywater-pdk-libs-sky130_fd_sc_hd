* File: sky130_fd_sc_hd__macro_sparecell.pxi.spice
* Created: Thu Aug 27 14:27:00 2020
* 
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_1/A
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1003_d
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1005_s
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1001_g
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1003_g
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n N_SKY130_FD_SC_HD__INV_2_1/A_c_242_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_259_p N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_265_p N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n N_SKY130_FD_SC_HD__INV_2_1/A_c_245_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_246_n N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n N_SKY130_FD_SC_HD__INV_2_1/A_c_249_n
+ N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_1/A
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__NOR2_2_1/B
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1003_s
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1000_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1005_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1001_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1002_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1003_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1004_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n N_SKY130_FD_SC_HD__NOR2_2_1/B_c_414_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_415_p N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_424_p N_SKY130_FD_SC_HD__NOR2_2_1/B_c_420_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_416_p N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_362_n N_SKY130_FD_SC_HD__NOR2_2_1/B_c_363_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_400_n N_SKY130_FD_SC_HD__NOR2_2_1/B_c_401_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_364_n N_SKY130_FD_SC_HD__NOR2_2_1/B_c_406_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_367_n N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_377_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__NOR2_2_1/B
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%LO N_LO_c_513_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1003_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g N_LO_c_514_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1004_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g N_LO_c_515_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1002_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g N_LO_c_516_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1007_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g N_LO_c_517_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1002_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g N_LO_c_518_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1007_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g N_LO_c_519_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1003_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g N_LO_c_520_n
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1004_g
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g N_LO_c_521_n N_LO_c_522_n
+ N_LO_c_523_n N_LO_c_583_n N_LO_c_524_n N_LO_c_525_n N_LO_c_526_n N_LO_c_527_n
+ N_LO_c_528_n N_LO_c_529_n N_LO_c_530_n N_LO_c_531_n LO
+ N_LO_Xsky130_fd_sc_hd__conb_1_0/R0_neg N_LO_c_532_n N_LO_c_533_n N_LO_c_534_n
+ N_LO_c_535_n N_LO_c_536_n N_LO_c_537_n N_LO_c_538_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%LO
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%VPWR
+ N_VPWR_Xsky130_fd_sc_hd__inv_2_1/M1000_d
+ N_VPWR_Xsky130_fd_sc_hd__inv_2_1/M1002_d
+ N_VPWR_Xsky130_fd_sc_hd__nor2_2_1/M1000_d
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1000_s
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1001_s
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1006_s
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1000_s
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1001_s
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1006_s
+ N_VPWR_Xsky130_fd_sc_hd__nor2_2_0/M1000_d
+ N_VPWR_Xsky130_fd_sc_hd__inv_2_0/M1000_d
+ N_VPWR_Xsky130_fd_sc_hd__inv_2_0/M1002_d N_VPWR_c_766_n N_VPWR_c_767_n
+ N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n
+ N_VPWR_c_773_n N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_764_n N_VPWR_c_777_n
+ N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n
+ N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n
+ N_VPWR_c_788_n N_VPWR_c_789_n VPWR N_VPWR_Xsky130_fd_sc_hd__conb_1_0/R1_neg
+ N_VPWR_c_790_n N_VPWR_c_791_n N_VPWR_c_792_n N_VPWR_c_793_n N_VPWR_c_794_n
+ N_VPWR_c_795_n N_VPWR_c_796_n N_VPWR_c_797_n N_VPWR_c_798_n N_VPWR_c_799_n
+ N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_804_n
+ N_VPWR_c_765_n PM_SKY130_FD_SC_HD__MACRO_SPARECELL%VPWR
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%VGND
+ N_VGND_Xsky130_fd_sc_hd__inv_2_1/M1001_s
+ N_VGND_Xsky130_fd_sc_hd__inv_2_1/M1003_s
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1001_s
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1002_s
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1004_s
+ N_VGND_Xsky130_fd_sc_hd__nand2_2_1/M1002_s
+ N_VGND_Xsky130_fd_sc_hd__nand2_2_0/M1002_s
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1001_s
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1002_s
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1004_s
+ N_VGND_Xsky130_fd_sc_hd__inv_2_0/M1001_s
+ N_VGND_Xsky130_fd_sc_hd__inv_2_0/M1003_s N_VGND_c_962_n N_VGND_c_963_n
+ N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n N_VGND_c_968_n
+ N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n
+ N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n
+ N_VGND_c_979_n N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n
+ N_VGND_c_984_n VGND N_VGND_Xsky130_fd_sc_hd__conb_1_0/R0_pos N_VGND_c_985_n
+ N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n
+ N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n
+ N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n
+ N_VGND_c_1001_n PM_SKY130_FD_SC_HD__MACRO_SPARECELL%VGND
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__NOR2_2_0/A
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1003_s
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1000_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1005_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1001_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1002_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1003_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1004_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1197_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1202_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1214_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1217_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1219_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1182_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1184_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1185_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1279_p N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1285_p
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1280_p N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1186_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1196_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__NOR2_2_0/A
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_0/A
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1003_d
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_s
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1001_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1003_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1375_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1383_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1418_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1343_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1344_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1346_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_0/A
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_1/Y
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1000_s
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1459_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1461_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1470_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1473_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_1/Y
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1005_d
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1006_d
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1007_s
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1483_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1484_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1485_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1524_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1488_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1000_s
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1007_s
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1006_d
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1532_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1534_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1547_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1536_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_0/Y
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1000_s
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1585_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1582_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1600_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1603_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_0/Y
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1003_d
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1004_d
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1007_d
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1622_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#
x_PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1002_d
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1007_d
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1004_d
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1670_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n
+ PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#
cc_1 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n 0.0209918f $X=-0.19 $Y=-0.24
+ $X2=0.48 $Y2=0.995
cc_2 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n 0.0198569f $X=-0.19 $Y=-0.24
+ $X2=0.9 $Y2=0.995
cc_3 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n 0.0011145f $X=-0.19 $Y=-0.24
+ $X2=1.975 $Y2=0.82
cc_4 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_242_n 0.00235966f $X=-0.19 $Y=-0.24
+ $X2=1.76 $Y2=0.82
cc_5 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n 0.00397808f $X=-0.19 $Y=-0.24
+ $X2=2.815 $Y2=0.815
cc_6 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n 0.00186749f $X=-0.19 $Y=-0.24
+ $X2=2.14 $Y2=0.815
cc_7 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_245_n 0.0011181f $X=-0.19 $Y=-0.24
+ $X2=1.15 $Y2=1.19
cc_8 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_246_n 0.0139471f $X=-0.19 $Y=-0.24
+ $X2=1.51 $Y2=1.19
cc_9 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n 0.00171731f $X=-0.19 $Y=-0.24
+ $X2=1.315 $Y2=1.19
cc_10 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n 0.00204182f $X=-0.19 $Y=-0.24
+ $X2=1.655 $Y2=1.19
cc_11 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_249_n 0.00830399f $X=-0.19 $Y=-0.24
+ $X2=1.655 $Y2=1.19
cc_12 VNB N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n 0.0646401f $X=-0.19 $Y=-0.24
+ $X2=1.11 $Y2=1.16
cc_13 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n 0.0191673f $X=-0.19 $Y=-0.24
+ $X2=0.48 $Y2=0.995
cc_14 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n 0.0157974f $X=-0.19 $Y=-0.24
+ $X2=0.9 $Y2=0.995
cc_15 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n 0.0158002f $X=-0.19 $Y=-0.24
+ $X2=1.975 $Y2=0.82
cc_16 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n 0.0196869f $X=-0.19 $Y=-0.24
+ $X2=2.305 $Y2=0.815
cc_17 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n 0.00394529f $X=-0.19 $Y=-0.24
+ $X2=2.14 $Y2=1.555
cc_18 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.00630293f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_19 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_362_n 0.00910986f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_20 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_363_n 0.00950816f $X=-0.19 $Y=-0.24
+ $X2=1.652 $Y2=1.19
cc_21 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_364_n 0.0119884f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_22 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n 0.0029375f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_23 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n 0.0340596f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_24 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_367_n 0.0345333f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_25 VNB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n 0.00513f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_26 VNB N_LO_c_513_n 0.0191995f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=0.235
cc_27 VNB N_LO_c_514_n 0.0158903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_LO_c_515_n 0.0159539f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.985
cc_29 VNB N_LO_c_516_n 0.0179842f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.985
cc_30 VNB N_LO_c_517_n 0.0179911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_LO_c_518_n 0.0159539f $X=-0.19 $Y=-0.24 $X2=1.652 $Y2=0.905
cc_32 VNB N_LO_c_519_n 0.0158903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_LO_c_520_n 0.0191995f $X=-0.19 $Y=-0.24 $X2=1.315 $Y2=1.19
cc_34 VNB N_LO_c_521_n 0.00204665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_LO_c_522_n 0.00339973f $X=-0.19 $Y=-0.24 $X2=1.652 $Y2=1.19
cc_36 VNB N_LO_c_523_n 0.00375524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_LO_c_524_n 0.00277937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_LO_c_525_n 0.0177343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_LO_c_526_n 0.00396254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_LO_c_527_n 0.0121303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_LO_c_528_n 0.00252956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_LO_c_529_n 7.38737e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_LO_c_530_n 0.00139603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_LO_c_531_n 0.00148871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_LO_c_532_n 0.00805225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_LO_c_533_n 0.0329092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_LO_c_534_n 0.0327227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_LO_c_535_n 0.0327566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_LO_c_536_n 0.00240457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_LO_c_537_n 0.0329092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_LO_c_538_n 0.00587963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB SKY130_FD_SC_HD__CONB_1_0/HI 0.117782f $X=-0.19 $Y=-0.24 $X2=2.005
+ $Y2=1.485
cc_53 VNB N_VPWR_c_764_n 0.00804647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_765_n 0.554392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_962_n 0.0108622f $X=-0.19 $Y=-0.24 $X2=1.652 $Y2=1.555
cc_56 VNB N_VGND_c_963_n 0.00872689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_964_n 0.0113508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_965_n 0.00821008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_966_n 0.00763157f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.19
cc_60 VNB N_VGND_c_967_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.19
cc_61 VNB N_VGND_c_968_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.655 $Y2=1.19
cc_62 VNB N_VGND_c_969_n 0.01493f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_63 VNB N_VGND_c_970_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.16
cc_64 VNB N_VGND_c_971_n 0.00554933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_972_n 0.105774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_973_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_974_n 0.01493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_975_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_976_n 0.00763157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_977_n 0.00821008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_978_n 0.0113508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_979_n 0.0108622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_980_n 0.00872689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_981_n 0.033536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_982_n 0.00452775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_983_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_984_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_985_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_986_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_987_n 0.0391719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_988_n 0.0222979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_989_n 0.0391719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_990_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_991_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_992_n 0.00442067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_993_n 0.00554706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_994_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_995_n 0.00528623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_996_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_997_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_998_n 0.00528623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_999_n 0.00554706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1000_n 0.00442067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1001_n 0.66454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n 0.0196869f $X=-0.19 $Y=-0.24
+ $X2=0.48 $Y2=0.995
cc_96 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n 0.0158002f $X=-0.19 $Y=-0.24
+ $X2=0.9 $Y2=0.995
cc_97 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n 0.0157974f $X=-0.19 $Y=-0.24
+ $X2=1.975 $Y2=0.82
cc_98 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n 0.0191673f $X=-0.19 $Y=-0.24
+ $X2=2.305 $Y2=0.815
cc_99 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n 0.00396855f $X=-0.19 $Y=-0.24
+ $X2=2.14 $Y2=0.815
cc_100 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n 0.00950816f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_101 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1182_n 0.00911045f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_102 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n 0.00630293f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_103 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1184_n 0.0123431f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_104 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1185_n 0.00274448f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_105 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1186_n 0.0345333f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_106 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n 0.0340596f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_107 VNB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n 0.00513f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_108 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n 0.0198569f $X=-0.19 $Y=-0.24
+ $X2=0.48 $Y2=0.995
cc_109 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n 0.0209918f $X=-0.19 $Y=-0.24
+ $X2=0.9 $Y2=0.995
cc_110 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00205847f $X=-0.19 $Y=-0.24
+ $X2=2.14 $Y2=0.39
cc_111 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00192043f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_112 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.00349083f $X=-0.19 $Y=-0.24
+ $X2=2.98 $Y2=0.39
cc_113 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n 0.00187633f $X=-0.19 $Y=-0.24
+ $X2=1.652 $Y2=0.905
cc_114 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1343_n 0.0011181f $X=-0.19 $Y=-0.24
+ $X2=0 $Y2=0
cc_115 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1344_n 0.0139471f $X=-0.19 $Y=-0.24
+ $X2=1.51 $Y2=1.19
cc_116 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n 0.00220609f $X=-0.19 $Y=-0.24
+ $X2=1.315 $Y2=1.19
cc_117 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1346_n 0.00830399f $X=-0.19 $Y=-0.24
+ $X2=1.17 $Y2=1.19
cc_118 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n 0.00153234f $X=-0.19 $Y=-0.24
+ $X2=1.655 $Y2=1.19
cc_119 VNB N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n 0.0646401f $X=-0.19 $Y=-0.24
+ $X2=1.11 $Y2=1.16
cc_120 VNB N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 9.8125e-19 $X=-0.19 $Y=-0.24
+ $X2=0.9 $Y2=1.325
cc_121 VNB N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 9.8125e-19 $X=-0.19 $Y=-0.24
+ $X2=0.9 $Y2=1.325
cc_122 VNB N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 0.00123987f $X=-0.19
+ $Y=-0.24 $X2=0.48 $Y2=1.325
cc_123 VNB N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.00334688f $X=-0.19
+ $Y=-0.24 $X2=0.48 $Y2=1.985
cc_124 VNB N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n 0.00400503f $X=-0.19
+ $Y=-0.24 $X2=0.9 $Y2=0.56
cc_125 VNB N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 0.00307565f $X=-0.19
+ $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n 0.00480403f $X=-0.19
+ $Y=-0.24 $X2=0.48 $Y2=0.56
cc_127 VNB N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n 0.00419179f $X=-0.19
+ $Y=-0.24 $X2=0.48 $Y2=1.985
cc_128 VNB N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 0.00124746f $X=-0.19
+ $Y=-0.24 $X2=0.9 $Y2=0.995
cc_129 VNB N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n 0.00307565f $X=-0.19
+ $Y=-0.24 $X2=1.76 $Y2=0.82
cc_130 VPB N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ 0.0253019f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_131 VPB N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ 0.0231079f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_132 VPB N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n 0.0067499f $X=-0.19 $Y=1.305
+ $X2=2.14 $Y2=1.62
cc_133 VPB N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n 0.00148865f $X=-0.19 $Y=1.305
+ $X2=1.315 $Y2=1.19
cc_134 VPB N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n 6.87247e-19 $X=-0.19 $Y=1.305
+ $X2=1.655 $Y2=1.19
cc_135 VPB N_SKY130_FD_SC_HD__INV_2_1/A_c_249_n 0.00439746f $X=-0.19 $Y=1.305
+ $X2=1.655 $Y2=1.19
cc_136 VPB N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n 0.0151211f $X=-0.19 $Y=1.305
+ $X2=1.11 $Y2=1.16
cc_137 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ 0.0219547f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_138 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ 0.0182972f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_139 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ 0.0179939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ 0.0225925f $X=-0.19 $Y=1.305 $X2=1.652 $Y2=0.905
cc_141 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_363_n 0.00561924f $X=-0.19 $Y=1.305
+ $X2=1.652 $Y2=1.19
cc_142 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n 2.60076e-19 $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_143 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n 0.00421086f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_144 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_367_n 0.00432833f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_145 VPB N_SKY130_FD_SC_HD__NOR2_2_1/B_c_377_n 0.00687837f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_146 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g 0.0219695f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_147 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g 0.0185026f $X=-0.19 $Y=1.305
+ $X2=0.48 $Y2=1.325
cc_148 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g 0.0185065f $X=-0.19 $Y=1.305
+ $X2=0.9 $Y2=1.325
cc_149 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g 0.0210045f $X=-0.19 $Y=1.305
+ $X2=2.14 $Y2=0.39
cc_150 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g 0.0208064f $X=-0.19 $Y=1.305
+ $X2=2.98 $Y2=0.39
cc_151 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g 0.0185065f $X=-0.19 $Y=1.305
+ $X2=2.14 $Y2=1.62
cc_152 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g 0.0185026f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_153 VPB N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g 0.0219695f $X=-0.19 $Y=1.305
+ $X2=1.655 $Y2=1.19
cc_154 VPB N_LO_c_521_n 0.00211564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_LO_c_522_n 0.0044275f $X=-0.19 $Y=1.305 $X2=1.652 $Y2=1.19
cc_156 VPB N_LO_c_523_n 0.00439189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_LO_c_524_n 2.9423e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_LO_c_526_n 0.00148865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_LO_c_528_n 0.00189803f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_LO_c_532_n 0.123209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_LO_c_533_n 0.00412859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_LO_c_534_n 0.00408514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_LO_c_535_n 0.00408639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_LO_c_536_n 0.00211564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_LO_c_537_n 0.00412859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_LO_c_538_n 0.0178775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB SKY130_FD_SC_HD__CONB_1_0/HI 0.00802111f $X=-0.19 $Y=1.305 $X2=2.005
+ $Y2=1.485
cc_168 VPB N_VPWR_c_766_n 0.0108363f $X=-0.19 $Y=1.305 $X2=1.652 $Y2=1.555
cc_169 VPB N_VPWR_c_767_n 0.00438892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_768_n 0.0149751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_769_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.19
cc_172 VPB N_VPWR_c_770_n 0.0193922f $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.19
cc_173 VPB N_VPWR_c_771_n 0.0120373f $X=-0.19 $Y=1.305 $X2=1.655 $Y2=1.19
cc_174 VPB N_VPWR_c_772_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_175 VPB N_VPWR_c_773_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.16
cc_176 VPB N_VPWR_c_774_n 0.0128121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_775_n 0.00584107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_764_n 0.127033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_777_n 0.0129905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_778_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_779_n 0.0120373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_780_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_781_n 0.0149751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_782_n 0.0108363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_783_n 0.00438892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_784_n 0.0103455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_785_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_786_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_787_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_788_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_789_n 0.00487564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_790_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_791_n 0.0375449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_792_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_793_n 0.0212654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_794_n 0.0193922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_795_n 0.0375449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_796_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_797_n 0.00439477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_798_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_799_n 0.00487564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_800_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_801_n 0.00497181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_802_n 0.00497181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_803_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_804_n 0.00439477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_765_n 0.116463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g
+ 0.0225925f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_209 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g
+ 0.0179939f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_210 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ 0.0182972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g
+ 0.0219547f $X=-0.19 $Y=1.305 $X2=1.652 $Y2=0.905
cc_212 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n 0.00561924f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_213 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1186_n 0.00432833f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_214 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n 0.00421086f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_215 VPB N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1196_n 0.00687837f $X=-0.19 $Y=1.305
+ $X2=0 $Y2=0
cc_216 VPB N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g
+ 0.0231079f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_217 VPB N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g
+ 0.0253019f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_218 VPB N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.00677654f $X=-0.19 $Y=1.305
+ $X2=2.14 $Y2=1.62
cc_219 VPB N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n 6.96869e-19 $X=-0.19 $Y=1.305
+ $X2=1.315 $Y2=1.19
cc_220 VPB N_SKY130_FD_SC_HD__INV_2_0/A_c_1346_n 0.00439746f $X=-0.19 $Y=1.305
+ $X2=1.17 $Y2=1.19
cc_221 VPB N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n 0.00130257f $X=-0.19 $Y=1.305
+ $X2=1.655 $Y2=1.19
cc_222 VPB N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n 0.0151211f $X=-0.19 $Y=1.305
+ $X2=1.11 $Y2=1.16
cc_223 VPB N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.00151227f $X=-0.19 $Y=1.305
+ $X2=0.9 $Y2=1.325
cc_224 VPB N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1483_n 0.00644428f $X=-0.19
+ $Y=1.305 $X2=0.48 $Y2=0.56
cc_225 VPB N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1484_n 0.0026524f $X=-0.19
+ $Y=1.305 $X2=0.48 $Y2=1.985
cc_226 VPB N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1485_n 0.00153792f $X=-0.19
+ $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.00265353f $X=-0.19
+ $Y=1.305 $X2=0.9 $Y2=0.56
cc_228 VPB N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n 0.00419803f $X=-0.19
+ $Y=1.305 $X2=0.9 $Y2=1.325
cc_229 VPB N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1488_n 0.00972405f $X=-0.19
+ $Y=1.305 $X2=0.9 $Y2=1.985
cc_230 VPB N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n 0.00419803f $X=-0.19
+ $Y=1.305 $X2=0.48 $Y2=0.995
cc_231 VPB N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1532_n 0.00972405f $X=-0.19
+ $Y=1.305 $X2=0.48 $Y2=0.56
cc_232 VPB N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00265432f $X=-0.19
+ $Y=1.305 $X2=0.48 $Y2=1.985
cc_233 VPB N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1534_n 0.00153792f $X=-0.19
+ $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.0026524f $X=-0.19
+ $Y=1.305 $X2=0.9 $Y2=0.56
cc_235 VPB N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1536_n 0.00652051f $X=-0.19
+ $Y=1.305 $X2=0.9 $Y2=1.985
cc_236 VPB N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.00151227f $X=-0.19 $Y=1.305
+ $X2=0.9 $Y2=1.325
cc_237 N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n 0.0108204f $X=1.975 $Y=0.82 $X2=0 $Y2=0
cc_238 N_SKY130_FD_SC_HD__INV_2_1/A_c_259_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n 0.0109314f $X=2.14 $Y=0.39 $X2=0 $Y2=0
cc_239 N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n 0.00158032f $X=2.14 $Y=0.815 $X2=0 $Y2=0
cc_240 N_SKY130_FD_SC_HD__INV_2_1/A_c_249_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n 0.0140806f $X=1.655 $Y=1.19 $X2=0 $Y2=0
cc_241 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g 0.0254664f
+ $X=2.14 $Y=1.62 $X2=0 $Y2=0
cc_242 N_SKY130_FD_SC_HD__INV_2_1/A_c_259_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n 0.00630972f $X=2.14 $Y=0.39 $X2=0 $Y2=0
cc_243 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n 0.00864955f $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_244 N_SKY130_FD_SC_HD__INV_2_1/A_c_265_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n 5.22228e-19 $X=2.98 $Y=0.39 $X2=0 $Y2=0
cc_245 N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n 0.00111672f $X=2.14 $Y=0.815 $X2=0 $Y2=0
cc_246 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g 0.00856424f
+ $X=2.14 $Y=1.62 $X2=0 $Y2=0
cc_247 N_SKY130_FD_SC_HD__INV_2_1/A_c_259_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n 5.22228e-19 $X=2.14 $Y=0.39 $X2=0 $Y2=0
cc_248 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n 0.0112985f $X=2.815 $Y=0.815 $X2=0 $Y2=0
cc_249 N_SKY130_FD_SC_HD__INV_2_1/A_c_265_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n 0.00630972f $X=2.98 $Y=0.39 $X2=0 $Y2=0
cc_250 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n 0.00261194f $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_251 N_SKY130_FD_SC_HD__INV_2_1/A_c_265_p
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n 0.00539651f $X=2.98 $Y=0.39 $X2=0 $Y2=0
cc_252 N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.00305484f $X=1.975 $Y=0.82 $X2=0 $Y2=0
cc_253 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.0266973f $X=2.815 $Y=0.815 $X2=0 $Y2=0
cc_254 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.0246539f $X=2.14 $Y=1.62 $X2=0 $Y2=0
cc_255 N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.023675f $X=2.14 $Y=0.815 $X2=0 $Y2=0
cc_256 N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.00178057f $X=1.655 $Y=1.19 $X2=0 $Y2=0
cc_257 N_SKY130_FD_SC_HD__INV_2_1/A_c_249_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n 0.0137365f $X=1.655 $Y=1.19 $X2=0 $Y2=0
cc_258 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_362_n 0.0193224f $X=2.815 $Y=0.815 $X2=0 $Y2=0
cc_259 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_400_n 0.00696298f $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_260 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_401_n 5.78068e-19 $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_261 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_401_n 0.00654189f $X=2.14 $Y=1.62 $X2=0 $Y2=0
cc_262 N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_401_n 0.00649173f $X=2.14 $Y=0.815 $X2=0 $Y2=0
cc_263 N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_401_n 0.0189613f $X=1.655 $Y=1.19 $X2=0 $Y2=0
cc_264 N_SKY130_FD_SC_HD__INV_2_1/A_c_249_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_401_n 3.75211e-19 $X=1.655 $Y=1.19 $X2=0 $Y2=0
cc_265 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_406_n 0.00600063f $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_266 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n 0.00215368f $X=2.14 $Y=1.62 $X2=0 $Y2=0
cc_267 N_SKY130_FD_SC_HD__INV_2_1/A_c_244_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n 0.00230339f $X=2.14 $Y=0.815 $X2=0 $Y2=0
cc_268 N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n 0.00234275f $X=1.655 $Y=1.19 $X2=0 $Y2=0
cc_269 N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_366_n 0.00478049f $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_270 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_c_367_n 0.00230339f $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_271 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_VPWR_c_767_n 0.0031902f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_272 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_VPWR_c_768_n 0.00320188f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_273 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n N_VPWR_c_768_n 0.0100425f $X=2.14
+ $Y=1.62 $X2=0 $Y2=0
cc_274 N_SKY130_FD_SC_HD__INV_2_1/A_c_245_n N_VPWR_c_768_n 0.0164326f $X=1.15
+ $Y=1.19 $X2=0 $Y2=0
cc_275 N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n N_VPWR_c_768_n 0.00184934f $X=1.315
+ $Y=1.19 $X2=0 $Y2=0
cc_276 N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n N_VPWR_c_768_n 0.00529313f $X=1.11
+ $Y=1.16 $X2=0 $Y2=0
cc_277 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_VPWR_c_790_n 0.00541359f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_278 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_VPWR_c_790_n 0.00541359f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_279 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1005_s
+ N_VPWR_c_765_n 0.00216833f $X=2.005 $Y=1.485 $X2=0 $Y2=0
cc_280 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_VPWR_c_765_n 0.0104652f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_281 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_VPWR_c_765_n 0.0108276f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_282 N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1001_s 3.93288e-19 $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_283 N_SKY130_FD_SC_HD__INV_2_1/A_c_242_n
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1001_s 0.00248165f $X=1.76 $Y=0.82 $X2=0
+ $Y2=0
cc_284 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1002_s 0.00162089f $X=2.815 $Y=0.815 $X2=0
+ $Y2=0
cc_285 N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n N_VGND_c_963_n 0.00363144f $X=0.48
+ $Y=0.995 $X2=0 $Y2=0
cc_286 N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n N_VGND_c_964_n 0.00366806f $X=0.9
+ $Y=0.995 $X2=0 $Y2=0
cc_287 N_SKY130_FD_SC_HD__INV_2_1/A_c_242_n N_VGND_c_964_n 0.0101019f $X=1.76
+ $Y=0.82 $X2=0 $Y2=0
cc_288 N_SKY130_FD_SC_HD__INV_2_1/A_c_245_n N_VGND_c_964_n 0.0161043f $X=1.15
+ $Y=1.19 $X2=0 $Y2=0
cc_289 N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n N_VGND_c_964_n 0.00560615f $X=1.315
+ $Y=1.19 $X2=0 $Y2=0
cc_290 N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n N_VGND_c_964_n 0.00585411f $X=1.11
+ $Y=1.16 $X2=0 $Y2=0
cc_291 N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n N_VGND_c_966_n 0.00268399f $X=1.975
+ $Y=0.82 $X2=0 $Y2=0
cc_292 N_SKY130_FD_SC_HD__INV_2_1/A_c_242_n N_VGND_c_966_n 0.0172644f $X=1.76
+ $Y=0.82 $X2=0 $Y2=0
cc_293 N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n N_VGND_c_966_n 0.00217186f $X=1.655
+ $Y=1.19 $X2=0 $Y2=0
cc_294 N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n N_VGND_c_967_n 0.00193763f $X=1.975
+ $Y=0.82 $X2=0 $Y2=0
cc_295 N_SKY130_FD_SC_HD__INV_2_1/A_c_259_p N_VGND_c_967_n 0.0188551f $X=2.14
+ $Y=0.39 $X2=0 $Y2=0
cc_296 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n N_VGND_c_967_n 0.00198695f $X=2.815
+ $Y=0.815 $X2=0 $Y2=0
cc_297 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n N_VGND_c_968_n 0.0118745f $X=2.815
+ $Y=0.815 $X2=0 $Y2=0
cc_298 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n N_VGND_c_969_n 0.00835456f $X=2.815
+ $Y=0.815 $X2=0 $Y2=0
cc_299 N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n N_VGND_c_985_n 0.00541359f $X=0.48
+ $Y=0.995 $X2=0 $Y2=0
cc_300 N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n N_VGND_c_985_n 0.00541359f $X=0.9
+ $Y=0.995 $X2=0 $Y2=0
cc_301 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n N_VGND_c_986_n 0.00198695f $X=2.815
+ $Y=0.815 $X2=0 $Y2=0
cc_302 N_SKY130_FD_SC_HD__INV_2_1/A_c_265_p N_VGND_c_986_n 0.0188551f $X=2.98
+ $Y=0.39 $X2=0 $Y2=0
cc_303 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1001_d
+ N_VGND_c_1001_n 0.00215201f $X=2.005 $Y=0.235 $X2=0 $Y2=0
cc_304 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1003_d
+ N_VGND_c_1001_n 0.00215201f $X=2.845 $Y=0.235 $X2=0 $Y2=0
cc_305 N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n N_VGND_c_1001_n 0.0104652f $X=0.48
+ $Y=0.995 $X2=0 $Y2=0
cc_306 N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n N_VGND_c_1001_n 0.0108276f $X=0.9
+ $Y=0.995 $X2=0 $Y2=0
cc_307 N_SKY130_FD_SC_HD__INV_2_1/A_c_241_n N_VGND_c_1001_n 0.00398137f $X=1.975
+ $Y=0.82 $X2=0 $Y2=0
cc_308 N_SKY130_FD_SC_HD__INV_2_1/A_c_242_n N_VGND_c_1001_n 9.4368e-19 $X=1.76
+ $Y=0.82 $X2=0 $Y2=0
cc_309 N_SKY130_FD_SC_HD__INV_2_1/A_c_259_p N_VGND_c_1001_n 0.0122069f $X=2.14
+ $Y=0.39 $X2=0 $Y2=0
cc_310 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n N_VGND_c_1001_n 0.00835832f $X=2.815
+ $Y=0.815 $X2=0 $Y2=0
cc_311 N_SKY130_FD_SC_HD__INV_2_1/A_c_265_p N_VGND_c_1001_n 0.0122069f $X=2.98
+ $Y=0.39 $X2=0 $Y2=0
cc_312 N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1459_n 0.00534153f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_313 N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1459_n 0.00534153f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_314 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1461_n 0.00918977f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_315 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1461_n 0.00918977f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_316 N_SKY130_FD_SC_HD__INV_2_1/A_c_239_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.00675111f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_317 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.00809641f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_318 N_SKY130_FD_SC_HD__INV_2_1/A_c_240_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.004954f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_319 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.00408533f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_320 N_SKY130_FD_SC_HD__INV_2_1/A_c_245_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.0156717f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_321 N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 3.89584e-19 $X=1.315 $Y=1.19 $X2=0 $Y2=0
cc_322 N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.0259992f $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_323 N_SKY130_FD_SC_HD__INV_2_1/A_c_245_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1470_n 0.00153058f $X=1.15 $Y=1.19 $X2=0 $Y2=0
cc_324 N_SKY130_FD_SC_HD__INV_2_1/A_c_247_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1470_n 0.0229882f $X=1.315 $Y=1.19 $X2=0 $Y2=0
cc_325 N_SKY130_FD_SC_HD__INV_2_1/A_c_250_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1470_n 0.0151782f $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_326 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1473_n 0.00214168f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_327 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_c_1473_n 0.00280787f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_328 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1005_d
+ 0.00296777f $X=2.14 $Y=1.62 $X2=-0.19 $Y2=-0.24
cc_329 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1483_n 0.0202286f $X=2.14 $Y=1.62
+ $X2=0 $Y2=0
cc_330 N_SKY130_FD_SC_HD__INV_2_1/A_c_248_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1483_n 0.00137335f $X=1.655 $Y=1.19
+ $X2=0 $Y2=0
cc_331 N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1005_s
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n 0.00312348f $X=2.005 $Y=1.485
+ $X2=0 $Y2=0
cc_332 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n 0.0183094f $X=2.14 $Y=1.62
+ $X2=0 $Y2=0
cc_333 N_SKY130_FD_SC_HD__INV_2_1/A_c_253_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1485_n 0.0102037f $X=2.14 $Y=1.62
+ $X2=0 $Y2=0
cc_334 N_SKY130_FD_SC_HD__INV_2_1/A_c_243_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.00202726f $X=2.815 $Y=0.815
+ $X2=0 $Y2=0
cc_335 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n N_LO_c_513_n 0.0137866f $X=4.46
+ $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_336 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_363_n N_LO_c_513_n 0.0198667f $X=3.905
+ $Y=0.835 $X2=-0.19 $Y2=-0.24
cc_337 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_414_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g 0.0129153f $X=4.295 $Y=1.58 $X2=0
+ $Y2=0
cc_338 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_415_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g 0.0145598f $X=4.46 $Y=2.34 $X2=0
+ $Y2=0
cc_339 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_416_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g 8.84614e-19 $X=4.46 $Y=1.66 $X2=0
+ $Y2=0
cc_340 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n N_LO_c_514_n 0.00382511f $X=4.46
+ $Y=0.74 $X2=0 $Y2=0
cc_341 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_415_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g 0.00975139f $X=4.46 $Y=2.34 $X2=0
+ $Y2=0
cc_342 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g 0.0107043f $X=5.135 $Y=1.58 $X2=0
+ $Y2=0
cc_343 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_420_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g 6.1949e-19 $X=5.3 $Y=2.34 $X2=0 $Y2=0
cc_344 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_416_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g 8.84614e-19 $X=4.46 $Y=1.66 $X2=0
+ $Y2=0
cc_345 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_415_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g 6.1949e-19 $X=4.46 $Y=2.34 $X2=0
+ $Y2=0
cc_346 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g 0.0120619f $X=5.135 $Y=1.58 $X2=0
+ $Y2=0
cc_347 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_424_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g 8.72449e-19 $X=5.3 $Y=1.665 $X2=0
+ $Y2=0
cc_348 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_420_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g 0.00975139f $X=5.3 $Y=2.34 $X2=0
+ $Y2=0
cc_349 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_424_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g 0.00224191f $X=5.3 $Y=1.665 $X2=0
+ $Y2=0
cc_350 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_420_p
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g 0.00882321f $X=5.3 $Y=2.34 $X2=0
+ $Y2=0
cc_351 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n N_LO_c_521_n 0.0305541f $X=4.46
+ $Y=0.74 $X2=0 $Y2=0
cc_352 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_414_p N_LO_c_521_n 0.00555408f $X=4.295
+ $Y=1.58 $X2=0 $Y2=0
cc_353 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p N_LO_c_521_n 0.0215822f $X=5.135
+ $Y=1.58 $X2=0 $Y2=0
cc_354 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_416_p N_LO_c_521_n 0.0213676f $X=4.46
+ $Y=1.66 $X2=0 $Y2=0
cc_355 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_363_n N_LO_c_521_n 0.0176457f $X=3.905
+ $Y=0.835 $X2=0 $Y2=0
cc_356 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n N_LO_c_521_n 0.00733902f $X=3.905
+ $Y=1.19 $X2=0 $Y2=0
cc_357 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_424_p N_LO_c_522_n 0.0198347f $X=5.3
+ $Y=1.665 $X2=0 $Y2=0
cc_358 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p N_LO_c_583_n 0.00311669f $X=5.135
+ $Y=1.58 $X2=0 $Y2=0
cc_359 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_424_p N_LO_c_583_n 0.00238622f $X=5.3
+ $Y=1.665 $X2=0 $Y2=0
cc_360 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p N_LO_c_524_n 0.00309698f $X=5.135
+ $Y=1.58 $X2=0 $Y2=0
cc_361 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n N_LO_c_533_n 0.00223984f $X=4.46
+ $Y=0.74 $X2=0 $Y2=0
cc_362 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_416_p N_LO_c_533_n 0.00209661f $X=4.46
+ $Y=1.66 $X2=0 $Y2=0
cc_363 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n N_LO_c_533_n 0.00753014f $X=3.905
+ $Y=1.19 $X2=0 $Y2=0
cc_364 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_424_p N_LO_c_534_n 0.00209661f $X=5.3
+ $Y=1.665 $X2=0 $Y2=0
cc_365 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_414_p
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1000_s 0.00202414f $X=4.295 $Y=1.58 $X2=0
+ $Y2=0
cc_366 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_377_n
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1000_s 0.00218031f $X=3.905 $Y=1.495 $X2=0
+ $Y2=0
cc_367 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1001_s 0.00317613f $X=5.135 $Y=1.58 $X2=0
+ $Y2=0
cc_368 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ N_VPWR_c_768_n 0.00680156f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_369 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_VPWR_c_769_n 0.00110007f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_370 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ N_VPWR_c_769_n 0.0122133f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_371 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_VPWR_c_769_n 0.0129672f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_372 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_VPWR_c_770_n 0.0046653f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_373 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_VPWR_c_771_n 0.00299545f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_374 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_414_p N_VPWR_c_771_n 0.00588864f $X=4.295
+ $Y=1.58 $X2=0 $Y2=0
cc_375 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n N_VPWR_c_771_n 7.43608e-19 $X=3.905
+ $Y=1.19 $X2=0 $Y2=0
cc_376 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_377_n N_VPWR_c_771_n 0.0153103f $X=3.905
+ $Y=1.495 $X2=0 $Y2=0
cc_377 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_415_p N_VPWR_c_772_n 0.0189039f $X=4.46
+ $Y=2.34 $X2=0 $Y2=0
cc_378 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p N_VPWR_c_773_n 0.0122533f $X=5.135
+ $Y=1.58 $X2=0 $Y2=0
cc_379 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ N_VPWR_c_791_n 0.00357877f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_380 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_VPWR_c_791_n 0.00357877f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_381 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ N_VPWR_c_791_n 0.0046653f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_382 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_420_p N_VPWR_c_792_n 0.0189039f $X=5.3
+ $Y=2.34 $X2=0 $Y2=0
cc_383 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1000_d
+ N_VPWR_c_765_n 0.00215201f $X=4.325 $Y=1.485 $X2=0 $Y2=0
cc_384 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1005_d
+ N_VPWR_c_765_n 0.00215201f $X=5.165 $Y=1.485 $X2=0 $Y2=0
cc_385 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ N_VPWR_c_765_n 0.00655123f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_386 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_VPWR_c_765_n 0.00522516f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_387 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ N_VPWR_c_765_n 0.00789179f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_388 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_VPWR_c_765_n 0.00921786f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_389 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_415_p N_VPWR_c_765_n 0.0122217f $X=4.46
+ $Y=2.34 $X2=0 $Y2=0
cc_390 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_420_p N_VPWR_c_765_n 0.0122217f $X=5.3
+ $Y=2.34 $X2=0 $Y2=0
cc_391 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n N_VGND_c_964_n 0.00503112f $X=1.93
+ $Y=0.995 $X2=0 $Y2=0
cc_392 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n N_VGND_c_966_n 0.0032322f $X=1.93
+ $Y=0.995 $X2=0 $Y2=0
cc_393 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n N_VGND_c_967_n 0.00424416f $X=1.93
+ $Y=0.995 $X2=0 $Y2=0
cc_394 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n N_VGND_c_967_n 0.00423334f $X=2.35
+ $Y=0.995 $X2=0 $Y2=0
cc_395 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n N_VGND_c_968_n 0.00146448f $X=2.35
+ $Y=0.995 $X2=0 $Y2=0
cc_396 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n N_VGND_c_968_n 0.00146448f $X=2.77
+ $Y=0.995 $X2=0 $Y2=0
cc_397 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n N_VGND_c_969_n 0.00366968f $X=3.19
+ $Y=0.995 $X2=0 $Y2=0
cc_398 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_362_n N_VGND_c_969_n 0.0211459f $X=2.985
+ $Y=1.19 $X2=0 $Y2=0
cc_399 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_364_n N_VGND_c_969_n 0.0021114f $X=3.76
+ $Y=1.19 $X2=0 $Y2=0
cc_400 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n N_VGND_c_969_n 0.0213859f $X=3.905
+ $Y=0.905 $X2=0 $Y2=0
cc_401 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n N_VGND_c_986_n 0.00423334f $X=2.77
+ $Y=0.995 $X2=0 $Y2=0
cc_402 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n N_VGND_c_986_n 0.00541359f $X=3.19
+ $Y=0.995 $X2=0 $Y2=0
cc_403 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n N_VGND_c_987_n 0.00214403f $X=3.905
+ $Y=0.905 $X2=0 $Y2=0
cc_404 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1003_s
+ N_VGND_c_1001_n 0.00216833f $X=4.325 $Y=0.235 $X2=0 $Y2=0
cc_405 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_356_n N_VGND_c_1001_n 0.00706214f $X=1.93
+ $Y=0.995 $X2=0 $Y2=0
cc_406 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_357_n N_VGND_c_1001_n 0.0057163f $X=2.35
+ $Y=0.995 $X2=0 $Y2=0
cc_407 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_358_n N_VGND_c_1001_n 0.0057163f $X=2.77
+ $Y=0.995 $X2=0 $Y2=0
cc_408 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_359_n N_VGND_c_1001_n 0.0108276f $X=3.19
+ $Y=0.995 $X2=0 $Y2=0
cc_409 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n N_VGND_c_1001_n 0.00368014f
+ $X=3.905 $Y=0.905 $X2=0 $Y2=0
cc_410 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n 0.00929492f $X=1.93 $Y=1.985
+ $X2=0 $Y2=0
cc_411 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n 0.0112436f $X=2.35 $Y=1.985
+ $X2=0 $Y2=0
cc_412 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1485_n 2.36323e-19 $X=2.35 $Y=1.985
+ $X2=0 $Y2=0
cc_413 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1485_n 0.0124486f $X=2.065 $Y=1.19
+ $X2=0 $Y2=0
cc_414 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_400_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1485_n 0.00142025f $X=2.9 $Y=1.19
+ $X2=0 $Y2=0
cc_415 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.0149365f $X=2.77 $Y=1.985
+ $X2=0 $Y2=0
cc_416 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.013736f $X=3.19 $Y=1.985
+ $X2=0 $Y2=0
cc_417 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_361_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.00362207f $X=2.065 $Y=1.19
+ $X2=0 $Y2=0
cc_418 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_362_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.0268321f $X=2.985 $Y=1.19
+ $X2=0 $Y2=0
cc_419 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_400_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.004896f $X=2.9 $Y=1.19 $X2=0
+ $Y2=0
cc_420 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_364_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 9.00165e-19 $X=3.76 $Y=1.19
+ $X2=0 $Y2=0
cc_421 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_406_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.00708673f $X=3.19 $Y=1.19
+ $X2=0 $Y2=0
cc_422 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_367_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.00213789f $X=3.19 $Y=1.16
+ $X2=0 $Y2=0
cc_423 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_362_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n 0.0201375f $X=2.985 $Y=1.19
+ $X2=0 $Y2=0
cc_424 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_363_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n 0.00338615f $X=3.905 $Y=0.835
+ $X2=0 $Y2=0
cc_425 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_364_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n 0.00229746f $X=3.76 $Y=1.19
+ $X2=0 $Y2=0
cc_426 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_377_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n 0.0156019f $X=3.905 $Y=1.495
+ $X2=0 $Y2=0
cc_427 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1003_d
+ 7.4958e-19 $X=4.46 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_428 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1003_d
+ 0.00241065f $X=3.905 $Y=0.905 $X2=-0.19 $Y2=-0.24
cc_429 N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1003_s
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n 0.00312175f $X=4.325 $Y=0.235
+ $X2=0 $Y2=0
cc_430 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n 0.0192847f $X=4.46 $Y=0.74
+ $X2=0 $Y2=0
cc_431 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 3.07688e-19 $X=5.135 $Y=1.58
+ $X2=0 $Y2=0
cc_432 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_419_p
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 8.34819e-19 $X=5.135 $Y=1.58
+ $X2=0 $Y2=0
cc_433 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_360_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 0.00727582f $X=4.46 $Y=0.74
+ $X2=0 $Y2=0
cc_434 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_365_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 6.02828e-19 $X=3.905 $Y=1.19
+ $X2=0 $Y2=0
cc_435 N_SKY130_FD_SC_HD__NOR2_2_1/B_c_368_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 0.0131928f $X=3.905 $Y=0.905
+ $X2=0 $Y2=0
cc_436 N_LO_c_516_n SKY130_FD_SC_HD__CONB_1_0/HI 0.0189792f $X=5.51 $Y=0.995
+ $X2=0 $Y2=0
cc_437 N_LO_c_522_n SKY130_FD_SC_HD__CONB_1_0/HI 0.0188372f $X=5.745 $Y=1.19
+ $X2=0 $Y2=0
cc_438 N_LO_c_525_n SKY130_FD_SC_HD__CONB_1_0/HI 0.0641014f $X=6.705 $Y=1.19
+ $X2=0 $Y2=0
cc_439 N_LO_c_526_n SKY130_FD_SC_HD__CONB_1_0/HI 0.00278662f $X=5.935 $Y=1.19
+ $X2=0 $Y2=0
cc_440 N_LO_c_528_n SKY130_FD_SC_HD__CONB_1_0/HI 0.00279426f $X=6.995 $Y=1.19
+ $X2=0 $Y2=0
cc_441 N_LO_c_532_n SKY130_FD_SC_HD__CONB_1_0/HI 0.00177247f $X=6.92 $Y=1.995
+ $X2=0 $Y2=0
cc_442 N_LO_c_534_n SKY130_FD_SC_HD__CONB_1_0/HI 0.00419262f $X=5.51 $Y=1.16
+ $X2=0 $Y2=0
cc_443 N_LO_c_538_n SKY130_FD_SC_HD__CONB_1_0/HI 0.0705118f $X=6.85 $Y=1.19
+ $X2=0 $Y2=0
cc_444 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g N_VPWR_c_771_n 0.00321527f
+ $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_445 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g N_VPWR_c_772_n 0.00541359f
+ $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_446 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g N_VPWR_c_772_n 0.00541359f
+ $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_447 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g N_VPWR_c_773_n 0.00146448f
+ $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_448 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g N_VPWR_c_773_n 0.00146448f
+ $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_449 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g N_VPWR_c_774_n 0.00183357f
+ $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_450 N_LO_c_522_n N_VPWR_c_774_n 0.0196879f $X=5.745 $Y=1.19 $X2=0 $Y2=0
cc_451 N_LO_c_526_n N_VPWR_c_774_n 0.00201967f $X=5.935 $Y=1.19 $X2=0 $Y2=0
cc_452 N_LO_c_532_n N_VPWR_c_775_n 0.00431607f $X=6.92 $Y=1.995 $X2=0 $Y2=0
cc_453 N_LO_c_538_n N_VPWR_c_775_n 0.0478402f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_454 N_LO_c_522_n N_VPWR_c_764_n 4.21998e-19 $X=5.745 $Y=1.19 $X2=0 $Y2=0
cc_455 N_LO_c_532_n N_VPWR_c_764_n 0.0921235f $X=6.92 $Y=1.995 $X2=0 $Y2=0
cc_456 N_LO_c_534_n N_VPWR_c_764_n 0.0179366f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_457 N_LO_c_538_n N_VPWR_c_764_n 0.00789999f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_458 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g N_VPWR_c_777_n 0.00183357f
+ $X=7.83 $Y=1.985 $X2=0 $Y2=0
cc_459 N_LO_c_523_n N_VPWR_c_777_n 0.0197828f $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_460 N_LO_c_527_n N_VPWR_c_777_n 8.71532e-19 $X=7.565 $Y=1.19 $X2=0 $Y2=0
cc_461 N_LO_c_530_n N_VPWR_c_777_n 0.00112745f $X=7.855 $Y=1.19 $X2=0 $Y2=0
cc_462 N_LO_c_532_n N_VPWR_c_777_n 0.00656332f $X=6.92 $Y=1.995 $X2=0 $Y2=0
cc_463 N_LO_c_538_n N_VPWR_c_777_n 0.0821969f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_464 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g N_VPWR_c_778_n 0.00146448f
+ $X=8.25 $Y=1.985 $X2=0 $Y2=0
cc_465 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g N_VPWR_c_778_n 0.00146448f
+ $X=8.67 $Y=1.985 $X2=0 $Y2=0
cc_466 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g N_VPWR_c_779_n 0.00321527f
+ $X=9.09 $Y=1.985 $X2=0 $Y2=0
cc_467 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g N_VPWR_c_786_n 0.00541359f
+ $X=7.83 $Y=1.985 $X2=0 $Y2=0
cc_468 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g N_VPWR_c_786_n 0.00541359f
+ $X=8.25 $Y=1.985 $X2=0 $Y2=0
cc_469 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g N_VPWR_c_788_n 0.00541359f
+ $X=8.67 $Y=1.985 $X2=0 $Y2=0
cc_470 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g N_VPWR_c_788_n 0.00541359f
+ $X=9.09 $Y=1.985 $X2=0 $Y2=0
cc_471 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g N_VPWR_c_792_n 0.00541359f
+ $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_472 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g N_VPWR_c_792_n 0.00541359f
+ $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_473 N_LO_c_532_n N_VPWR_c_793_n 0.0114454f $X=6.92 $Y=1.995 $X2=0 $Y2=0
cc_474 N_LO_c_538_n N_VPWR_c_793_n 0.0354508f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_475 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g N_VPWR_c_765_n 0.0108276f
+ $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_476 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g N_VPWR_c_765_n 0.00950154f
+ $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_477 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g N_VPWR_c_765_n 0.00950154f
+ $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_478 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g N_VPWR_c_765_n 0.00999367f
+ $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_479 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g N_VPWR_c_765_n 0.00999669f
+ $X=7.83 $Y=1.985 $X2=0 $Y2=0
cc_480 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g N_VPWR_c_765_n 0.00950154f
+ $X=8.25 $Y=1.985 $X2=0 $Y2=0
cc_481 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g N_VPWR_c_765_n 0.00950154f
+ $X=8.67 $Y=1.985 $X2=0 $Y2=0
cc_482 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g N_VPWR_c_765_n 0.0108276f
+ $X=9.09 $Y=1.985 $X2=0 $Y2=0
cc_483 N_LO_c_532_n N_VPWR_c_765_n 0.0137178f $X=6.92 $Y=1.995 $X2=0 $Y2=0
cc_484 N_LO_c_538_n N_VPWR_c_765_n 0.017754f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_485 N_LO_c_513_n N_VGND_c_969_n 0.00581848f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_486 N_LO_c_515_n N_VGND_c_970_n 0.00268723f $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_487 N_LO_c_516_n N_VGND_c_970_n 0.00268723f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_488 N_LO_c_517_n N_VGND_c_971_n 7.40199e-19 $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_489 N_LO_c_527_n N_VGND_c_971_n 4.96106e-19 $X=7.565 $Y=1.19 $X2=0 $Y2=0
cc_490 N_LO_c_528_n N_VGND_c_971_n 0.00130139f $X=6.995 $Y=1.19 $X2=0 $Y2=0
cc_491 N_LO_c_538_n N_VGND_c_971_n 0.0270844f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_492 N_LO_c_517_n N_VGND_c_972_n 0.0151826f $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_493 N_LO_c_523_n N_VGND_c_972_n 3.2733e-19 $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_494 N_LO_c_538_n N_VGND_c_972_n 0.0262939f $X=6.85 $Y=1.19 $X2=0 $Y2=0
cc_495 N_LO_c_517_n N_VGND_c_973_n 0.00268723f $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_496 N_LO_c_518_n N_VGND_c_973_n 0.00268723f $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_497 N_LO_c_520_n N_VGND_c_974_n 0.00581848f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_498 N_LO_c_516_n N_VGND_c_981_n 0.00422241f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_499 N_LO_c_513_n N_VGND_c_987_n 0.00357877f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_500 N_LO_c_514_n N_VGND_c_987_n 0.00357877f $X=4.67 $Y=0.995 $X2=0 $Y2=0
cc_501 N_LO_c_515_n N_VGND_c_987_n 0.00420723f $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_502 N_LO_c_517_n N_VGND_c_988_n 0.00422241f $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_503 N_LO_c_518_n N_VGND_c_989_n 0.00420723f $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_504 N_LO_c_519_n N_VGND_c_989_n 0.00357877f $X=8.67 $Y=0.995 $X2=0 $Y2=0
cc_505 N_LO_c_520_n N_VGND_c_989_n 0.00357877f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_506 N_LO_c_513_n N_VGND_c_1001_n 0.00655123f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_507 N_LO_c_514_n N_VGND_c_1001_n 0.00522516f $X=4.67 $Y=0.995 $X2=0 $Y2=0
cc_508 N_LO_c_515_n N_VGND_c_1001_n 0.00570563f $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_509 N_LO_c_516_n N_VGND_c_1001_n 0.00618869f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_510 N_LO_c_517_n N_VGND_c_1001_n 0.00618869f $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_511 N_LO_c_518_n N_VGND_c_1001_n 0.00570563f $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_512 N_LO_c_519_n N_VGND_c_1001_n 0.00522516f $X=8.67 $Y=0.995 $X2=0 $Y2=0
cc_513 N_LO_c_520_n N_VGND_c_1001_n 0.00655123f $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_514 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1197_n 0.00224191f $X=7.83 $Y=1.985 $X2=0
+ $Y2=0
cc_515 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1197_n 8.72449e-19 $X=8.25 $Y=1.985 $X2=0
+ $Y2=0
cc_516 N_LO_c_523_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1197_n 0.0198347f $X=8.055
+ $Y=1.19 $X2=0 $Y2=0
cc_517 N_LO_c_529_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1197_n 0.00238622f $X=8.425
+ $Y=1.19 $X2=0 $Y2=0
cc_518 N_LO_c_535_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1197_n 0.00209661f $X=8.25
+ $Y=1.16 $X2=0 $Y2=0
cc_519 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1202_n 0.00882321f $X=7.83 $Y=1.985 $X2=0
+ $Y2=0
cc_520 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1202_n 0.00975139f $X=8.25 $Y=1.985 $X2=0
+ $Y2=0
cc_521 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1202_n 6.1949e-19 $X=8.67 $Y=1.985 $X2=0 $Y2=0
cc_522 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.0120619f $X=8.25 $Y=1.985 $X2=0 $Y2=0
cc_523 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.0106611f $X=8.67 $Y=1.985 $X2=0 $Y2=0
cc_524 N_LO_c_529_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.00461219f $X=8.425
+ $Y=1.19 $X2=0 $Y2=0
cc_525 N_LO_c_531_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.00203861f $X=8.57
+ $Y=1.19 $X2=0 $Y2=0
cc_526 N_LO_c_536_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.0210625f $X=8.88
+ $Y=1.16 $X2=0 $Y2=0
cc_527 N_LO_c_519_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n 0.00382511f $X=8.67
+ $Y=0.995 $X2=0 $Y2=0
cc_528 N_LO_c_520_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n 0.0137866f $X=9.09
+ $Y=0.995 $X2=0 $Y2=0
cc_529 N_LO_c_536_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n 0.0305541f $X=8.88
+ $Y=1.16 $X2=0 $Y2=0
cc_530 N_LO_c_537_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n 0.00223984f $X=9.09
+ $Y=1.16 $X2=0 $Y2=0
cc_531 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1214_n 6.1949e-19 $X=8.25 $Y=1.985 $X2=0 $Y2=0
cc_532 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1214_n 0.00975139f $X=8.67 $Y=1.985 $X2=0
+ $Y2=0
cc_533 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1214_n 0.0145598f $X=9.09 $Y=1.985 $X2=0 $Y2=0
cc_534 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1217_n 0.0129153f $X=9.09 $Y=1.985 $X2=0 $Y2=0
cc_535 N_LO_c_536_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1217_n 0.00555408f $X=8.88
+ $Y=1.16 $X2=0 $Y2=0
cc_536 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1219_n 8.84614e-19 $X=8.67 $Y=1.985 $X2=0
+ $Y2=0
cc_537 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1219_n 8.84614e-19 $X=9.09 $Y=1.985 $X2=0
+ $Y2=0
cc_538 N_LO_c_536_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1219_n 0.0213676f $X=8.88
+ $Y=1.16 $X2=0 $Y2=0
cc_539 N_LO_c_537_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1219_n 0.00209661f $X=9.09
+ $Y=1.16 $X2=0 $Y2=0
cc_540 N_LO_c_520_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n 0.0198667f $X=9.09
+ $Y=0.995 $X2=0 $Y2=0
cc_541 N_LO_c_531_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n 4.62104e-19 $X=8.57
+ $Y=1.19 $X2=0 $Y2=0
cc_542 N_LO_c_536_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n 0.0176283f $X=8.88
+ $Y=1.16 $X2=0 $Y2=0
cc_543 N_LO_c_536_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1185_n 0.00738035f $X=8.88
+ $Y=1.16 $X2=0 $Y2=0
cc_544 N_LO_c_537_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1185_n 0.00755246f $X=9.09
+ $Y=1.16 $X2=0 $Y2=0
cc_545 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1487_n 6.56838e-19 $X=4.25 $Y=1.985
+ $X2=0 $Y2=0
cc_546 N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1488_n 0.00482016f $X=4.25 $Y=1.985
+ $X2=0 $Y2=0
cc_547 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n 6.56838e-19 $X=9.09 $Y=1.985
+ $X2=0 $Y2=0
cc_548 N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1532_n 0.00482016f $X=9.09 $Y=1.985
+ $X2=0 $Y2=0
cc_549 N_LO_c_513_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n 0.00750429f
+ $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_550 N_LO_c_514_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n 0.0103415f
+ $X=4.67 $Y=0.995 $X2=0 $Y2=0
cc_551 N_LO_c_521_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n 0.00299901f
+ $X=4.825 $Y=1.19 $X2=0 $Y2=0
cc_552 N_LO_c_524_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1611_n 0.00151741f
+ $X=5.005 $Y=1.19 $X2=0 $Y2=0
cc_553 N_LO_c_515_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1622_n 0.00244813f
+ $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_554 N_LO_c_515_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 0.0049983f
+ $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_555 N_LO_c_516_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 4.58193e-19
+ $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_556 N_LO_c_521_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 0.0104608f
+ $X=4.825 $Y=1.19 $X2=0 $Y2=0
cc_557 N_LO_c_583_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 0.00105162f
+ $X=5.645 $Y=1.19 $X2=0 $Y2=0
cc_558 N_LO_c_524_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1605_n 0.00618556f
+ $X=5.005 $Y=1.19 $X2=0 $Y2=0
cc_559 N_LO_c_515_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.00945687f
+ $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_560 N_LO_c_516_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.00931947f
+ $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_561 N_LO_c_522_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0420214f
+ $X=5.745 $Y=1.19 $X2=0 $Y2=0
cc_562 N_LO_c_583_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0055921f
+ $X=5.645 $Y=1.19 $X2=0 $Y2=0
cc_563 N_LO_c_526_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.00703017f
+ $X=5.935 $Y=1.19 $X2=0 $Y2=0
cc_564 N_LO_c_534_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.00218981f
+ $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_565 N_LO_c_515_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n 5.19117e-19
+ $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_566 N_LO_c_516_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n 0.00620543f
+ $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_567 N_LO_c_513_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 0.00157861f
+ $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_568 N_LO_c_517_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n 0.00620543f
+ $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_569 N_LO_c_518_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n 5.19117e-19
+ $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_570 N_LO_c_517_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.00843297f
+ $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_571 N_LO_c_518_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.00945687f
+ $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_572 N_LO_c_523_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.0213774f
+ $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_573 N_LO_c_529_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.00448318f
+ $X=8.425 $Y=1.19 $X2=0 $Y2=0
cc_574 N_LO_c_530_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.0015981f
+ $X=7.855 $Y=1.19 $X2=0 $Y2=0
cc_575 N_LO_c_535_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.00218981f
+ $X=8.25 $Y=1.16 $X2=0 $Y2=0
cc_576 N_LO_c_517_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n 8.76612e-19
+ $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_577 N_LO_c_523_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n 0.0205585f
+ $X=8.055 $Y=1.19 $X2=0 $Y2=0
cc_578 N_LO_c_527_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n 9.16516e-19
+ $X=7.565 $Y=1.19 $X2=0 $Y2=0
cc_579 N_LO_c_530_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n 0.00604792f
+ $X=7.855 $Y=1.19 $X2=0 $Y2=0
cc_580 N_LO_c_518_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1670_n 0.00244813f
+ $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_581 N_LO_c_517_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 4.58193e-19
+ $X=7.83 $Y=0.995 $X2=0 $Y2=0
cc_582 N_LO_c_518_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 0.0049983f
+ $X=8.25 $Y=0.995 $X2=0 $Y2=0
cc_583 N_LO_c_529_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 0.00269701f
+ $X=8.425 $Y=1.19 $X2=0 $Y2=0
cc_584 N_LO_c_531_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 0.00337445f
+ $X=8.57 $Y=1.19 $X2=0 $Y2=0
cc_585 N_LO_c_536_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 0.0107404f
+ $X=8.88 $Y=1.16 $X2=0 $Y2=0
cc_586 N_LO_c_520_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n 0.00157861f
+ $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_587 N_LO_c_519_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.0102965f
+ $X=8.67 $Y=0.995 $X2=0 $Y2=0
cc_588 N_LO_c_520_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.00750429f
+ $X=9.09 $Y=0.995 $X2=0 $Y2=0
cc_589 N_LO_c_531_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.00298747f
+ $X=8.57 $Y=1.19 $X2=0 $Y2=0
cc_590 N_LO_c_536_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.00187885f
+ $X=8.88 $Y=1.16 $X2=0 $Y2=0
cc_591 SKY130_FD_SC_HD__CONB_1_0/HI N_VPWR_c_774_n 0.0207611f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_592 SKY130_FD_SC_HD__CONB_1_0/HI N_VPWR_c_775_n 0.0279374f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_593 SKY130_FD_SC_HD__CONB_1_0/HI N_VPWR_c_764_n 0.0425229f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_594 SKY130_FD_SC_HD__CONB_1_0/HI N_VGND_c_971_n 0.0464596f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_595 SKY130_FD_SC_HD__CONB_1_0/HI N_VGND_c_972_n 0.0757432f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_596 SKY130_FD_SC_HD__CONB_1_0/HI N_VGND_c_981_n 0.0468962f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_597 SKY130_FD_SC_HD__CONB_1_0/HI N_VGND_c_1001_n 0.031487f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_598 SKY130_FD_SC_HD__CONB_1_0/HI
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0162853f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_599 SKY130_FD_SC_HD__CONB_1_0/HI
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n 0.0415033f $X=6.325 $Y=1.16
+ $X2=0 $Y2=0
cc_600 N_VPWR_c_767_n N_VGND_c_963_n 0.00765463f $X=0.27 $Y=1.66 $X2=0 $Y2=0
cc_601 N_VPWR_c_783_n N_VGND_c_980_n 0.00765463f $X=13.07 $Y=1.66 $X2=0 $Y2=0
cc_602 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1000_d 0.00215201f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_603 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1005_d 0.00215201f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_604 N_VPWR_c_779_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g 0.00299545f
+ $X=9.3 $Y=2 $X2=0 $Y2=0
cc_605 N_VPWR_c_780_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g 0.0129672f
+ $X=10.36 $Y=2 $X2=0 $Y2=0
cc_606 N_VPWR_c_794_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g 0.0046653f
+ $X=10.195 $Y=2.72 $X2=0 $Y2=0
cc_607 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g 0.00921786f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_608 N_VPWR_c_780_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g 0.0122133f
+ $X=10.36 $Y=2 $X2=0 $Y2=0
cc_609 N_VPWR_c_795_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g 0.0046653f
+ $X=12.085 $Y=2.72 $X2=0 $Y2=0
cc_610 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g 0.00789179f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_611 N_VPWR_c_780_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g 0.00110007f
+ $X=10.36 $Y=2 $X2=0 $Y2=0
cc_612 N_VPWR_c_795_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g 0.00357877f
+ $X=12.085 $Y=2.72 $X2=0 $Y2=0
cc_613 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g 0.00522516f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_614 N_VPWR_c_781_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g 0.00680156f
+ $X=12.23 $Y=1.66 $X2=0 $Y2=0
cc_615 N_VPWR_c_795_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g 0.00357877f
+ $X=12.085 $Y=2.72 $X2=0 $Y2=0
cc_616 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g 0.00655123f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_617 N_VPWR_c_786_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1202_n 0.0189039f $X=8.375
+ $Y=2.72 $X2=0 $Y2=0
cc_618 N_VPWR_c_765_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1202_n 0.0122217f $X=13.11
+ $Y=2.72 $X2=0 $Y2=0
cc_619 N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1001_s
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.00318167f $X=8.325 $Y=1.485 $X2=0
+ $Y2=0
cc_620 N_VPWR_c_778_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n 0.012272f $X=8.46
+ $Y=2 $X2=0 $Y2=0
cc_621 N_VPWR_c_788_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1214_n 0.0189039f $X=9.215
+ $Y=2.72 $X2=0 $Y2=0
cc_622 N_VPWR_c_765_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1214_n 0.0122217f $X=13.11
+ $Y=2.72 $X2=0 $Y2=0
cc_623 N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1006_s
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1217_n 0.00207121f $X=9.165 $Y=1.485 $X2=0
+ $Y2=0
cc_624 N_VPWR_c_779_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1217_n 0.00587458f $X=9.3
+ $Y=2 $X2=0 $Y2=0
cc_625 N_VPWR_c_779_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1185_n 7.53817e-19 $X=9.3
+ $Y=2 $X2=0 $Y2=0
cc_626 N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1006_s
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1196_n 0.00218031f $X=9.165 $Y=1.485 $X2=0
+ $Y2=0
cc_627 N_VPWR_c_779_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1196_n 0.0153103f $X=9.3
+ $Y=2 $X2=0 $Y2=0
cc_628 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_s 0.00216833f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_629 N_VPWR_c_781_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g 0.00320188f
+ $X=12.23 $Y=1.66 $X2=0 $Y2=0
cc_630 N_VPWR_c_796_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g 0.00541359f
+ $X=12.985 $Y=2.72 $X2=0 $Y2=0
cc_631 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g 0.0108276f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_632 N_VPWR_c_783_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g 0.0031902f
+ $X=13.07 $Y=1.66 $X2=0 $Y2=0
cc_633 N_VPWR_c_796_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g 0.00541359f
+ $X=12.985 $Y=2.72 $X2=0 $Y2=0
cc_634 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g 0.0104652f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_635 N_VPWR_c_781_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.0100425f $X=12.23
+ $Y=1.66 $X2=0 $Y2=0
cc_636 N_VPWR_c_781_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1343_n 0.0164326f $X=12.23
+ $Y=1.66 $X2=0 $Y2=0
cc_637 N_VPWR_c_781_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n 0.00184934f $X=12.23
+ $Y=1.66 $X2=0 $Y2=0
cc_638 N_VPWR_c_781_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n 0.00529313f $X=12.23
+ $Y=1.66 $X2=0 $Y2=0
cc_639 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1000_s 0.00215201f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_640 N_VPWR_c_790_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1461_n 0.0189039f $X=1.025
+ $Y=2.72 $X2=0 $Y2=0
cc_641 N_VPWR_c_765_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1461_n 0.0122217f $X=13.11
+ $Y=2.72 $X2=0 $Y2=0
cc_642 N_VPWR_c_765_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1005_d
+ 0.00209324f $X=13.11 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_643 N_VPWR_c_765_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1006_d
+ 0.00385313f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_644 N_VPWR_c_765_n
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1007_s
+ 0.00399293f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_645 N_VPWR_c_768_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1483_n 0.0282587f
+ $X=1.11 $Y=1.66 $X2=0 $Y2=0
cc_646 N_VPWR_c_791_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n 0.0358391f
+ $X=2.815 $Y=2.72 $X2=0 $Y2=0
cc_647 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1492_n 0.0234424f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_648 N_VPWR_c_768_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1484_n 0.0111901f
+ $X=1.11 $Y=1.66 $X2=0 $Y2=0
cc_649 N_VPWR_c_791_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1484_n 0.0208596f
+ $X=2.815 $Y=2.72 $X2=0 $Y2=0
cc_650 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1484_n 0.0115253f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_651 N_VPWR_c_791_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1524_n 0.0114668f
+ $X=2.815 $Y=2.72 $X2=0 $Y2=0
cc_652 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1524_n
+ 0.00653655f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_653 N_VPWR_Xsky130_fd_sc_hd__nor2_2_1/M1000_d
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.00166915f $X=2.845 $Y=1.485
+ $X2=0 $Y2=0
cc_654 N_VPWR_c_769_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1486_n 0.0166992f
+ $X=2.98 $Y=2 $X2=0 $Y2=0
cc_655 N_VPWR_c_770_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1488_n 0.019049f
+ $X=3.87 $Y=2.72 $X2=0 $Y2=0
cc_656 N_VPWR_c_771_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1488_n 0.0358806f
+ $X=4.04 $Y=2 $X2=0 $Y2=0
cc_657 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_c_1488_n 0.0105137f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_658 N_VPWR_c_765_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1000_s
+ 0.00399293f $X=13.11 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_659 N_VPWR_c_765_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1007_s
+ 0.00385313f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_660 N_VPWR_c_765_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1006_d
+ 0.00209324f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_661 N_VPWR_c_779_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1532_n 0.0358806f
+ $X=9.3 $Y=2 $X2=0 $Y2=0
cc_662 N_VPWR_c_794_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1532_n 0.019049f
+ $X=10.195 $Y=2.72 $X2=0 $Y2=0
cc_663 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1532_n 0.0105137f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_664 N_VPWR_Xsky130_fd_sc_hd__nor2_2_0/M1000_d
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00166915f $X=10.225 $Y=1.485
+ $X2=0 $Y2=0
cc_665 N_VPWR_c_780_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.0167005f
+ $X=10.36 $Y=2 $X2=0 $Y2=0
cc_666 N_VPWR_c_795_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1547_n 0.0114668f
+ $X=12.085 $Y=2.72 $X2=0 $Y2=0
cc_667 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1547_n
+ 0.00653655f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_668 N_VPWR_c_781_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.0111901f
+ $X=12.23 $Y=1.66 $X2=0 $Y2=0
cc_669 N_VPWR_c_795_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.0566987f
+ $X=12.085 $Y=2.72 $X2=0 $Y2=0
cc_670 N_VPWR_c_765_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.0349677f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_671 N_VPWR_c_781_n N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1536_n 0.0282587f
+ $X=12.23 $Y=1.66 $X2=0 $Y2=0
cc_672 N_VPWR_c_765_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1000_s 0.00215201f
+ $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_673 N_VPWR_c_796_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1582_n 0.0189039f $X=12.985
+ $Y=2.72 $X2=0 $Y2=0
cc_674 N_VPWR_c_765_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1582_n 0.0122217f $X=13.11
+ $Y=2.72 $X2=0 $Y2=0
cc_675 N_VGND_c_1001_n
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1003_s 0.00216833f
+ $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_676 N_VGND_c_974_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n 0.00366968f $X=9.94
+ $Y=0.39 $X2=0 $Y2=0
cc_677 N_VGND_c_983_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n 0.00541359f
+ $X=10.695 $Y=0 $X2=0 $Y2=0
cc_678 N_VGND_c_1001_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n 0.0108276f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_975_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n 0.00146448f
+ $X=10.78 $Y=0.39 $X2=0 $Y2=0
cc_680 N_VGND_c_983_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n 0.00423334f
+ $X=10.695 $Y=0 $X2=0 $Y2=0
cc_681 N_VGND_c_1001_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n 0.0057163f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_975_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n 0.00146448f
+ $X=10.78 $Y=0.39 $X2=0 $Y2=0
cc_683 N_VGND_c_990_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n 0.00423334f
+ $X=11.535 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1001_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n 0.0057163f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_685 N_VGND_c_976_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n 0.0032322f $X=11.62
+ $Y=0.39 $X2=0 $Y2=0
cc_686 N_VGND_c_978_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n 0.00503112f
+ $X=12.23 $Y=0.38 $X2=0 $Y2=0
cc_687 N_VGND_c_990_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n 0.00424416f
+ $X=11.535 $Y=0 $X2=0 $Y2=0
cc_688 N_VGND_c_1001_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n 0.00706214f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_689 N_VGND_c_974_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1182_n 0.0211459f $X=9.94
+ $Y=0.39 $X2=0 $Y2=0
cc_690 N_VGND_c_974_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1184_n 0.0021114f $X=9.94
+ $Y=0.39 $X2=0 $Y2=0
cc_691 N_VGND_c_974_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n 0.0213859f $X=9.94
+ $Y=0.39 $X2=0 $Y2=0
cc_692 N_VGND_c_989_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n 0.00214403f $X=9.75
+ $Y=0 $X2=0 $Y2=0
cc_693 N_VGND_c_1001_n N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n 0.00368014f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_694 N_VGND_c_1001_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1001_d 0.00215201f
+ $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_695 N_VGND_c_1001_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1003_d 0.00215201f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_696 N_VGND_c_978_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n 0.00366806f $X=12.23
+ $Y=0.38 $X2=0 $Y2=0
cc_697 N_VGND_c_991_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n 0.00541359f
+ $X=12.985 $Y=0 $X2=0 $Y2=0
cc_698 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n 0.0108276f $X=13.11
+ $Y=0 $X2=0 $Y2=0
cc_699 N_VGND_c_980_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n 0.00363144f $X=13.07
+ $Y=0.38 $X2=0 $Y2=0
cc_700 N_VGND_c_991_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n 0.00541359f
+ $X=12.985 $Y=0 $X2=0 $Y2=0
cc_701 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n 0.0104652f $X=13.11
+ $Y=0 $X2=0 $Y2=0
cc_702 N_VGND_c_983_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1375_n 0.0188551f $X=10.695
+ $Y=0 $X2=0 $Y2=0
cc_703 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1375_n 0.0122069f $X=13.11
+ $Y=0 $X2=0 $Y2=0
cc_704 N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1002_s
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00162089f $X=10.645 $Y=0.235 $X2=0
+ $Y2=0
cc_705 N_VGND_c_975_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.0118745f $X=10.78
+ $Y=0.39 $X2=0 $Y2=0
cc_706 N_VGND_c_983_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00198695f
+ $X=10.695 $Y=0 $X2=0 $Y2=0
cc_707 N_VGND_c_990_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00198695f
+ $X=11.535 $Y=0 $X2=0 $Y2=0
cc_708 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00835832f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_709 N_VGND_c_974_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00835456f $X=9.94
+ $Y=0.39 $X2=0 $Y2=0
cc_710 N_VGND_c_990_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1383_n 0.0188551f $X=11.535
+ $Y=0 $X2=0 $Y2=0
cc_711 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1383_n 0.0122069f $X=13.11
+ $Y=0 $X2=0 $Y2=0
cc_712 N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1004_s
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.00287493f $X=11.485 $Y=0.235 $X2=0
+ $Y2=0
cc_713 N_VGND_c_976_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.0199581f $X=11.62
+ $Y=0.39 $X2=0 $Y2=0
cc_714 N_VGND_c_978_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.0101019f $X=12.23
+ $Y=0.38 $X2=0 $Y2=0
cc_715 N_VGND_c_990_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.00193763f
+ $X=11.535 $Y=0 $X2=0 $Y2=0
cc_716 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.00492504f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_717 N_VGND_c_978_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1343_n 0.0161043f $X=12.23
+ $Y=0.38 $X2=0 $Y2=0
cc_718 N_VGND_c_976_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n 0.00216104f $X=11.62
+ $Y=0.39 $X2=0 $Y2=0
cc_719 N_VGND_c_978_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n 0.00560615f $X=12.23
+ $Y=0.38 $X2=0 $Y2=0
cc_720 N_VGND_c_978_n N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n 0.00585411f $X=12.23
+ $Y=0.38 $X2=0 $Y2=0
cc_721 N_VGND_c_1001_n
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1001_d 0.00215201f
+ $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_722 N_VGND_c_963_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1459_n 0.025023f $X=0.27
+ $Y=0.38 $X2=0 $Y2=0
cc_723 N_VGND_c_985_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1459_n 0.0188933f $X=1.025
+ $Y=0 $X2=0 $Y2=0
cc_724 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1459_n 0.0122158f $X=13.11
+ $Y=0 $X2=0 $Y2=0
cc_725 N_VGND_c_964_n N_SKY130_FD_SC_HD__INV_2_1/Y_c_1457_n 0.00115029f $X=1.11
+ $Y=0.38 $X2=0 $Y2=0
cc_726 N_VGND_c_1001_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1001_d 0.00215201f
+ $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_727 N_VGND_c_980_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1585_n 0.025023f $X=13.07
+ $Y=0.38 $X2=0 $Y2=0
cc_728 N_VGND_c_991_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1585_n 0.0188933f $X=12.985
+ $Y=0 $X2=0 $Y2=0
cc_729 N_VGND_c_1001_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1585_n 0.0122158f $X=13.11
+ $Y=0 $X2=0 $Y2=0
cc_730 N_VGND_c_978_n N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.00115029f $X=12.23
+ $Y=0.38 $X2=0 $Y2=0
cc_731 N_VGND_c_1001_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1003_d
+ 0.00209344f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_732 N_VGND_c_1001_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1004_d
+ 0.00215206f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_733 N_VGND_c_1001_n
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1007_d
+ 0.00209319f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_734 N_VGND_c_987_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1622_n 0.0151813f
+ $X=5.215 $Y=0 $X2=0 $Y2=0
cc_735 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1622_n
+ 0.0093992f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_736 N_VGND_Xsky130_fd_sc_hd__nand2_2_1/M1002_s
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0030073f $X=5.165 $Y=0.235
+ $X2=0 $Y2=0
cc_737 N_VGND_c_970_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0118126f
+ $X=5.3 $Y=0.38 $X2=0 $Y2=0
cc_738 N_VGND_c_981_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0020257f
+ $X=6.755 $Y=0 $X2=0 $Y2=0
cc_739 N_VGND_c_987_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n 0.0020257f
+ $X=5.215 $Y=0 $X2=0 $Y2=0
cc_740 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1606_n
+ 0.00841425f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_741 N_VGND_c_981_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n 0.0216446f
+ $X=6.755 $Y=0 $X2=0 $Y2=0
cc_742 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1607_n 0.012786f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_743 N_VGND_c_969_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 0.0138207f
+ $X=3.4 $Y=0.39 $X2=0 $Y2=0
cc_744 N_VGND_c_987_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n 0.0522346f
+ $X=5.215 $Y=0 $X2=0 $Y2=0
cc_745 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_c_1608_n
+ 0.0329318f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_746 N_VGND_c_1001_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1002_d
+ 0.00209319f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_747 N_VGND_c_1001_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1007_d
+ 0.00215206f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_748 N_VGND_c_1001_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1004_d
+ 0.00209344f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_749 N_VGND_c_971_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n 0.0213372f
+ $X=6.92 $Y=0.32 $X2=0 $Y2=0
cc_750 N_VGND_c_972_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n
+ 0.00534646f $X=6.92 $Y=0.32 $X2=0 $Y2=0
cc_751 N_VGND_c_988_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n 0.0216446f
+ $X=7.955 $Y=0 $X2=0 $Y2=0
cc_752 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1654_n 0.012786f
+ $X=13.11 $Y=0 $X2=0 $Y2=0
cc_753 N_VGND_Xsky130_fd_sc_hd__nand2_2_0/M1002_s
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.0030073f $X=7.905 $Y=0.235
+ $X2=0 $Y2=0
cc_754 N_VGND_c_973_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.0118126f
+ $X=8.04 $Y=0.38 $X2=0 $Y2=0
cc_755 N_VGND_c_988_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.0020257f
+ $X=7.955 $Y=0 $X2=0 $Y2=0
cc_756 N_VGND_c_989_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 0.0020257f
+ $X=9.75 $Y=0 $X2=0 $Y2=0
cc_757 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n
+ 0.00841425f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_758 N_VGND_c_971_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n
+ 0.00148053f $X=6.92 $Y=0.32 $X2=0 $Y2=0
cc_759 N_VGND_c_972_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1655_n
+ 0.00465853f $X=6.92 $Y=0.32 $X2=0 $Y2=0
cc_760 N_VGND_c_989_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1670_n 0.0151813f
+ $X=9.75 $Y=0 $X2=0 $Y2=0
cc_761 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1670_n
+ 0.0093992f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_762 N_VGND_c_974_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n 0.0138207f
+ $X=9.94 $Y=0.39 $X2=0 $Y2=0
cc_763 N_VGND_c_989_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.0522346f
+ $X=9.75 $Y=0 $X2=0 $Y2=0
cc_764 N_VGND_c_1001_n N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n
+ 0.0329318f $X=13.11 $Y=0 $X2=0 $Y2=0
cc_765 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1375_n 0.00539651f $X=10.15 $Y=0.995 $X2=0
+ $Y2=0
cc_766 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1375_n 0.00630972f $X=10.57 $Y=0.995 $X2=0
+ $Y2=0
cc_767 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1375_n 5.22228e-19 $X=10.99 $Y=0.995 $X2=0
+ $Y2=0
cc_768 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.009853f $X=10.57 $Y=0.995 $X2=0 $Y2=0
cc_769 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00864909f $X=10.99 $Y=0.995 $X2=0
+ $Y2=0
cc_770 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.026683f $X=11.275 $Y=1.19 $X2=0 $Y2=0
cc_771 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1279_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 0.00523428f $X=11.005 $Y=1.19 $X2=0
+ $Y2=0
cc_772 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1280_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n 6.94178e-19 $X=11.15 $Y=1.19 $X2=0 $Y2=0
cc_773 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1176_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00261194f $X=10.15 $Y=0.995 $X2=0
+ $Y2=0
cc_774 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00144547f $X=10.57 $Y=0.995 $X2=0
+ $Y2=0
cc_775 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1182_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.0193374f $X=10.355 $Y=1.19 $X2=0 $Y2=0
cc_776 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1279_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00173485f $X=11.005 $Y=1.19 $X2=0
+ $Y2=0
cc_777 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1285_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00587785f $X=10.435 $Y=1.19 $X2=0
+ $Y2=0
cc_778 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1186_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n 0.00230339f $X=10.57 $Y=1.16 $X2=0 $Y2=0
cc_779 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1177_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1383_n 5.22228e-19 $X=10.57 $Y=0.995 $X2=0
+ $Y2=0
cc_780 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1383_n 0.00630972f $X=10.99 $Y=0.995 $X2=0
+ $Y2=0
cc_781 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1383_n 0.0109314f $X=11.41 $Y=0.995 $X2=0 $Y2=0
cc_782 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.0108204f $X=11.41 $Y=0.995 $X2=0 $Y2=0
cc_783 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1341_n 0.00305484f $X=11.275 $Y=1.19 $X2=0
+ $Y2=0
cc_784 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1178_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n 0.00111672f $X=10.99 $Y=0.995 $X2=0
+ $Y2=0
cc_785 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n 0.00158032f $X=11.41 $Y=0.995 $X2=0
+ $Y2=0
cc_786 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n 0.0237296f $X=11.275 $Y=1.19 $X2=0 $Y2=0
cc_787 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1280_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n 0.00636895f $X=11.15 $Y=1.19 $X2=0 $Y2=0
cc_788 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1342_n 0.00230339f $X=11.41 $Y=1.16 $X2=0 $Y2=0
cc_789 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1418_n 0.00527847f $X=10.99 $Y=1.985 $X2=0
+ $Y2=0
cc_790 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1418_n 0.0111068f $X=11.41 $Y=1.985 $X2=0 $Y2=0
cc_791 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.00328577f $X=10.99 $Y=1.985 $X2=0
+ $Y2=0
cc_792 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.0143596f $X=11.41 $Y=1.985 $X2=0 $Y2=0
cc_793 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.0247043f $X=11.275 $Y=1.19 $X2=0 $Y2=0
cc_794 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1280_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.00641818f $X=11.15 $Y=1.19 $X2=0 $Y2=0
cc_795 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n 0.00215368f $X=11.41 $Y=1.16 $X2=0 $Y2=0
cc_796 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n 0.00180246f $X=11.275 $Y=1.19 $X2=0
+ $Y2=0
cc_797 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1280_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n 0.0185691f $X=11.15 $Y=1.19 $X2=0 $Y2=0
cc_798 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n 0.00235288f $X=11.41 $Y=1.16 $X2=0 $Y2=0
cc_799 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1179_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1346_n 0.0140806f $X=11.41 $Y=0.995 $X2=0 $Y2=0
cc_800 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1346_n 0.0137498f $X=11.275 $Y=1.19 $X2=0 $Y2=0
cc_801 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1280_p
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1346_n 3.77336e-19 $X=11.15 $Y=1.19 $X2=0 $Y2=0
cc_802 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1187_n
+ N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n 0.00478049f $X=11.41 $Y=1.16 $X2=0 $Y2=0
cc_803 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1181_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n 0.00338615f $X=9.435 $Y=0.835
+ $X2=0 $Y2=0
cc_804 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1182_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n 0.0201375f $X=10.355 $Y=1.19
+ $X2=0 $Y2=0
cc_805 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1184_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n 0.00229746f $X=10.145 $Y=1.19
+ $X2=0 $Y2=0
cc_806 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1196_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1531_n 0.0156019f $X=9.435 $Y=1.495
+ $X2=0 $Y2=0
cc_807 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.0137355f $X=10.15 $Y=1.985
+ $X2=0 $Y2=0
cc_808 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.0149365f $X=10.57 $Y=1.985
+ $X2=0 $Y2=0
cc_809 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1182_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.0268324f $X=10.355 $Y=1.19
+ $X2=0 $Y2=0
cc_810 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00362207f $X=11.275 $Y=1.19
+ $X2=0 $Y2=0
cc_811 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1184_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 8.64843e-19 $X=10.145 $Y=1.19
+ $X2=0 $Y2=0
cc_812 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1279_p
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00493378f $X=11.005 $Y=1.19
+ $X2=0 $Y2=0
cc_813 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1285_p
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00708414f $X=10.435 $Y=1.19
+ $X2=0 $Y2=0
cc_814 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1186_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00213789f $X=10.57 $Y=1.16
+ $X2=0 $Y2=0
cc_815 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1534_n 2.36323e-19 $X=10.99 $Y=1.985
+ $X2=0 $Y2=0
cc_816 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1183_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1534_n 0.0124486f $X=11.275 $Y=1.19
+ $X2=0 $Y2=0
cc_817 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1279_p
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1534_n 0.00142025f $X=11.005 $Y=1.19
+ $X2=0 $Y2=0
cc_818 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.0112436f $X=10.99 $Y=1.985
+ $X2=0 $Y2=0
cc_819 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.00929492f $X=11.41 $Y=1.985
+ $X2=0 $Y2=0
cc_820 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1004_d
+ 7.4958e-19 $X=9.295 $Y=0.78 $X2=0 $Y2=0
cc_821 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1004_d
+ 0.00241065f $X=9.435 $Y=0.905 $X2=0 $Y2=0
cc_822 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1660_n 8.34819e-19 $X=8.715 $Y=1.58
+ $X2=0 $Y2=0
cc_823 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1205_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1656_n 3.07688e-19 $X=8.715 $Y=1.58
+ $X2=0 $Y2=0
cc_824 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n 0.00726619f $X=9.295 $Y=0.78
+ $X2=0 $Y2=0
cc_825 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1185_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n 6.10376e-19 $X=9.575 $Y=1.19
+ $X2=0 $Y2=0
cc_826 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1188_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1657_n 0.0131928f $X=9.435 $Y=0.905
+ $X2=0 $Y2=0
cc_827 N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1003_s
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.00312175f $X=8.745 $Y=0.235
+ $X2=0 $Y2=0
cc_828 N_SKY130_FD_SC_HD__NOR2_2_0/A_c_1180_n
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_c_1677_n 0.0192847f $X=9.295 $Y=0.78
+ $X2=0 $Y2=0
cc_829 N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1006_d
+ 0.00296777f $X=11.687 $Y=1.555 $X2=0 $Y2=0
cc_830 N_SKY130_FD_SC_HD__INV_2_0/A_c_1339_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 0.00126399f $X=11.035 $Y=0.815
+ $X2=0 $Y2=0
cc_831 N_SKY130_FD_SC_HD__INV_2_0/A_c_1340_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1533_n 7.6328e-19 $X=10.525 $Y=0.815
+ $X2=0 $Y2=0
cc_832 N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1534_n 0.0102037f $X=11.687 $Y=1.555
+ $X2=0 $Y2=0
cc_833 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_s
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.00312348f $X=11.065 $Y=1.485
+ $X2=0 $Y2=0
cc_834 N_SKY130_FD_SC_HD__INV_2_0/A_c_1418_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.0154795f $X=11.2 $Y=1.62
+ $X2=0 $Y2=0
cc_835 N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1535_n 0.00282992f $X=11.687 $Y=1.555
+ $X2=0 $Y2=0
cc_836 N_SKY130_FD_SC_HD__INV_2_0/A_c_1351_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1536_n 0.0202369f $X=11.687 $Y=1.555
+ $X2=0 $Y2=0
cc_837 N_SKY130_FD_SC_HD__INV_2_0/A_c_1345_n
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_c_1536_n 0.00152808f $X=11.835 $Y=1.19
+ $X2=0 $Y2=0
cc_838 N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1585_n 0.00534153f $X=12.44 $Y=0.995 $X2=0
+ $Y2=0
cc_839 N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1585_n 0.00534153f $X=12.86 $Y=0.995 $X2=0
+ $Y2=0
cc_840 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1582_n 0.00918977f $X=12.44 $Y=1.985 $X2=0
+ $Y2=0
cc_841 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1582_n 0.00918977f $X=12.86 $Y=1.985 $X2=0
+ $Y2=0
cc_842 N_SKY130_FD_SC_HD__INV_2_0/A_c_1337_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.004954f $X=12.44 $Y=0.995 $X2=0 $Y2=0
cc_843 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.00408533f $X=12.44 $Y=1.985 $X2=0
+ $Y2=0
cc_844 N_SKY130_FD_SC_HD__INV_2_0/A_c_1338_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.00675111f $X=12.86 $Y=0.995 $X2=0
+ $Y2=0
cc_845 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.00809641f $X=12.86 $Y=1.985 $X2=0
+ $Y2=0
cc_846 N_SKY130_FD_SC_HD__INV_2_0/A_c_1343_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.0156803f $X=12.19 $Y=1.19 $X2=0 $Y2=0
cc_847 N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 3.94596e-19 $X=12.175 $Y=1.19 $X2=0
+ $Y2=0
cc_848 N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1579_n 0.0259992f $X=12.86 $Y=1.16 $X2=0 $Y2=0
cc_849 N_SKY130_FD_SC_HD__INV_2_0/A_c_1343_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1600_n 0.00151169f $X=12.19 $Y=1.19 $X2=0 $Y2=0
cc_850 N_SKY130_FD_SC_HD__INV_2_0/A_c_1347_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1600_n 0.0229696f $X=12.175 $Y=1.19 $X2=0 $Y2=0
cc_851 N_SKY130_FD_SC_HD__INV_2_0/A_c_1348_n
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1600_n 0.0147405f $X=12.86 $Y=1.16 $X2=0 $Y2=0
cc_852 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1603_n 0.00280787f $X=12.44 $Y=1.985 $X2=0
+ $Y2=0
cc_853 N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_c_1603_n 0.00214168f $X=12.86 $Y=1.985 $X2=0
+ $Y2=0

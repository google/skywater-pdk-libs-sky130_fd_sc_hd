* File: sky130_fd_sc_hd__and3b_2.pxi.spice
* Created: Thu Aug 27 14:08:05 2020
* 
x_PM_SKY130_FD_SC_HD__AND3B_2%A_N N_A_N_M1005_g N_A_N_M1006_g A_N A_N
+ N_A_N_c_71_n PM_SKY130_FD_SC_HD__AND3B_2%A_N
x_PM_SKY130_FD_SC_HD__AND3B_2%A_109_53# N_A_109_53#_M1005_d N_A_109_53#_M1006_d
+ N_A_109_53#_M1010_g N_A_109_53#_M1002_g N_A_109_53#_c_96_n N_A_109_53#_c_97_n
+ N_A_109_53#_c_98_n N_A_109_53#_c_99_n N_A_109_53#_c_100_n
+ PM_SKY130_FD_SC_HD__AND3B_2%A_109_53#
x_PM_SKY130_FD_SC_HD__AND3B_2%B N_B_M1003_g N_B_M1007_g N_B_c_139_n B
+ N_B_c_142_n PM_SKY130_FD_SC_HD__AND3B_2%B
x_PM_SKY130_FD_SC_HD__AND3B_2%C N_C_M1004_g N_C_M1008_g C C N_C_c_178_n
+ PM_SKY130_FD_SC_HD__AND3B_2%C
x_PM_SKY130_FD_SC_HD__AND3B_2%A_215_311# N_A_215_311#_M1002_s
+ N_A_215_311#_M1010_s N_A_215_311#_M1007_d N_A_215_311#_c_221_n
+ N_A_215_311#_M1009_g N_A_215_311#_M1000_g N_A_215_311#_c_222_n
+ N_A_215_311#_M1011_g N_A_215_311#_M1001_g N_A_215_311#_c_229_n
+ N_A_215_311#_c_223_n N_A_215_311#_c_230_n N_A_215_311#_c_231_n
+ N_A_215_311#_c_224_n N_A_215_311#_c_257_n N_A_215_311#_c_233_n
+ N_A_215_311#_c_234_n N_A_215_311#_c_225_n N_A_215_311#_c_226_n
+ PM_SKY130_FD_SC_HD__AND3B_2%A_215_311#
x_PM_SKY130_FD_SC_HD__AND3B_2%VPWR N_VPWR_M1006_s N_VPWR_M1010_d N_VPWR_M1008_d
+ N_VPWR_M1001_d N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n
+ N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_347_n VPWR N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_330_n
+ PM_SKY130_FD_SC_HD__AND3B_2%VPWR
x_PM_SKY130_FD_SC_HD__AND3B_2%X N_X_M1009_d N_X_M1000_s N_X_c_387_n N_X_c_396_n
+ N_X_c_389_n X X X N_X_c_411_n X N_X_c_412_n PM_SKY130_FD_SC_HD__AND3B_2%X
x_PM_SKY130_FD_SC_HD__AND3B_2%VGND N_VGND_M1005_s N_VGND_M1004_d N_VGND_M1011_s
+ N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n
+ VGND N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n
+ PM_SKY130_FD_SC_HD__AND3B_2%VGND
cc_1 VNB N_A_N_M1005_g 0.0374011f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB A_N 0.0116594f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A_N_c_71_n 0.0482177f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_109_53#_M1002_g 0.0320842f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_5 VNB N_A_109_53#_c_96_n 0.013992f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=0.85
cc_6 VNB N_A_109_53#_c_97_n 0.00154999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_109_53#_c_98_n 0.0151677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_109_53#_c_99_n 0.00361993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_109_53#_c_100_n 0.0340277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_M1003_g 0.0249958f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_11 VNB N_B_M1007_g 0.00462644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_139_n 0.0120087f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_13 VNB N_C_M1004_g 0.0266067f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_14 VNB C 4.7131e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_15 VNB C 0.0107095f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_C_c_178_n 0.0194923f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_17 VNB N_A_215_311#_c_221_n 0.0176302f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_A_215_311#_c_222_n 0.0202418f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=0.85
cc_19 VNB N_A_215_311#_c_223_n 0.0032547f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_215_311#_c_224_n 0.00510463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_215_311#_c_225_n 0.00382265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_215_311#_c_226_n 0.0402727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_330_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_387_n 7.23192e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.0224173f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_26 VNB N_VGND_c_421_n 0.010079f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_27 VNB N_VGND_c_422_n 0.0199104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_423_n 0.00311252f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_29 VNB N_VGND_c_424_n 0.0100062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_425_n 0.0243823f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_426_n 0.0543489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_427_n 0.015254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_428_n 0.00510766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_429_n 0.222608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_N_M1006_g 0.0378397f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.765
cc_36 VPB A_N 0.0026867f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_37 VPB N_A_N_c_71_n 0.0097152f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_38 VPB N_A_109_53#_M1010_g 0.0287481f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_39 VPB N_A_109_53#_c_97_n 0.0115132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_109_53#_c_100_n 0.00815536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B_M1007_g 0.0211481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB B 0.00971454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B_c_142_n 0.0414351f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_44 VPB N_C_M1008_g 0.0205363f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.765
cc_45 VPB N_C_c_178_n 0.00425601f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_46 VPB N_A_215_311#_M1000_g 0.0207234f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_47 VPB N_A_215_311#_M1001_g 0.0231128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_215_311#_c_229_n 0.00352671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_215_311#_c_230_n 0.00319006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_215_311#_c_231_n 0.00337561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_215_311#_c_224_n 0.00164465f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_215_311#_c_233_n 0.00634289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_215_311#_c_234_n 0.00558352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_215_311#_c_225_n 0.00121877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_215_311#_c_226_n 0.00810712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_331_n 0.0109454f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_57 VPB N_VPWR_c_332_n 0.0494594f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_58 VPB N_VPWR_c_333_n 0.0212745f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.16
cc_59 VPB N_VPWR_c_334_n 0.00444413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_335_n 0.00998035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_336_n 0.0377907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_337_n 0.0563065f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_338_n 0.0179932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_339_n 0.00141883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_340_n 0.00410958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_330_n 0.0650786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_X_c_389_n 5.95156e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB X 0.0116895f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_69 N_A_N_M1005_g N_A_109_53#_c_96_n 0.00882834f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_70 A_N N_A_109_53#_c_96_n 0.020647f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_71 A_N N_A_109_53#_c_97_n 0.00609989f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_72 N_A_N_c_71_n N_A_109_53#_c_97_n 0.0106502f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_73 A_N N_A_109_53#_c_99_n 0.019107f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_74 N_A_N_c_71_n N_A_109_53#_c_99_n 0.00315652f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_N_c_71_n N_A_109_53#_c_100_n 0.00518656f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_N_M1006_g N_A_215_311#_c_229_n 9.76835e-19 $X=0.47 $Y=1.765 $X2=0
+ $Y2=0
cc_77 N_A_N_M1006_g N_VPWR_c_332_n 0.014987f $X=0.47 $Y=1.765 $X2=0 $Y2=0
cc_78 A_N N_VPWR_c_332_n 0.0142442f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_N_c_71_n N_VPWR_c_332_n 0.00326847f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_N_M1006_g N_VPWR_c_337_n 0.00353352f $X=0.47 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_N_M1006_g N_VPWR_c_330_n 0.00428307f $X=0.47 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_N_M1005_g N_VGND_c_422_n 0.00470487f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_83 A_N N_VGND_c_422_n 0.0174883f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_84 N_A_N_c_71_n N_VGND_c_422_n 0.00223068f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_N_M1005_g N_VGND_c_426_n 0.00542149f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_86 A_N N_VGND_c_426_n 8.36374e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_87 N_A_N_M1005_g N_VGND_c_429_n 0.0117518f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_88 A_N N_VGND_c_429_n 0.00231313f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_109_53#_M1002_g N_B_M1003_g 0.0330914f $X=1.43 $Y=0.475 $X2=0 $Y2=0
cc_90 N_A_109_53#_M1010_g N_B_M1007_g 0.0211943f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_109_53#_c_100_n N_B_M1007_g 0.00622468f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_109_53#_c_100_n N_B_c_139_n 0.0330914f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_109_53#_c_97_n N_A_215_311#_c_229_n 0.0224984f $X=0.68 $Y=1.74 $X2=0
+ $Y2=0
cc_94 N_A_109_53#_M1002_g N_A_215_311#_c_223_n 0.0131578f $X=1.43 $Y=0.475 $X2=0
+ $Y2=0
cc_95 N_A_109_53#_c_96_n N_A_215_311#_c_223_n 0.0204758f $X=0.7 $Y=0.47 $X2=0
+ $Y2=0
cc_96 N_A_109_53#_c_98_n N_A_215_311#_c_223_n 0.0116666f $X=1.22 $Y=1.16 $X2=0
+ $Y2=0
cc_97 N_A_109_53#_c_100_n N_A_215_311#_c_223_n 0.00499852f $X=1.43 $Y=1.16 $X2=0
+ $Y2=0
cc_98 N_A_109_53#_M1010_g N_A_215_311#_c_230_n 0.0144635f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_99 N_A_109_53#_c_98_n N_A_215_311#_c_230_n 0.00876907f $X=1.22 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_109_53#_c_100_n N_A_215_311#_c_230_n 0.00211758f $X=1.43 $Y=1.16
+ $X2=0 $Y2=0
cc_101 N_A_109_53#_c_97_n N_A_215_311#_c_231_n 0.0134726f $X=0.68 $Y=1.74 $X2=0
+ $Y2=0
cc_102 N_A_109_53#_c_98_n N_A_215_311#_c_231_n 0.0182953f $X=1.22 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_109_53#_c_100_n N_A_215_311#_c_231_n 0.00506215f $X=1.43 $Y=1.16
+ $X2=0 $Y2=0
cc_104 N_A_109_53#_M1010_g N_A_215_311#_c_224_n 0.0024221f $X=1.41 $Y=1.765
+ $X2=0 $Y2=0
cc_105 N_A_109_53#_M1002_g N_A_215_311#_c_224_n 0.014381f $X=1.43 $Y=0.475 $X2=0
+ $Y2=0
cc_106 N_A_109_53#_c_98_n N_A_215_311#_c_224_n 0.0187659f $X=1.22 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_109_53#_M1010_g N_VPWR_c_347_n 0.00256209f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_109_53#_M1010_g N_VPWR_c_337_n 0.00483317f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_109_53#_M1010_g N_VPWR_c_339_n 0.00874185f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_109_53#_c_97_n N_VPWR_c_330_n 0.0109339f $X=0.68 $Y=1.74 $X2=0 $Y2=0
cc_111 N_A_109_53#_M1002_g N_VGND_c_426_n 0.00347765f $X=1.43 $Y=0.475 $X2=0
+ $Y2=0
cc_112 N_A_109_53#_c_96_n N_VGND_c_426_n 0.0140092f $X=0.7 $Y=0.47 $X2=0 $Y2=0
cc_113 N_A_109_53#_M1002_g N_VGND_c_429_n 0.0059338f $X=1.43 $Y=0.475 $X2=0
+ $Y2=0
cc_114 N_A_109_53#_c_96_n N_VGND_c_429_n 0.0102507f $X=0.7 $Y=0.47 $X2=0 $Y2=0
cc_115 N_B_M1003_g N_C_M1004_g 0.0416246f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_C_M1008_g 0.0122184f $X=1.83 $Y=1.765 $X2=0 $Y2=0
cc_117 B N_C_M1008_g 0.00206749f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_118 N_B_M1003_g C 0.00410142f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_119 N_B_c_139_n C 0.0014215f $X=1.81 $Y=1.2 $X2=0 $Y2=0
cc_120 N_B_c_139_n N_C_c_178_n 0.0180091f $X=1.81 $Y=1.2 $X2=0 $Y2=0
cc_121 N_B_c_142_n N_A_215_311#_M1000_g 0.00208029f $X=1.9 $Y=2.3 $X2=0 $Y2=0
cc_122 N_B_M1003_g N_A_215_311#_c_223_n 0.00808008f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_123 N_B_M1003_g N_A_215_311#_c_224_n 0.0096969f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_124 N_B_M1007_g N_A_215_311#_c_224_n 0.00656763f $X=1.83 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B_c_139_n N_A_215_311#_c_224_n 0.00500625f $X=1.81 $Y=1.2 $X2=0 $Y2=0
cc_126 B N_A_215_311#_c_257_n 0.0107664f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_127 N_B_M1007_g N_A_215_311#_c_234_n 0.0130234f $X=1.83 $Y=1.765 $X2=0 $Y2=0
cc_128 B N_A_215_311#_c_234_n 0.00781453f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_129 N_B_c_142_n N_A_215_311#_c_234_n 3.77868e-19 $X=1.9 $Y=2.3 $X2=0 $Y2=0
cc_130 B N_VPWR_c_333_n 0.0314336f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_131 N_B_c_142_n N_VPWR_c_333_n 0.00596674f $X=1.9 $Y=2.3 $X2=0 $Y2=0
cc_132 N_B_M1007_g N_VPWR_c_334_n 0.00239172f $X=1.83 $Y=1.765 $X2=0 $Y2=0
cc_133 B N_VPWR_c_334_n 0.0277107f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_134 N_B_c_142_n N_VPWR_c_334_n 0.00132062f $X=1.9 $Y=2.3 $X2=0 $Y2=0
cc_135 N_B_M1007_g N_VPWR_c_347_n 0.00379873f $X=1.83 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B_c_142_n N_VPWR_c_337_n 0.00665957f $X=1.9 $Y=2.3 $X2=0 $Y2=0
cc_137 N_B_M1007_g N_VPWR_c_339_n 0.00665957f $X=1.83 $Y=1.765 $X2=0 $Y2=0
cc_138 B N_VPWR_c_339_n 0.0288888f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_139 B N_VPWR_c_330_n 0.0169635f $X=2.01 $Y=2.125 $X2=0 $Y2=0
cc_140 N_B_c_142_n N_VPWR_c_330_n 0.00834174f $X=1.9 $Y=2.3 $X2=0 $Y2=0
cc_141 N_B_M1003_g N_VGND_c_426_n 0.00382191f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_142 N_B_M1003_g N_VGND_c_429_n 0.00577482f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_143 N_C_M1004_g N_A_215_311#_c_221_n 0.0147418f $X=2.195 $Y=0.475 $X2=0 $Y2=0
cc_144 C N_A_215_311#_c_221_n 6.38142e-19 $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_145 C N_A_215_311#_c_221_n 0.00232992f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_146 N_C_M1008_g N_A_215_311#_M1000_g 0.0187411f $X=2.305 $Y=1.695 $X2=0 $Y2=0
cc_147 N_C_M1004_g N_A_215_311#_c_223_n 2.65899e-19 $X=2.195 $Y=0.475 $X2=0
+ $Y2=0
cc_148 C N_A_215_311#_c_223_n 0.0211398f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_149 N_C_M1004_g N_A_215_311#_c_224_n 6.6184e-19 $X=2.195 $Y=0.475 $X2=0 $Y2=0
cc_150 N_C_M1008_g N_A_215_311#_c_224_n 5.32924e-19 $X=2.305 $Y=1.695 $X2=0
+ $Y2=0
cc_151 C N_A_215_311#_c_224_n 0.052259f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_152 N_C_c_178_n N_A_215_311#_c_224_n 4.81118e-19 $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_153 N_C_M1008_g N_A_215_311#_c_233_n 0.013148f $X=2.305 $Y=1.695 $X2=0 $Y2=0
cc_154 N_C_c_178_n N_A_215_311#_c_233_n 2.44767e-19 $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_155 C N_A_215_311#_c_234_n 0.0308291f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_156 N_C_c_178_n N_A_215_311#_c_234_n 0.00315743f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_157 N_C_M1008_g N_A_215_311#_c_225_n 0.00212173f $X=2.305 $Y=1.695 $X2=0
+ $Y2=0
cc_158 C N_A_215_311#_c_225_n 0.020603f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_159 N_C_c_178_n N_A_215_311#_c_225_n 0.00238051f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_160 C N_A_215_311#_c_226_n 8.32628e-19 $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_161 N_C_c_178_n N_A_215_311#_c_226_n 0.0212377f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_162 N_C_M1008_g N_VPWR_c_333_n 0.00200243f $X=2.305 $Y=1.695 $X2=0 $Y2=0
cc_163 N_C_M1008_g N_VPWR_c_334_n 0.0037598f $X=2.305 $Y=1.695 $X2=0 $Y2=0
cc_164 N_C_M1008_g N_VPWR_c_347_n 2.09407e-19 $X=2.305 $Y=1.695 $X2=0 $Y2=0
cc_165 N_C_M1008_g N_VPWR_c_330_n 0.00250493f $X=2.305 $Y=1.695 $X2=0 $Y2=0
cc_166 C N_X_c_387_n 0.00535475f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_167 C X 0.00262087f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_168 N_C_M1004_g N_VGND_c_423_n 0.00607028f $X=2.195 $Y=0.475 $X2=0 $Y2=0
cc_169 C N_VGND_c_423_n 0.0189612f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_170 C N_VGND_c_423_n 6.45863e-19 $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_171 N_C_M1004_g N_VGND_c_426_n 0.00418186f $X=2.195 $Y=0.475 $X2=0 $Y2=0
cc_172 C N_VGND_c_426_n 0.00940062f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_173 N_C_M1004_g N_VGND_c_429_n 0.0055742f $X=2.195 $Y=0.475 $X2=0 $Y2=0
cc_174 C N_VGND_c_429_n 0.0073435f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_175 C N_VGND_c_429_n 0.0073758f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_176 C A_373_53# 0.00371982f $X=2.01 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_177 N_A_215_311#_c_230_n N_VPWR_M1010_d 4.47557e-19 $X=1.585 $Y=1.51 $X2=0
+ $Y2=0
cc_178 N_A_215_311#_c_234_n N_VPWR_M1010_d 0.00120414f $X=2.2 $Y=1.51 $X2=0
+ $Y2=0
cc_179 N_A_215_311#_c_233_n N_VPWR_M1008_d 0.00314201f $X=2.59 $Y=1.51 $X2=0
+ $Y2=0
cc_180 N_A_215_311#_c_229_n N_VPWR_c_332_n 0.00152152f $X=1.2 $Y=1.76 $X2=0
+ $Y2=0
cc_181 N_A_215_311#_M1000_g N_VPWR_c_334_n 0.00310368f $X=2.79 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_215_311#_c_233_n N_VPWR_c_334_n 0.0149225f $X=2.59 $Y=1.51 $X2=0
+ $Y2=0
cc_183 N_A_215_311#_c_226_n N_VPWR_c_334_n 2.9535e-19 $X=3.21 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_215_311#_M1001_g N_VPWR_c_336_n 0.00594697f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_215_311#_c_230_n N_VPWR_c_347_n 0.0154228f $X=1.585 $Y=1.51 $X2=0
+ $Y2=0
cc_186 N_A_215_311#_c_257_n N_VPWR_c_347_n 0.0074696f $X=2.095 $Y=1.725 $X2=0
+ $Y2=0
cc_187 N_A_215_311#_c_229_n N_VPWR_c_337_n 0.0201855f $X=1.2 $Y=1.76 $X2=0 $Y2=0
cc_188 N_A_215_311#_c_230_n N_VPWR_c_337_n 0.00511706f $X=1.585 $Y=1.51 $X2=0
+ $Y2=0
cc_189 N_A_215_311#_M1000_g N_VPWR_c_338_n 0.00585385f $X=2.79 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_215_311#_M1001_g N_VPWR_c_338_n 0.0054895f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_215_311#_M1000_g N_VPWR_c_330_n 0.0117707f $X=2.79 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_215_311#_M1001_g N_VPWR_c_330_n 0.0106281f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_215_311#_c_229_n N_VPWR_c_330_n 9.29713e-19 $X=1.2 $Y=1.76 $X2=0
+ $Y2=0
cc_194 N_A_215_311#_c_221_n N_X_c_387_n 0.00269233f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_215_311#_c_222_n N_X_c_387_n 0.00905919f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_215_311#_c_226_n N_X_c_387_n 4.25328e-19 $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_215_311#_M1001_g N_X_c_396_n 0.00151268f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_215_311#_c_226_n N_X_c_396_n 0.00112447f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_215_311#_M1000_g N_X_c_389_n 0.00505627f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_215_311#_M1001_g N_X_c_389_n 0.0114063f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_215_311#_c_233_n N_X_c_389_n 0.0118423f $X=2.59 $Y=1.51 $X2=0 $Y2=0
cc_202 N_A_215_311#_c_226_n N_X_c_389_n 3.21959e-19 $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_215_311#_c_222_n X 0.00129962f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_215_311#_c_226_n X 0.00130953f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_215_311#_c_221_n X 8.72726e-19 $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_215_311#_M1000_g X 7.99116e-19 $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_215_311#_c_222_n X 0.00923584f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_215_311#_M1001_g X 0.0113091f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_215_311#_c_233_n X 0.00167834f $X=2.59 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_215_311#_c_225_n X 0.0335046f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_215_311#_c_226_n X 0.0222013f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_215_311#_c_222_n N_X_c_411_n 0.00450041f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_215_311#_M1001_g N_X_c_412_n 0.00581098f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_215_311#_c_221_n N_VGND_c_423_n 0.00933971f $X=2.79 $Y=0.995 $X2=0
+ $Y2=0
cc_215 N_A_215_311#_c_222_n N_VGND_c_423_n 6.46241e-19 $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_216 N_A_215_311#_c_225_n N_VGND_c_423_n 0.00503735f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_217 N_A_215_311#_c_226_n N_VGND_c_423_n 5.53235e-19 $X=3.21 $Y=1.16 $X2=0
+ $Y2=0
cc_218 N_A_215_311#_c_222_n N_VGND_c_425_n 0.00546769f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_215_311#_c_223_n N_VGND_c_426_n 0.0353135f $X=1.585 $Y=0.437 $X2=0
+ $Y2=0
cc_220 N_A_215_311#_c_221_n N_VGND_c_427_n 0.00486043f $X=2.79 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_215_311#_c_222_n N_VGND_c_427_n 0.0054895f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_215_311#_c_221_n N_VGND_c_429_n 0.0082748f $X=2.79 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_215_311#_c_222_n N_VGND_c_429_n 0.0107794f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_215_311#_c_223_n N_VGND_c_429_n 0.0276241f $X=1.585 $Y=0.437 $X2=0
+ $Y2=0
cc_225 N_A_215_311#_c_223_n A_301_53# 0.00191292f $X=1.585 $Y=0.437 $X2=-0.19
+ $Y2=-0.24
cc_226 N_A_215_311#_c_224_n A_301_53# 0.00132529f $X=1.712 $Y=1.425 $X2=-0.19
+ $Y2=-0.24
cc_227 N_VPWR_c_330_n N_X_M1000_s 0.00249917f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_336_n X 0.0222348f $X=3.42 $Y=1.96 $X2=0 $Y2=0
cc_229 N_VPWR_c_338_n N_X_c_412_n 0.016223f $X=3.33 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_330_n N_X_c_412_n 0.0107149f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_231 X N_VGND_c_425_n 0.0222348f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_232 N_X_c_411_n N_VGND_c_427_n 0.0146998f $X=3.037 $Y=0.593 $X2=0 $Y2=0
cc_233 N_X_M1009_d N_VGND_c_429_n 0.00393857f $X=2.865 $Y=0.235 $X2=0 $Y2=0
cc_234 N_X_c_411_n N_VGND_c_429_n 0.00921777f $X=3.037 $Y=0.593 $X2=0 $Y2=0

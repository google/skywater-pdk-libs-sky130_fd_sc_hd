* File: sky130_fd_sc_hd__a31oi_1.pxi.spice
* Created: Tue Sep  1 18:55:19 2020
* 
x_PM_SKY130_FD_SC_HD__A31OI_1%A3 N_A3_c_43_n N_A3_M1007_g N_A3_M1006_g A3
+ N_A3_c_45_n PM_SKY130_FD_SC_HD__A31OI_1%A3
x_PM_SKY130_FD_SC_HD__A31OI_1%A2 N_A2_M1003_g N_A2_M1002_g A2 A2 A2 N_A2_c_67_n
+ N_A2_c_68_n PM_SKY130_FD_SC_HD__A31OI_1%A2
x_PM_SKY130_FD_SC_HD__A31OI_1%A1 N_A1_M1004_g N_A1_M1005_g N_A1_c_105_n
+ N_A1_c_106_n A1 N_A1_c_107_n N_A1_c_111_n PM_SKY130_FD_SC_HD__A31OI_1%A1
x_PM_SKY130_FD_SC_HD__A31OI_1%B1 N_B1_c_147_n N_B1_M1000_g N_B1_M1001_g B1
+ N_B1_c_149_n PM_SKY130_FD_SC_HD__A31OI_1%B1
x_PM_SKY130_FD_SC_HD__A31OI_1%VPWR N_VPWR_M1006_s N_VPWR_M1002_d N_VPWR_c_176_n
+ N_VPWR_c_177_n N_VPWR_c_178_n VPWR N_VPWR_c_179_n N_VPWR_c_180_n
+ N_VPWR_c_175_n N_VPWR_c_182_n PM_SKY130_FD_SC_HD__A31OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A31OI_1%A_109_297# N_A_109_297#_M1006_d
+ N_A_109_297#_M1005_d N_A_109_297#_c_224_n N_A_109_297#_c_215_n
+ N_A_109_297#_c_218_n N_A_109_297#_c_231_n
+ PM_SKY130_FD_SC_HD__A31OI_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A31OI_1%Y N_Y_M1004_d N_Y_M1001_d N_Y_c_240_n N_Y_c_236_n
+ N_Y_c_249_n N_Y_c_238_n Y Y PM_SKY130_FD_SC_HD__A31OI_1%Y
x_PM_SKY130_FD_SC_HD__A31OI_1%VGND N_VGND_M1007_s N_VGND_M1000_d N_VGND_c_275_n
+ N_VGND_c_276_n N_VGND_c_277_n N_VGND_c_278_n VGND N_VGND_c_279_n
+ N_VGND_c_280_n PM_SKY130_FD_SC_HD__A31OI_1%VGND
cc_1 VNB N_A3_c_43_n 0.0206809f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A3 0.0140863f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A3_c_45_n 0.0366615f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB A2 0.00863844f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_5 VNB N_A2_c_67_n 0.0190055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A2_c_68_n 0.0153872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A1_c_105_n 3.16405e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_8 VNB N_A1_c_106_n 0.0234644f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_9 VNB N_A1_c_107_n 0.0177526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_147_n 0.0220799f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB B1 0.014545f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_12 VNB N_B1_c_149_n 0.0372046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_175_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_236_n 0.0028679f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_15 VNB N_VGND_c_275_n 0.0103393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_276_n 0.0256844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_277_n 0.00988631f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_18 VNB N_VGND_c_278_n 0.0182011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_279_n 0.0403011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_280_n 0.141241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_A3_M1006_g 0.0254473f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_22 VPB A3 0.00344411f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_23 VPB N_A3_c_45_n 0.00999597f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_24 VPB N_A2_M1002_g 0.019233f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_25 VPB N_A2_c_67_n 0.00508691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A1_M1005_g 0.0189637f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_27 VPB N_A1_c_105_n 8.65482e-19 $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_28 VPB N_A1_c_106_n 0.00462679f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_29 VPB N_A1_c_111_n 0.00691897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_B1_M1001_g 0.0259703f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_31 VPB B1 0.00297428f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_B1_c_149_n 0.010021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_176_n 0.0100778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_177_n 0.041437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_178_n 0.00271083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_179_n 0.0121021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_180_n 0.0293422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_175_n 0.0431118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_182_n 0.00507625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_Y_c_236_n 0.00108863f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_41 VPB N_Y_c_238_n 0.00742573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB Y 0.0308277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 N_A3_M1006_g N_A2_M1002_g 0.0416173f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_44 N_A3_c_43_n A2 0.0106428f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_45 A3 A2 0.0170893f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_46 A3 N_A2_c_67_n 4.53948e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A3_c_45_n N_A2_c_67_n 0.0373407f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_48 N_A3_c_43_n N_A2_c_68_n 0.0373407f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A3_M1006_g N_VPWR_c_177_n 0.0187768f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_50 A3 N_VPWR_c_177_n 0.0216203f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_51 N_A3_c_45_n N_VPWR_c_177_n 0.00197112f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A3_M1006_g N_VPWR_c_178_n 6.41967e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_53 N_A3_M1006_g N_VPWR_c_179_n 0.00486043f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_54 N_A3_M1006_g N_VPWR_c_175_n 0.00830305f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_55 N_A3_c_43_n N_VGND_c_276_n 0.0144105f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_56 A3 N_VGND_c_276_n 0.0206839f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_57 N_A3_c_45_n N_VGND_c_276_n 0.0019532f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A3_c_43_n N_VGND_c_279_n 0.00447018f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A3_c_43_n N_VGND_c_280_n 0.00752597f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A2_M1002_g N_A1_M1005_g 0.038494f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A2_M1002_g N_A1_c_105_n 7.37482e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_62 A2 N_A1_c_105_n 0.0183076f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_63 N_A2_c_67_n N_A1_c_105_n 6.42974e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_64 A2 N_A1_c_106_n 0.0017393f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_65 N_A2_c_67_n N_A1_c_106_n 0.020558f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_66 A2 N_A1_c_107_n 0.00598194f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_67 N_A2_c_68_n N_A1_c_107_n 0.0273278f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A2_M1002_g N_A1_c_111_n 0.00360124f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A2_M1002_g N_VPWR_c_177_n 0.00217006f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A2_M1002_g N_VPWR_c_178_n 0.00776704f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A2_M1002_g N_VPWR_c_179_n 0.00348405f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A2_M1002_g N_VPWR_c_175_n 0.00417382f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A2_M1002_g N_A_109_297#_c_215_n 0.0133089f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_74 A2 N_A_109_297#_c_215_n 0.00707668f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_75 N_A2_c_67_n N_A_109_297#_c_215_n 8.60234e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_76 A2 N_A_109_297#_c_218_n 0.00573994f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_77 A2 N_Y_c_240_n 0.024034f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_78 N_A2_c_68_n N_Y_c_240_n 6.36618e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_79 A2 N_Y_c_236_n 0.00570474f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_80 A2 N_VGND_c_276_n 0.0365714f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_81 N_A2_c_68_n N_VGND_c_276_n 0.00204042f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_82 A2 N_VGND_c_279_n 0.0177213f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_83 N_A2_c_68_n N_VGND_c_279_n 0.00373852f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_84 A2 N_VGND_c_280_n 0.0156373f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_85 N_A2_c_68_n N_VGND_c_280_n 0.00542691f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_86 A2 A_109_47# 0.00598676f $X=0.61 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_87 A2 A_181_47# 0.0075528f $X=0.61 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_88 N_A1_c_107_n N_B1_c_147_n 0.00918239f $X=1.37 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_89 N_A1_M1005_g N_B1_M1001_g 0.0333343f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A1_c_105_n N_B1_M1001_g 2.99028e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A1_c_105_n N_B1_c_149_n 3.09473e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A1_c_106_n N_B1_c_149_n 0.0170403f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A1_c_111_n N_VPWR_M1002_d 0.00433069f $X=1.362 $Y=1.555 $X2=0 $Y2=0
cc_94 N_A1_c_111_n N_VPWR_c_177_n 0.0045841f $X=1.362 $Y=1.555 $X2=0 $Y2=0
cc_95 N_A1_M1005_g N_VPWR_c_178_n 0.00319712f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A1_M1005_g N_VPWR_c_180_n 0.00436487f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A1_M1005_g N_VPWR_c_175_n 0.00606729f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A1_M1005_g N_A_109_297#_c_215_n 0.0121031f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A1_c_106_n N_A_109_297#_c_215_n 9.47875e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A1_c_111_n N_A_109_297#_c_215_n 0.0208947f $X=1.362 $Y=1.555 $X2=0
+ $Y2=0
cc_101 N_A1_c_107_n N_Y_c_240_n 0.00685888f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A1_M1005_g N_Y_c_236_n 5.08735e-19 $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A1_c_105_n N_Y_c_236_n 0.0328402f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A1_c_106_n N_Y_c_236_n 0.00201257f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A1_c_107_n N_Y_c_236_n 0.00138377f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A1_c_111_n N_Y_c_236_n 0.00346597f $X=1.362 $Y=1.555 $X2=0 $Y2=0
cc_107 N_A1_c_105_n N_Y_c_249_n 0.00445013f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A1_c_106_n N_Y_c_249_n 0.00166435f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A1_c_107_n N_Y_c_249_n 0.00217538f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A1_M1005_g N_Y_c_238_n 6.17011e-19 $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A1_M1005_g Y 0.00106135f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A1_c_107_n N_VGND_c_279_n 0.00528321f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A1_c_107_n N_VGND_c_280_n 0.00974305f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B1_M1001_g N_VPWR_c_180_n 0.00557067f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B1_M1001_g N_VPWR_c_175_n 0.011197f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_c_147_n N_Y_c_240_n 0.0103332f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B1_c_147_n N_Y_c_236_n 0.00794198f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_M1001_g N_Y_c_236_n 0.00860214f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_119 B1 N_Y_c_236_n 0.0230504f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B1_c_149_n N_Y_c_236_n 0.00790497f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B1_c_147_n N_Y_c_249_n 0.00533806f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B1_M1001_g N_Y_c_238_n 0.0140715f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_123 B1 N_Y_c_238_n 0.0182285f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B1_c_149_n N_Y_c_238_n 0.00329318f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B1_M1001_g Y 0.00976569f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_c_147_n N_VGND_c_278_n 0.00648481f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_127 B1 N_VGND_c_278_n 0.0101625f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_c_149_n N_VGND_c_278_n 0.00190009f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B1_c_147_n N_VGND_c_279_n 0.00519379f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_147_n N_VGND_c_280_n 0.00995033f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_131 N_VPWR_c_175_n N_A_109_297#_M1006_d 0.00401945f $X=2.07 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_132 N_VPWR_c_175_n N_A_109_297#_M1005_d 0.00464084f $X=2.07 $Y=2.72 $X2=0
+ $Y2=0
cc_133 N_VPWR_c_179_n N_A_109_297#_c_224_n 0.00866598f $X=0.935 $Y=2.72 $X2=0
+ $Y2=0
cc_134 N_VPWR_c_175_n N_A_109_297#_c_224_n 0.00646445f $X=2.07 $Y=2.72 $X2=0
+ $Y2=0
cc_135 N_VPWR_M1002_d N_A_109_297#_c_215_n 0.00466875f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_136 N_VPWR_c_178_n N_A_109_297#_c_215_n 0.0169895f $X=1.1 $Y=2.34 $X2=0 $Y2=0
cc_137 N_VPWR_c_179_n N_A_109_297#_c_215_n 0.00203142f $X=0.935 $Y=2.72 $X2=0
+ $Y2=0
cc_138 N_VPWR_c_180_n N_A_109_297#_c_215_n 0.00247588f $X=2.07 $Y=2.72 $X2=0
+ $Y2=0
cc_139 N_VPWR_c_175_n N_A_109_297#_c_215_n 0.00987224f $X=2.07 $Y=2.72 $X2=0
+ $Y2=0
cc_140 N_VPWR_c_180_n N_A_109_297#_c_231_n 0.011419f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_141 N_VPWR_c_175_n N_A_109_297#_c_231_n 0.00833279f $X=2.07 $Y=2.72 $X2=0
+ $Y2=0
cc_142 N_VPWR_c_175_n N_Y_M1001_d 0.00218354f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_143 N_VPWR_c_180_n Y 0.0189982f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_144 N_VPWR_c_175_n Y 0.0125416f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_145 N_VPWR_c_177_n N_VGND_c_276_n 6.05903e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_146 N_A_109_297#_M1005_d N_Y_c_236_n 2.67876e-19 $X=1.42 $Y=1.485 $X2=0 $Y2=0
cc_147 N_A_109_297#_M1005_d N_Y_c_238_n 0.0023141f $X=1.42 $Y=1.485 $X2=0.832
+ $Y2=0.51
cc_148 N_A_109_297#_c_215_n N_Y_c_238_n 0.00502319f $X=1.47 $Y=1.92 $X2=0.832
+ $Y2=0.51
cc_149 N_Y_c_240_n N_VGND_c_278_n 0.0209024f $X=1.555 $Y=0.38 $X2=0 $Y2=0
cc_150 N_Y_c_240_n N_VGND_c_279_n 0.0190489f $X=1.555 $Y=0.38 $X2=0 $Y2=0
cc_151 N_Y_M1004_d N_VGND_c_280_n 0.00262165f $X=1.42 $Y=0.235 $X2=0 $Y2=0
cc_152 N_Y_c_240_n N_VGND_c_280_n 0.0146397f $X=1.555 $Y=0.38 $X2=0 $Y2=0
cc_153 N_Y_c_249_n N_VGND_c_280_n 2.08993e-19 $X=1.587 $Y=0.825 $X2=0 $Y2=0
cc_154 N_VGND_c_280_n A_109_47# 0.00401615f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
cc_155 N_VGND_c_280_n A_181_47# 0.0104695f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a31oi_2.pxi.spice
* Created: Tue Sep  1 18:55:24 2020
* 
x_PM_SKY130_FD_SC_HD__A31OI_2%A3 N_A3_c_70_n N_A3_M1002_g N_A3_M1001_g
+ N_A3_c_71_n N_A3_M1014_g N_A3_M1007_g A3 A3 N_A3_c_72_n
+ PM_SKY130_FD_SC_HD__A31OI_2%A3
x_PM_SKY130_FD_SC_HD__A31OI_2%A2 N_A2_c_110_n N_A2_M1004_g N_A2_M1000_g
+ N_A2_c_111_n N_A2_M1005_g N_A2_M1013_g A2 A2 N_A2_c_112_n N_A2_c_113_n
+ PM_SKY130_FD_SC_HD__A31OI_2%A2
x_PM_SKY130_FD_SC_HD__A31OI_2%A1 N_A1_M1010_g N_A1_c_156_n N_A1_M1003_g
+ N_A1_c_157_n N_A1_M1008_g N_A1_M1012_g N_A1_c_158_n N_A1_c_159_n A1 A1
+ N_A1_c_160_n N_A1_c_161_n N_A1_c_162_n PM_SKY130_FD_SC_HD__A31OI_2%A1
x_PM_SKY130_FD_SC_HD__A31OI_2%B1 N_B1_c_220_n N_B1_M1006_g N_B1_M1009_g
+ N_B1_c_221_n N_B1_c_222_n N_B1_M1011_g N_B1_M1015_g N_B1_c_223_n B1 B1 B1
+ N_B1_c_225_n N_B1_c_251_p PM_SKY130_FD_SC_HD__A31OI_2%B1
x_PM_SKY130_FD_SC_HD__A31OI_2%A_27_297# N_A_27_297#_M1001_d N_A_27_297#_M1007_d
+ N_A_27_297#_M1013_s N_A_27_297#_M1012_s N_A_27_297#_M1015_s
+ N_A_27_297#_c_276_n N_A_27_297#_c_283_n N_A_27_297#_c_289_n
+ N_A_27_297#_c_333_p N_A_27_297#_c_295_n N_A_27_297#_c_299_n
+ N_A_27_297#_c_296_n N_A_27_297#_c_301_n N_A_27_297#_c_280_n
+ N_A_27_297#_c_287_n N_A_27_297#_c_297_n PM_SKY130_FD_SC_HD__A31OI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__A31OI_2%VPWR N_VPWR_M1001_s N_VPWR_M1000_d N_VPWR_M1010_d
+ N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n VPWR
+ N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_334_n N_VPWR_c_343_n
+ N_VPWR_c_344_n PM_SKY130_FD_SC_HD__A31OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A31OI_2%Y N_Y_M1003_s N_Y_M1008_s N_Y_M1011_d N_Y_M1009_d
+ N_Y_c_400_n N_Y_c_418_n N_Y_c_401_n N_Y_c_404_n N_Y_c_430_n N_Y_c_402_n Y Y Y
+ Y PM_SKY130_FD_SC_HD__A31OI_2%Y
x_PM_SKY130_FD_SC_HD__A31OI_2%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1014_d
+ N_A_27_47#_M1005_d N_A_27_47#_c_470_n PM_SKY130_FD_SC_HD__A31OI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__A31OI_2%VGND N_VGND_M1002_s N_VGND_M1006_s N_VGND_c_493_n
+ N_VGND_c_494_n VGND N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n
+ N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n PM_SKY130_FD_SC_HD__A31OI_2%VGND
x_PM_SKY130_FD_SC_HD__A31OI_2%A_277_47# N_A_277_47#_M1004_s N_A_277_47#_M1003_d
+ N_A_277_47#_c_553_n PM_SKY130_FD_SC_HD__A31OI_2%A_277_47#
cc_1 VNB N_A3_c_70_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A3_c_71_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A3_c_72_n 0.0595485f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_4 VNB N_A2_c_110_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_A2_c_111_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_6 VNB N_A2_c_112_n 0.00319969f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_7 VNB N_A2_c_113_n 0.0327026f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_8 VNB N_A1_c_156_n 0.0222717f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_9 VNB N_A1_c_157_n 0.0172785f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_10 VNB N_A1_c_158_n 0.0163416f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_A1_c_159_n 4.54479e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_160_n 0.0217081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A1_c_161_n 0.00254047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_162_n 0.0298391f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.305
cc_15 VNB N_B1_c_220_n 0.0169195f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_B1_c_221_n 0.0155576f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_17 VNB N_B1_c_222_n 0.0227273f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_18 VNB N_B1_c_223_n 0.00997566f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_19 VNB B1 0.00804951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B1_c_225_n 0.0329828f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_21 VNB N_VPWR_c_334_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_400_n 0.00208743f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_23 VNB N_Y_c_401_n 0.00790145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_402_n 0.0142007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Y 0.00424886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_470_n 0.0104497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_493_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_28 VNB N_VGND_c_494_n 0.00276998f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_29 VNB N_VGND_c_495_n 0.0156958f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_30 VNB N_VGND_c_496_n 0.0673517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_497_n 0.0174893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_498_n 0.240835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_499_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_500_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_277_47#_c_553_n 0.00646116f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_36 VPB N_A3_M1001_g 0.0221004f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A3_M1007_g 0.0178811f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_38 VPB A3 0.00651054f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_39 VPB N_A3_c_72_n 0.0147647f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_40 VPB N_A2_M1000_g 0.0169734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_41 VPB N_A2_M1013_g 0.0178783f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_42 VPB N_A2_c_112_n 0.00117989f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_43 VPB N_A2_c_113_n 0.00616604f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_44 VPB N_A1_M1010_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_45 VPB N_A1_M1012_g 0.0238063f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_46 VPB N_A1_c_158_n 0.00236409f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_A1_c_159_n 6.90647e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A1_c_160_n 0.00875738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A1_c_161_n 0.00291486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A1_c_162_n 0.0127098f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.305
cc_51 VPB N_B1_M1009_g 0.0195598f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_52 VPB N_B1_c_221_n 0.00474242f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_53 VPB N_B1_M1015_g 0.0225981f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_54 VPB N_B1_c_223_n 6.43591e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_55 VPB B1 0.0130867f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_B1_c_225_n 0.0113063f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_57 VPB N_VPWR_c_335_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_58 VPB N_VPWR_c_336_n 3.21049e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_337_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_338_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_339_n 0.0159043f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_62 VPB N_VPWR_c_340_n 0.0172297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_341_n 0.0431879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_334_n 0.0469402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_343_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_344_n 0.0198531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_Y_c_404_n 0.0032006f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_68 VPB Y 5.51301e-19 $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.305
cc_69 VPB Y 0.00182448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 N_A3_c_71_n N_A2_c_110_n 0.0267608f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_71 N_A3_M1007_g N_A2_M1000_g 0.0263282f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_72 A3 N_A2_M1000_g 2.26074e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_73 A3 N_A2_c_112_n 0.0436822f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A3_c_72_n N_A2_c_112_n 0.00547121f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 A3 N_A2_c_113_n 2.65639e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A3_c_72_n N_A2_c_113_n 0.0217198f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_77 A3 N_A_27_297#_M1001_d 0.00937732f $X=0.61 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_78 N_A3_M1001_g N_A_27_297#_c_276_n 0.00936448f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A3_M1007_g N_A_27_297#_c_276_n 0.0137183f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_80 A3 N_A_27_297#_c_276_n 0.0241617f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A3_c_72_n N_A_27_297#_c_276_n 3.35338e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_82 A3 N_A_27_297#_c_280_n 0.0145285f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A3_c_72_n N_A_27_297#_c_280_n 7.02443e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_84 A3 N_VPWR_M1001_s 0.00172977f $X=0.61 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_85 N_A3_M1001_g N_VPWR_c_335_n 0.0107254f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A3_M1007_g N_VPWR_c_335_n 0.00889062f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A3_M1007_g N_VPWR_c_336_n 5.47116e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A3_M1007_g N_VPWR_c_337_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A3_M1001_g N_VPWR_c_339_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A3_M1001_g N_VPWR_c_334_n 0.00515525f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A3_M1007_g N_VPWR_c_334_n 0.00422825f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A3_c_70_n N_A_27_47#_c_470_n 0.00954728f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A3_c_71_n N_A_27_47#_c_470_n 0.0139452f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_94 A3 N_A_27_47#_c_470_n 0.0457839f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A3_c_72_n N_A_27_47#_c_470_n 0.00881276f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A3_c_70_n N_VGND_c_493_n 0.0152492f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A3_c_71_n N_VGND_c_493_n 0.00930495f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A3_c_70_n N_VGND_c_495_n 0.00341689f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A3_c_71_n N_VGND_c_496_n 0.00341689f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A3_c_70_n N_VGND_c_498_n 0.0050171f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A3_c_71_n N_VGND_c_498_n 0.00405445f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A3_c_71_n N_A_277_47#_c_553_n 4.913e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A2_M1013_g N_A1_M1010_g 0.0264319f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A2_c_112_n N_A1_M1010_g 2.79246e-19 $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A2_c_112_n N_A1_c_158_n 3.33588e-19 $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A2_c_113_n N_A1_c_158_n 0.0216834f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A2_c_112_n N_A1_c_161_n 0.0487326f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A2_c_113_n N_A1_c_161_n 0.004454f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A2_c_112_n N_A_27_297#_M1007_d 0.00268034f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A2_M1000_g N_A_27_297#_c_283_n 0.00936448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A2_M1013_g N_A_27_297#_c_283_n 0.010861f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A2_c_112_n N_A_27_297#_c_283_n 0.0313067f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A2_c_113_n N_A_27_297#_c_283_n 3.35338e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A2_c_112_n N_A_27_297#_c_287_n 0.0114089f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A2_c_112_n N_VPWR_M1000_d 0.00172977f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A2_M1000_g N_VPWR_c_335_n 5.47116e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A2_M1000_g N_VPWR_c_336_n 0.00894861f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A2_M1013_g N_VPWR_c_336_n 0.00921012f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A2_M1000_g N_VPWR_c_337_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A2_M1013_g N_VPWR_c_340_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A2_M1000_g N_VPWR_c_334_n 0.00422825f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A2_M1013_g N_VPWR_c_334_n 0.00422825f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A2_c_110_n N_A_27_47#_c_470_n 0.00956275f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A2_c_111_n N_A_27_47#_c_470_n 0.00997392f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A2_c_112_n N_A_27_47#_c_470_n 0.0484422f $X=1.67 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A2_c_113_n N_A_27_47#_c_470_n 0.00323803f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A2_c_110_n N_VGND_c_493_n 0.0018398f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A2_c_110_n N_VGND_c_496_n 0.00415639f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_111_n N_VGND_c_496_n 0.00366111f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_110_n N_VGND_c_498_n 0.00578549f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_c_111_n N_VGND_c_498_n 0.00661716f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A2_c_110_n N_A_277_47#_c_553_n 0.00365451f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_111_n N_A_277_47#_c_553_n 0.0101156f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A1_c_157_n N_B1_c_220_n 0.0185071f $X=3.12 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_135 N_A1_M1012_g N_B1_M1009_g 0.0185071f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A1_c_159_n N_B1_c_223_n 2.31662e-19 $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_c_162_n N_B1_c_223_n 0.0185071f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_c_161_n N_A_27_297#_M1013_s 0.00188529f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A1_M1010_g N_A_27_297#_c_289_n 0.0117091f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_M1012_g N_A_27_297#_c_289_n 0.0178105f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_c_159_n N_A_27_297#_c_289_n 0.00468836f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A1_c_160_n N_A_27_297#_c_289_n 0.00129833f $X=2.595 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A1_c_161_n N_A_27_297#_c_289_n 0.0420303f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A1_c_162_n N_A_27_297#_c_289_n 0.00743936f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A1_M1012_g N_A_27_297#_c_295_n 0.00528901f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1012_g N_A_27_297#_c_296_n 0.0018177f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_c_161_n N_A_27_297#_c_297_n 0.00561531f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A1_c_161_n N_VPWR_M1010_d 0.00791891f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A1_M1010_g N_VPWR_c_336_n 5.93951e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A1_M1010_g N_VPWR_c_340_n 0.00585385f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A1_M1012_g N_VPWR_c_341_n 0.00585385f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1010_g N_VPWR_c_334_n 0.00752222f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A1_M1012_g N_VPWR_c_334_n 0.00773145f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A1_M1010_g N_VPWR_c_344_n 0.0118402f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A1_M1012_g N_VPWR_c_344_n 0.0143674f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A1_c_156_n N_Y_c_400_n 0.0109066f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A1_c_157_n N_Y_c_400_n 0.013409f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A1_c_159_n N_Y_c_400_n 0.010318f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_c_160_n N_Y_c_400_n 0.00665969f $X=2.595 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_c_161_n N_Y_c_400_n 0.0264627f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A1_c_162_n N_Y_c_400_n 0.00301263f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A1_M1012_g Y 0.00277982f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A1_c_161_n Y 0.00611586f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A1_c_157_n Y 0.00962256f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_159_n Y 0.0237769f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_c_161_n Y 0.00439959f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A1_c_158_n N_A_27_47#_c_470_n 0.00213605f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A1_c_161_n N_A_27_47#_c_470_n 0.0119666f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A1_c_157_n N_VGND_c_494_n 0.00104176f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_156_n N_VGND_c_496_n 0.00366111f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_157_n N_VGND_c_496_n 0.00415639f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A1_c_156_n N_VGND_c_498_n 0.0066948f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_157_n N_VGND_c_498_n 0.00602414f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_156_n N_A_277_47#_c_553_n 0.0101156f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A1_c_157_n N_A_277_47#_c_553_n 0.00253136f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A1_c_158_n N_A_277_47#_c_553_n 0.00415574f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A1_c_161_n N_A_277_47#_c_553_n 0.00632968f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_178 B1 N_A_27_297#_M1015_s 0.00602613f $X=4.28 $Y=1.445 $X2=0 $Y2=0
cc_179 N_B1_M1009_g N_A_27_297#_c_299_n 0.0126304f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1015_g N_A_27_297#_c_299_n 0.0117554f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_181 B1 N_A_27_297#_c_301_n 0.0140093f $X=4.28 $Y=1.445 $X2=0 $Y2=0
cc_182 N_B1_c_225_n N_A_27_297#_c_301_n 8.29256e-19 $X=4.325 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B1_M1009_g N_VPWR_c_341_n 0.00357877f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1015_g N_VPWR_c_341_n 0.00357877f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1009_g N_VPWR_c_334_n 0.00566282f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_M1015_g N_VPWR_c_334_n 0.00638447f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B1_c_220_n N_Y_c_418_n 0.00593249f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_220_n N_Y_c_401_n 0.011021f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_221_n N_Y_c_401_n 0.00405806f $X=4.055 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B1_c_222_n N_Y_c_401_n 0.0100337f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_191 B1 N_Y_c_401_n 0.0141344f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_192 N_B1_c_225_n N_Y_c_401_n 0.00668981f $X=4.325 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B1_c_251_p N_Y_c_401_n 0.0201082f $X=4.265 $Y=1.175 $X2=0 $Y2=0
cc_194 N_B1_M1009_g N_Y_c_404_n 0.0140932f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_c_221_n N_Y_c_404_n 0.00436748f $X=4.055 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B1_M1015_g N_Y_c_404_n 0.00290127f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_197 B1 N_Y_c_404_n 0.0130906f $X=4.28 $Y=1.445 $X2=0 $Y2=0
cc_198 N_B1_c_251_p N_Y_c_404_n 0.0214133f $X=4.265 $Y=1.175 $X2=0 $Y2=0
cc_199 N_B1_M1015_g N_Y_c_430_n 0.0115884f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_200 B1 N_Y_c_430_n 6.85526e-19 $X=4.28 $Y=1.445 $X2=0 $Y2=0
cc_201 N_B1_c_220_n N_Y_c_402_n 6.43414e-19 $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_222_n N_Y_c_402_n 0.00580295f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B1_c_220_n Y 0.00300792f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B1_M1009_g Y 0.00303095f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B1_c_220_n Y 0.00515573f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B1_M1009_g Y 0.00362128f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_c_222_n Y 7.82988e-19 $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B1_M1015_g Y 5.50641e-19 $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_c_223_n Y 0.0141203f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B1_c_251_p Y 0.0115438f $X=4.265 $Y=1.175 $X2=0 $Y2=0
cc_211 N_B1_c_220_n N_VGND_c_494_n 0.00835481f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_222_n N_VGND_c_494_n 0.00417809f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_220_n N_VGND_c_496_n 0.00341675f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_222_n N_VGND_c_497_n 0.00417062f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_220_n N_VGND_c_498_n 0.00426746f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_222_n N_VGND_c_498_n 0.00678426f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_27_297#_c_276_n N_VPWR_M1001_s 0.00317012f $X=1.015 $Y=1.87 $X2=0.47
+ $Y2=0.995
cc_218 N_A_27_297#_c_283_n N_VPWR_M1000_d 0.00317012f $X=1.855 $Y=1.87 $X2=0.47
+ $Y2=0.56
cc_219 N_A_27_297#_c_289_n N_VPWR_M1010_d 0.0204381f $X=3.335 $Y=1.87 $X2=0.47
+ $Y2=0.56
cc_220 N_A_27_297#_c_276_n N_VPWR_c_335_n 0.0165384f $X=1.015 $Y=1.87 $X2=0.89
+ $Y2=1.985
cc_221 N_A_27_297#_c_283_n N_VPWR_c_336_n 0.0165384f $X=1.855 $Y=1.87 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_c_287_n N_VPWR_c_337_n 0.0113958f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_223 N_A_27_297#_c_280_n N_VPWR_c_339_n 0.0116048f $X=0.26 $Y=1.95 $X2=0.47
+ $Y2=1.16
cc_224 N_A_27_297#_c_297_n N_VPWR_c_340_n 0.0113958f $X=1.94 $Y=1.95 $X2=0 $Y2=0
cc_225 N_A_27_297#_c_299_n N_VPWR_c_341_n 0.0526088f $X=4.255 $Y=2.38 $X2=0
+ $Y2=0
cc_226 N_A_27_297#_c_296_n N_VPWR_c_341_n 0.0117106f $X=3.505 $Y=2.38 $X2=0
+ $Y2=0
cc_227 N_A_27_297#_M1001_d N_VPWR_c_334_n 0.00378138f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_228 N_A_27_297#_M1007_d N_VPWR_c_334_n 0.00268171f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_229 N_A_27_297#_M1013_s N_VPWR_c_334_n 0.00268171f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_A_27_297#_M1012_s N_VPWR_c_334_n 0.00366244f $X=3.195 $Y=1.485 $X2=0
+ $Y2=0
cc_231 N_A_27_297#_M1015_s N_VPWR_c_334_n 0.00348186f $X=4.205 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_27_297#_c_276_n N_VPWR_c_334_n 0.0117708f $X=1.015 $Y=1.87 $X2=0
+ $Y2=0
cc_233 N_A_27_297#_c_283_n N_VPWR_c_334_n 0.0117708f $X=1.855 $Y=1.87 $X2=0
+ $Y2=0
cc_234 N_A_27_297#_c_289_n N_VPWR_c_334_n 0.0236525f $X=3.335 $Y=1.87 $X2=0
+ $Y2=0
cc_235 N_A_27_297#_c_299_n N_VPWR_c_334_n 0.0329665f $X=4.255 $Y=2.38 $X2=0
+ $Y2=0
cc_236 N_A_27_297#_c_296_n N_VPWR_c_334_n 0.006547f $X=3.505 $Y=2.38 $X2=0 $Y2=0
cc_237 N_A_27_297#_c_280_n N_VPWR_c_334_n 0.00646998f $X=0.26 $Y=1.95 $X2=0
+ $Y2=0
cc_238 N_A_27_297#_c_287_n N_VPWR_c_334_n 0.00646998f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_239 N_A_27_297#_c_297_n N_VPWR_c_334_n 0.00646998f $X=1.94 $Y=1.95 $X2=0
+ $Y2=0
cc_240 N_A_27_297#_c_289_n N_VPWR_c_344_n 0.0527982f $X=3.335 $Y=1.87 $X2=0
+ $Y2=0
cc_241 N_A_27_297#_c_295_n N_VPWR_c_344_n 0.00797239f $X=3.42 $Y=2.295 $X2=0
+ $Y2=0
cc_242 N_A_27_297#_c_296_n N_VPWR_c_344_n 0.00883915f $X=3.505 $Y=2.38 $X2=0
+ $Y2=0
cc_243 N_A_27_297#_c_299_n N_Y_M1009_d 0.00478617f $X=4.255 $Y=2.38 $X2=0.47
+ $Y2=1.325
cc_244 N_A_27_297#_c_299_n N_Y_c_430_n 0.0190265f $X=4.255 $Y=2.38 $X2=0.605
+ $Y2=1.16
cc_245 N_A_27_297#_M1012_s Y 0.00533555f $X=3.195 $Y=1.485 $X2=0.695 $Y2=1.305
cc_246 N_A_27_297#_c_289_n Y 0.00647221f $X=3.335 $Y=1.87 $X2=0.695 $Y2=1.305
cc_247 N_A_27_297#_c_333_p Y 0.0146964f $X=3.42 $Y=1.955 $X2=0.695 $Y2=1.305
cc_248 N_VPWR_c_334_n N_Y_M1009_d 0.0028108f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_249 N_Y_c_400_n N_A_27_47#_c_470_n 0.0145425f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_250 N_Y_c_401_n N_VGND_M1006_s 0.00533383f $X=4.175 $Y=0.74 $X2=0 $Y2=0
cc_251 N_Y_c_418_n N_VGND_c_494_n 0.0115284f $X=3.34 $Y=0.42 $X2=0 $Y2=0
cc_252 N_Y_c_401_n N_VGND_c_494_n 0.0182521f $X=4.175 $Y=0.74 $X2=0 $Y2=0
cc_253 N_Y_c_400_n N_VGND_c_496_n 0.0024261f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_254 N_Y_c_418_n N_VGND_c_496_n 0.0118139f $X=3.34 $Y=0.42 $X2=0 $Y2=0
cc_255 N_Y_c_401_n N_VGND_c_496_n 0.00162524f $X=4.175 $Y=0.74 $X2=0 $Y2=0
cc_256 Y N_VGND_c_496_n 0.00213984f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_257 N_Y_c_401_n N_VGND_c_497_n 0.00232396f $X=4.175 $Y=0.74 $X2=0 $Y2=0
cc_258 N_Y_c_402_n N_VGND_c_497_n 0.0164902f $X=4.34 $Y=0.38 $X2=0 $Y2=0
cc_259 N_Y_M1003_s N_VGND_c_498_n 0.00212464f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_260 N_Y_M1008_s N_VGND_c_498_n 0.00360908f $X=3.195 $Y=0.235 $X2=0 $Y2=0
cc_261 N_Y_M1011_d N_VGND_c_498_n 0.00211564f $X=4.205 $Y=0.235 $X2=0 $Y2=0
cc_262 N_Y_c_400_n N_VGND_c_498_n 0.00590784f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_263 N_Y_c_418_n N_VGND_c_498_n 0.00646998f $X=3.34 $Y=0.42 $X2=0 $Y2=0
cc_264 N_Y_c_401_n N_VGND_c_498_n 0.00802915f $X=4.175 $Y=0.74 $X2=0 $Y2=0
cc_265 N_Y_c_402_n N_VGND_c_498_n 0.0120857f $X=4.34 $Y=0.38 $X2=0 $Y2=0
cc_266 Y N_VGND_c_498_n 0.00422206f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_267 N_Y_c_400_n N_A_277_47#_M1003_d 0.00484436f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_268 N_Y_M1003_s N_A_277_47#_c_553_n 0.0048485f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_269 N_Y_c_400_n N_A_277_47#_c_553_n 0.0374379f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_270 N_Y_c_418_n N_A_277_47#_c_553_n 0.012629f $X=3.34 $Y=0.42 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_470_n N_VGND_M1002_s 0.00313177f $X=1.94 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_272 N_A_27_47#_c_470_n N_VGND_c_493_n 0.0145262f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_470_n N_VGND_c_495_n 0.00649125f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_470_n N_VGND_c_496_n 0.00740101f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_27_47#_M1002_d N_VGND_c_498_n 0.00312512f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1014_d N_VGND_c_498_n 0.00323135f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_M1005_d N_VGND_c_498_n 0.00212464f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_470_n N_VGND_c_498_n 0.027121f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_470_n N_A_277_47#_M1004_s 0.00313543f $X=1.94 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_280 N_A_27_47#_M1005_d N_A_277_47#_c_553_n 0.00502908f $X=1.805 $Y=0.235
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_470_n N_A_277_47#_c_553_n 0.0355537f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_VGND_c_498_n N_A_277_47#_M1004_s 0.00217615f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_283 N_VGND_c_498_n N_A_277_47#_M1003_d 0.00241975f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_493_n N_A_277_47#_c_553_n 0.00545039f $X=0.68 $Y=0.38 $X2=0
+ $Y2=0
cc_285 N_VGND_c_496_n N_A_277_47#_c_553_n 0.0790384f $X=3.675 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_498_n N_A_277_47#_c_553_n 0.060558f $X=4.37 $Y=0 $X2=0 $Y2=0

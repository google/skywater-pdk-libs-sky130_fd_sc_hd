* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_461_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=2.7e+11p ps=2.54e+06u
M1001 a_461_297# A2 a_333_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=4.9e+11p ps=2.98e+06u
M1002 Y B2 a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=6.1e+11p pd=3.22e+06u as=2.1e+11p ps=2.42e+06u
M1003 VGND A3 a_27_47# VNB nshort w=650000u l=150000u
+  ad=6.7275e+11p pd=4.67e+06u as=5.46e+11p ps=5.58e+06u
M1004 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_109_297# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_333_297# A3 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.1125e+11p pd=1.95e+06u as=0p ps=0u
M1009 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__o311ai_1.pxi.spice
* Created: Tue Sep  1 19:24:45 2020
* 
x_PM_SKY130_FD_SC_HD__O311AI_1%A1 N_A1_c_50_n N_A1_M1006_g N_A1_M1009_g A1 A1
+ N_A1_c_52_n PM_SKY130_FD_SC_HD__O311AI_1%A1
x_PM_SKY130_FD_SC_HD__O311AI_1%A2 N_A2_c_73_n N_A2_M1000_g N_A2_M1002_g A2
+ N_A2_c_75_n PM_SKY130_FD_SC_HD__O311AI_1%A2
x_PM_SKY130_FD_SC_HD__O311AI_1%A3 N_A3_M1003_g N_A3_M1001_g A3 N_A3_c_110_n
+ N_A3_c_111_n PM_SKY130_FD_SC_HD__O311AI_1%A3
x_PM_SKY130_FD_SC_HD__O311AI_1%B1 N_B1_M1004_g N_B1_M1008_g B1 N_B1_c_141_n
+ N_B1_c_142_n PM_SKY130_FD_SC_HD__O311AI_1%B1
x_PM_SKY130_FD_SC_HD__O311AI_1%C1 N_C1_c_175_n N_C1_M1007_g N_C1_M1005_g C1
+ N_C1_c_177_n PM_SKY130_FD_SC_HD__O311AI_1%C1
x_PM_SKY130_FD_SC_HD__O311AI_1%VPWR N_VPWR_M1009_s N_VPWR_M1004_d N_VPWR_c_201_n
+ N_VPWR_c_202_n N_VPWR_c_203_n N_VPWR_c_204_n N_VPWR_c_205_n VPWR
+ N_VPWR_c_206_n N_VPWR_c_200_n PM_SKY130_FD_SC_HD__O311AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O311AI_1%Y N_Y_M1007_d N_Y_M1001_d N_Y_M1005_d N_Y_c_244_n
+ Y Y Y Y Y Y Y Y Y PM_SKY130_FD_SC_HD__O311AI_1%Y
x_PM_SKY130_FD_SC_HD__O311AI_1%VGND N_VGND_M1006_s N_VGND_M1000_d N_VGND_c_279_n
+ N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n VGND N_VGND_c_283_n
+ N_VGND_c_284_n N_VGND_c_285_n PM_SKY130_FD_SC_HD__O311AI_1%VGND
x_PM_SKY130_FD_SC_HD__O311AI_1%A_138_47# N_A_138_47#_M1006_d N_A_138_47#_M1003_d
+ N_A_138_47#_c_335_n N_A_138_47#_c_321_n N_A_138_47#_c_320_n
+ N_A_138_47#_c_331_n PM_SKY130_FD_SC_HD__O311AI_1%A_138_47#
cc_1 VNB N_A1_c_50_n 0.0213312f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.995
cc_2 VNB A1 0.0184734f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_3 VNB N_A1_c_52_n 0.0323103f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.16
cc_4 VNB N_A2_c_73_n 0.0162214f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.995
cc_5 VNB A2 0.00267852f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_A2_c_75_n 0.0200136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB A3 0.00405923f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A3_c_110_n 0.021583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A3_c_111_n 0.0186451f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_10 VNB B1 0.00139441f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_11 VNB N_B1_c_141_n 0.0265384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_142_n 0.0175573f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_13 VNB N_C1_c_175_n 0.0188874f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.995
cc_14 VNB C1 0.0122044f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_C1_c_177_n 0.0397748f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_16 VNB N_VPWR_c_200_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB Y 0.0304446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.00667466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_279_n 0.0129985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_280_n 0.0318775f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_21 VNB N_VGND_c_281_n 0.0117571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_282_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_283_n 0.0479725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_284_n 0.181396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_285_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A1_M1009_g 0.0246762f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_27 VPB A1 0.00342191f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_28 VPB N_A1_c_52_n 0.00814889f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.16
cc_29 VPB N_A2_M1002_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_30 VPB A2 0.00348948f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_31 VPB N_A2_c_75_n 0.00563225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A3_M1001_g 0.0209139f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_33 VPB A3 0.00132946f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_34 VPB N_A3_c_110_n 0.00407411f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_B1_M1004_g 0.0219765f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.56
cc_36 VPB N_B1_c_141_n 0.00554115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_C1_M1005_g 0.0234627f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_38 VPB C1 0.00149016f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_39 VPB N_C1_c_177_n 0.01158f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_40 VPB N_VPWR_c_201_n 0.0157691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_202_n 0.0535914f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_42 VPB N_VPWR_c_203_n 0.00561515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_204_n 0.0346647f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_44 VPB N_VPWR_c_205_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_206_n 0.0211221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_200_n 0.0441037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB Y 0.00931654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB Y 0.0376231f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_49 VPB Y 0.00751936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 N_A1_c_50_n N_A2_c_73_n 0.0236382f $X=0.615 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_51 N_A1_M1009_g N_A2_M1002_g 0.0603914f $X=0.615 $Y=1.985 $X2=0 $Y2=0
cc_52 N_A1_M1009_g A2 0.00334254f $X=0.615 $Y=1.985 $X2=0 $Y2=0
cc_53 A1 A2 0.027727f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A1_c_52_n A2 3.14876e-19 $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_55 A1 N_A2_c_75_n 0.00215956f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A1_c_52_n N_A2_c_75_n 0.0202495f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A1_M1009_g N_VPWR_c_202_n 0.0296774f $X=0.615 $Y=1.985 $X2=0 $Y2=0
cc_58 A1 N_VPWR_c_202_n 0.0530866f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A1_c_52_n N_VPWR_c_202_n 0.00611614f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A1_c_50_n N_VGND_c_280_n 0.0117393f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_61 A1 N_VGND_c_280_n 0.0382706f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A1_c_52_n N_VGND_c_280_n 0.00611614f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A1_c_50_n N_VGND_c_281_n 0.0046653f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A1_c_50_n N_VGND_c_282_n 5.54209e-19 $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A1_c_50_n N_VGND_c_284_n 0.00799591f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_66 A1 N_A_138_47#_c_320_n 0.0031152f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A2_M1002_g N_A3_M1001_g 0.0559324f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_68 A2 A3 0.0261953f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A2_c_75_n A3 3.1636e-19 $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_70 A2 N_A3_c_110_n 0.012346f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A2_c_75_n N_A3_c_110_n 0.0201852f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A2_c_73_n N_A3_c_111_n 0.0273838f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A2_M1002_g N_VPWR_c_202_n 0.00665426f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A2_M1002_g N_VPWR_c_204_n 0.00357877f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_75 A2 N_VPWR_c_204_n 0.0190217f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A2_M1002_g N_VPWR_c_200_n 0.00532055f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_77 A2 N_VPWR_c_200_n 0.0112467f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_78 A2 A_222_297# 0.0091484f $X=1.065 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_79 A2 N_Y_c_244_n 0.0140159f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A2_M1002_g Y 7.29289e-19 $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_81 A2 Y 0.0644441f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A2_c_73_n N_VGND_c_280_n 6.99357e-19 $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A2_c_73_n N_VGND_c_281_n 0.00341689f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A2_c_73_n N_VGND_c_282_n 0.00681952f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A2_c_73_n N_VGND_c_284_n 0.00405445f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A2_c_73_n N_A_138_47#_c_321_n 0.0102357f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_87 A2 N_A_138_47#_c_321_n 0.0218658f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_88 N_A2_c_75_n N_A_138_47#_c_321_n 0.00122018f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A2_c_75_n N_A_138_47#_c_320_n 2.71297e-19 $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A3_M1001_g N_B1_M1004_g 0.0297906f $X=1.455 $Y=1.985 $X2=0 $Y2=0
cc_91 A3 B1 0.0221833f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A3_c_110_n B1 3.42843e-19 $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A3_c_111_n B1 0.00335495f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_94 A3 N_B1_c_141_n 0.00235967f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A3_c_110_n N_B1_c_141_n 0.0113895f $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A3_c_111_n N_B1_c_142_n 0.00990207f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A3_M1001_g N_VPWR_c_204_n 0.00435091f $X=1.455 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A3_M1001_g N_VPWR_c_200_n 0.00760094f $X=1.455 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A3_M1001_g N_Y_c_244_n 0.00683987f $X=1.455 $Y=1.985 $X2=0 $Y2=0
cc_100 A3 N_Y_c_244_n 0.0266038f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A3_c_110_n N_Y_c_244_n 0.00262179f $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A3_M1001_g Y 0.025506f $X=1.455 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A3_c_111_n N_VGND_c_282_n 0.00853411f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A3_c_111_n N_VGND_c_283_n 0.00341689f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A3_c_111_n N_VGND_c_284_n 0.00470573f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_106 A3 N_A_138_47#_c_321_n 0.0229651f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A3_c_110_n N_A_138_47#_c_321_n 0.0015994f $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A3_c_111_n N_A_138_47#_c_321_n 0.0122513f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_109 B1 N_C1_c_175_n 0.00101088f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_110 N_B1_c_142_n N_C1_c_175_n 0.0371541f $X=2.135 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_111 N_B1_M1004_g N_C1_M1005_g 0.017839f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B1_c_141_n N_C1_c_177_n 0.0371541f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B1_M1004_g N_VPWR_c_203_n 0.00320532f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B1_M1004_g N_VPWR_c_204_n 0.00585385f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B1_M1004_g N_VPWR_c_200_n 0.0112137f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_M1004_g N_Y_c_244_n 0.00280657f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B1_M1004_g Y 0.0133675f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_118 B1 Y 0.0144001f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B1_c_141_n Y 0.00541634f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_M1004_g Y 0.00304359f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_121 B1 Y 0.0263972f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B1_c_142_n Y 0.00295127f $X=2.135 $Y=0.995 $X2=0 $Y2=0
cc_123 B1 N_VGND_c_283_n 0.00913452f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B1_c_142_n N_VGND_c_283_n 0.00499673f $X=2.135 $Y=0.995 $X2=0 $Y2=0
cc_125 B1 N_VGND_c_284_n 0.00771639f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B1_c_142_n N_VGND_c_284_n 0.00915061f $X=2.135 $Y=0.995 $X2=0 $Y2=0
cc_127 B1 N_A_138_47#_M1003_d 0.00738627f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_128 B1 N_A_138_47#_c_321_n 0.0110939f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B1_c_142_n N_A_138_47#_c_321_n 6.18624e-19 $X=2.135 $Y=0.995 $X2=0
+ $Y2=0
cc_130 B1 N_A_138_47#_c_331_n 0.0194914f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B1_c_142_n N_A_138_47#_c_331_n 0.00215332f $X=2.135 $Y=0.995 $X2=0
+ $Y2=0
cc_132 N_C1_M1005_g N_VPWR_c_203_n 0.00320532f $X=2.575 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C1_M1005_g N_VPWR_c_206_n 0.00585385f $X=2.575 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C1_M1005_g N_VPWR_c_200_n 0.0118001f $X=2.575 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C1_M1005_g Y 0.0125849f $X=2.575 $Y=1.985 $X2=0 $Y2=0
cc_136 C1 Y 0.0258447f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_137 N_C1_c_177_n Y 0.00978841f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_138 N_C1_c_175_n Y 0.0114181f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_139 C1 Y 0.0254119f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_140 N_C1_c_177_n Y 0.0097006f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_141 N_C1_c_175_n Y 0.00485784f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C1_M1005_g Y 0.00569102f $X=2.575 $Y=1.985 $X2=0 $Y2=0
cc_143 C1 Y 0.0238092f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_144 N_C1_c_177_n Y 0.0108162f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_145 N_C1_c_175_n N_VGND_c_283_n 0.00357877f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_146 N_C1_c_175_n N_VGND_c_284_n 0.00617552f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_147 N_VPWR_c_202_n A_138_297# 0.00912644f $X=0.405 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_148 N_VPWR_c_200_n A_138_297# 0.0073898f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_149 N_VPWR_c_200_n A_222_297# 0.0063341f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_150 N_VPWR_c_200_n N_Y_M1001_d 0.00362055f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_151 N_VPWR_c_200_n N_Y_M1005_d 0.00250309f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_152 N_VPWR_c_204_n Y 0.0343869f $X=2.15 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_200_n Y 0.0206517f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_M1004_d Y 0.00980034f $X=2.13 $Y=1.485 $X2=0 $Y2=0
cc_155 N_VPWR_c_203_n Y 0.0208278f $X=2.315 $Y=1.96 $X2=0 $Y2=0
cc_156 N_VPWR_c_206_n Y 0.032253f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_200_n Y 0.0185907f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_158 Y N_VGND_c_283_n 0.0437346f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_159 N_Y_M1007_d N_VGND_c_284_n 0.00225742f $X=2.65 $Y=0.235 $X2=0 $Y2=0
cc_160 Y N_VGND_c_284_n 0.0256781f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_161 N_VGND_c_284_n N_A_138_47#_M1006_d 0.00412745f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_162 N_VGND_c_284_n N_A_138_47#_M1003_d 0.0133522f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_163 N_VGND_c_281_n N_A_138_47#_c_335_n 0.0112554f $X=1.08 $Y=0 $X2=0 $Y2=0
cc_164 N_VGND_c_284_n N_A_138_47#_c_335_n 0.00644035f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_165 N_VGND_M1000_d N_A_138_47#_c_321_n 0.004964f $X=1.11 $Y=0.235 $X2=0 $Y2=0
cc_166 N_VGND_c_281_n N_A_138_47#_c_321_n 0.00232396f $X=1.08 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_c_282_n N_A_138_47#_c_321_n 0.0160613f $X=1.245 $Y=0.36 $X2=0
+ $Y2=0
cc_168 N_VGND_c_283_n N_A_138_47#_c_321_n 0.00232396f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_169 N_VGND_c_284_n N_A_138_47#_c_321_n 0.00970544f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_c_283_n N_A_138_47#_c_331_n 0.011459f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_171 N_VGND_c_284_n N_A_138_47#_c_331_n 0.00644035f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_172 N_VGND_c_284_n A_458_47# 0.00705923f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

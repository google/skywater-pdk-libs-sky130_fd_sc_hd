* File: sky130_fd_sc_hd__dlxbn_1.pxi.spice
* Created: Thu Aug 27 14:17:49 2020
* 
x_PM_SKY130_FD_SC_HD__DLXBN_1%GATE_N N_GATE_N_c_158_n N_GATE_N_c_153_n
+ N_GATE_N_M1018_g N_GATE_N_c_159_n N_GATE_N_M1009_g N_GATE_N_c_154_n
+ N_GATE_N_c_160_n GATE_N GATE_N N_GATE_N_c_156_n N_GATE_N_c_157_n
+ PM_SKY130_FD_SC_HD__DLXBN_1%GATE_N
x_PM_SKY130_FD_SC_HD__DLXBN_1%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1009_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_c_197_n N_A_27_47#_M1016_g
+ N_A_27_47#_M1021_g N_A_27_47#_c_341_p N_A_27_47#_c_199_n N_A_27_47#_c_200_n
+ N_A_27_47#_c_208_n N_A_27_47#_c_201_n N_A_27_47#_c_209_n N_A_27_47#_c_202_n
+ N_A_27_47#_c_203_n N_A_27_47#_c_211_n N_A_27_47#_c_212_n N_A_27_47#_c_213_n
+ N_A_27_47#_c_214_n N_A_27_47#_c_215_n N_A_27_47#_c_204_n N_A_27_47#_c_217_n
+ N_A_27_47#_c_205_n PM_SKY130_FD_SC_HD__DLXBN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLXBN_1%D N_D_c_353_n N_D_c_354_n N_D_M1003_g N_D_M1004_g
+ N_D_c_355_n N_D_c_359_n D N_D_c_356_n PM_SKY130_FD_SC_HD__DLXBN_1%D
x_PM_SKY130_FD_SC_HD__DLXBN_1%A_299_47# N_A_299_47#_M1003_s N_A_299_47#_M1004_s
+ N_A_299_47#_M1007_g N_A_299_47#_c_403_n N_A_299_47#_M1001_g
+ N_A_299_47#_c_410_n N_A_299_47#_c_405_n N_A_299_47#_c_411_n
+ N_A_299_47#_c_412_n N_A_299_47#_c_406_n N_A_299_47#_c_407_n
+ N_A_299_47#_c_408_n PM_SKY130_FD_SC_HD__DLXBN_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLXBN_1%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1012_g N_A_193_47#_c_493_n N_A_193_47#_M1013_g
+ N_A_193_47#_c_494_n N_A_193_47#_c_495_n N_A_193_47#_c_499_n
+ N_A_193_47#_c_500_n N_A_193_47#_c_501_n N_A_193_47#_c_502_n
+ N_A_193_47#_c_503_n N_A_193_47#_c_504_n N_A_193_47#_c_496_n
+ PM_SKY130_FD_SC_HD__DLXBN_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLXBN_1%A_716_21# N_A_716_21#_M1020_s N_A_716_21#_M1019_s
+ N_A_716_21#_M1006_g N_A_716_21#_M1002_g N_A_716_21#_c_599_n
+ N_A_716_21#_M1017_g N_A_716_21#_M1008_g N_A_716_21#_c_600_n
+ N_A_716_21#_c_601_n N_A_716_21#_c_602_n N_A_716_21#_M1005_g
+ N_A_716_21#_M1014_g N_A_716_21#_c_611_n N_A_716_21#_c_612_n
+ N_A_716_21#_c_613_n N_A_716_21#_c_614_n N_A_716_21#_c_630_p
+ N_A_716_21#_c_626_p N_A_716_21#_c_603_n N_A_716_21#_c_615_n
+ N_A_716_21#_c_604_n N_A_716_21#_c_605_n N_A_716_21#_c_632_p
+ N_A_716_21#_c_638_p PM_SKY130_FD_SC_HD__DLXBN_1%A_716_21#
x_PM_SKY130_FD_SC_HD__DLXBN_1%A_560_47# N_A_560_47#_M1016_d N_A_560_47#_M1012_d
+ N_A_560_47#_c_710_n N_A_560_47#_M1020_g N_A_560_47#_M1019_g
+ N_A_560_47#_c_711_n N_A_560_47#_c_712_n N_A_560_47#_c_722_n
+ N_A_560_47#_c_719_n N_A_560_47#_c_713_n N_A_560_47#_c_720_n
+ N_A_560_47#_c_714_n N_A_560_47#_c_715_n PM_SKY130_FD_SC_HD__DLXBN_1%A_560_47#
x_PM_SKY130_FD_SC_HD__DLXBN_1%A_1124_47# N_A_1124_47#_M1005_s
+ N_A_1124_47#_M1014_s N_A_1124_47#_M1015_g N_A_1124_47#_M1011_g
+ N_A_1124_47#_c_797_n N_A_1124_47#_c_802_n N_A_1124_47#_c_798_n
+ N_A_1124_47#_c_799_n N_A_1124_47#_c_814_n N_A_1124_47#_c_800_n
+ PM_SKY130_FD_SC_HD__DLXBN_1%A_1124_47#
x_PM_SKY130_FD_SC_HD__DLXBN_1%VPWR N_VPWR_M1009_d N_VPWR_M1004_d N_VPWR_M1002_d
+ N_VPWR_M1019_d N_VPWR_M1014_d N_VPWR_c_843_n N_VPWR_c_844_n N_VPWR_c_845_n
+ N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_848_n N_VPWR_c_849_n VPWR
+ N_VPWR_c_850_n N_VPWR_c_851_n N_VPWR_c_852_n N_VPWR_c_853_n N_VPWR_c_854_n
+ N_VPWR_c_842_n N_VPWR_c_856_n N_VPWR_c_857_n N_VPWR_c_858_n N_VPWR_c_859_n
+ PM_SKY130_FD_SC_HD__DLXBN_1%VPWR
x_PM_SKY130_FD_SC_HD__DLXBN_1%Q N_Q_M1017_d N_Q_M1008_d Q Q Q Q N_Q_c_954_n
+ N_Q_c_955_n PM_SKY130_FD_SC_HD__DLXBN_1%Q
x_PM_SKY130_FD_SC_HD__DLXBN_1%Q_N N_Q_N_M1015_d N_Q_N_M1011_d N_Q_N_c_979_n
+ N_Q_N_c_982_n N_Q_N_c_980_n Q_N Q_N Q_N PM_SKY130_FD_SC_HD__DLXBN_1%Q_N
x_PM_SKY130_FD_SC_HD__DLXBN_1%VGND N_VGND_M1018_d N_VGND_M1003_d N_VGND_M1006_d
+ N_VGND_M1020_d N_VGND_M1005_d N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n
+ N_VGND_c_996_n N_VGND_c_997_n VGND N_VGND_c_998_n N_VGND_c_999_n
+ N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n
+ N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n
+ N_VGND_c_1008_n N_VGND_c_1009_n PM_SKY130_FD_SC_HD__DLXBN_1%VGND
cc_1 VNB N_GATE_N_c_153_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_154_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0153903f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_156_n 0.0210048f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_157_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0397112f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_197_n 0.030401f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_8 VNB N_A_27_47#_M1016_g 0.0184067f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_9 VNB N_A_27_47#_c_199_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_200_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_201_n 0.00834675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_202_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_203_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_204_n 0.023029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_205_n 0.0035432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_c_353_n 0.0520733f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_17 VNB N_D_c_354_n 0.0171218f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_18 VNB N_D_c_355_n 0.00634062f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_19 VNB N_D_c_356_n 0.00399698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_299_47#_M1007_g 0.0238123f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_21 VNB N_A_299_47#_c_403_n 0.0263114f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_22 VNB N_A_299_47#_M1001_g 0.00401758f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_23 VNB N_A_299_47#_c_405_n 0.00348116f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB N_A_299_47#_c_406_n 0.0117658f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_25 VNB N_A_299_47#_c_407_n 0.0010594f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_26 VNB N_A_299_47#_c_408_n 0.00247806f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_27 VNB N_A_193_47#_c_493_n 0.0230679f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_28 VNB N_A_193_47#_c_494_n 0.0206359f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_29 VNB N_A_193_47#_c_495_n 0.0139441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_496_n 0.0206501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_716_21#_M1006_g 0.0491883f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_716_21#_c_599_n 0.0193171f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_33 VNB N_A_716_21#_c_600_n 0.0467082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_716_21#_c_601_n 0.0257075f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_35 VNB N_A_716_21#_c_602_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_36 VNB N_A_716_21#_c_603_n 0.00162539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_716_21#_c_604_n 0.00367214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_716_21#_c_605_n 0.00991944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_560_47#_c_710_n 0.019906f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_40 VNB N_A_560_47#_c_711_n 0.0397654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_560_47#_c_712_n 0.00865064f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_42 VNB N_A_560_47#_c_713_n 0.0064658f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_560_47#_c_714_n 0.00443274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_560_47#_c_715_n 0.0086097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_1124_47#_c_797_n 0.00276448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1124_47#_c_798_n 0.00433139f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_47 VNB N_A_1124_47#_c_799_n 0.0227253f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_48 VNB N_A_1124_47#_c_800_n 0.0197028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_842_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Q_c_954_n 0.0053609f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_51 VNB N_Q_c_955_n 0.00350417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Q_N_c_979_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_53 VNB N_Q_N_c_980_n 0.0224379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB Q_N 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_55 VNB N_VGND_c_993_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_994_n 4.89433e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_995_n 0.0105294f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_58 VNB N_VGND_c_996_n 4.01796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_997_n 0.00262354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_998_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_999_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1000_n 0.0412999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1001_n 0.0145977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1002_n 0.0297283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1003_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1004_n 0.359548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1005_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1006_n 0.00469257f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1007_n 0.00632231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1008_n 0.00436333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1009_n 0.00440331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VPB N_GATE_N_c_158_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_73 VPB N_GATE_N_c_159_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_74 VPB N_GATE_N_c_160_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_75 VPB GATE_N 0.0153801f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_76 VPB N_GATE_N_c_156_n 0.0106763f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_77 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_78 VPB N_A_27_47#_M1021_g 0.0208628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_208_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.53
cc_80 VPB N_A_27_47#_c_209_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_202_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_211_n 0.0301745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_212_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_213_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_214_n 0.00264253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_215_n 0.00787946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_204_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_217_n 0.0284794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_D_M1004_g 0.0212065f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_90 VPB N_D_c_355_n 0.0165744f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_91 VPB N_D_c_359_n 0.0136433f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_92 VPB N_D_c_356_n 0.00229947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_299_47#_M1001_g 0.0372975f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_94 VPB N_A_299_47#_c_410_n 0.00699215f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_95 VPB N_A_299_47#_c_411_n 0.00498318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_299_47#_c_412_n 0.00230079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_299_47#_c_407_n 0.00339586f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_98 VPB N_A_193_47#_M1012_g 0.0310778f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_99 VPB N_A_193_47#_c_495_n 0.00802625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_193_47#_c_499_n 0.00297711f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_101 VPB N_A_193_47#_c_500_n 0.00550346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_193_47#_c_501_n 0.00240335f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_103 VPB N_A_193_47#_c_502_n 0.00738175f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_104 VPB N_A_193_47#_c_503_n 0.00114133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_193_47#_c_504_n 0.00897778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_193_47#_c_496_n 0.0447984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_716_21#_M1006_g 0.0152367f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_108 VPB N_A_716_21#_M1002_g 0.0239967f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_109 VPB N_A_716_21#_M1008_g 0.0221973f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_110 VPB N_A_716_21#_c_600_n 0.0228215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_716_21#_c_601_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_112 VPB N_A_716_21#_c_611_n 0.0192026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_716_21#_c_612_n 0.0285551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_716_21#_c_613_n 0.00702551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_716_21#_c_614_n 0.0430898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_716_21#_c_615_n 0.00237098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_716_21#_c_604_n 0.00483831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_716_21#_c_605_n 0.00120305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_560_47#_M1019_g 0.0233445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_560_47#_c_711_n 0.0144191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_560_47#_c_712_n 5.46857e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_122 VPB N_A_560_47#_c_719_n 0.00345844f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_123 VPB N_A_560_47#_c_720_n 0.00463497f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_124 VPB N_A_560_47#_c_714_n 0.00210713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_1124_47#_M1011_g 0.022632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_1124_47#_c_802_n 0.00436529f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_127 VPB N_A_1124_47#_c_798_n 0.0044672f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_128 VPB N_A_1124_47#_c_799_n 0.00492386f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_129 VPB N_VPWR_c_843_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_844_n 0.00329003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_845_n 0.00472845f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_132 VPB N_VPWR_c_846_n 0.00232137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_847_n 0.00289402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_848_n 0.0405103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_849_n 0.0032427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_850_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_851_n 0.0303088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_852_n 0.0222391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_853_n 0.0288878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_854_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_842_n 0.0671165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_856_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_857_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_858_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_859_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB Q 0.00200009f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_147 VPB Q 0.00828788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_Q_c_955_n 0.00475021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_Q_N_c_982_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_150 VPB N_Q_N_c_980_n 0.00978899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB Q_N 0.0318651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 N_GATE_N_c_153_n N_A_27_47#_M1010_g 0.0187834f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_153 N_GATE_N_c_157_n N_A_27_47#_M1010_g 0.00419721f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_154 N_GATE_N_c_160_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_155 N_GATE_N_c_156_n N_A_27_47#_M1000_g 0.00527139f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_156 N_GATE_N_c_153_n N_A_27_47#_c_199_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_157 N_GATE_N_c_154_n N_A_27_47#_c_199_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_158 N_GATE_N_c_154_n N_A_27_47#_c_200_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_159 GATE_N N_A_27_47#_c_200_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_160 N_GATE_N_c_156_n N_A_27_47#_c_200_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_161 N_GATE_N_c_159_n N_A_27_47#_c_208_n 0.0135489f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_162 N_GATE_N_c_160_n N_A_27_47#_c_208_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_163 N_GATE_N_c_159_n N_A_27_47#_c_209_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_164 N_GATE_N_c_160_n N_A_27_47#_c_209_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_165 GATE_N N_A_27_47#_c_209_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_166 N_GATE_N_c_156_n N_A_27_47#_c_209_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_167 N_GATE_N_c_156_n N_A_27_47#_c_202_n 0.00319349f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_168 N_GATE_N_c_154_n N_A_27_47#_c_203_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_169 GATE_N N_A_27_47#_c_203_n 0.0288278f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_170 N_GATE_N_c_157_n N_A_27_47#_c_203_n 0.00151818f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_171 N_GATE_N_c_158_n N_A_27_47#_c_212_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_172 N_GATE_N_c_160_n N_A_27_47#_c_212_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_173 GATE_N N_A_27_47#_c_212_n 0.00653562f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_174 N_GATE_N_c_158_n N_A_27_47#_c_213_n 7.602e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_175 N_GATE_N_c_160_n N_A_27_47#_c_213_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_176 GATE_N N_A_27_47#_c_204_n 9.06856e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_177 N_GATE_N_c_156_n N_A_27_47#_c_204_n 0.0165768f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_178 N_GATE_N_c_159_n N_VPWR_c_843_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_179 N_GATE_N_c_159_n N_VPWR_c_850_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_180 N_GATE_N_c_159_n N_VPWR_c_842_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_181 N_GATE_N_c_153_n N_VGND_c_993_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_182 N_GATE_N_c_153_n N_VGND_c_998_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_183 N_GATE_N_c_154_n N_VGND_c_998_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_184 N_GATE_N_c_153_n N_VGND_c_1004_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1010_g N_D_c_353_n 0.0054595f $X=0.89 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_186 N_A_27_47#_c_211_n N_D_c_353_n 3.18903e-19 $X=2.895 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_27_47#_c_211_n N_D_c_355_n 0.00474321f $X=2.895 $Y=1.53 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_211_n N_D_c_356_n 0.00957673f $X=2.895 $Y=1.53 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_197_n N_A_299_47#_M1007_g 0.00880707f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1016_g N_A_299_47#_M1007_g 0.0247945f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_201_n N_A_299_47#_M1007_g 8.2645e-19 $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_197_n N_A_299_47#_c_403_n 0.00879426f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_205_n N_A_299_47#_c_403_n 8.75667e-19 $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_211_n N_A_299_47#_M1001_g 0.00476495f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_205_n N_A_299_47#_M1001_g 6.68536e-19 $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_211_n N_A_299_47#_c_411_n 0.0120631f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_211_n N_A_299_47#_c_412_n 0.0118176f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_197_n N_A_299_47#_c_406_n 5.80475e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_201_n N_A_299_47#_c_406_n 0.0181483f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_211_n N_A_299_47#_c_406_n 0.00621587f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_205_n N_A_299_47#_c_406_n 0.00677094f $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_211_n N_A_299_47#_c_407_n 0.00907512f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1021_g N_A_193_47#_M1012_g 0.0180503f $X=3.295 $Y=2.275 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_197_n N_A_193_47#_c_493_n 0.0019914f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1016_g N_A_193_47#_c_493_n 0.0129628f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_201_n N_A_193_47#_c_493_n 0.00185589f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_197_n N_A_193_47#_c_494_n 0.0137064f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_201_n N_A_193_47#_c_494_n 0.00224918f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_205_n N_A_193_47#_c_494_n 0.00317732f $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_M1010_g N_A_193_47#_c_495_n 0.00778071f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_199_n N_A_193_47#_c_495_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_202_n N_A_193_47#_c_495_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_203_n N_A_193_47#_c_495_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_211_n N_A_193_47#_c_495_n 0.0185577f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_212_n N_A_193_47#_c_495_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_213_n N_A_193_47#_c_495_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_208_n N_A_193_47#_c_499_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_211_n N_A_193_47#_c_499_n 0.00195186f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_204_n N_A_193_47#_c_499_n 0.00778071f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_211_n N_A_193_47#_c_500_n 0.0891962f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_M1000_g N_A_193_47#_c_501_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_208_n N_A_193_47#_c_501_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_211_n N_A_193_47#_c_501_n 0.0259095f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_213_n N_A_193_47#_c_501_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_M1000_g N_A_193_47#_c_502_n 0.00778071f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_211_n N_A_193_47#_c_503_n 0.0255946f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_215_n N_A_193_47#_c_503_n 0.00104402f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_197_n N_A_193_47#_c_504_n 8.22516e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1021_g N_A_193_47#_c_504_n 5.26344e-19 $X=3.295 $Y=2.275
+ $X2=0 $Y2=0
cc_230 N_A_27_47#_c_201_n N_A_193_47#_c_504_n 0.0088829f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_211_n N_A_193_47#_c_504_n 0.0200219f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_214_n N_A_193_47#_c_504_n 0.00262555f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_217_n N_A_193_47#_c_504_n 2.60208e-19 $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_234 N_A_27_47#_c_205_n N_A_193_47#_c_504_n 0.0393616f $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_197_n N_A_193_47#_c_496_n 0.0204307f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_201_n N_A_193_47#_c_496_n 0.00281201f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_211_n N_A_193_47#_c_496_n 0.00576745f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_214_n N_A_193_47#_c_496_n 0.00289277f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_215_n N_A_193_47#_c_496_n 0.00983293f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_217_n N_A_193_47#_c_496_n 0.0316651f $X=3.205 $Y=1.745 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_205_n N_A_193_47#_c_496_n 0.0157456f $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_215_n N_A_716_21#_M1006_g 9.47199e-19 $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_205_n N_A_716_21#_M1006_g 2.55699e-19 $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1021_g N_A_716_21#_M1002_g 0.0314861f $X=3.295 $Y=2.275 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_215_n N_A_716_21#_c_614_n 2.60641e-19 $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_217_n N_A_716_21#_c_614_n 0.0314861f $X=3.205 $Y=1.745 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_197_n N_A_560_47#_c_722_n 5.71128e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1016_g N_A_560_47#_c_722_n 0.00332918f $X=2.725 $Y=0.415
+ $X2=0 $Y2=0
cc_249 N_A_27_47#_c_201_n N_A_560_47#_c_722_n 0.0210242f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1021_g N_A_560_47#_c_719_n 0.0127001f $X=3.295 $Y=2.275 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_214_n N_A_560_47#_c_719_n 0.0021292f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_215_n N_A_560_47#_c_719_n 0.020881f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_217_n N_A_560_47#_c_719_n 0.00101654f $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_254 N_A_27_47#_c_201_n N_A_560_47#_c_713_n 0.0188625f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_214_n N_A_560_47#_c_720_n 0.00130177f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_215_n N_A_560_47#_c_720_n 0.0367792f $X=3.04 $Y=1.53 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_217_n N_A_560_47#_c_720_n 0.00412397f $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_258 N_A_27_47#_c_205_n N_A_560_47#_c_720_n 0.00387408f $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_201_n N_A_560_47#_c_715_n 0.00293434f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_217_n N_A_560_47#_c_715_n 5.43103e-19 $X=3.205 $Y=1.745
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_205_n N_A_560_47#_c_715_n 0.0164606f $X=3.12 $Y=1.415 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_208_n N_VPWR_M1009_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_263 N_A_27_47#_M1000_g N_VPWR_c_843_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_208_n N_VPWR_c_843_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_209_n N_VPWR_c_843_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_212_n N_VPWR_c_843_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_211_n N_VPWR_c_844_n 0.00101715f $X=2.895 $Y=1.53 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1021_g N_VPWR_c_848_n 0.00394409f $X=3.295 $Y=2.275 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_208_n N_VPWR_c_850_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_209_n N_VPWR_c_850_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_271 N_A_27_47#_M1000_g N_VPWR_c_851_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1000_g N_VPWR_c_842_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1021_g N_VPWR_c_842_n 0.00563532f $X=3.295 $Y=2.275 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_208_n N_VPWR_c_842_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_209_n N_VPWR_c_842_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_199_n N_VGND_M1018_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_277 N_A_27_47#_M1010_g N_VGND_c_993_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_199_n N_VGND_c_993_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_202_n N_VGND_c_993_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_204_n N_VGND_c_993_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_M1016_g N_VGND_c_994_n 0.00193219f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_341_p N_VGND_c_998_n 0.00713694f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_199_n N_VGND_c_998_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_284 N_A_27_47#_M1010_g N_VGND_c_999_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_197_n N_VGND_c_1000_n 2.95456e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1016_g N_VGND_c_1000_n 0.00431421f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_201_n N_VGND_c_1000_n 0.00346042f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1018_s N_VGND_c_1004_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_M1010_g N_VGND_c_1004_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1016_g N_VGND_c_1004_n 0.00627964f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_341_p N_VGND_c_1004_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_199_n N_VGND_c_1004_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_201_n N_VGND_c_1004_n 0.00581168f $X=2.95 $Y=0.87 $X2=0
+ $Y2=0
cc_294 N_D_c_353_n N_A_299_47#_M1007_g 0.00386645f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_295 N_D_c_354_n N_A_299_47#_M1007_g 0.0161181f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_296 N_D_c_353_n N_A_299_47#_c_403_n 0.0199316f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_297 N_D_c_356_n N_A_299_47#_c_403_n 2.66716e-19 $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_298 N_D_c_355_n N_A_299_47#_M1001_g 0.0102066f $X=1.822 $Y=1.565 $X2=0 $Y2=0
cc_299 N_D_c_359_n N_A_299_47#_M1001_g 0.0192108f $X=1.822 $Y=1.715 $X2=0 $Y2=0
cc_300 N_D_M1004_g N_A_299_47#_c_410_n 0.0109158f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_301 N_D_c_359_n N_A_299_47#_c_410_n 0.00368967f $X=1.822 $Y=1.715 $X2=0 $Y2=0
cc_302 N_D_c_353_n N_A_299_47#_c_405_n 0.00913816f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_303 N_D_c_354_n N_A_299_47#_c_405_n 0.00680452f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_304 N_D_c_356_n N_A_299_47#_c_405_n 0.00576082f $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_305 N_D_c_353_n N_A_299_47#_c_411_n 5.96048e-19 $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_306 N_D_c_355_n N_A_299_47#_c_411_n 0.00243526f $X=1.822 $Y=1.565 $X2=0 $Y2=0
cc_307 N_D_c_359_n N_A_299_47#_c_411_n 0.00481255f $X=1.822 $Y=1.715 $X2=0 $Y2=0
cc_308 N_D_c_353_n N_A_299_47#_c_412_n 0.00116923f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_309 N_D_c_355_n N_A_299_47#_c_412_n 0.00306233f $X=1.822 $Y=1.565 $X2=0 $Y2=0
cc_310 N_D_c_359_n N_A_299_47#_c_412_n 0.00279839f $X=1.822 $Y=1.715 $X2=0 $Y2=0
cc_311 N_D_c_356_n N_A_299_47#_c_412_n 0.0212479f $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_312 N_D_c_353_n N_A_299_47#_c_406_n 0.00590642f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_313 N_D_c_356_n N_A_299_47#_c_406_n 0.0191772f $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_314 N_D_c_355_n N_A_299_47#_c_407_n 0.00427242f $X=1.822 $Y=1.565 $X2=0 $Y2=0
cc_315 N_D_c_356_n N_A_299_47#_c_407_n 0.00575207f $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_316 N_D_c_353_n N_A_299_47#_c_408_n 0.00526279f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_317 N_D_c_354_n N_A_299_47#_c_408_n 6.93286e-19 $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_318 N_D_c_356_n N_A_299_47#_c_408_n 0.0138491f $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_319 N_D_c_353_n N_A_193_47#_c_495_n 0.00471466f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_320 N_D_c_355_n N_A_193_47#_c_495_n 0.00484352f $X=1.822 $Y=1.565 $X2=0 $Y2=0
cc_321 N_D_c_356_n N_A_193_47#_c_495_n 0.0218739f $X=1.61 $Y=1.04 $X2=0 $Y2=0
cc_322 N_D_M1004_g N_A_193_47#_c_499_n 0.00127046f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_323 N_D_M1004_g N_A_193_47#_c_500_n 0.00296602f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_324 N_D_M1004_g N_VPWR_c_844_n 0.00304701f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_325 N_D_M1004_g N_VPWR_c_851_n 0.00543342f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_326 N_D_M1004_g N_VPWR_c_842_n 0.00734866f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_327 N_D_c_354_n N_VGND_c_994_n 0.0109478f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_328 N_D_c_354_n N_VGND_c_999_n 0.00337001f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_329 N_D_c_353_n N_VGND_c_1004_n 0.00136965f $X=1.79 $Y=1.205 $X2=0 $Y2=0
cc_330 N_D_c_354_n N_VGND_c_1004_n 0.0053254f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_331 N_A_299_47#_M1001_g N_A_193_47#_M1012_g 0.0342233f $X=2.275 $Y=2.165
+ $X2=0 $Y2=0
cc_332 N_A_299_47#_c_410_n N_A_193_47#_c_495_n 0.00102774f $X=1.645 $Y=1.99
+ $X2=0 $Y2=0
cc_333 N_A_299_47#_c_412_n N_A_193_47#_c_495_n 0.00816005f $X=1.81 $Y=1.58 $X2=0
+ $Y2=0
cc_334 N_A_299_47#_c_408_n N_A_193_47#_c_495_n 0.0191832f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_410_n N_A_193_47#_c_499_n 0.0432762f $X=1.645 $Y=1.99 $X2=0
+ $Y2=0
cc_336 N_A_299_47#_M1001_g N_A_193_47#_c_500_n 0.00334905f $X=2.275 $Y=2.165
+ $X2=0 $Y2=0
cc_337 N_A_299_47#_c_410_n N_A_193_47#_c_500_n 0.0228554f $X=1.645 $Y=1.99 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_411_n N_A_193_47#_c_500_n 0.00551435f $X=1.995 $Y=1.58
+ $X2=0 $Y2=0
cc_339 N_A_299_47#_c_410_n N_A_193_47#_c_501_n 0.0026925f $X=1.645 $Y=1.99 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_M1001_g N_A_193_47#_c_503_n 0.00149195f $X=2.275 $Y=2.165
+ $X2=0 $Y2=0
cc_341 N_A_299_47#_M1001_g N_A_193_47#_c_504_n 0.00673436f $X=2.275 $Y=2.165
+ $X2=0 $Y2=0
cc_342 N_A_299_47#_c_411_n N_A_193_47#_c_504_n 0.00754519f $X=1.995 $Y=1.58
+ $X2=0 $Y2=0
cc_343 N_A_299_47#_c_407_n N_A_193_47#_c_504_n 0.00645446f $X=2.08 $Y=1.495
+ $X2=0 $Y2=0
cc_344 N_A_299_47#_c_403_n N_A_193_47#_c_496_n 5.83528e-19 $X=2.275 $Y=1.235
+ $X2=0 $Y2=0
cc_345 N_A_299_47#_M1001_g N_A_193_47#_c_496_n 0.0247492f $X=2.275 $Y=2.165
+ $X2=0 $Y2=0
cc_346 N_A_299_47#_M1007_g N_A_560_47#_c_722_n 6.41898e-19 $X=2.25 $Y=0.445
+ $X2=0 $Y2=0
cc_347 N_A_299_47#_c_403_n N_VPWR_c_844_n 3.65226e-19 $X=2.275 $Y=1.235 $X2=0
+ $Y2=0
cc_348 N_A_299_47#_M1001_g N_VPWR_c_844_n 0.0219486f $X=2.275 $Y=2.165 $X2=0
+ $Y2=0
cc_349 N_A_299_47#_c_410_n N_VPWR_c_844_n 0.0232987f $X=1.645 $Y=1.99 $X2=0
+ $Y2=0
cc_350 N_A_299_47#_c_411_n N_VPWR_c_844_n 0.013562f $X=1.995 $Y=1.58 $X2=0 $Y2=0
cc_351 N_A_299_47#_c_406_n N_VPWR_c_844_n 0.00151378f $X=2.08 $Y=1.235 $X2=0
+ $Y2=0
cc_352 N_A_299_47#_M1001_g N_VPWR_c_848_n 0.00212864f $X=2.275 $Y=2.165 $X2=0
+ $Y2=0
cc_353 N_A_299_47#_c_410_n N_VPWR_c_851_n 0.0159418f $X=1.645 $Y=1.99 $X2=0
+ $Y2=0
cc_354 N_A_299_47#_M1004_s N_VPWR_c_842_n 0.00174533f $X=1.52 $Y=1.845 $X2=0
+ $Y2=0
cc_355 N_A_299_47#_M1001_g N_VPWR_c_842_n 0.00262666f $X=2.275 $Y=2.165 $X2=0
+ $Y2=0
cc_356 N_A_299_47#_c_410_n N_VPWR_c_842_n 0.00576627f $X=1.645 $Y=1.99 $X2=0
+ $Y2=0
cc_357 N_A_299_47#_c_405_n N_VGND_M1003_d 3.25986e-19 $X=1.995 $Y=0.7 $X2=0
+ $Y2=0
cc_358 N_A_299_47#_c_406_n N_VGND_M1003_d 0.00135909f $X=2.08 $Y=1.235 $X2=0
+ $Y2=0
cc_359 N_A_299_47#_M1007_g N_VGND_c_994_n 0.0112495f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_360 N_A_299_47#_c_403_n N_VGND_c_994_n 2.69913e-19 $X=2.275 $Y=1.235 $X2=0
+ $Y2=0
cc_361 N_A_299_47#_c_405_n N_VGND_c_994_n 0.00448601f $X=1.995 $Y=0.7 $X2=0
+ $Y2=0
cc_362 N_A_299_47#_c_406_n N_VGND_c_994_n 0.012332f $X=2.08 $Y=1.235 $X2=0 $Y2=0
cc_363 N_A_299_47#_c_405_n N_VGND_c_999_n 0.00255672f $X=1.995 $Y=0.7 $X2=0
+ $Y2=0
cc_364 N_A_299_47#_c_408_n N_VGND_c_999_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_365 N_A_299_47#_M1007_g N_VGND_c_1000_n 0.00368966f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_A_299_47#_M1003_s N_VGND_c_1004_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_299_47#_M1007_g N_VGND_c_1004_n 0.00660474f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_368 N_A_299_47#_c_405_n N_VGND_c_1004_n 0.00484661f $X=1.995 $Y=0.7 $X2=0
+ $Y2=0
cc_369 N_A_299_47#_c_406_n N_VGND_c_1004_n 8.89004e-19 $X=2.08 $Y=1.235 $X2=0
+ $Y2=0
cc_370 N_A_299_47#_c_408_n N_VGND_c_1004_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_493_n N_A_716_21#_M1006_g 0.0467823f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_496_n N_A_716_21#_M1006_g 9.79947e-19 $X=2.755 $Y=1.42
+ $X2=0 $Y2=0
cc_373 N_A_193_47#_c_493_n N_A_560_47#_c_722_n 0.0118198f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_496_n N_A_560_47#_c_722_n 2.13332e-19 $X=2.755 $Y=1.42
+ $X2=0 $Y2=0
cc_375 N_A_193_47#_M1012_g N_A_560_47#_c_719_n 0.00283345f $X=2.755 $Y=2.275
+ $X2=0 $Y2=0
cc_376 N_A_193_47#_c_496_n N_A_560_47#_c_719_n 4.93948e-19 $X=2.755 $Y=1.42
+ $X2=0 $Y2=0
cc_377 N_A_193_47#_c_493_n N_A_560_47#_c_713_n 0.00619431f $X=3.18 $Y=0.685
+ $X2=0 $Y2=0
cc_378 N_A_193_47#_M1012_g N_A_560_47#_c_720_n 3.20592e-19 $X=2.755 $Y=2.275
+ $X2=0 $Y2=0
cc_379 N_A_193_47#_c_496_n N_A_560_47#_c_720_n 6.6801e-19 $X=2.755 $Y=1.42 $X2=0
+ $Y2=0
cc_380 N_A_193_47#_c_494_n N_A_560_47#_c_715_n 0.00317352f $X=3.215 $Y=1.175
+ $X2=0 $Y2=0
cc_381 N_A_193_47#_c_500_n N_VPWR_M1004_d 6.81311e-19 $X=2.435 $Y=1.87 $X2=0
+ $Y2=0
cc_382 N_A_193_47#_c_502_n N_VPWR_c_843_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_M1012_g N_VPWR_c_844_n 0.00357312f $X=2.755 $Y=2.275 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_c_500_n N_VPWR_c_844_n 0.0165674f $X=2.435 $Y=1.87 $X2=0
+ $Y2=0
cc_385 N_A_193_47#_c_503_n N_VPWR_c_844_n 0.0013481f $X=2.58 $Y=1.87 $X2=0 $Y2=0
cc_386 N_A_193_47#_c_504_n N_VPWR_c_844_n 0.00972665f $X=2.695 $Y=1.52 $X2=0
+ $Y2=0
cc_387 N_A_193_47#_M1012_g N_VPWR_c_848_n 0.00487021f $X=2.755 $Y=2.275 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_c_504_n N_VPWR_c_848_n 0.00456724f $X=2.695 $Y=1.52 $X2=0
+ $Y2=0
cc_389 N_A_193_47#_c_502_n N_VPWR_c_851_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_390 N_A_193_47#_M1012_g N_VPWR_c_842_n 0.00803197f $X=2.755 $Y=2.275 $X2=0
+ $Y2=0
cc_391 N_A_193_47#_c_500_n N_VPWR_c_842_n 0.0530141f $X=2.435 $Y=1.87 $X2=0
+ $Y2=0
cc_392 N_A_193_47#_c_501_n N_VPWR_c_842_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_393 N_A_193_47#_c_502_n N_VPWR_c_842_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_394 N_A_193_47#_c_503_n N_VPWR_c_842_n 0.0151013f $X=2.58 $Y=1.87 $X2=0 $Y2=0
cc_395 N_A_193_47#_c_504_n N_VPWR_c_842_n 0.00403974f $X=2.695 $Y=1.52 $X2=0
+ $Y2=0
cc_396 N_A_193_47#_c_500_n A_470_369# 0.00119229f $X=2.435 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_397 N_A_193_47#_c_503_n A_470_369# 0.00120144f $X=2.58 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_398 N_A_193_47#_c_504_n A_470_369# 0.0030615f $X=2.695 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_399 N_A_193_47#_c_495_n N_VGND_c_999_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_400 N_A_193_47#_c_493_n N_VGND_c_1000_n 0.00378965f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_401 N_A_193_47#_M1010_d N_VGND_c_1004_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_402 N_A_193_47#_c_493_n N_VGND_c_1004_n 0.00558598f $X=3.18 $Y=0.685 $X2=0
+ $Y2=0
cc_403 N_A_193_47#_c_495_n N_VGND_c_1004_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_404 N_A_716_21#_c_599_n N_A_560_47#_c_710_n 0.0243964f $X=5.015 $Y=0.995
+ $X2=0 $Y2=0
cc_405 N_A_716_21#_c_626_p N_A_560_47#_c_710_n 0.00629098f $X=4.487 $Y=0.84
+ $X2=0 $Y2=0
cc_406 N_A_716_21#_c_603_n N_A_560_47#_c_710_n 0.00560518f $X=4.487 $Y=0.995
+ $X2=0 $Y2=0
cc_407 N_A_716_21#_M1008_g N_A_560_47#_M1019_g 0.0271706f $X=5.015 $Y=1.985
+ $X2=0 $Y2=0
cc_408 N_A_716_21#_c_614_n N_A_560_47#_M1019_g 0.00346217f $X=3.885 $Y=1.7 $X2=0
+ $Y2=0
cc_409 N_A_716_21#_c_630_p N_A_560_47#_M1019_g 0.00856694f $X=4.385 $Y=2.27
+ $X2=0 $Y2=0
cc_410 N_A_716_21#_c_615_n N_A_560_47#_M1019_g 0.00762012f $X=4.487 $Y=1.535
+ $X2=0 $Y2=0
cc_411 N_A_716_21#_c_632_p N_A_560_47#_M1019_g 0.00819586f $X=4.385 $Y=1.755
+ $X2=0 $Y2=0
cc_412 N_A_716_21#_M1006_g N_A_560_47#_c_711_n 0.0153386f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_413 N_A_716_21#_c_613_n N_A_560_47#_c_711_n 0.0074966f $X=4.3 $Y=1.7 $X2=0
+ $Y2=0
cc_414 N_A_716_21#_c_614_n N_A_560_47#_c_711_n 9.14109e-19 $X=3.885 $Y=1.7 $X2=0
+ $Y2=0
cc_415 N_A_716_21#_c_626_p N_A_560_47#_c_711_n 0.00402633f $X=4.487 $Y=0.84
+ $X2=0 $Y2=0
cc_416 N_A_716_21#_c_632_p N_A_560_47#_c_711_n 0.0040439f $X=4.385 $Y=1.755
+ $X2=0 $Y2=0
cc_417 N_A_716_21#_c_638_p N_A_560_47#_c_711_n 0.0142491f $X=4.487 $Y=1.16 $X2=0
+ $Y2=0
cc_418 N_A_716_21#_c_604_n N_A_560_47#_c_712_n 0.014151f $X=5.055 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_716_21#_c_605_n N_A_560_47#_c_712_n 0.0174257f $X=5.055 $Y=1.16 $X2=0
+ $Y2=0
cc_420 N_A_716_21#_c_638_p N_A_560_47#_c_712_n 0.00186446f $X=4.487 $Y=1.16
+ $X2=0 $Y2=0
cc_421 N_A_716_21#_M1002_g N_A_560_47#_c_719_n 0.00953172f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_422 N_A_716_21#_c_630_p N_A_560_47#_c_719_n 0.00225108f $X=4.385 $Y=2.27
+ $X2=0 $Y2=0
cc_423 N_A_716_21#_M1006_g N_A_560_47#_c_713_n 0.00871786f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_424 N_A_716_21#_M1006_g N_A_560_47#_c_720_n 0.0113092f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_425 N_A_716_21#_M1002_g N_A_560_47#_c_720_n 0.00430059f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_426 N_A_716_21#_c_613_n N_A_560_47#_c_720_n 0.0247769f $X=4.3 $Y=1.7 $X2=0
+ $Y2=0
cc_427 N_A_716_21#_c_614_n N_A_560_47#_c_720_n 0.00849091f $X=3.885 $Y=1.7 $X2=0
+ $Y2=0
cc_428 N_A_716_21#_c_630_p N_A_560_47#_c_720_n 0.00363279f $X=4.385 $Y=2.27
+ $X2=0 $Y2=0
cc_429 N_A_716_21#_M1006_g N_A_560_47#_c_714_n 0.0162815f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_430 N_A_716_21#_c_613_n N_A_560_47#_c_714_n 0.0286551f $X=4.3 $Y=1.7 $X2=0
+ $Y2=0
cc_431 N_A_716_21#_c_614_n N_A_560_47#_c_714_n 0.00732235f $X=3.885 $Y=1.7 $X2=0
+ $Y2=0
cc_432 N_A_716_21#_c_638_p N_A_560_47#_c_714_n 0.0277655f $X=4.487 $Y=1.16 $X2=0
+ $Y2=0
cc_433 N_A_716_21#_M1006_g N_A_560_47#_c_715_n 0.00683303f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_434 N_A_716_21#_c_611_n N_A_1124_47#_M1011_g 0.0100318f $X=5.952 $Y=1.62
+ $X2=0 $Y2=0
cc_435 N_A_716_21#_c_612_n N_A_1124_47#_M1011_g 0.01223f $X=5.952 $Y=1.77 $X2=0
+ $Y2=0
cc_436 N_A_716_21#_c_599_n N_A_1124_47#_c_797_n 0.00417556f $X=5.015 $Y=0.995
+ $X2=0 $Y2=0
cc_437 N_A_716_21#_c_601_n N_A_1124_47#_c_797_n 0.0102162f $X=5.95 $Y=1.325
+ $X2=0 $Y2=0
cc_438 N_A_716_21#_c_602_n N_A_1124_47#_c_797_n 0.00951761f $X=5.955 $Y=0.73
+ $X2=0 $Y2=0
cc_439 N_A_716_21#_c_611_n N_A_1124_47#_c_802_n 0.011231f $X=5.952 $Y=1.62 $X2=0
+ $Y2=0
cc_440 N_A_716_21#_c_612_n N_A_1124_47#_c_802_n 0.019991f $X=5.952 $Y=1.77 $X2=0
+ $Y2=0
cc_441 N_A_716_21#_c_601_n N_A_1124_47#_c_798_n 0.017655f $X=5.95 $Y=1.325 $X2=0
+ $Y2=0
cc_442 N_A_716_21#_c_601_n N_A_1124_47#_c_799_n 0.0214963f $X=5.95 $Y=1.325
+ $X2=0 $Y2=0
cc_443 N_A_716_21#_c_600_n N_A_1124_47#_c_814_n 0.0177004f $X=5.875 $Y=1.16
+ $X2=0 $Y2=0
cc_444 N_A_716_21#_c_601_n N_A_1124_47#_c_814_n 0.0010876f $X=5.95 $Y=1.325
+ $X2=0 $Y2=0
cc_445 N_A_716_21#_c_601_n N_A_1124_47#_c_800_n 0.00393897f $X=5.95 $Y=1.325
+ $X2=0 $Y2=0
cc_446 N_A_716_21#_c_602_n N_A_1124_47#_c_800_n 0.0157324f $X=5.955 $Y=0.73
+ $X2=0 $Y2=0
cc_447 N_A_716_21#_M1002_g N_VPWR_c_845_n 0.00438629f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_448 N_A_716_21#_c_613_n N_VPWR_c_845_n 0.00707659f $X=4.3 $Y=1.7 $X2=0 $Y2=0
cc_449 N_A_716_21#_c_614_n N_VPWR_c_845_n 0.00377554f $X=3.885 $Y=1.7 $X2=0
+ $Y2=0
cc_450 N_A_716_21#_c_630_p N_VPWR_c_845_n 0.011437f $X=4.385 $Y=2.27 $X2=0 $Y2=0
cc_451 N_A_716_21#_M1008_g N_VPWR_c_846_n 0.0129712f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_452 N_A_716_21#_c_604_n N_VPWR_c_846_n 0.00826346f $X=5.055 $Y=1.16 $X2=0
+ $Y2=0
cc_453 N_A_716_21#_c_612_n N_VPWR_c_847_n 0.00537515f $X=5.952 $Y=1.77 $X2=0
+ $Y2=0
cc_454 N_A_716_21#_M1002_g N_VPWR_c_848_n 0.00525264f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_455 N_A_716_21#_c_630_p N_VPWR_c_852_n 0.0128916f $X=4.385 $Y=2.27 $X2=0
+ $Y2=0
cc_456 N_A_716_21#_M1008_g N_VPWR_c_853_n 0.0046653f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_457 N_A_716_21#_c_612_n N_VPWR_c_853_n 0.00541359f $X=5.952 $Y=1.77 $X2=0
+ $Y2=0
cc_458 N_A_716_21#_M1019_s N_VPWR_c_842_n 0.00238199f $X=4.26 $Y=1.485 $X2=0
+ $Y2=0
cc_459 N_A_716_21#_M1002_g N_VPWR_c_842_n 0.0100685f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_460 N_A_716_21#_M1008_g N_VPWR_c_842_n 0.00921786f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_461 N_A_716_21#_c_612_n N_VPWR_c_842_n 0.0110992f $X=5.952 $Y=1.77 $X2=0
+ $Y2=0
cc_462 N_A_716_21#_c_613_n N_VPWR_c_842_n 0.0129435f $X=4.3 $Y=1.7 $X2=0 $Y2=0
cc_463 N_A_716_21#_c_614_n N_VPWR_c_842_n 0.00269099f $X=3.885 $Y=1.7 $X2=0
+ $Y2=0
cc_464 N_A_716_21#_c_630_p N_VPWR_c_842_n 0.00926541f $X=4.385 $Y=2.27 $X2=0
+ $Y2=0
cc_465 N_A_716_21#_c_600_n Q 0.0047956f $X=5.875 $Y=1.16 $X2=0 $Y2=0
cc_466 N_A_716_21#_c_612_n Q 0.00304486f $X=5.952 $Y=1.77 $X2=0 $Y2=0
cc_467 N_A_716_21#_c_600_n N_Q_c_954_n 0.00550705f $X=5.875 $Y=1.16 $X2=0 $Y2=0
cc_468 N_A_716_21#_c_602_n N_Q_c_954_n 7.5837e-19 $X=5.955 $Y=0.73 $X2=0 $Y2=0
cc_469 N_A_716_21#_c_599_n N_Q_c_955_n 0.0076145f $X=5.015 $Y=0.995 $X2=0 $Y2=0
cc_470 N_A_716_21#_M1008_g N_Q_c_955_n 0.0106802f $X=5.015 $Y=1.985 $X2=0 $Y2=0
cc_471 N_A_716_21#_c_600_n N_Q_c_955_n 0.0215882f $X=5.875 $Y=1.16 $X2=0 $Y2=0
cc_472 N_A_716_21#_c_601_n N_Q_c_955_n 0.00109445f $X=5.95 $Y=1.325 $X2=0 $Y2=0
cc_473 N_A_716_21#_c_611_n N_Q_c_955_n 9.74328e-19 $X=5.952 $Y=1.62 $X2=0 $Y2=0
cc_474 N_A_716_21#_c_604_n N_Q_c_955_n 0.0249855f $X=5.055 $Y=1.16 $X2=0 $Y2=0
cc_475 N_A_716_21#_M1006_g N_VGND_c_995_n 0.00498076f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_476 N_A_716_21#_c_626_p N_VGND_c_995_n 0.0133418f $X=4.487 $Y=0.84 $X2=0
+ $Y2=0
cc_477 N_A_716_21#_c_599_n N_VGND_c_996_n 0.0142448f $X=5.015 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_716_21#_c_604_n N_VGND_c_996_n 0.0101778f $X=5.055 $Y=1.16 $X2=0
+ $Y2=0
cc_479 N_A_716_21#_c_602_n N_VGND_c_997_n 0.00420958f $X=5.955 $Y=0.73 $X2=0
+ $Y2=0
cc_480 N_A_716_21#_M1006_g N_VGND_c_1000_n 0.00585385f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_481 N_A_716_21#_c_626_p N_VGND_c_1001_n 0.00708699f $X=4.487 $Y=0.84 $X2=0
+ $Y2=0
cc_482 N_A_716_21#_c_599_n N_VGND_c_1002_n 0.0046653f $X=5.015 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_716_21#_c_602_n N_VGND_c_1002_n 0.00541359f $X=5.955 $Y=0.73 $X2=0
+ $Y2=0
cc_484 N_A_716_21#_M1020_s N_VGND_c_1004_n 0.00383951f $X=4.26 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_716_21#_M1006_g N_VGND_c_1004_n 0.0121908f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_A_716_21#_c_599_n N_VGND_c_1004_n 0.00934473f $X=5.015 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_A_716_21#_c_602_n N_VGND_c_1004_n 0.0110992f $X=5.955 $Y=0.73 $X2=0
+ $Y2=0
cc_488 N_A_716_21#_c_626_p N_VGND_c_1004_n 0.00884264f $X=4.487 $Y=0.84 $X2=0
+ $Y2=0
cc_489 N_A_560_47#_c_719_n N_VPWR_c_844_n 0.00493731f $X=3.36 $Y=2.19 $X2=0
+ $Y2=0
cc_490 N_A_560_47#_M1019_g N_VPWR_c_845_n 0.00248972f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_A_560_47#_M1019_g N_VPWR_c_846_n 0.00279634f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_492 N_A_560_47#_c_719_n N_VPWR_c_848_n 0.0179866f $X=3.36 $Y=2.19 $X2=0 $Y2=0
cc_493 N_A_560_47#_M1019_g N_VPWR_c_852_n 0.0054256f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A_560_47#_M1012_d N_VPWR_c_842_n 0.00661403f $X=2.83 $Y=2.065 $X2=0
+ $Y2=0
cc_495 N_A_560_47#_M1019_g N_VPWR_c_842_n 0.0109465f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_560_47#_c_719_n N_VPWR_c_842_n 0.0224794f $X=3.36 $Y=2.19 $X2=0 $Y2=0
cc_497 N_A_560_47#_c_719_n A_674_413# 0.00129169f $X=3.36 $Y=2.19 $X2=-0.19
+ $Y2=-0.24
cc_498 N_A_560_47#_c_722_n N_VGND_c_994_n 0.00237054f $X=3.355 $Y=0.45 $X2=0
+ $Y2=0
cc_499 N_A_560_47#_c_710_n N_VGND_c_995_n 0.00455513f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_500 N_A_560_47#_c_711_n N_VGND_c_995_n 0.00181231f $X=4.52 $Y=1.16 $X2=0
+ $Y2=0
cc_501 N_A_560_47#_c_714_n N_VGND_c_995_n 0.015157f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_502 N_A_560_47#_c_710_n N_VGND_c_996_n 0.00896856f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_503 N_A_560_47#_c_722_n N_VGND_c_1000_n 0.0250007f $X=3.355 $Y=0.45 $X2=0
+ $Y2=0
cc_504 N_A_560_47#_c_710_n N_VGND_c_1001_n 0.00403817f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_560_47#_M1016_d N_VGND_c_1004_n 0.00259228f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_506 N_A_560_47#_c_710_n N_VGND_c_1004_n 0.00739419f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_507 N_A_560_47#_c_722_n N_VGND_c_1004_n 0.0249534f $X=3.355 $Y=0.45 $X2=0
+ $Y2=0
cc_508 N_A_560_47#_c_722_n A_651_47# 0.00497444f $X=3.355 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_509 N_A_560_47#_c_713_n A_651_47# 0.00190728f $X=3.44 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_510 N_A_1124_47#_M1011_g N_VPWR_c_847_n 0.0132029f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_A_1124_47#_c_802_n N_VPWR_c_847_n 0.0454653f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_512 N_A_1124_47#_c_798_n N_VPWR_c_847_n 0.00970026f $X=6.37 $Y=1.16 $X2=0
+ $Y2=0
cc_513 N_A_1124_47#_c_799_n N_VPWR_c_847_n 0.00197978f $X=6.37 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_A_1124_47#_c_802_n N_VPWR_c_853_n 0.0153916f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_515 N_A_1124_47#_M1011_g N_VPWR_c_854_n 0.0046653f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_516 N_A_1124_47#_M1014_s N_VPWR_c_842_n 0.00352456f $X=5.62 $Y=1.845 $X2=0
+ $Y2=0
cc_517 N_A_1124_47#_M1011_g N_VPWR_c_842_n 0.00895857f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_518 N_A_1124_47#_c_802_n N_VPWR_c_842_n 0.00941829f $X=5.745 $Y=2.165 $X2=0
+ $Y2=0
cc_519 N_A_1124_47#_c_797_n N_Q_c_954_n 0.0255149f $X=5.745 $Y=0.51 $X2=0 $Y2=0
cc_520 N_A_1124_47#_c_797_n N_Q_c_955_n 0.0185881f $X=5.745 $Y=0.51 $X2=0 $Y2=0
cc_521 N_A_1124_47#_c_802_n N_Q_c_955_n 0.0870977f $X=5.745 $Y=2.165 $X2=0 $Y2=0
cc_522 N_A_1124_47#_c_814_n N_Q_c_955_n 0.024005f $X=5.785 $Y=1.16 $X2=0 $Y2=0
cc_523 N_A_1124_47#_c_798_n N_Q_N_c_980_n 0.0264222f $X=6.37 $Y=1.16 $X2=0 $Y2=0
cc_524 N_A_1124_47#_c_800_n N_Q_N_c_980_n 0.0203256f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_525 N_A_1124_47#_c_797_n N_VGND_c_997_n 0.0209216f $X=5.745 $Y=0.51 $X2=0
+ $Y2=0
cc_526 N_A_1124_47#_c_798_n N_VGND_c_997_n 0.0106046f $X=6.37 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_A_1124_47#_c_799_n N_VGND_c_997_n 0.00207666f $X=6.37 $Y=1.16 $X2=0
+ $Y2=0
cc_528 N_A_1124_47#_c_800_n N_VGND_c_997_n 0.00941229f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_529 N_A_1124_47#_c_797_n N_VGND_c_1002_n 0.0153916f $X=5.745 $Y=0.51 $X2=0
+ $Y2=0
cc_530 N_A_1124_47#_c_800_n N_VGND_c_1003_n 0.0046653f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_1124_47#_M1005_s N_VGND_c_1004_n 0.00352456f $X=5.62 $Y=0.235 $X2=0
+ $Y2=0
cc_532 N_A_1124_47#_c_797_n N_VGND_c_1004_n 0.0094183f $X=5.745 $Y=0.51 $X2=0
+ $Y2=0
cc_533 N_A_1124_47#_c_800_n N_VGND_c_1004_n 0.00895857f $X=6.37 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_842_n A_470_369# 0.00373974f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_535 N_VPWR_c_842_n A_674_413# 0.00193462f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_536 N_VPWR_c_842_n N_Q_M1008_d 0.00382897f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_537 N_VPWR_c_853_n Q 0.0237367f $X=6.09 $Y=2.72 $X2=0 $Y2=0
cc_538 N_VPWR_c_842_n Q 0.013017f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_c_842_n N_Q_N_M1011_d 0.00387172f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_540 N_VPWR_c_854_n Q_N 0.018001f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_541 N_VPWR_c_842_n Q_N 0.00993603f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_542 N_Q_c_954_n N_VGND_c_1002_n 0.0110946f $X=5.395 $Y=0.58 $X2=0 $Y2=0
cc_543 N_Q_M1017_d N_VGND_c_1004_n 0.00402409f $X=5.09 $Y=0.235 $X2=0 $Y2=0
cc_544 N_Q_c_954_n N_VGND_c_1004_n 0.0116259f $X=5.395 $Y=0.58 $X2=0 $Y2=0
cc_545 Q_N N_VGND_c_1003_n 0.0179443f $X=6.595 $Y=0.425 $X2=0 $Y2=0
cc_546 N_Q_N_M1015_d N_VGND_c_1004_n 0.00387172f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_547 Q_N N_VGND_c_1004_n 0.00992387f $X=6.595 $Y=0.425 $X2=0 $Y2=0
cc_548 N_VGND_c_1004_n A_465_47# 0.0113625f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_549 N_VGND_c_1004_n A_651_47# 0.00464458f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24

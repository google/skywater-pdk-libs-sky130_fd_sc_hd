* File: sky130_fd_sc_hd__mux2_4.pxi.spice
* Created: Tue Sep  1 19:14:30 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2_4%S N_S_M1017_g N_S_M1015_g N_S_c_87_n N_S_M1011_g
+ N_S_M1016_g N_S_c_88_n N_S_c_111_p N_S_c_167_p N_S_c_89_n N_S_c_90_n
+ N_S_c_91_n N_S_c_92_n S N_S_c_93_n N_S_c_94_n N_S_c_137_p
+ PM_SKY130_FD_SC_HD__MUX2_4%S
x_PM_SKY130_FD_SC_HD__MUX2_4%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1015_s
+ N_A_27_47#_M1000_g N_A_27_47#_M1005_g N_A_27_47#_c_184_n N_A_27_47#_c_191_n
+ N_A_27_47#_c_201_n N_A_27_47#_c_185_n N_A_27_47#_c_186_n N_A_27_47#_c_187_n
+ N_A_27_47#_c_194_n N_A_27_47#_c_188_n PM_SKY130_FD_SC_HD__MUX2_4%A_27_47#
x_PM_SKY130_FD_SC_HD__MUX2_4%A0 N_A0_c_238_n N_A0_M1007_g N_A0_M1004_g A0 A0
+ N_A0_c_240_n PM_SKY130_FD_SC_HD__MUX2_4%A0
x_PM_SKY130_FD_SC_HD__MUX2_4%A1 N_A1_M1002_g N_A1_M1001_g A1 N_A1_c_272_n
+ N_A1_c_273_n N_A1_c_274_n PM_SKY130_FD_SC_HD__MUX2_4%A1
x_PM_SKY130_FD_SC_HD__MUX2_4%A_396_47# N_A_396_47#_M1007_d N_A_396_47#_M1004_d
+ N_A_396_47#_c_306_n N_A_396_47#_M1008_g N_A_396_47#_M1003_g
+ N_A_396_47#_c_307_n N_A_396_47#_M1009_g N_A_396_47#_M1006_g
+ N_A_396_47#_c_308_n N_A_396_47#_M1012_g N_A_396_47#_M1010_g
+ N_A_396_47#_c_309_n N_A_396_47#_M1014_g N_A_396_47#_M1013_g
+ N_A_396_47#_c_324_n N_A_396_47#_c_318_n N_A_396_47#_c_332_n
+ N_A_396_47#_c_334_n N_A_396_47#_c_337_n N_A_396_47#_c_310_n
+ N_A_396_47#_c_311_n N_A_396_47#_c_384_p N_A_396_47#_c_312_n
+ N_A_396_47#_c_313_n PM_SKY130_FD_SC_HD__MUX2_4%A_396_47#
x_PM_SKY130_FD_SC_HD__MUX2_4%VPWR N_VPWR_M1015_d N_VPWR_M1016_d N_VPWR_M1006_s
+ N_VPWR_M1013_s N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n
+ N_VPWR_c_438_n VPWR N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_433_n
+ PM_SKY130_FD_SC_HD__MUX2_4%VPWR
x_PM_SKY130_FD_SC_HD__MUX2_4%A_204_297# N_A_204_297#_M1000_d
+ N_A_204_297#_M1001_d N_A_204_297#_c_510_n N_A_204_297#_c_511_n
+ PM_SKY130_FD_SC_HD__MUX2_4%A_204_297#
x_PM_SKY130_FD_SC_HD__MUX2_4%A_314_297# N_A_314_297#_M1004_s
+ N_A_314_297#_M1016_s N_A_314_297#_c_533_n N_A_314_297#_c_540_n
+ PM_SKY130_FD_SC_HD__MUX2_4%A_314_297#
x_PM_SKY130_FD_SC_HD__MUX2_4%X N_X_M1008_d N_X_M1012_d N_X_M1003_d N_X_M1010_d
+ N_X_c_601_p N_X_c_583_n N_X_c_559_n N_X_c_563_n N_X_c_565_n N_X_c_569_n
+ N_X_c_604_p N_X_c_587_n N_X_c_571_n N_X_c_573_n X X X N_X_c_555_n N_X_c_557_n
+ X X PM_SKY130_FD_SC_HD__MUX2_4%X
x_PM_SKY130_FD_SC_HD__MUX2_4%VGND N_VGND_M1017_d N_VGND_M1011_d N_VGND_M1009_s
+ N_VGND_M1014_s N_VGND_c_613_n N_VGND_c_614_n N_VGND_c_615_n N_VGND_c_616_n
+ N_VGND_c_617_n VGND N_VGND_c_618_n N_VGND_c_619_n N_VGND_c_620_n
+ N_VGND_c_621_n N_VGND_c_622_n N_VGND_c_623_n N_VGND_c_624_n N_VGND_c_625_n
+ PM_SKY130_FD_SC_HD__MUX2_4%VGND
cc_1 VNB N_S_c_87_n 0.019748f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=0.995
cc_2 VNB N_S_c_88_n 0.00205824f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.995
cc_3 VNB N_S_c_89_n 0.00242396f $X=-0.19 $Y=-0.24 $X2=2.765 $Y2=0.995
cc_4 VNB N_S_c_90_n 0.0230207f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_5 VNB N_S_c_91_n 0.00208902f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_6 VNB N_S_c_92_n 0.00216163f $X=-0.19 $Y=-0.24 $X2=2.85 $Y2=1.16
cc_7 VNB N_S_c_93_n 0.0197405f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_8 VNB N_S_c_94_n 0.0431691f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=1.16
cc_9 VNB N_A_27_47#_c_184_n 0.0288307f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=1.985
cc_10 VNB N_A_27_47#_c_185_n 4.78091e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_11 VNB N_A_27_47#_c_186_n 0.0244297f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_12 VNB N_A_27_47#_c_187_n 0.0127969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_188_n 0.0227662f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_14 VNB N_A0_c_238_n 0.022682f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_15 VNB A0 0.0054184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A0_c_240_n 0.0319948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A1_c_272_n 0.0220634f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=0.56
cc_18 VNB N_A1_c_273_n 0.00226885f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=0.56
cc_19 VNB N_A1_c_274_n 0.0200732f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=1.325
cc_20 VNB N_A_396_47#_c_306_n 0.0153255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_396_47#_c_307_n 0.0157706f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=1.985
cc_22 VNB N_A_396_47#_c_308_n 0.0157741f $X=-0.19 $Y=-0.24 $X2=2.765 $Y2=0.805
cc_23 VNB N_A_396_47#_c_309_n 0.0182854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_396_47#_c_310_n 0.00149244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_396_47#_c_311_n 3.46824e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_396_47#_c_312_n 0.00102135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_396_47#_c_313_n 0.0673175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_433_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_555_n 0.00760135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.0243437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_613_n 0.00280471f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=1.985
cc_32 VNB N_VGND_c_614_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=2.68 $Y2=0.72
cc_33 VNB N_VGND_c_615_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_34 VNB N_VGND_c_616_n 0.0102807f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_35 VNB N_VGND_c_617_n 0.0118704f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_36 VNB N_VGND_c_618_n 0.0152837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_619_n 0.0639701f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=1.16
cc_38 VNB N_VGND_c_620_n 0.0117278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_621_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_622_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_623_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_624_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_625_n 0.27659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VPB N_S_M1015_g 0.022619f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB N_S_M1016_g 0.0259973f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.985
cc_46 VPB N_S_c_90_n 0.00412822f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_47 VPB N_S_c_91_n 9.49139e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_48 VPB N_S_c_92_n 0.00203566f $X=-0.19 $Y=1.305 $X2=2.85 $Y2=1.16
cc_49 VPB N_S_c_94_n 0.0138692f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=1.16
cc_50 VPB N_A_27_47#_M1000_g 0.0239397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_184_n 0.00884863f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.985
cc_52 VPB N_A_27_47#_c_191_n 0.0304719f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.995
cc_53 VPB N_A_27_47#_c_185_n 0.00208145f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_54 VPB N_A_27_47#_c_186_n 0.00496299f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_55 VPB N_A_27_47#_c_194_n 0.00720662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A0_M1004_g 0.0227834f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_57 VPB A0 0.00621422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A0_c_240_n 0.0104496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A1_M1001_g 0.0268584f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_60 VPB N_A1_c_272_n 0.00432076f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=0.56
cc_61 VPB N_A1_c_273_n 0.00259849f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=0.56
cc_62 VPB N_A_396_47#_M1003_g 0.0176213f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=0.56
cc_63 VPB N_A_396_47#_M1006_g 0.0182683f $X=-0.19 $Y=1.305 $X2=2.68 $Y2=0.72
cc_64 VPB N_A_396_47#_M1010_g 0.0182735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_396_47#_M1013_g 0.0210031f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_66 VPB N_A_396_47#_c_318_n 0.00678936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_396_47#_c_311_n 0.00161135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_396_47#_c_313_n 0.0106066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_434_n 0.00262493f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.985
cc_70 VPB N_VPWR_c_435_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=2.68 $Y2=0.72
cc_71 VPB N_VPWR_c_436_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_72 VPB N_VPWR_c_437_n 0.0102077f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_73 VPB N_VPWR_c_438_n 0.0250335f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_74 VPB N_VPWR_c_439_n 0.0151047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_440_n 0.062391f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=1.16
cc_76 VPB N_VPWR_c_441_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_442_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_443_n 0.00459796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_444_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_445_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_433_n 0.0497334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_204_297#_c_510_n 0.01149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_204_297#_c_511_n 0.00658858f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=0.56
cc_84 VPB N_A_314_297#_c_533_n 0.00978395f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_X_c_557_n 0.00777576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB X 0.012588f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 N_S_M1015_g N_A_27_47#_M1000_g 0.0228985f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_88 N_S_M1015_g N_A_27_47#_c_184_n 0.00421983f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_89 N_S_c_88_n N_A_27_47#_c_184_n 0.00729016f $X=0.655 $Y=0.995 $X2=0 $Y2=0
cc_90 N_S_c_90_n N_A_27_47#_c_184_n 0.00753857f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_91 N_S_c_91_n N_A_27_47#_c_184_n 0.0246541f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_92 N_S_c_93_n N_A_27_47#_c_184_n 0.00756436f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_93 N_S_M1015_g N_A_27_47#_c_201_n 0.0168485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_94 N_S_c_90_n N_A_27_47#_c_201_n 0.00222911f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_95 N_S_c_91_n N_A_27_47#_c_201_n 0.0209111f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_96 N_S_M1015_g N_A_27_47#_c_185_n 6.24468e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_97 N_S_c_111_p N_A_27_47#_c_185_n 0.0101604f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_98 N_S_c_90_n N_A_27_47#_c_185_n 3.18713e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_99 N_S_c_91_n N_A_27_47#_c_185_n 0.0247586f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_100 N_S_c_111_p N_A_27_47#_c_186_n 0.00173923f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_101 N_S_c_90_n N_A_27_47#_c_186_n 0.020191f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_102 N_S_c_91_n N_A_27_47#_c_186_n 0.00198104f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_103 N_S_c_88_n N_A_27_47#_c_188_n 0.00416964f $X=0.655 $Y=0.995 $X2=0 $Y2=0
cc_104 N_S_c_111_p N_A_27_47#_c_188_n 0.0149247f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_105 N_S_c_93_n N_A_27_47#_c_188_n 0.0227395f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_106 N_S_c_111_p N_A0_c_238_n 0.0181794f $X=2.68 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_107 N_S_c_111_p A0 0.0193968f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_108 N_S_c_111_p N_A0_c_240_n 0.00351787f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_109 N_S_c_111_p N_A1_c_272_n 0.00174798f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_110 N_S_c_92_n N_A1_c_272_n 0.00283577f $X=2.85 $Y=1.16 $X2=0 $Y2=0
cc_111 N_S_c_94_n N_A1_c_272_n 0.0103875f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_112 N_S_c_111_p N_A1_c_273_n 0.0286526f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_113 N_S_c_92_n N_A1_c_273_n 0.0217291f $X=2.85 $Y=1.16 $X2=0 $Y2=0
cc_114 N_S_c_94_n N_A1_c_273_n 3.08871e-19 $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_115 N_S_c_111_p N_A1_c_274_n 0.0128194f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_116 N_S_c_89_n N_A1_c_274_n 0.00605028f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_117 N_S_c_111_p N_A_396_47#_M1007_d 0.00434603f $X=2.68 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_118 N_S_c_87_n N_A_396_47#_c_306_n 0.0130972f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_119 N_S_M1016_g N_A_396_47#_M1003_g 0.0220635f $X=3.37 $Y=1.985 $X2=0 $Y2=0
cc_120 N_S_c_87_n N_A_396_47#_c_324_n 0.00391863f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_121 N_S_c_111_p N_A_396_47#_c_324_n 0.0490692f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_122 N_S_c_94_n N_A_396_47#_c_324_n 0.00362358f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_123 N_S_c_137_p N_A_396_47#_c_324_n 0.00635313f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_124 N_S_M1016_g N_A_396_47#_c_318_n 0.018787f $X=3.37 $Y=1.985 $X2=0 $Y2=0
cc_125 N_S_c_92_n N_A_396_47#_c_318_n 0.0102322f $X=2.85 $Y=1.16 $X2=0 $Y2=0
cc_126 N_S_c_94_n N_A_396_47#_c_318_n 0.00923449f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_127 N_S_c_137_p N_A_396_47#_c_318_n 0.0267106f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_128 N_S_c_87_n N_A_396_47#_c_332_n 0.0072547f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_129 N_S_c_111_p N_A_396_47#_c_332_n 0.00135923f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_130 N_S_c_87_n N_A_396_47#_c_334_n 0.0142816f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_131 N_S_c_94_n N_A_396_47#_c_334_n 0.00130986f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_132 N_S_c_137_p N_A_396_47#_c_334_n 0.00979689f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_133 N_S_c_111_p N_A_396_47#_c_337_n 0.0115397f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_134 N_S_c_89_n N_A_396_47#_c_337_n 0.00135839f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_135 N_S_c_94_n N_A_396_47#_c_337_n 0.00392529f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_136 N_S_c_137_p N_A_396_47#_c_337_n 0.0137618f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_137 N_S_c_87_n N_A_396_47#_c_310_n 0.00426797f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_138 N_S_c_137_p N_A_396_47#_c_310_n 0.00630069f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_139 N_S_c_94_n N_A_396_47#_c_311_n 0.00645554f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_140 N_S_c_137_p N_A_396_47#_c_311_n 0.00630069f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_141 N_S_c_94_n N_A_396_47#_c_312_n 0.001309f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_142 N_S_c_137_p N_A_396_47#_c_312_n 0.0152104f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_143 N_S_c_94_n N_A_396_47#_c_313_n 0.050404f $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_144 N_S_c_137_p N_A_396_47#_c_313_n 3.06175e-19 $X=3.31 $Y=1.16 $X2=0 $Y2=0
cc_145 N_S_M1015_g N_VPWR_c_434_n 0.0128878f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_146 N_S_M1016_g N_VPWR_c_435_n 0.00863421f $X=3.37 $Y=1.985 $X2=0 $Y2=0
cc_147 N_S_M1015_g N_VPWR_c_439_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_148 N_S_M1016_g N_VPWR_c_440_n 0.0046653f $X=3.37 $Y=1.985 $X2=0 $Y2=0
cc_149 N_S_M1015_g N_VPWR_c_433_n 0.008846f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_150 N_S_M1016_g N_VPWR_c_433_n 0.00921786f $X=3.37 $Y=1.985 $X2=0 $Y2=0
cc_151 N_S_c_88_n N_VGND_M1017_d 9.53637e-19 $X=0.655 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_152 N_S_c_111_p N_VGND_M1017_d 0.00396736f $X=2.68 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_153 N_S_c_167_p N_VGND_M1017_d 0.0022983f $X=0.74 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_154 N_S_c_111_p N_VGND_c_613_n 0.00629984f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_155 N_S_c_167_p N_VGND_c_613_n 0.0111292f $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_156 N_S_c_90_n N_VGND_c_613_n 2.41877e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_157 N_S_c_91_n N_VGND_c_613_n 0.0012826f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_158 N_S_c_93_n N_VGND_c_613_n 0.0100153f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_159 N_S_c_87_n N_VGND_c_614_n 0.00970925f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_160 N_S_c_93_n N_VGND_c_618_n 0.0046653f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_161 N_S_c_87_n N_VGND_c_619_n 0.00341689f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_162 N_S_c_111_p N_VGND_c_619_n 0.0182828f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_163 N_S_c_87_n N_VGND_c_625_n 0.00540327f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_164 N_S_c_111_p N_VGND_c_625_n 0.0323092f $X=2.68 $Y=0.72 $X2=0 $Y2=0
cc_165 N_S_c_167_p N_VGND_c_625_n 8.07506e-19 $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_166 N_S_c_93_n N_VGND_c_625_n 0.00895857f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_167 N_S_c_111_p A_206_47# 0.0327043f $X=2.68 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_168 N_S_c_111_p A_490_47# 0.0139742f $X=2.68 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_169 N_S_c_89_n A_490_47# 0.00210306f $X=2.765 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_170 N_A_27_47#_M1000_g A0 0.00163071f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_201_n A0 0.00554875f $X=0.91 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_185_n A0 0.0202926f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_186_n A0 0.00247512f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_185_n N_A0_c_240_n 3.62599e-19 $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_186_n N_A0_c_240_n 0.00891269f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_201_n N_VPWR_M1015_d 0.00637844f $X=0.91 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_27_47#_M1000_g N_VPWR_c_434_n 0.00293578f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_201_n N_VPWR_c_434_n 0.0193336f $X=0.91 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_191_n N_VPWR_c_439_n 0.0176426f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1000_g N_VPWR_c_440_n 0.00542163f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1015_s N_VPWR_c_433_n 0.00382897f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1000_g N_VPWR_c_433_n 0.0109852f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_191_n N_VPWR_c_433_n 0.00974347f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_201_n N_A_204_297#_M1000_d 0.00426876f $X=0.91 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_185 N_A_27_47#_M1000_g N_A_204_297#_c_511_n 0.00614498f $X=0.945 $Y=1.985
+ $X2=0 $Y2=0
cc_186 N_A_27_47#_c_201_n N_A_204_297#_c_511_n 0.0016549f $X=0.91 $Y=1.58 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_186_n N_A_204_297#_c_511_n 0.00136468f $X=0.995 $Y=1.16
+ $X2=0 $Y2=0
cc_188 N_A_27_47#_c_188_n N_VGND_c_613_n 0.00423719f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_187_n N_VGND_c_618_n 0.0138219f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_188_n N_VGND_c_619_n 0.00425094f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1017_s N_VGND_c_625_n 0.00388984f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_187_n N_VGND_c_625_n 0.00948668f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_188_n N_VGND_c_625_n 0.00727912f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A0_M1004_g N_A1_M1001_g 0.037163f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_195 A0 N_A1_c_272_n 2.0566e-19 $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_196 N_A0_c_240_n N_A1_c_272_n 0.0186624f $X=1.905 $Y=1.16 $X2=0 $Y2=0
cc_197 A0 N_A1_c_273_n 0.0207423f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A0_c_240_n N_A1_c_273_n 0.00974287f $X=1.905 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A0_c_238_n N_A1_c_274_n 0.0233056f $X=1.905 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A0_c_238_n N_A_396_47#_c_324_n 0.00763795f $X=1.905 $Y=0.995 $X2=0
+ $Y2=0
cc_201 A0 N_A_396_47#_c_318_n 0.0013102f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A0_M1004_g N_VPWR_c_440_n 0.00362032f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A0_M1004_g N_VPWR_c_433_n 0.00679758f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A0_M1004_g N_A_204_297#_c_510_n 0.0118076f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_205 A0 N_A_204_297#_c_510_n 0.00158857f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_206 N_A0_M1004_g N_A_204_297#_c_511_n 0.00365238f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_207 A0 N_A_314_297#_M1004_s 0.00522984f $X=1.52 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_208 N_A0_M1004_g N_A_314_297#_c_533_n 0.0128949f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_209 A0 N_A_314_297#_c_533_n 0.0112202f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_210 N_A0_c_240_n N_A_314_297#_c_533_n 0.00210677f $X=1.905 $Y=1.16 $X2=0
+ $Y2=0
cc_211 N_A0_c_238_n N_VGND_c_619_n 0.00423128f $X=1.905 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A0_c_238_n N_VGND_c_625_n 0.00730383f $X=1.905 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A1_c_274_n N_A_396_47#_c_324_n 0.00999448f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A1_M1001_g N_A_396_47#_c_318_n 0.0114591f $X=2.375 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A1_c_272_n N_A_396_47#_c_318_n 0.00162184f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A1_c_273_n N_A_396_47#_c_318_n 0.0212577f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A1_c_274_n N_A_396_47#_c_332_n 0.00374734f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A1_c_274_n N_A_396_47#_c_337_n 5.79924e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A1_M1001_g N_VPWR_c_440_n 0.00362032f $X=2.375 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A1_M1001_g N_VPWR_c_433_n 0.00670766f $X=2.375 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A1_M1001_g N_A_204_297#_c_510_n 0.00800006f $X=2.375 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A1_M1001_g N_A_314_297#_c_533_n 0.0126849f $X=2.375 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A1_c_273_n N_A_314_297#_c_533_n 3.7176e-19 $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A1_M1001_g N_A_314_297#_c_540_n 0.0024733f $X=2.375 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A1_c_274_n N_VGND_c_619_n 0.00366111f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A1_c_274_n N_VGND_c_625_n 0.00676258f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_396_47#_c_318_n N_VPWR_M1016_d 0.00537906f $X=3.565 $Y=1.68 $X2=0
+ $Y2=0
cc_228 N_A_396_47#_c_311_n N_VPWR_M1016_d 0.00122758f $X=3.65 $Y=1.595 $X2=0
+ $Y2=0
cc_229 N_A_396_47#_M1003_g N_VPWR_c_435_n 0.00711767f $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_396_47#_M1006_g N_VPWR_c_435_n 5.08801e-19 $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_396_47#_c_318_n N_VPWR_c_435_n 0.0077152f $X=3.565 $Y=1.68 $X2=0
+ $Y2=0
cc_232 N_A_396_47#_M1003_g N_VPWR_c_436_n 6.0901e-19 $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_396_47#_M1006_g N_VPWR_c_436_n 0.0101939f $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_396_47#_M1010_g N_VPWR_c_436_n 0.0101939f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_396_47#_M1013_g N_VPWR_c_436_n 6.0901e-19 $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_396_47#_M1010_g N_VPWR_c_438_n 6.0901e-19 $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_396_47#_M1013_g N_VPWR_c_438_n 0.0112954f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_396_47#_M1003_g N_VPWR_c_441_n 0.0046653f $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A_396_47#_M1006_g N_VPWR_c_441_n 0.0046653f $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_396_47#_M1010_g N_VPWR_c_442_n 0.0046653f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_396_47#_M1013_g N_VPWR_c_442_n 0.0046653f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_396_47#_M1004_d N_VPWR_c_433_n 0.00258022f $X=1.98 $Y=1.485 $X2=0
+ $Y2=0
cc_243 N_A_396_47#_M1003_g N_VPWR_c_433_n 0.00789179f $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_A_396_47#_M1006_g N_VPWR_c_433_n 0.00789179f $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_A_396_47#_M1010_g N_VPWR_c_433_n 0.00789179f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_A_396_47#_M1013_g N_VPWR_c_433_n 0.00789179f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_396_47#_c_318_n N_A_204_297#_M1001_d 0.011224f $X=3.565 $Y=1.68 $X2=0
+ $Y2=0
cc_248 N_A_396_47#_M1004_d N_A_204_297#_c_510_n 0.00421632f $X=1.98 $Y=1.485
+ $X2=0 $Y2=0
cc_249 N_A_396_47#_c_318_n N_A_314_297#_M1016_s 0.00503149f $X=3.565 $Y=1.68
+ $X2=0 $Y2=0
cc_250 N_A_396_47#_M1004_d N_A_314_297#_c_533_n 0.00427371f $X=1.98 $Y=1.485
+ $X2=0 $Y2=0
cc_251 N_A_396_47#_c_318_n N_A_314_297#_c_533_n 0.0800729f $X=3.565 $Y=1.68
+ $X2=0 $Y2=0
cc_252 N_A_396_47#_c_307_n N_X_c_559_n 0.0115547f $X=4.21 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_396_47#_c_308_n N_X_c_559_n 0.0119869f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_396_47#_c_384_p N_X_c_559_n 0.026745f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_396_47#_c_313_n N_X_c_559_n 0.00207061f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_396_47#_c_384_p N_X_c_563_n 0.00881067f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_396_47#_c_313_n N_X_c_563_n 0.00216182f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_396_47#_M1006_g N_X_c_565_n 0.0144787f $X=4.21 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A_396_47#_M1010_g N_X_c_565_n 0.014911f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_396_47#_c_384_p N_X_c_565_n 0.0228036f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_396_47#_c_313_n N_X_c_565_n 0.00197867f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_396_47#_c_384_p N_X_c_569_n 0.00768518f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_396_47#_c_313_n N_X_c_569_n 0.00210139f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_396_47#_c_384_p N_X_c_571_n 0.00881067f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_396_47#_c_313_n N_X_c_571_n 0.00216182f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_396_47#_c_384_p N_X_c_573_n 0.00768518f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_396_47#_c_313_n N_X_c_573_n 0.00210139f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_396_47#_c_309_n X 0.0160156f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_396_47#_c_384_p X 0.00374684f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_396_47#_M1013_g X 0.0187409f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_396_47#_c_384_p X 0.0031876f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_396_47#_c_309_n X 0.029899f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_396_47#_c_384_p X 0.0137226f $X=4.865 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_396_47#_c_334_n N_VGND_M1011_d 0.00407149f $X=3.565 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_396_47#_c_310_n N_VGND_M1011_d 6.64472e-19 $X=3.65 $Y=1.075 $X2=0
+ $Y2=0
cc_276 N_A_396_47#_c_306_n N_VGND_c_614_n 0.00675799f $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_396_47#_c_307_n N_VGND_c_614_n 5.08801e-19 $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_396_47#_c_324_n N_VGND_c_614_n 0.0131487f $X=3.06 $Y=0.38 $X2=0 $Y2=0
cc_279 N_A_396_47#_c_334_n N_VGND_c_614_n 0.0147155f $X=3.565 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_396_47#_c_384_p N_VGND_c_614_n 2.21221e-19 $X=4.865 $Y=1.16 $X2=0
+ $Y2=0
cc_281 N_A_396_47#_c_306_n N_VGND_c_615_n 5.08801e-19 $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_396_47#_c_307_n N_VGND_c_615_n 0.00664421f $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_396_47#_c_308_n N_VGND_c_615_n 0.00664421f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_396_47#_c_309_n N_VGND_c_615_n 5.08801e-19 $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A_396_47#_c_308_n N_VGND_c_617_n 5.08801e-19 $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_396_47#_c_309_n N_VGND_c_617_n 0.00774571f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_396_47#_c_324_n N_VGND_c_619_n 0.0601177f $X=3.06 $Y=0.38 $X2=0 $Y2=0
cc_288 N_A_396_47#_c_334_n N_VGND_c_619_n 0.00252187f $X=3.565 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_396_47#_c_306_n N_VGND_c_620_n 0.0046653f $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_396_47#_c_307_n N_VGND_c_620_n 0.00339367f $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_396_47#_c_308_n N_VGND_c_621_n 0.00339367f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_396_47#_c_309_n N_VGND_c_621_n 0.00339367f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_396_47#_M1007_d N_VGND_c_625_n 0.00258215f $X=1.98 $Y=0.235 $X2=0
+ $Y2=0
cc_294 N_A_396_47#_c_306_n N_VGND_c_625_n 0.00789179f $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A_396_47#_c_307_n N_VGND_c_625_n 0.00394406f $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_396_47#_c_308_n N_VGND_c_625_n 0.00394406f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_396_47#_c_309_n N_VGND_c_625_n 0.00394406f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_396_47#_c_324_n N_VGND_c_625_n 0.0449378f $X=3.06 $Y=0.38 $X2=0 $Y2=0
cc_299 N_A_396_47#_c_334_n N_VGND_c_625_n 0.00610827f $X=3.565 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_396_47#_c_324_n A_490_47# 0.0214455f $X=3.06 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_301 N_A_396_47#_c_332_n A_490_47# 0.00574357f $X=3.145 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_302 N_A_396_47#_c_337_n A_490_47# 0.00383072f $X=3.23 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_303 N_VPWR_c_433_n N_A_204_297#_M1000_d 0.00226583f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_304 N_VPWR_c_433_n N_A_204_297#_M1001_d 0.00243107f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_440_n N_A_204_297#_c_510_n 0.0745259f $X=3.415 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_433_n N_A_204_297#_c_510_n 0.0511724f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_440_n N_A_204_297#_c_511_n 0.0194754f $X=3.415 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_433_n N_A_204_297#_c_511_n 0.0129525f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_433_n N_A_314_297#_M1004_s 0.00210988f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_310 N_VPWR_c_433_n N_A_314_297#_M1016_s 0.00395542f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_440_n N_A_314_297#_c_533_n 0.00578029f $X=3.415 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_433_n N_A_314_297#_c_533_n 0.0111513f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_440_n N_A_314_297#_c_540_n 0.0114f $X=3.415 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_433_n N_A_314_297#_c_540_n 0.00642843f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_433_n N_X_M1003_d 0.00562358f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_c_433_n N_X_M1010_d 0.00562358f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_317 N_VPWR_c_441_n N_X_c_583_n 0.0113958f $X=4.255 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_433_n N_X_c_583_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_M1006_s N_X_c_565_n 0.00363759f $X=4.285 $Y=1.485 $X2=0 $Y2=0
cc_320 N_VPWR_c_436_n N_X_c_565_n 0.0170259f $X=4.42 $Y=2 $X2=0 $Y2=0
cc_321 N_VPWR_c_442_n N_X_c_587_n 0.0113958f $X=5.095 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_c_433_n N_X_c_587_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_323 N_VPWR_M1013_s X 8.29358e-19 $X=5.125 $Y=1.485 $X2=0 $Y2=0
cc_324 N_VPWR_c_438_n X 0.00359494f $X=5.26 $Y=2 $X2=0 $Y2=0
cc_325 N_VPWR_M1013_s N_X_c_557_n 0.00278895f $X=5.125 $Y=1.485 $X2=0 $Y2=0
cc_326 N_VPWR_c_438_n N_X_c_557_n 0.0202891f $X=5.26 $Y=2 $X2=0 $Y2=0
cc_327 N_VPWR_M1013_s X 0.00141418f $X=5.125 $Y=1.485 $X2=0 $Y2=0
cc_328 N_A_204_297#_c_510_n N_A_314_297#_M1004_s 0.00489883f $X=2.605 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_329 N_A_204_297#_M1001_d N_A_314_297#_c_533_n 0.00618651f $X=2.45 $Y=1.485
+ $X2=0 $Y2=0
cc_330 N_A_204_297#_c_510_n N_A_314_297#_c_533_n 0.0682125f $X=2.605 $Y=2.36
+ $X2=0 $Y2=0
cc_331 N_A_204_297#_c_511_n N_A_314_297#_c_533_n 0.0137945f $X=1.175 $Y=2.02
+ $X2=0 $Y2=0
cc_332 N_A_204_297#_c_510_n N_A_314_297#_c_540_n 0.00919603f $X=2.605 $Y=2.36
+ $X2=0 $Y2=0
cc_333 N_X_c_559_n N_VGND_M1009_s 0.00337587f $X=4.755 $Y=0.72 $X2=0 $Y2=0
cc_334 X N_VGND_M1014_s 8.22501e-19 $X=5.2 $Y=0.765 $X2=0 $Y2=0
cc_335 N_X_c_555_n N_VGND_M1014_s 0.00272217f $X=5.315 $Y=0.805 $X2=0 $Y2=0
cc_336 X N_VGND_M1014_s 0.00125528f $X=5.285 $Y=0.85 $X2=0 $Y2=0
cc_337 N_X_c_559_n N_VGND_c_615_n 0.0159625f $X=4.755 $Y=0.72 $X2=0 $Y2=0
cc_338 X N_VGND_c_617_n 0.00337064f $X=5.2 $Y=0.765 $X2=0 $Y2=0
cc_339 N_X_c_555_n N_VGND_c_617_n 0.0190055f $X=5.315 $Y=0.805 $X2=0 $Y2=0
cc_340 N_X_c_601_p N_VGND_c_620_n 0.0112274f $X=4 $Y=0.42 $X2=0 $Y2=0
cc_341 N_X_c_559_n N_VGND_c_620_n 0.00244309f $X=4.755 $Y=0.72 $X2=0 $Y2=0
cc_342 N_X_c_559_n N_VGND_c_621_n 0.00244309f $X=4.755 $Y=0.72 $X2=0 $Y2=0
cc_343 N_X_c_604_p N_VGND_c_621_n 0.0112274f $X=4.84 $Y=0.42 $X2=0 $Y2=0
cc_344 X N_VGND_c_621_n 0.00244309f $X=5.2 $Y=0.765 $X2=0 $Y2=0
cc_345 N_X_M1008_d N_VGND_c_625_n 0.00405853f $X=3.865 $Y=0.235 $X2=0 $Y2=0
cc_346 N_X_M1012_d N_VGND_c_625_n 0.00249348f $X=4.705 $Y=0.235 $X2=0 $Y2=0
cc_347 N_X_c_601_p N_VGND_c_625_n 0.00643448f $X=4 $Y=0.42 $X2=0 $Y2=0
cc_348 N_X_c_559_n N_VGND_c_625_n 0.00984256f $X=4.755 $Y=0.72 $X2=0 $Y2=0
cc_349 N_X_c_604_p N_VGND_c_625_n 0.00643448f $X=4.84 $Y=0.42 $X2=0 $Y2=0
cc_350 X N_VGND_c_625_n 0.00465289f $X=5.2 $Y=0.765 $X2=0 $Y2=0
cc_351 N_X_c_555_n N_VGND_c_625_n 0.00132683f $X=5.315 $Y=0.805 $X2=0 $Y2=0
cc_352 N_VGND_c_625_n A_206_47# 0.00941645f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
cc_353 N_VGND_c_625_n A_490_47# 0.00719245f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__and4bb_4.spice
* Created: Thu Aug 27 14:09:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4bb_4.pex.spice"
.subckt sky130_fd_sc_hd__and4bb_4  VNB VPB B_N D C A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_B_N_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_174_21#_M1001_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11785 PD=0.92 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1001_d N_A_174_21#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_174_21#_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.3
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1019 N_X_M1007_d N_A_174_21#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75001.7
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1004 A_556_47# N_D_M1004_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.11375 PD=0.98 PS=1 NRD=20.304 NRS=10.152 M=1 R=4.33333 SA=75002.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1008 A_652_47# N_C_M1008_g A_556_47# VNB NSHORT L=0.15 W=0.65 AD=0.1365
+ AS=0.10725 PD=1.07 PS=0.98 NRD=28.608 NRS=20.304 M=1 R=4.33333 SA=75002.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1013 A_766_47# N_A_27_47#_M1013_g A_652_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.1365 PD=0.98 PS=1.07 NRD=20.304 NRS=28.608 M=1 R=4.33333
+ SA=75003.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1018 N_A_174_21#_M1018_d N_A_832_21#_M1018_g A_766_47# VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333
+ SA=75003.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_832_21#_M1014_d N_A_N_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1764 PD=1.36 PS=1.68 NRD=0 NRS=44.28 M=1 R=2.8 SA=75000.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_B_N_M1009_g N_A_27_47#_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75005.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1009_d N_A_174_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.198239 AS=0.135 PD=1.8662 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.4 SB=75004 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_174_21#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1002_d N_A_174_21#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A_174_21#_M1012_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.135 PD=1.35 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1016 N_A_174_21#_M1016_d N_D_M1016_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.175 PD=1.33 PS=1.35 NRD=10.8153 NRS=14.7553 M=1 R=6.66667
+ SA=75002.1 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g N_A_174_21#_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.165 PD=1.42 PS=1.33 NRD=18.715 NRS=0 M=1 R=6.66667 SA=75002.6
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1005 N_A_174_21#_M1005_d N_A_27_47#_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=1 AD=0.165 AS=0.21 PD=1.33 PS=1.42 NRD=2.9353 NRS=8.8453 M=1 R=6.66667
+ SA=75003.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_832_21#_M1015_g N_A_174_21#_M1005_d VPB PHIGHVT L=0.15
+ W=1 AD=0.438944 AS=0.165 PD=2.99296 PS=1.33 NRD=14.7553 NRS=6.8753 M=1
+ R=6.66667 SA=75003.7 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1006 N_A_832_21#_M1006_d N_A_N_M1006_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.184356 PD=1.36 PS=1.25704 NRD=0 NRS=42.1974 M=1 R=2.8
+ SA=75005.2 SB=75000.2 A=0.063 P=1.14 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__and4bb_4.pxi.spice"
*
.ends
*
*

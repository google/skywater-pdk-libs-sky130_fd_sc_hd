* File: sky130_fd_sc_hd__and3_4.spice
* Created: Thu Aug 27 14:07:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and3_4.pex.spice"
.subckt sky130_fd_sc_hd__and3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 A_185_47# N_A_M1006_g N_A_94_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128375 AS=0.19825 PD=1.045 PS=1.91 NRD=26.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003 A=0.0975 P=1.6 MULT=1
MM1005 A_294_47# N_B_M1005_g A_185_47# VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.128375 PD=0.86 PS=1.045 NRD=9.228 NRS=26.304 M=1 R=4.33333 SA=75000.8
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g A_294_47# VNB NSHORT L=0.15 W=0.65 AD=0.138125
+ AS=0.06825 PD=1.075 PS=0.86 NRD=18.456 NRS=9.228 M=1 R=4.33333 SA=75001.1
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1000 N_X_M1000_d N_A_94_47#_M1000_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.138125 PD=0.93 PS=1.075 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1000_d N_A_94_47#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1010_d N_A_94_47#_M1010_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1010_d N_A_94_47#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.18525 PD=0.93 PS=1.87 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_94_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1975 AS=0.305 PD=1.395 PS=2.61 NRD=12.7853 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003 A=0.15 P=2.3 MULT=1
MM1009 N_A_94_47#_M1009_d N_B_M1009_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1975 PD=1.28 PS=1.395 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75000.8
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_C_M1013_g N_A_94_47#_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1775 AS=0.14 PD=1.355 PS=1.28 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_94_47#_M1001_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1775 PD=1.28 PS=1.355 NRD=0 NRS=7.8603 M=1 R=6.66667 SA=75001.7
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1001_d N_A_94_47#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.1
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1008_d N_A_94_47#_M1008_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_X_M1008_d N_A_94_47#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75003 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__and3_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__fa_4.spice.SKY130_FD_SC_HD__FA_4.pxi
* Created: Thu Aug 27 14:21:17 2020
* 
x_PM_SKY130_FD_SC_HD__FA_4%A_79_21# N_A_79_21#_M1010_d N_A_79_21#_M1006_d
+ N_A_79_21#_c_212_n N_A_79_21#_M1020_g N_A_79_21#_M1005_g N_A_79_21#_c_213_n
+ N_A_79_21#_M1028_g N_A_79_21#_M1011_g N_A_79_21#_c_214_n N_A_79_21#_M1029_g
+ N_A_79_21#_M1031_g N_A_79_21#_c_215_n N_A_79_21#_M1036_g N_A_79_21#_M1035_g
+ N_A_79_21#_M1017_g N_A_79_21#_M1016_g N_A_79_21#_c_380_p N_A_79_21#_c_218_n
+ N_A_79_21#_c_219_n N_A_79_21#_c_220_n N_A_79_21#_c_390_p N_A_79_21#_c_235_n
+ N_A_79_21#_c_236_n N_A_79_21#_c_254_p N_A_79_21#_c_248_p N_A_79_21#_c_221_n
+ N_A_79_21#_c_222_n N_A_79_21#_c_223_n N_A_79_21#_c_224_n N_A_79_21#_c_225_n
+ N_A_79_21#_c_226_n N_A_79_21#_c_227_n N_A_79_21#_c_228_n
+ PM_SKY130_FD_SC_HD__FA_4%A_79_21#
x_PM_SKY130_FD_SC_HD__FA_4%A N_A_c_468_n N_A_M1034_g N_A_M1024_g N_A_M1018_g
+ N_A_M1019_g N_A_M1039_g N_A_M1004_g N_A_M1003_g N_A_M1026_g N_A_c_474_n A
+ N_A_c_476_n N_A_c_477_n N_A_c_478_n N_A_c_479_n N_A_c_480_n N_A_c_481_n
+ N_A_c_482_n N_A_c_483_n N_A_c_484_n N_A_c_485_n N_A_c_486_n N_A_c_487_n
+ N_A_c_488_n PM_SKY130_FD_SC_HD__FA_4%A
x_PM_SKY130_FD_SC_HD__FA_4%B N_B_M1006_g N_B_M1010_g N_B_c_737_n N_B_M1014_g
+ N_B_c_746_n N_B_M1038_g N_B_c_738_n N_B_c_739_n N_B_c_747_n N_B_c_748_n
+ N_B_c_740_n N_B_M1000_g N_B_M1023_g N_B_M1030_g N_B_M1007_g N_B_c_742_n B
+ N_B_c_752_n N_B_c_753_n N_B_c_754_n N_B_c_821_n N_B_c_755_n N_B_c_756_n
+ N_B_c_757_n N_B_c_758_n N_B_c_759_n N_B_c_743_n N_B_c_761_n N_B_c_762_n
+ PM_SKY130_FD_SC_HD__FA_4%B
x_PM_SKY130_FD_SC_HD__FA_4%CIN N_CIN_M1021_g N_CIN_M1032_g N_CIN_M1001_g
+ N_CIN_M1013_g N_CIN_M1009_g N_CIN_M1037_g N_CIN_c_969_n N_CIN_c_970_n
+ N_CIN_c_971_n N_CIN_c_984_n N_CIN_c_985_n N_CIN_c_972_n N_CIN_c_973_n
+ N_CIN_c_974_n N_CIN_c_975_n N_CIN_c_988_n N_CIN_c_976_n N_CIN_c_977_n
+ N_CIN_c_990_n N_CIN_c_991_n CIN N_CIN_c_978_n N_CIN_c_993_n N_CIN_c_994_n
+ PM_SKY130_FD_SC_HD__FA_4%CIN
x_PM_SKY130_FD_SC_HD__FA_4%A_1271_47# N_A_1271_47#_M1017_d N_A_1271_47#_M1016_d
+ N_A_1271_47#_c_1195_n N_A_1271_47#_M1015_g N_A_1271_47#_M1002_g
+ N_A_1271_47#_M1008_g N_A_1271_47#_c_1196_n N_A_1271_47#_M1022_g
+ N_A_1271_47#_c_1197_n N_A_1271_47#_M1027_g N_A_1271_47#_M1012_g
+ N_A_1271_47#_c_1198_n N_A_1271_47#_M1033_g N_A_1271_47#_M1025_g
+ N_A_1271_47#_c_1246_n N_A_1271_47#_c_1212_n N_A_1271_47#_c_1225_n
+ N_A_1271_47#_c_1199_n N_A_1271_47#_c_1200_n N_A_1271_47#_c_1230_n
+ N_A_1271_47#_c_1233_n N_A_1271_47#_c_1201_n N_A_1271_47#_c_1202_n
+ N_A_1271_47#_c_1300_p N_A_1271_47#_c_1216_n N_A_1271_47#_c_1257_n
+ N_A_1271_47#_c_1210_n N_A_1271_47#_c_1203_n N_A_1271_47#_c_1204_n
+ PM_SKY130_FD_SC_HD__FA_4%A_1271_47#
x_PM_SKY130_FD_SC_HD__FA_4%VPWR N_VPWR_M1005_s N_VPWR_M1011_s N_VPWR_M1035_s
+ N_VPWR_M1019_d N_VPWR_M1023_s N_VPWR_M1013_d N_VPWR_M1026_d N_VPWR_M1008_d
+ N_VPWR_M1025_d N_VPWR_c_1374_n N_VPWR_c_1375_n N_VPWR_c_1376_n N_VPWR_c_1377_n
+ N_VPWR_c_1378_n N_VPWR_c_1379_n N_VPWR_c_1380_n N_VPWR_c_1381_n
+ N_VPWR_c_1382_n N_VPWR_c_1383_n N_VPWR_c_1384_n N_VPWR_c_1385_n
+ N_VPWR_c_1386_n N_VPWR_c_1387_n VPWR VPWR N_VPWR_c_1389_n N_VPWR_c_1390_n
+ N_VPWR_c_1391_n N_VPWR_c_1392_n N_VPWR_c_1393_n N_VPWR_c_1394_n
+ N_VPWR_c_1373_n N_VPWR_c_1396_n N_VPWR_c_1397_n N_VPWR_c_1398_n
+ N_VPWR_c_1399_n N_VPWR_c_1400_n N_VPWR_c_1401_n PM_SKY130_FD_SC_HD__FA_4%VPWR
x_PM_SKY130_FD_SC_HD__FA_4%COUT N_COUT_M1020_s N_COUT_M1029_s N_COUT_M1005_d
+ N_COUT_M1031_d N_COUT_c_1538_n N_COUT_c_1550_n N_COUT_c_1539_n N_COUT_c_1540_n
+ N_COUT_c_1542_n N_COUT_c_1543_n N_COUT_c_1574_n N_COUT_c_1595_n
+ N_COUT_c_1578_n N_COUT_c_1582_n N_COUT_c_1585_n COUT N_COUT_c_1586_n
+ PM_SKY130_FD_SC_HD__FA_4%COUT
x_PM_SKY130_FD_SC_HD__FA_4%A_658_369# N_A_658_369#_M1032_d N_A_658_369#_M1038_d
+ N_A_658_369#_c_1629_n N_A_658_369#_c_1617_n N_A_658_369#_c_1623_n
+ N_A_658_369#_c_1618_n PM_SKY130_FD_SC_HD__FA_4%A_658_369#
x_PM_SKY130_FD_SC_HD__FA_4%A_1014_369# N_A_1014_369#_M1023_d
+ N_A_1014_369#_M1004_d N_A_1014_369#_c_1651_n N_A_1014_369#_c_1640_n
+ N_A_1014_369#_c_1643_n N_A_1014_369#_c_1658_n
+ PM_SKY130_FD_SC_HD__FA_4%A_1014_369#
x_PM_SKY130_FD_SC_HD__FA_4%SUM N_SUM_M1015_s N_SUM_M1027_s N_SUM_M1002_s
+ N_SUM_M1012_s N_SUM_c_1666_n N_SUM_c_1671_n N_SUM_c_1672_n N_SUM_c_1667_n
+ N_SUM_c_1696_n N_SUM_c_1699_n N_SUM_c_1668_n N_SUM_c_1673_n N_SUM_c_1704_n
+ N_SUM_c_1708_n N_SUM_c_1711_n N_SUM_c_1669_n N_SUM_c_1674_n SUM
+ PM_SKY130_FD_SC_HD__FA_4%SUM
x_PM_SKY130_FD_SC_HD__FA_4%VGND N_VGND_M1020_d N_VGND_M1028_d N_VGND_M1036_d
+ N_VGND_M1018_d N_VGND_M1000_s N_VGND_M1001_d N_VGND_M1003_d N_VGND_M1022_d
+ N_VGND_M1033_d N_VGND_c_1752_n N_VGND_c_1753_n N_VGND_c_1754_n N_VGND_c_1755_n
+ N_VGND_c_1756_n N_VGND_c_1757_n N_VGND_c_1758_n N_VGND_c_1759_n
+ N_VGND_c_1760_n N_VGND_c_1761_n N_VGND_c_1762_n N_VGND_c_1763_n
+ N_VGND_c_1764_n N_VGND_c_1765_n N_VGND_c_1766_n N_VGND_c_1767_n VGND VGND
+ N_VGND_c_1769_n N_VGND_c_1770_n N_VGND_c_1771_n N_VGND_c_1772_n
+ N_VGND_c_1773_n N_VGND_c_1774_n N_VGND_c_1775_n N_VGND_c_1776_n
+ N_VGND_c_1777_n N_VGND_c_1778_n N_VGND_c_1779_n PM_SKY130_FD_SC_HD__FA_4%VGND
x_PM_SKY130_FD_SC_HD__FA_4%A_658_47# N_A_658_47#_M1021_d N_A_658_47#_M1014_d
+ N_A_658_47#_c_1962_n N_A_658_47#_c_1937_n N_A_658_47#_c_1938_n
+ N_A_658_47#_c_1954_n PM_SKY130_FD_SC_HD__FA_4%A_658_47#
x_PM_SKY130_FD_SC_HD__FA_4%A_1014_47# N_A_1014_47#_M1000_d N_A_1014_47#_M1039_d
+ N_A_1014_47#_c_1995_n N_A_1014_47#_c_1972_n N_A_1014_47#_c_1973_n
+ N_A_1014_47#_c_1992_n PM_SKY130_FD_SC_HD__FA_4%A_1014_47#
cc_1 VNB N_A_79_21#_c_212_n 0.0198049f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_213_n 0.0157804f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_214_n 0.0157921f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_215_n 0.0163085f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_M1017_g 0.0230444f $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=0.445
cc_6 VNB N_A_79_21#_M1016_g 0.00523751f $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=2.165
cc_7 VNB N_A_79_21#_c_218_n 0.00157651f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.075
cc_8 VNB N_A_79_21#_c_219_n 3.20669e-19 $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.43
cc_9 VNB N_A_79_21#_c_220_n 0.00279192f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.74
cc_10 VNB N_A_79_21#_c_221_n 9.44169e-19 $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.16
cc_11 VNB N_A_79_21#_c_222_n 0.0123286f $X=-0.19 $Y=-0.24 $X2=6.55 $Y2=0.85
cc_12 VNB N_A_79_21#_c_223_n 0.00402697f $X=-0.19 $Y=-0.24 $X2=3.14 $Y2=0.85
cc_13 VNB N_A_79_21#_c_224_n 0.00994223f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=0.85
cc_14 VNB N_A_79_21#_c_225_n 0.00132437f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=0.85
cc_15 VNB N_A_79_21#_c_226_n 0.0651633f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_16 VNB N_A_79_21#_c_227_n 0.0252305f $X=-0.19 $Y=-0.24 $X2=6.34 $Y2=1.04
cc_17 VNB N_A_79_21#_c_228_n 0.00649189f $X=-0.19 $Y=-0.24 $X2=6.34 $Y2=1.04
cc_18 VNB N_A_c_468_n 0.022157f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=0.235
cc_19 VNB N_A_M1024_g 0.0288159f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A_M1018_g 0.0299029f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_21 VNB N_A_M1039_g 0.0198556f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_22 VNB N_A_M1004_g 0.00424732f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_23 VNB N_A_M1003_g 0.0294745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_c_474_n 4.23616e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB A 0.00481396f $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=1.205
cc_26 VNB N_A_c_476_n 0.00432352f $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=2.165
cc_27 VNB N_A_c_477_n 2.01406e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_c_478_n 0.00614383f $X=-0.19 $Y=-0.24 $X2=1.74 $Y2=1.16
cc_29 VNB N_A_c_479_n 8.64789e-19 $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_30 VNB N_A_c_480_n 0.00558474f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_31 VNB N_A_c_481_n 0.00124236f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_32 VNB N_A_c_482_n 0.00253456f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.245
cc_33 VNB N_A_c_483_n 0.00170256f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.58
cc_34 VNB N_A_c_484_n 0.0224949f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.16
cc_35 VNB N_A_c_485_n 0.0244928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_c_486_n 0.00666652f $X=-0.19 $Y=-0.24 $X2=6.55 $Y2=0.85
cc_37 VNB N_A_c_487_n 0.0209216f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=0.85
cc_38 VNB N_A_c_488_n 0.012294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_B_M1010_g 0.0444388f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_40 VNB N_B_c_737_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_41 VNB N_B_c_738_n 0.0530718f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_42 VNB N_B_c_739_n 0.00947258f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_43 VNB N_B_c_740_n 0.0171497f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_44 VNB N_B_M1030_g 0.0415238f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_45 VNB N_B_c_742_n 0.00469281f $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=0.875
cc_46 VNB N_B_c_743_n 0.0213523f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=1.995
cc_47 VNB N_CIN_M1021_g 0.0299955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_CIN_M1037_g 0.0416782f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_49 VNB N_CIN_c_969_n 0.0134432f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_50 VNB N_CIN_c_970_n 0.00664345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_CIN_c_971_n 3.21027e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_52 VNB N_CIN_c_972_n 0.00215826f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_53 VNB N_CIN_c_973_n 0.0152367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_CIN_c_974_n 0.00451859f $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=0.875
cc_55 VNB N_CIN_c_975_n 5.41591e-19 $X=-0.19 $Y=-0.24 $X2=6.28 $Y2=0.445
cc_56 VNB N_CIN_c_976_n 0.020086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_CIN_c_977_n 0.00304308f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_58 VNB N_CIN_c_978_n 0.0187439f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=0.74
cc_59 VNB N_A_1271_47#_c_1195_n 0.0173318f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_60 VNB N_A_1271_47#_c_1196_n 0.0165379f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_61 VNB N_A_1271_47#_c_1197_n 0.0157973f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_62 VNB N_A_1271_47#_c_1198_n 0.019164f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_63 VNB N_A_1271_47#_c_1199_n 0.00364909f $X=-0.19 $Y=-0.24 $X2=1.74 $Y2=1.16
cc_64 VNB N_A_1271_47#_c_1200_n 0.0033791f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_65 VNB N_A_1271_47#_c_1201_n 0.001669f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.16
cc_66 VNB N_A_1271_47#_c_1202_n 4.74296e-19 $X=-0.19 $Y=-0.24 $X2=1.825
+ $Y2=1.075
cc_67 VNB N_A_1271_47#_c_1203_n 0.00105672f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=0.85
cc_68 VNB N_A_1271_47#_c_1204_n 0.0693337f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_69 VNB N_VPWR_c_1373_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_COUT_c_1538_n 0.017806f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_71 VNB N_COUT_c_1539_n 0.00343673f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_72 VNB N_COUT_c_1540_n 0.0112067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_SUM_c_1666_n 0.00175519f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_74 VNB N_SUM_c_1667_n 0.00217862f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_75 VNB N_SUM_c_1668_n 0.0110037f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_76 VNB N_SUM_c_1669_n 0.0022746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB SUM 0.0224348f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=0.825
cc_78 VNB N_VGND_c_1752_n 0.00360014f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_79 VNB N_VGND_c_1753_n 0.0022431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1754_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1755_n 0.0049662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1756_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_83 VNB N_VGND_c_1757_n 0.00281836f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.16
cc_84 VNB N_VGND_c_1758_n 0.00410953f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.43
cc_85 VNB N_VGND_c_1759_n 0.00416643f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.58
cc_86 VNB N_VGND_c_1760_n 0.0167116f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=1.995
cc_87 VNB N_VGND_c_1761_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=2.31 $Y2=1.995
cc_88 VNB N_VGND_c_1762_n 0.0456861f $X=-0.19 $Y=-0.24 $X2=1.842 $Y2=1.58
cc_89 VNB N_VGND_c_1763_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1764_n 0.0202688f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.995
cc_91 VNB N_VGND_c_1765_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1766_n 0.0170047f $X=-0.19 $Y=-0.24 $X2=3.14 $Y2=0.85
cc_93 VNB N_VGND_c_1767_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=0.85
cc_94 VNB VGND 0.0106949f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=0.85
cc_95 VNB N_VGND_c_1769_n 0.0173944f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.16
cc_96 VNB N_VGND_c_1770_n 0.0353132f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_97 VNB N_VGND_c_1771_n 0.0159136f $X=-0.19 $Y=-0.24 $X2=3.005 $Y2=0.595
cc_98 VNB N_VGND_c_1772_n 0.0116974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1773_n 0.0106277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1774_n 0.469755f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1775_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1776_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1777_n 0.00507318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1778_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1779_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_A_658_47#_c_1937_n 0.00310751f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_107 VNB N_A_658_47#_c_1938_n 0.00259269f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_108 VNB N_A_1014_47#_c_1972_n 0.00540238f $X=-0.19 $Y=-0.24 $X2=0.47
+ $Y2=1.985
cc_109 VNB N_A_1014_47#_c_1973_n 0.00218811f $X=-0.19 $Y=-0.24 $X2=0.47
+ $Y2=1.985
cc_110 VPB N_A_79_21#_M1005_g 0.022676f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_111 VPB N_A_79_21#_M1011_g 0.0178626f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_112 VPB N_A_79_21#_M1031_g 0.0178784f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_113 VPB N_A_79_21#_M1035_g 0.0184713f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_114 VPB N_A_79_21#_M1016_g 0.0378103f $X=-0.19 $Y=1.305 $X2=6.28 $Y2=2.165
cc_115 VPB N_A_79_21#_c_219_n 0.00216187f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.43
cc_116 VPB N_A_79_21#_c_235_n 0.00292419f $X=-0.19 $Y=1.305 $X2=2.14 $Y2=1.58
cc_117 VPB N_A_79_21#_c_236_n 0.00184251f $X=-0.19 $Y=1.305 $X2=2.225 $Y2=1.91
cc_118 VPB N_A_79_21#_c_226_n 0.010057f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_119 VPB N_A_c_468_n 0.00414423f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=0.235
cc_120 VPB N_A_M1034_g 0.0367825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_M1019_g 0.0369395f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_122 VPB N_A_M1004_g 0.0364185f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_123 VPB N_A_M1026_g 0.0396698f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_124 VPB N_A_c_474_n 7.8182e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_c_477_n 0.00213469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_c_479_n 2.32744e-19 $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.16
cc_127 VPB N_A_c_481_n 5.14832e-19 $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.16
cc_128 VPB N_A_c_482_n 0.00178219f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.245
cc_129 VPB N_A_c_483_n 7.64837e-19 $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.58
cc_130 VPB N_A_c_484_n 0.00700974f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.16
cc_131 VPB N_A_c_487_n 0.00485547f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=0.85
cc_132 VPB N_B_M1006_g 0.0208944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_B_M1010_g 0.00337255f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_134 VPB N_B_c_746_n 0.0190907f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_135 VPB N_B_c_747_n 0.0399721f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_136 VPB N_B_c_748_n 0.00881125f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_137 VPB N_B_M1030_g 0.00322479f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_138 VPB N_B_M1007_g 0.0205486f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_139 VPB B 0.00966646f $X=-0.19 $Y=1.305 $X2=6.28 $Y2=0.445
cc_140 VPB N_B_c_752_n 0.00733903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_B_c_753_n 0.00220153f $X=-0.19 $Y=1.305 $X2=6.28 $Y2=1.205
cc_142 VPB N_B_c_754_n 0.0105272f $X=-0.19 $Y=1.305 $X2=6.28 $Y2=2.165
cc_143 VPB N_B_c_755_n 0.00168228f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.16
cc_144 VPB N_B_c_756_n 0.00813082f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=0.825
cc_145 VPB N_B_c_757_n 0.0255568f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.43
cc_146 VPB N_B_c_758_n 0.0389846f $X=-0.19 $Y=1.305 $X2=2.225 $Y2=1.665
cc_147 VPB N_B_c_759_n 0.00182223f $X=-0.19 $Y=1.305 $X2=2.225 $Y2=1.91
cc_148 VPB N_B_c_743_n 0.00173871f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=1.995
cc_149 VPB N_B_c_761_n 0.0184685f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.16
cc_150 VPB N_B_c_762_n 0.0243326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_CIN_M1032_g 0.0358736f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_152 VPB N_CIN_M1013_g 0.0188895f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_153 VPB N_CIN_M1009_g 0.0179457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_CIN_M1037_g 0.00271333f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_155 VPB N_CIN_c_971_n 0.00267764f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_156 VPB N_CIN_c_984_n 0.00934831f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_157 VPB N_CIN_c_985_n 0.00271596f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_158 VPB N_CIN_c_972_n 0.0069689f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_159 VPB N_CIN_c_975_n 0.00124245f $X=-0.19 $Y=1.305 $X2=6.28 $Y2=0.445
cc_160 VPB N_CIN_c_988_n 0.0171474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_CIN_c_976_n 0.00657573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_CIN_c_990_n 0.0233104f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.16
cc_163 VPB N_CIN_c_991_n 0.00366471f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=0.825
cc_164 VPB N_CIN_c_978_n 0.00233543f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=0.74
cc_165 VPB N_CIN_c_993_n 0.0253827f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.58
cc_166 VPB N_CIN_c_994_n 0.00644752f $X=-0.19 $Y=1.305 $X2=2.225 $Y2=1.665
cc_167 VPB N_A_1271_47#_M1002_g 0.0182277f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_168 VPB N_A_1271_47#_M1008_g 0.0187642f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_169 VPB N_A_1271_47#_M1012_g 0.0187844f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_170 VPB N_A_1271_47#_M1025_g 0.022035f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_171 VPB N_A_1271_47#_c_1202_n 0.00157521f $X=-0.19 $Y=1.305 $X2=1.825
+ $Y2=1.075
cc_172 VPB N_A_1271_47#_c_1210_n 0.00203197f $X=-0.19 $Y=1.305 $X2=2.995
+ $Y2=0.85
cc_173 VPB N_A_1271_47#_c_1204_n 0.0124904f $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.16
cc_174 VPB N_VPWR_c_1374_n 0.00359124f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_175 VPB N_VPWR_c_1375_n 0.00231272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1376_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1377_n 0.00765493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1378_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.16
cc_179 VPB N_VPWR_c_1379_n 0.0027527f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.16
cc_180 VPB N_VPWR_c_1380_n 0.00412306f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.43
cc_181 VPB N_VPWR_c_1381_n 0.00469317f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.58
cc_182 VPB N_VPWR_c_1382_n 0.0182896f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=1.995
cc_183 VPB N_VPWR_c_1383_n 0.00324402f $X=-0.19 $Y=1.305 $X2=2.31 $Y2=1.995
cc_184 VPB N_VPWR_c_1384_n 0.0159536f $X=-0.19 $Y=1.305 $X2=1.842 $Y2=1.58
cc_185 VPB N_VPWR_c_1385_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1386_n 0.0209492f $X=-0.19 $Y=1.305 $X2=2.94 $Y2=1.995
cc_187 VPB N_VPWR_c_1387_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB VPWR 0.0110272f $X=-0.19 $Y=1.305 $X2=6.55 $Y2=0.85
cc_189 VPB N_VPWR_c_1389_n 0.0180274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1390_n 0.0375067f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_191 VPB N_VPWR_c_1391_n 0.0153149f $X=-0.19 $Y=1.305 $X2=6.34 $Y2=1.04
cc_192 VPB N_VPWR_c_1392_n 0.0116974f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=0.595
cc_193 VPB N_VPWR_c_1393_n 0.0484432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1394_n 0.0113717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1373_n 0.0595624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1396_n 0.0051592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1397_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1398_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1399_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1400_n 0.00510002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1401_n 0.00416791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_COUT_c_1538_n 0.00553627f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_203 VPB N_COUT_c_1542_n 0.00400074f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_204 VPB N_COUT_c_1543_n 0.0123158f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_205 VPB N_A_658_369#_c_1617_n 0.00158421f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.325
cc_206 VPB N_A_658_369#_c_1618_n 0.0032459f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_207 VPB N_SUM_c_1671_n 0.00264533f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_208 VPB N_SUM_c_1672_n 0.00156186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_SUM_c_1673_n 0.0144284f $X=-0.19 $Y=1.305 $X2=6.28 $Y2=0.875
cc_210 VPB N_SUM_c_1674_n 0.00227704f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.16
cc_211 VPB SUM 0.00614182f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=0.825
cc_212 N_A_79_21#_c_218_n N_A_c_468_n 4.84784e-19 $X=1.825 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_213 N_A_79_21#_c_219_n N_A_c_468_n 4.83622e-19 $X=1.825 $Y=1.43 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_79_21#_c_220_n N_A_c_468_n 0.00314729f $X=2.37 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_215 N_A_79_21#_c_235_n N_A_c_468_n 0.00305547f $X=2.14 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_216 N_A_79_21#_c_221_n N_A_c_468_n 0.00116088f $X=1.825 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_79_21#_c_226_n N_A_c_468_n 0.0185821f $X=1.73 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_79_21#_M1035_g N_A_M1034_g 0.0343293f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_219_n N_A_M1034_g 0.00289362f $X=1.825 $Y=1.43 $X2=0 $Y2=0
cc_220 N_A_79_21#_c_235_n N_A_M1034_g 0.00743643f $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A_79_21#_c_236_n N_A_M1034_g 0.00710889f $X=2.225 $Y=1.91 $X2=0 $Y2=0
cc_222 N_A_79_21#_c_248_p N_A_M1034_g 0.00932588f $X=2.31 $Y=1.995 $X2=0 $Y2=0
cc_223 N_A_79_21#_c_215_n N_A_M1024_g 0.0229188f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_79_21#_c_218_n N_A_M1024_g 0.00329971f $X=1.825 $Y=1.075 $X2=0 $Y2=0
cc_225 N_A_79_21#_c_220_n N_A_M1024_g 0.0122069f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_79_21#_c_224_n N_A_M1024_g 0.00789386f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_227 N_A_79_21#_c_222_n N_A_M1018_g 0.00338905f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_228 N_A_79_21#_c_254_p N_A_M1019_g 2.03713e-19 $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_229 N_A_79_21#_M1017_g N_A_M1039_g 0.0165256f $X=6.28 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_79_21#_c_222_n N_A_M1039_g 0.00113591f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_231 N_A_79_21#_c_228_n N_A_M1039_g 7.05654e-19 $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_232 N_A_79_21#_M1016_g N_A_M1004_g 0.044851f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_233 N_A_79_21#_c_218_n N_A_c_474_n 0.00621239f $X=1.825 $Y=1.075 $X2=0 $Y2=0
cc_234 N_A_79_21#_c_219_n N_A_c_474_n 0.00580417f $X=1.825 $Y=1.43 $X2=0 $Y2=0
cc_235 N_A_79_21#_c_220_n N_A_c_474_n 0.0213932f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_79_21#_c_235_n N_A_c_474_n 0.01802f $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A_79_21#_c_254_p N_A_c_474_n 5.72713e-19 $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_238 N_A_79_21#_c_221_n N_A_c_474_n 0.01443f $X=1.825 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_79_21#_c_226_n N_A_c_474_n 3.11849e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_79_21#_c_254_p A 0.00286887f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_241 N_A_79_21#_c_224_n A 0.0242805f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_242 N_A_79_21#_c_222_n N_A_c_476_n 0.0499403f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_243 N_A_79_21#_c_223_n N_A_c_476_n 0.0274738f $X=3.14 $Y=0.85 $X2=0 $Y2=0
cc_244 N_A_79_21#_c_224_n N_A_c_476_n 0.00520722f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_245 N_A_79_21#_c_254_p N_A_c_477_n 0.00219144f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_246 N_A_79_21#_c_221_n N_A_c_477_n 7.37443e-19 $X=1.825 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_79_21#_c_224_n N_A_c_477_n 0.00196475f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_248 N_A_79_21#_c_222_n N_A_c_478_n 0.124008f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_249 N_A_79_21#_c_222_n N_A_c_479_n 0.0266325f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_250 N_A_79_21#_M1016_g N_A_c_480_n 0.00200174f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_251 N_A_79_21#_c_222_n N_A_c_480_n 0.0490684f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_252 N_A_79_21#_c_225_n N_A_c_480_n 0.0249445f $X=6.695 $Y=0.85 $X2=0 $Y2=0
cc_253 N_A_79_21#_c_227_n N_A_c_480_n 0.00198965f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_254 N_A_79_21#_c_228_n N_A_c_480_n 0.0168241f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_255 N_A_79_21#_M1016_g N_A_c_481_n 4.24426e-19 $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_256 N_A_79_21#_c_222_n N_A_c_481_n 0.0261862f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_257 N_A_79_21#_c_228_n N_A_c_481_n 3.07492e-19 $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_258 N_A_79_21#_c_222_n N_A_c_482_n 0.00306165f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_259 N_A_79_21#_c_228_n N_A_c_483_n 0.00133594f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_260 N_A_79_21#_c_222_n N_A_c_484_n 0.00187757f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_261 N_A_79_21#_c_222_n N_A_c_485_n 0.00347599f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_262 N_A_79_21#_c_227_n N_A_c_485_n 0.0196997f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_263 N_A_79_21#_c_228_n N_A_c_485_n 0.00115543f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_264 N_A_79_21#_c_222_n N_A_c_486_n 0.00253419f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_265 N_A_79_21#_c_227_n N_A_c_486_n 0.00311574f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_266 N_A_79_21#_c_228_n N_A_c_486_n 0.014709f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_267 N_A_79_21#_c_228_n N_A_c_488_n 0.0106157f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_268 N_A_79_21#_c_236_n N_B_M1006_g 0.00311481f $X=2.225 $Y=1.91 $X2=0 $Y2=0
cc_269 N_A_79_21#_c_254_p N_B_M1006_g 0.0112199f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_270 N_A_79_21#_c_223_n N_B_M1010_g 5.09542e-19 $X=3.14 $Y=0.85 $X2=0 $Y2=0
cc_271 N_A_79_21#_c_224_n N_B_M1010_g 0.0287112f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_272 N_A_79_21#_c_222_n N_B_c_738_n 0.0124329f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_273 N_A_79_21#_c_222_n N_B_c_739_n 0.00188483f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_274 N_A_79_21#_c_228_n N_B_M1030_g 0.00137141f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_275 N_A_79_21#_c_222_n N_B_c_742_n 0.00336351f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_276 N_A_79_21#_c_219_n B 0.00184322f $X=1.825 $Y=1.43 $X2=0 $Y2=0
cc_277 N_A_79_21#_c_235_n B 0.0151331f $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_278 N_A_79_21#_c_236_n B 0.00196768f $X=2.225 $Y=1.91 $X2=0 $Y2=0
cc_279 N_A_79_21#_c_254_p B 0.0325517f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_280 N_A_79_21#_c_224_n B 0.00649937f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_281 N_A_79_21#_c_254_p N_B_c_752_n 6.65518e-19 $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_282 N_A_79_21#_c_235_n N_B_c_753_n 5.80777e-19 $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_283 N_A_79_21#_c_254_p N_B_c_753_n 0.00363907f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_284 N_A_79_21#_M1016_g N_B_c_754_n 0.00173774f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_285 N_A_79_21#_c_227_n N_B_c_754_n 5.89663e-19 $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_286 N_A_79_21#_c_228_n N_B_c_754_n 0.00221477f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_287 N_A_79_21#_c_235_n N_B_c_757_n 5.79882e-19 $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_288 N_A_79_21#_c_254_p N_B_c_757_n 0.00127292f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_289 N_A_79_21#_c_222_n N_B_c_743_n 0.00135025f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_290 N_A_79_21#_c_222_n N_CIN_M1021_g 0.00462124f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_291 N_A_79_21#_c_223_n N_CIN_M1021_g 0.00221673f $X=3.14 $Y=0.85 $X2=0 $Y2=0
cc_292 N_A_79_21#_c_224_n N_CIN_M1021_g 0.00480374f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_293 N_A_79_21#_c_254_p N_CIN_M1032_g 0.0151768f $X=2.735 $Y=1.995 $X2=0 $Y2=0
cc_294 N_A_79_21#_M1016_g N_CIN_M1009_g 0.0251353f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_295 N_A_79_21#_M1017_g N_CIN_M1037_g 0.0126f $X=6.28 $Y=0.445 $X2=0 $Y2=0
cc_296 N_A_79_21#_M1016_g N_CIN_M1037_g 0.00538209f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_297 N_A_79_21#_c_225_n N_CIN_M1037_g 0.00134755f $X=6.695 $Y=0.85 $X2=0 $Y2=0
cc_298 N_A_79_21#_c_227_n N_CIN_M1037_g 0.0160461f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_299 N_A_79_21#_c_228_n N_CIN_M1037_g 0.0149352f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_300 N_A_79_21#_c_222_n N_CIN_c_970_n 0.00117521f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_301 N_A_79_21#_c_222_n N_CIN_c_973_n 0.021158f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_302 N_A_79_21#_c_222_n N_CIN_c_974_n 0.00158362f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_303 N_A_79_21#_M1016_g N_CIN_c_988_n 0.0148758f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_304 N_A_79_21#_c_227_n N_CIN_c_988_n 0.00169335f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_305 N_A_79_21#_c_228_n N_CIN_c_988_n 0.0114048f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_306 N_A_79_21#_c_254_p N_CIN_c_976_n 8.27068e-19 $X=2.735 $Y=1.995 $X2=0
+ $Y2=0
cc_307 N_A_79_21#_c_222_n N_CIN_c_976_n 9.52651e-19 $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_308 N_A_79_21#_c_223_n N_CIN_c_976_n 9.74524e-19 $X=3.14 $Y=0.85 $X2=0 $Y2=0
cc_309 N_A_79_21#_c_224_n N_CIN_c_976_n 2.46291e-19 $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_310 N_A_79_21#_c_254_p N_CIN_c_977_n 5.46291e-19 $X=2.735 $Y=1.995 $X2=0
+ $Y2=0
cc_311 N_A_79_21#_c_222_n N_CIN_c_977_n 0.00500146f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_312 N_A_79_21#_c_223_n N_CIN_c_977_n 0.0013906f $X=3.14 $Y=0.85 $X2=0 $Y2=0
cc_313 N_A_79_21#_c_224_n N_CIN_c_977_n 0.00266523f $X=2.995 $Y=0.85 $X2=0 $Y2=0
cc_314 N_A_79_21#_c_222_n N_CIN_c_978_n 0.00174757f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_315 N_A_79_21#_M1016_g N_CIN_c_993_n 0.0153265f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_316 N_A_79_21#_c_228_n N_CIN_c_993_n 7.33058e-19 $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_317 N_A_79_21#_M1016_g N_CIN_c_994_n 0.00668536f $X=6.28 $Y=2.165 $X2=0 $Y2=0
cc_318 N_A_79_21#_c_228_n N_CIN_c_994_n 0.0119833f $X=6.34 $Y=1.04 $X2=0 $Y2=0
cc_319 N_A_79_21#_c_225_n N_A_1271_47#_c_1212_n 0.00212136f $X=6.695 $Y=0.85
+ $X2=0 $Y2=0
cc_320 N_A_79_21#_c_228_n N_A_1271_47#_c_1212_n 0.00815626f $X=6.34 $Y=1.04
+ $X2=0 $Y2=0
cc_321 N_A_79_21#_c_225_n N_A_1271_47#_c_1200_n 0.00161347f $X=6.695 $Y=0.85
+ $X2=0 $Y2=0
cc_322 N_A_79_21#_c_228_n N_A_1271_47#_c_1200_n 0.00199818f $X=6.34 $Y=1.04
+ $X2=0 $Y2=0
cc_323 N_A_79_21#_c_222_n N_A_1271_47#_c_1216_n 4.08874e-19 $X=6.55 $Y=0.85
+ $X2=0 $Y2=0
cc_324 N_A_79_21#_c_225_n N_A_1271_47#_c_1216_n 0.00101125f $X=6.695 $Y=0.85
+ $X2=0 $Y2=0
cc_325 N_A_79_21#_c_228_n N_A_1271_47#_c_1216_n 0.0120345f $X=6.34 $Y=1.04 $X2=0
+ $Y2=0
cc_326 N_A_79_21#_c_219_n N_VPWR_M1035_s 0.00185736f $X=1.825 $Y=1.43 $X2=0
+ $Y2=0
cc_327 N_A_79_21#_c_235_n N_VPWR_M1035_s 0.00422101f $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_328 N_A_79_21#_M1011_g N_VPWR_c_1374_n 0.00146448f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A_79_21#_M1031_g N_VPWR_c_1374_n 0.00142012f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_A_79_21#_M1035_g N_VPWR_c_1375_n 0.00176026f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_331 N_A_79_21#_c_219_n N_VPWR_c_1375_n 0.00271926f $X=1.825 $Y=1.43 $X2=0
+ $Y2=0
cc_332 N_A_79_21#_c_235_n N_VPWR_c_1375_n 0.0050401f $X=2.14 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A_79_21#_M1016_g N_VPWR_c_1378_n 0.00114511f $X=6.28 $Y=2.165 $X2=0
+ $Y2=0
cc_334 N_A_79_21#_M1005_g N_VPWR_c_1382_n 0.00542163f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_79_21#_M1011_g N_VPWR_c_1382_n 0.00542163f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_79_21#_M1031_g N_VPWR_c_1389_n 0.00585385f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A_79_21#_M1035_g N_VPWR_c_1389_n 0.00585385f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_79_21#_c_254_p N_VPWR_c_1390_n 0.0329257f $X=2.735 $Y=1.995 $X2=0
+ $Y2=0
cc_339 N_A_79_21#_c_248_p N_VPWR_c_1390_n 0.00265378f $X=2.31 $Y=1.995 $X2=0
+ $Y2=0
cc_340 N_A_79_21#_M1016_g N_VPWR_c_1393_n 0.00585385f $X=6.28 $Y=2.165 $X2=0
+ $Y2=0
cc_341 N_A_79_21#_M1006_d N_VPWR_c_1373_n 0.00337082f $X=2.725 $Y=1.855 $X2=0
+ $Y2=0
cc_342 N_A_79_21#_M1005_g N_VPWR_c_1373_n 0.0104567f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_79_21#_M1011_g N_VPWR_c_1373_n 0.00950252f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_79_21#_M1031_g N_VPWR_c_1373_n 0.0105371f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_345 N_A_79_21#_M1035_g N_VPWR_c_1373_n 0.0105934f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_79_21#_M1016_g N_VPWR_c_1373_n 0.0108663f $X=6.28 $Y=2.165 $X2=0
+ $Y2=0
cc_347 N_A_79_21#_c_254_p N_VPWR_c_1373_n 0.0276946f $X=2.735 $Y=1.995 $X2=0
+ $Y2=0
cc_348 N_A_79_21#_c_248_p N_VPWR_c_1373_n 0.00425201f $X=2.31 $Y=1.995 $X2=0
+ $Y2=0
cc_349 N_A_79_21#_M1005_g N_VPWR_c_1401_n 0.00316354f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A_79_21#_c_212_n N_COUT_c_1538_n 0.00365765f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_79_21#_M1005_g N_COUT_c_1538_n 0.00365765f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_79_21#_c_213_n N_COUT_c_1538_n 4.4806e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A_79_21#_M1011_g N_COUT_c_1538_n 4.4806e-19 $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_79_21#_c_380_p N_COUT_c_1538_n 0.0134679f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_355 N_A_79_21#_c_226_n N_COUT_c_1538_n 0.0180538f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A_79_21#_c_212_n N_COUT_c_1550_n 0.0111734f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_79_21#_c_213_n N_COUT_c_1550_n 0.0065119f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_79_21#_c_214_n N_COUT_c_1550_n 5.25965e-19 $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_359 N_A_79_21#_c_213_n N_COUT_c_1539_n 0.00845772f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_360 N_A_79_21#_c_214_n N_COUT_c_1539_n 0.0105731f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_79_21#_c_215_n N_COUT_c_1539_n 0.00129105f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_362 N_A_79_21#_c_380_p N_COUT_c_1539_n 0.0130429f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_363 N_A_79_21#_c_218_n N_COUT_c_1539_n 0.00527838f $X=1.825 $Y=1.075 $X2=0
+ $Y2=0
cc_364 N_A_79_21#_c_390_p N_COUT_c_1539_n 0.00655392f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_365 N_A_79_21#_c_226_n N_COUT_c_1539_n 0.00348171f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_366 N_A_79_21#_c_212_n N_COUT_c_1540_n 0.0120485f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_367 N_A_79_21#_c_213_n N_COUT_c_1540_n 0.00124227f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_368 N_A_79_21#_c_380_p N_COUT_c_1540_n 0.0525681f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A_79_21#_c_226_n N_COUT_c_1540_n 0.00221825f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_370 N_A_79_21#_M1011_g N_COUT_c_1542_n 0.0106747f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_A_79_21#_M1031_g N_COUT_c_1542_n 0.0143489f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_372 N_A_79_21#_M1035_g N_COUT_c_1542_n 0.00126569f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_373 N_A_79_21#_c_380_p N_COUT_c_1542_n 0.0136608f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_79_21#_c_219_n N_COUT_c_1542_n 0.0142595f $X=1.825 $Y=1.43 $X2=0
+ $Y2=0
cc_375 N_A_79_21#_c_226_n N_COUT_c_1542_n 0.00452908f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_376 N_A_79_21#_M1005_g N_COUT_c_1543_n 0.0148116f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_377 N_A_79_21#_M1011_g N_COUT_c_1543_n 0.00175109f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_378 N_A_79_21#_c_380_p N_COUT_c_1543_n 0.0556709f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_79_21#_c_226_n N_COUT_c_1543_n 0.00221825f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_380 N_A_79_21#_c_213_n N_COUT_c_1574_n 4.60039e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A_79_21#_c_214_n N_COUT_c_1574_n 0.00491662f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A_79_21#_c_215_n N_COUT_c_1574_n 0.0038f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_383 N_A_79_21#_c_390_p N_COUT_c_1574_n 0.00520964f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_79_21#_c_214_n N_COUT_c_1578_n 0.0021751f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_385 N_A_79_21#_c_215_n N_COUT_c_1578_n 0.00306707f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_386 N_A_79_21#_c_380_p N_COUT_c_1578_n 0.0033652f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A_79_21#_c_226_n N_COUT_c_1578_n 7.13848e-19 $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_388 N_A_79_21#_M1035_g N_COUT_c_1582_n 0.00176697f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_389 N_A_79_21#_c_219_n N_COUT_c_1582_n 0.00545866f $X=1.825 $Y=1.43 $X2=0
+ $Y2=0
cc_390 N_A_79_21#_c_236_n N_COUT_c_1582_n 0.00309381f $X=2.225 $Y=1.91 $X2=0
+ $Y2=0
cc_391 N_A_79_21#_c_380_p N_COUT_c_1585_n 0.00151726f $X=1.74 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_A_79_21#_M1005_g N_COUT_c_1586_n 0.0166869f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_393 N_A_79_21#_M1011_g N_COUT_c_1586_n 0.0109416f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_394 N_A_79_21#_M1031_g N_COUT_c_1586_n 7.55688e-19 $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_395 N_A_79_21#_c_254_p A_456_371# 0.00639507f $X=2.735 $Y=1.995 $X2=-0.19
+ $Y2=-0.24
cc_396 N_A_79_21#_M1016_g N_A_1014_369#_c_1640_n 0.0048174f $X=6.28 $Y=2.165
+ $X2=0 $Y2=0
cc_397 N_A_79_21#_c_218_n N_VGND_M1036_d 7.2386e-19 $X=1.825 $Y=1.075 $X2=0
+ $Y2=0
cc_398 N_A_79_21#_c_220_n N_VGND_M1036_d 0.00448661f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A_79_21#_c_390_p N_VGND_M1036_d 5.36799e-19 $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A_79_21#_c_213_n N_VGND_c_1752_n 0.00146448f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_401 N_A_79_21#_c_214_n N_VGND_c_1752_n 0.00146448f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_402 N_A_79_21#_c_215_n N_VGND_c_1753_n 0.00285054f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_403 N_A_79_21#_c_220_n N_VGND_c_1753_n 0.016676f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A_79_21#_c_390_p N_VGND_c_1753_n 0.00368134f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_405 N_A_79_21#_c_224_n N_VGND_c_1753_n 0.0163179f $X=2.995 $Y=0.85 $X2=0
+ $Y2=0
cc_406 N_A_79_21#_c_222_n N_VGND_c_1754_n 0.00115864f $X=6.55 $Y=0.85 $X2=0
+ $Y2=0
cc_407 N_A_79_21#_c_222_n N_VGND_c_1755_n 0.00407154f $X=6.55 $Y=0.85 $X2=0
+ $Y2=0
cc_408 N_A_79_21#_M1017_g N_VGND_c_1756_n 0.00114511f $X=6.28 $Y=0.445 $X2=0
+ $Y2=0
cc_409 N_A_79_21#_c_222_n N_VGND_c_1756_n 0.00115864f $X=6.55 $Y=0.85 $X2=0
+ $Y2=0
cc_410 N_A_79_21#_c_212_n N_VGND_c_1760_n 0.00423442f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_411 N_A_79_21#_c_213_n N_VGND_c_1760_n 0.00423442f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_412 N_A_79_21#_M1017_g N_VGND_c_1762_n 0.00585385f $X=6.28 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_79_21#_c_214_n N_VGND_c_1769_n 0.00425388f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_414 N_A_79_21#_c_215_n N_VGND_c_1769_n 0.00474077f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_415 N_A_79_21#_c_390_p N_VGND_c_1769_n 0.0015722f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A_79_21#_c_220_n N_VGND_c_1770_n 0.00299685f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_A_79_21#_c_224_n N_VGND_c_1770_n 0.0457698f $X=2.995 $Y=0.85 $X2=0
+ $Y2=0
cc_418 N_A_79_21#_M1010_d N_VGND_c_1774_n 0.00277879f $X=2.78 $Y=0.235 $X2=0
+ $Y2=0
cc_419 N_A_79_21#_c_212_n N_VGND_c_1774_n 0.00670508f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A_79_21#_c_213_n N_VGND_c_1774_n 0.00575087f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_A_79_21#_c_214_n N_VGND_c_1774_n 0.00574144f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_422 N_A_79_21#_c_215_n N_VGND_c_1774_n 0.00764688f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_423 N_A_79_21#_M1017_g N_VGND_c_1774_n 0.00673586f $X=6.28 $Y=0.445 $X2=0
+ $Y2=0
cc_424 N_A_79_21#_c_220_n N_VGND_c_1774_n 0.00580564f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_425 N_A_79_21#_c_390_p N_VGND_c_1774_n 0.00335468f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_426 N_A_79_21#_c_222_n N_VGND_c_1774_n 0.156698f $X=6.55 $Y=0.85 $X2=0 $Y2=0
cc_427 N_A_79_21#_c_223_n N_VGND_c_1774_n 0.0149244f $X=3.14 $Y=0.85 $X2=0 $Y2=0
cc_428 N_A_79_21#_c_224_n N_VGND_c_1774_n 0.0219117f $X=2.995 $Y=0.85 $X2=0
+ $Y2=0
cc_429 N_A_79_21#_c_225_n N_VGND_c_1774_n 0.015806f $X=6.695 $Y=0.85 $X2=0 $Y2=0
cc_430 N_A_79_21#_c_228_n N_VGND_c_1774_n 0.00304902f $X=6.34 $Y=1.04 $X2=0
+ $Y2=0
cc_431 N_A_79_21#_c_212_n N_VGND_c_1779_n 0.00316354f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_A_79_21#_c_224_n A_461_47# 0.00728689f $X=2.995 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_433 N_A_79_21#_c_222_n N_A_658_47#_c_1937_n 0.0271275f $X=6.55 $Y=0.85 $X2=0
+ $Y2=0
cc_434 N_A_79_21#_c_222_n N_A_658_47#_c_1938_n 0.00797006f $X=6.55 $Y=0.85 $X2=0
+ $Y2=0
cc_435 N_A_79_21#_c_223_n N_A_658_47#_c_1938_n 0.00117968f $X=3.14 $Y=0.85 $X2=0
+ $Y2=0
cc_436 N_A_79_21#_c_224_n N_A_658_47#_c_1938_n 0.0081472f $X=2.995 $Y=0.85 $X2=0
+ $Y2=0
cc_437 N_A_79_21#_M1017_g N_A_1014_47#_c_1972_n 0.00472067f $X=6.28 $Y=0.445
+ $X2=0 $Y2=0
cc_438 N_A_79_21#_c_222_n N_A_1014_47#_c_1972_n 0.0286552f $X=6.55 $Y=0.85 $X2=0
+ $Y2=0
cc_439 N_A_79_21#_c_225_n N_A_1014_47#_c_1972_n 0.00140299f $X=6.695 $Y=0.85
+ $X2=0 $Y2=0
cc_440 N_A_79_21#_c_228_n N_A_1014_47#_c_1972_n 0.00128307f $X=6.34 $Y=1.04
+ $X2=0 $Y2=0
cc_441 N_A_79_21#_c_222_n N_A_1014_47#_c_1973_n 0.00610599f $X=6.55 $Y=0.85
+ $X2=0 $Y2=0
cc_442 N_A_M1034_g N_B_M1006_g 0.0383136f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_443 N_A_c_468_n N_B_M1010_g 0.00660104f $X=2.205 $Y=1.325 $X2=0 $Y2=0
cc_444 N_A_M1034_g N_B_M1010_g 0.00161938f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_445 N_A_M1024_g N_B_M1010_g 0.0382754f $X=2.23 $Y=0.445 $X2=0 $Y2=0
cc_446 N_A_c_474_n N_B_M1010_g 9.5302e-19 $X=2.34 $Y=1.16 $X2=0 $Y2=0
cc_447 A N_B_M1010_g 0.00925882f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_448 N_A_c_476_n N_B_M1010_g 0.00281072f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_449 N_A_c_477_n N_B_M1010_g 0.0017855f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_450 N_A_M1018_g N_B_c_737_n 0.0218633f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_451 N_A_c_478_n N_B_c_739_n 5.6387e-19 $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_452 N_A_c_479_n N_B_c_739_n 3.21623e-19 $X=4.06 $Y=1.19 $X2=0 $Y2=0
cc_453 N_A_c_482_n N_B_c_739_n 4.12248e-19 $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_454 N_A_M1019_g N_B_c_748_n 0.0329021f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_455 N_A_M1003_g N_B_M1030_g 0.043667f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_456 N_A_M1026_g N_B_M1030_g 0.00146789f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_457 N_A_c_483_n N_B_M1030_g 8.60102e-19 $X=7.155 $Y=1.19 $X2=0 $Y2=0
cc_458 N_A_c_488_n N_B_M1030_g 0.0135237f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_459 N_A_M1026_g N_B_M1007_g 0.0262997f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_460 N_A_M1034_g B 0.0011743f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_461 A B 0.0128348f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_462 N_A_c_476_n B 0.00561395f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_463 N_A_c_477_n B 0.00545311f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_464 N_A_M1019_g N_B_c_752_n 0.00360106f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_465 N_A_c_476_n N_B_c_752_n 0.0492111f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_466 N_A_c_478_n N_B_c_752_n 0.0518636f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_467 N_A_c_479_n N_B_c_752_n 0.0266263f $X=4.06 $Y=1.19 $X2=0 $Y2=0
cc_468 N_A_c_482_n N_B_c_752_n 0.00287761f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_469 N_A_c_484_n N_B_c_752_n 0.00189048f $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_470 N_A_c_476_n N_B_c_753_n 0.0274741f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_471 N_A_M1004_g N_B_c_754_n 0.00147663f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_472 N_A_c_478_n N_B_c_754_n 0.049641f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_473 N_A_c_480_n N_B_c_754_n 0.0886059f $X=7.01 $Y=1.19 $X2=0 $Y2=0
cc_474 N_A_c_481_n N_B_c_754_n 0.0275415f $X=5.92 $Y=1.19 $X2=0 $Y2=0
cc_475 N_A_c_483_n N_B_c_754_n 0.0266188f $X=7.155 $Y=1.19 $X2=0 $Y2=0
cc_476 N_A_c_486_n N_B_c_754_n 0.00168577f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_477 N_A_c_488_n N_B_c_754_n 0.00203106f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_478 N_A_c_478_n N_B_c_821_n 0.0274198f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_479 N_A_M1026_g N_B_c_755_n 0.00308106f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_480 N_A_c_487_n N_B_c_755_n 0.00186167f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_481 N_A_c_488_n N_B_c_755_n 0.00780453f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_482 N_A_M1026_g N_B_c_756_n 0.0100188f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_483 N_A_c_483_n N_B_c_756_n 0.00127994f $X=7.155 $Y=1.19 $X2=0 $Y2=0
cc_484 N_A_c_487_n N_B_c_756_n 0.00165748f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_485 N_A_c_488_n N_B_c_756_n 0.0454517f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_486 N_A_M1034_g N_B_c_757_n 0.018974f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_487 A N_B_c_757_n 0.00315799f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_488 N_A_c_477_n N_B_c_757_n 0.00353207f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_489 N_A_c_478_n N_B_c_758_n 0.00153932f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_490 N_A_c_478_n N_B_c_759_n 0.00207379f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_491 N_A_c_478_n N_B_c_743_n 0.00138637f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_492 N_A_M1026_g N_B_c_762_n 0.0159725f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_493 N_A_c_483_n N_B_c_762_n 7.30893e-19 $X=7.155 $Y=1.19 $X2=0 $Y2=0
cc_494 N_A_c_488_n N_B_c_762_n 0.00296771f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_495 N_A_M1018_g N_CIN_M1021_g 0.0261054f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_496 N_A_c_484_n N_CIN_M1032_g 0.0412793f $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_497 N_A_M1004_g N_CIN_M1013_g 0.0298654f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_498 N_A_c_480_n N_CIN_M1037_g 0.00347129f $X=7.01 $Y=1.19 $X2=0 $Y2=0
cc_499 N_A_c_483_n N_CIN_M1037_g 0.00137964f $X=7.155 $Y=1.19 $X2=0 $Y2=0
cc_500 N_A_c_488_n N_CIN_M1037_g 0.0036571f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_501 N_A_M1039_g N_CIN_c_969_n 0.0141455f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_502 N_A_M1039_g N_CIN_c_970_n 0.00744646f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_503 N_A_c_485_n N_CIN_c_970_n 0.0209378f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_504 N_A_c_476_n N_CIN_c_971_n 6.22985e-19 $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_505 N_A_c_477_n N_CIN_c_971_n 7.92681e-19 $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_506 N_A_c_482_n N_CIN_c_971_n 0.00575336f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_507 N_A_c_484_n N_CIN_c_971_n 0.00450847f $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_508 N_A_M1019_g N_CIN_c_984_n 0.0111093f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_509 N_A_c_476_n N_CIN_c_984_n 0.00162254f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_510 N_A_c_478_n N_CIN_c_984_n 6.24857e-19 $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_511 N_A_c_479_n N_CIN_c_984_n 5.60263e-19 $X=4.06 $Y=1.19 $X2=0 $Y2=0
cc_512 N_A_c_482_n N_CIN_c_984_n 0.0202345f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_513 N_A_c_484_n N_CIN_c_984_n 0.00255109f $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_514 N_A_M1019_g N_CIN_c_972_n 0.00429073f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_515 N_A_c_478_n N_CIN_c_972_n 0.00318872f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_516 N_A_c_479_n N_CIN_c_972_n 0.00137624f $X=4.06 $Y=1.19 $X2=0 $Y2=0
cc_517 N_A_c_482_n N_CIN_c_972_n 0.00802988f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_518 N_A_c_484_n N_CIN_c_972_n 5.0579e-19 $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_519 N_A_c_478_n N_CIN_c_973_n 0.0373123f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_520 N_A_c_481_n N_CIN_c_973_n 0.00126698f $X=5.92 $Y=1.19 $X2=0 $Y2=0
cc_521 N_A_c_485_n N_CIN_c_973_n 2.96853e-19 $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_522 N_A_c_486_n N_CIN_c_973_n 0.0147988f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_523 N_A_M1018_g N_CIN_c_974_n 0.00195651f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_524 N_A_c_478_n N_CIN_c_974_n 0.00560548f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_525 N_A_c_479_n N_CIN_c_974_n 0.00142282f $X=4.06 $Y=1.19 $X2=0 $Y2=0
cc_526 N_A_c_482_n N_CIN_c_974_n 0.0168914f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_527 N_A_c_484_n N_CIN_c_974_n 0.0010498f $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_528 N_A_M1004_g N_CIN_c_975_n 7.9432e-19 $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_529 N_A_c_478_n N_CIN_c_975_n 0.00235868f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_530 N_A_c_481_n N_CIN_c_975_n 0.00166046f $X=5.92 $Y=1.19 $X2=0 $Y2=0
cc_531 N_A_c_486_n N_CIN_c_975_n 0.00105124f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_532 N_A_M1004_g N_CIN_c_988_n 0.0100247f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_533 N_A_c_478_n N_CIN_c_988_n 3.16966e-19 $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_534 N_A_c_480_n N_CIN_c_988_n 0.00292909f $X=7.01 $Y=1.19 $X2=0 $Y2=0
cc_535 N_A_c_481_n N_CIN_c_988_n 0.00113336f $X=5.92 $Y=1.19 $X2=0 $Y2=0
cc_536 N_A_c_485_n N_CIN_c_988_n 5.94361e-19 $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_537 N_A_c_486_n N_CIN_c_988_n 0.0170478f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_538 N_A_M1018_g N_CIN_c_976_n 0.0215001f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_539 A N_CIN_c_976_n 8.76754e-19 $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_540 N_A_c_482_n N_CIN_c_976_n 7.99315e-19 $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_541 A N_CIN_c_977_n 0.00494488f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_542 N_A_c_476_n N_CIN_c_977_n 0.0143043f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_543 N_A_c_477_n N_CIN_c_977_n 2.10722e-19 $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_544 N_A_c_482_n N_CIN_c_977_n 0.0106105f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_545 N_A_c_484_n N_CIN_c_977_n 8.25882e-19 $X=3.695 $Y=1.195 $X2=0 $Y2=0
cc_546 N_A_M1004_g N_CIN_c_990_n 0.0213309f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_547 N_A_c_478_n N_CIN_c_990_n 8.79356e-19 $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_548 N_A_M1004_g N_CIN_c_991_n 0.00147223f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_549 N_A_c_478_n N_CIN_c_991_n 0.00232417f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_550 N_A_M1004_g N_CIN_c_978_n 0.00733914f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_551 N_A_c_478_n N_CIN_c_978_n 0.00214774f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_552 N_A_c_481_n N_CIN_c_978_n 0.00137864f $X=5.92 $Y=1.19 $X2=0 $Y2=0
cc_553 N_A_c_486_n N_CIN_c_978_n 0.00203847f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_554 N_A_c_480_n N_CIN_c_994_n 0.00212697f $X=7.01 $Y=1.19 $X2=0 $Y2=0
cc_555 N_A_M1003_g N_A_1271_47#_c_1195_n 0.020681f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_556 N_A_M1026_g N_A_1271_47#_M1002_g 0.0316775f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_557 N_A_M1003_g N_A_1271_47#_c_1212_n 0.00349977f $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_558 N_A_c_480_n N_A_1271_47#_c_1212_n 0.00451776f $X=7.01 $Y=1.19 $X2=0 $Y2=0
cc_559 N_A_c_483_n N_A_1271_47#_c_1212_n 0.00220053f $X=7.155 $Y=1.19 $X2=0
+ $Y2=0
cc_560 N_A_c_488_n N_A_1271_47#_c_1212_n 0.00641421f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_561 N_A_M1003_g N_A_1271_47#_c_1225_n 0.00339087f $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_562 N_A_M1003_g N_A_1271_47#_c_1199_n 0.0120577f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_563 N_A_c_487_n N_A_1271_47#_c_1199_n 0.00292686f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_564 N_A_c_488_n N_A_1271_47#_c_1199_n 0.0297985f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_565 N_A_c_488_n N_A_1271_47#_c_1200_n 0.0146449f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_566 N_A_M1026_g N_A_1271_47#_c_1230_n 0.011406f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_567 N_A_c_487_n N_A_1271_47#_c_1230_n 7.79054e-19 $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_568 N_A_c_488_n N_A_1271_47#_c_1230_n 0.00240743f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_569 N_A_M1026_g N_A_1271_47#_c_1233_n 0.00499834f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_570 N_A_M1003_g N_A_1271_47#_c_1201_n 0.00306196f $X=7.66 $Y=0.445 $X2=0
+ $Y2=0
cc_571 N_A_c_487_n N_A_1271_47#_c_1201_n 2.24683e-19 $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_572 N_A_c_488_n N_A_1271_47#_c_1201_n 0.00663255f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_573 N_A_M1026_g N_A_1271_47#_c_1202_n 0.00244048f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_574 N_A_c_487_n N_A_1271_47#_c_1202_n 0.00111224f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_575 N_A_c_488_n N_A_1271_47#_c_1202_n 0.00241081f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_576 N_A_M1026_g N_A_1271_47#_c_1210_n 0.00113171f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_577 N_A_c_487_n N_A_1271_47#_c_1203_n 6.24375e-19 $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_578 N_A_c_488_n N_A_1271_47#_c_1203_n 0.0159237f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_579 N_A_c_487_n N_A_1271_47#_c_1204_n 0.0159689f $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_580 N_A_c_488_n N_A_1271_47#_c_1204_n 9.44274e-19 $X=7.72 $Y=1.16 $X2=0 $Y2=0
cc_581 N_A_M1034_g N_VPWR_c_1375_n 0.00846964f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_582 N_A_M1019_g N_VPWR_c_1376_n 0.00760687f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_583 N_A_M1004_g N_VPWR_c_1378_n 0.00761262f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_584 N_A_M1026_g N_VPWR_c_1379_n 0.00313672f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_585 N_A_M1034_g N_VPWR_c_1390_n 0.00382403f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_586 N_A_M1019_g N_VPWR_c_1390_n 0.00337001f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_587 N_A_M1004_g N_VPWR_c_1393_n 0.00337001f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_588 N_A_M1026_g N_VPWR_c_1393_n 0.00422112f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_589 N_A_M1034_g N_VPWR_c_1373_n 0.00451477f $X=2.205 $Y=2.17 $X2=0 $Y2=0
cc_590 N_A_M1019_g N_VPWR_c_1373_n 0.00397658f $X=3.635 $Y=2.165 $X2=0 $Y2=0
cc_591 N_A_M1004_g N_VPWR_c_1373_n 0.00403935f $X=5.835 $Y=2.165 $X2=0 $Y2=0
cc_592 N_A_M1026_g N_VPWR_c_1373_n 0.00605013f $X=7.72 $Y=2.17 $X2=0 $Y2=0
cc_593 N_A_M1019_g N_A_658_369#_c_1617_n 0.0100291f $X=3.635 $Y=2.165 $X2=0
+ $Y2=0
cc_594 N_A_M1004_g N_A_1014_369#_c_1640_n 0.0111197f $X=5.835 $Y=2.165 $X2=0
+ $Y2=0
cc_595 N_A_M1024_g N_VGND_c_1753_n 0.00801931f $X=2.23 $Y=0.445 $X2=0 $Y2=0
cc_596 N_A_M1018_g N_VGND_c_1754_n 0.00760016f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_597 N_A_M1039_g N_VGND_c_1756_n 0.00760591f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_598 N_A_M1003_g N_VGND_c_1757_n 0.00810631f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_599 N_A_M1039_g N_VGND_c_1762_n 0.00337001f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_600 N_A_M1003_g N_VGND_c_1762_n 0.00341689f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_601 N_A_M1024_g N_VGND_c_1770_n 0.00341689f $X=2.23 $Y=0.445 $X2=0 $Y2=0
cc_602 N_A_M1018_g N_VGND_c_1770_n 0.00337001f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_603 N_A_M1024_g N_VGND_c_1774_n 0.00418888f $X=2.23 $Y=0.445 $X2=0 $Y2=0
cc_604 N_A_M1018_g N_VGND_c_1774_n 0.00377406f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_605 N_A_M1039_g N_VGND_c_1774_n 0.00383683f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_606 N_A_M1003_g N_VGND_c_1774_n 0.00420045f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_607 N_A_M1018_g N_A_658_47#_c_1937_n 0.0108136f $X=3.635 $Y=0.445 $X2=0 $Y2=0
cc_608 N_A_c_476_n N_A_658_47#_c_1937_n 0.00108134f $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_609 N_A_c_478_n N_A_658_47#_c_1937_n 0.00161385f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_610 N_A_c_479_n N_A_658_47#_c_1937_n 9.66928e-19 $X=4.06 $Y=1.19 $X2=0 $Y2=0
cc_611 N_A_c_482_n N_A_658_47#_c_1937_n 0.0169746f $X=3.915 $Y=1.19 $X2=0 $Y2=0
cc_612 N_A_c_484_n N_A_658_47#_c_1937_n 0.00247695f $X=3.695 $Y=1.195 $X2=0
+ $Y2=0
cc_613 N_A_c_476_n N_A_658_47#_c_1938_n 5.45312e-19 $X=3.77 $Y=1.19 $X2=0 $Y2=0
cc_614 N_A_M1039_g N_A_1014_47#_c_1972_n 0.00973522f $X=5.835 $Y=0.445 $X2=0
+ $Y2=0
cc_615 N_A_c_478_n N_A_1014_47#_c_1972_n 0.00124068f $X=5.63 $Y=1.19 $X2=0 $Y2=0
cc_616 N_A_c_480_n N_A_1014_47#_c_1972_n 7.16872e-19 $X=7.01 $Y=1.19 $X2=0 $Y2=0
cc_617 N_A_c_481_n N_A_1014_47#_c_1972_n 4.03515e-19 $X=5.92 $Y=1.19 $X2=0 $Y2=0
cc_618 N_A_c_485_n N_A_1014_47#_c_1972_n 0.00230741f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_619 N_A_c_486_n N_A_1014_47#_c_1972_n 0.0230574f $X=5.84 $Y=1.04 $X2=0 $Y2=0
cc_620 N_B_M1010_g N_CIN_M1021_g 0.0244199f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_621 N_B_M1006_g N_CIN_M1032_g 0.0254422f $X=2.65 $Y=2.17 $X2=0 $Y2=0
cc_622 N_B_M1010_g N_CIN_M1032_g 0.0117014f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_623 B N_CIN_M1032_g 0.00181415f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_624 N_B_c_752_n N_CIN_M1032_g 0.00429611f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_625 N_B_c_753_n N_CIN_M1032_g 0.00221673f $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_626 N_B_c_758_n N_CIN_M1013_g 0.0268107f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_627 N_B_c_759_n N_CIN_M1013_g 3.15588e-19 $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_628 N_B_c_762_n N_CIN_M1009_g 0.0352431f $X=7.24 $Y=1.53 $X2=0 $Y2=0
cc_629 N_B_M1030_g N_CIN_M1037_g 0.0500916f $X=7.18 $Y=0.445 $X2=0 $Y2=0
cc_630 N_B_c_740_n N_CIN_c_969_n 0.00946436f $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_631 N_B_c_742_n N_CIN_c_970_n 0.00946436f $X=4.995 $Y=0.805 $X2=0 $Y2=0
cc_632 N_B_M1010_g N_CIN_c_971_n 8.26322e-19 $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_633 B N_CIN_c_971_n 0.00851593f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_634 N_B_c_752_n N_CIN_c_971_n 0.0085825f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_635 N_B_c_753_n N_CIN_c_971_n 0.00173655f $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_636 N_B_c_739_n N_CIN_c_984_n 0.00203699f $X=4.13 $Y=0.805 $X2=0 $Y2=0
cc_637 N_B_c_747_n N_CIN_c_984_n 0.0111006f $X=4.695 $Y=1.695 $X2=0 $Y2=0
cc_638 N_B_c_748_n N_CIN_c_984_n 0.00751562f $X=4.13 $Y=1.695 $X2=0 $Y2=0
cc_639 N_B_c_752_n N_CIN_c_984_n 0.0266023f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_640 N_B_c_821_n N_CIN_c_984_n 2.72288e-19 $X=5 $Y=1.53 $X2=0 $Y2=0
cc_641 N_B_c_758_n N_CIN_c_984_n 2.61162e-19 $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_642 N_B_c_759_n N_CIN_c_984_n 0.0100882f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_643 N_B_M1006_g N_CIN_c_985_n 2.07028e-19 $X=2.65 $Y=2.17 $X2=0 $Y2=0
cc_644 B N_CIN_c_985_n 0.00918003f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_645 N_B_c_752_n N_CIN_c_985_n 0.00591938f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_646 N_B_c_753_n N_CIN_c_985_n 0.00122285f $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_647 N_B_c_752_n N_CIN_c_972_n 0.00984268f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_648 N_B_c_821_n N_CIN_c_972_n 8.96072e-19 $X=5 $Y=1.53 $X2=0 $Y2=0
cc_649 N_B_c_758_n N_CIN_c_972_n 0.00315065f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_650 N_B_c_759_n N_CIN_c_972_n 0.00699272f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_651 N_B_c_743_n N_CIN_c_972_n 2.3672e-19 $X=4.882 $Y=1.355 $X2=0 $Y2=0
cc_652 N_B_c_738_n N_CIN_c_973_n 0.0147995f $X=4.92 $Y=0.805 $X2=0 $Y2=0
cc_653 N_B_c_747_n N_CIN_c_973_n 0.0061986f $X=4.695 $Y=1.695 $X2=0 $Y2=0
cc_654 N_B_c_752_n N_CIN_c_973_n 0.00184237f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_655 N_B_c_754_n N_CIN_c_973_n 0.00209743f $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_656 N_B_c_821_n N_CIN_c_973_n 0.00103879f $X=5 $Y=1.53 $X2=0 $Y2=0
cc_657 N_B_c_758_n N_CIN_c_973_n 0.00231696f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_658 N_B_c_759_n N_CIN_c_973_n 0.0258113f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_659 N_B_c_743_n N_CIN_c_973_n 0.0188183f $X=4.882 $Y=1.355 $X2=0 $Y2=0
cc_660 N_B_c_738_n N_CIN_c_974_n 0.00347447f $X=4.92 $Y=0.805 $X2=0 $Y2=0
cc_661 N_B_c_754_n N_CIN_c_975_n 4.57159e-19 $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_662 N_B_c_821_n N_CIN_c_975_n 8.51268e-19 $X=5 $Y=1.53 $X2=0 $Y2=0
cc_663 N_B_c_743_n N_CIN_c_975_n 0.00397174f $X=4.882 $Y=1.355 $X2=0 $Y2=0
cc_664 N_B_c_754_n N_CIN_c_988_n 0.0425084f $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_665 N_B_M1010_g N_CIN_c_976_n 0.0143765f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_666 N_B_c_753_n N_CIN_c_976_n 9.74524e-19 $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_667 N_B_M1010_g N_CIN_c_977_n 9.22498e-19 $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_668 B N_CIN_c_977_n 0.00197411f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_669 N_B_c_752_n N_CIN_c_977_n 0.00217963f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_670 N_B_c_753_n N_CIN_c_977_n 8.46704e-19 $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_671 N_B_c_758_n N_CIN_c_990_n 0.0216836f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_672 N_B_c_759_n N_CIN_c_990_n 3.87164e-19 $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_673 N_B_c_754_n N_CIN_c_991_n 0.0164483f $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_674 N_B_c_821_n N_CIN_c_991_n 0.00171886f $X=5 $Y=1.53 $X2=0 $Y2=0
cc_675 N_B_c_758_n N_CIN_c_991_n 0.00153667f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_676 N_B_c_759_n N_CIN_c_991_n 0.0135944f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_677 N_B_c_743_n N_CIN_c_978_n 0.0225963f $X=4.882 $Y=1.355 $X2=0 $Y2=0
cc_678 N_B_c_754_n N_CIN_c_993_n 0.00175799f $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_679 N_B_c_756_n N_CIN_c_993_n 0.00134146f $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_680 N_B_c_762_n N_CIN_c_993_n 0.0500916f $X=7.24 $Y=1.53 $X2=0 $Y2=0
cc_681 N_B_M1030_g N_CIN_c_994_n 5.62374e-19 $X=7.18 $Y=0.445 $X2=0 $Y2=0
cc_682 N_B_M1007_g N_CIN_c_994_n 0.00428927f $X=7.18 $Y=2.17 $X2=0 $Y2=0
cc_683 N_B_c_754_n N_CIN_c_994_n 0.0141879f $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_684 N_B_c_756_n N_CIN_c_994_n 0.017102f $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_685 N_B_c_762_n N_CIN_c_994_n 5.23813e-19 $X=7.24 $Y=1.53 $X2=0 $Y2=0
cc_686 N_B_c_756_n N_A_1271_47#_M1002_g 3.1636e-19 $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_687 N_B_M1007_g N_A_1271_47#_c_1246_n 0.0173719f $X=7.18 $Y=2.17 $X2=0 $Y2=0
cc_688 N_B_c_754_n N_A_1271_47#_c_1246_n 0.0120753f $X=7.47 $Y=1.53 $X2=0 $Y2=0
cc_689 N_B_c_756_n N_A_1271_47#_c_1246_n 0.011759f $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_690 N_B_c_762_n N_A_1271_47#_c_1246_n 5.22774e-19 $X=7.24 $Y=1.53 $X2=0 $Y2=0
cc_691 N_B_M1030_g N_A_1271_47#_c_1212_n 0.0132015f $X=7.18 $Y=0.445 $X2=0 $Y2=0
cc_692 N_B_M1030_g N_A_1271_47#_c_1200_n 0.00438384f $X=7.18 $Y=0.445 $X2=0
+ $Y2=0
cc_693 N_B_c_755_n N_A_1271_47#_c_1230_n 8.48123e-19 $X=7.615 $Y=1.53 $X2=0
+ $Y2=0
cc_694 N_B_c_756_n N_A_1271_47#_c_1230_n 0.00776504f $X=7.615 $Y=1.53 $X2=0
+ $Y2=0
cc_695 N_B_c_756_n N_A_1271_47#_c_1233_n 0.0071466f $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_696 N_B_c_755_n N_A_1271_47#_c_1202_n 0.00138572f $X=7.615 $Y=1.53 $X2=0
+ $Y2=0
cc_697 N_B_c_756_n N_A_1271_47#_c_1202_n 8.41183e-19 $X=7.615 $Y=1.53 $X2=0
+ $Y2=0
cc_698 N_B_M1007_g N_A_1271_47#_c_1257_n 0.00429324f $X=7.18 $Y=2.17 $X2=0 $Y2=0
cc_699 N_B_c_755_n N_A_1271_47#_c_1257_n 9.31973e-19 $X=7.615 $Y=1.53 $X2=0
+ $Y2=0
cc_700 N_B_c_756_n N_A_1271_47#_c_1257_n 0.0107388f $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_701 N_B_c_755_n N_A_1271_47#_c_1210_n 0.00128946f $X=7.615 $Y=1.53 $X2=0
+ $Y2=0
cc_702 N_B_c_756_n N_A_1271_47#_c_1210_n 0.0106926f $X=7.615 $Y=1.53 $X2=0 $Y2=0
cc_703 N_B_M1006_g N_VPWR_c_1375_n 0.00163718f $X=2.65 $Y=2.17 $X2=0 $Y2=0
cc_704 N_B_c_746_n N_VPWR_c_1376_n 0.00677587f $X=4.055 $Y=1.77 $X2=0 $Y2=0
cc_705 N_B_c_746_n N_VPWR_c_1377_n 0.00321545f $X=4.055 $Y=1.77 $X2=0 $Y2=0
cc_706 N_B_c_747_n N_VPWR_c_1377_n 0.00489764f $X=4.695 $Y=1.695 $X2=0 $Y2=0
cc_707 N_B_c_752_n N_VPWR_c_1377_n 5.45078e-19 $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_708 N_B_c_821_n N_VPWR_c_1377_n 0.00157163f $X=5 $Y=1.53 $X2=0 $Y2=0
cc_709 N_B_c_759_n N_VPWR_c_1377_n 0.0225991f $X=4.83 $Y=1.52 $X2=0 $Y2=0
cc_710 N_B_c_761_n N_VPWR_c_1377_n 0.0114275f $X=4.882 $Y=1.77 $X2=0 $Y2=0
cc_711 N_B_c_761_n N_VPWR_c_1378_n 5.31689e-19 $X=4.882 $Y=1.77 $X2=0 $Y2=0
cc_712 N_B_M1006_g N_VPWR_c_1390_n 0.00425831f $X=2.65 $Y=2.17 $X2=0 $Y2=0
cc_713 N_B_c_746_n N_VPWR_c_1391_n 0.00337001f $X=4.055 $Y=1.77 $X2=0 $Y2=0
cc_714 N_B_c_761_n N_VPWR_c_1392_n 0.0046653f $X=4.882 $Y=1.77 $X2=0 $Y2=0
cc_715 N_B_M1007_g N_VPWR_c_1393_n 0.00357877f $X=7.18 $Y=2.17 $X2=0 $Y2=0
cc_716 N_B_M1006_g N_VPWR_c_1373_n 0.00633573f $X=2.65 $Y=2.17 $X2=0 $Y2=0
cc_717 N_B_c_746_n N_VPWR_c_1373_n 0.0053254f $X=4.055 $Y=1.77 $X2=0 $Y2=0
cc_718 N_B_M1007_g N_VPWR_c_1373_n 0.00573192f $X=7.18 $Y=2.17 $X2=0 $Y2=0
cc_719 N_B_c_761_n N_VPWR_c_1373_n 0.00799591f $X=4.882 $Y=1.77 $X2=0 $Y2=0
cc_720 N_B_c_746_n N_A_658_369#_c_1617_n 0.0107429f $X=4.055 $Y=1.77 $X2=0 $Y2=0
cc_721 N_B_c_747_n N_A_658_369#_c_1617_n 0.00540826f $X=4.695 $Y=1.695 $X2=0
+ $Y2=0
cc_722 N_B_c_752_n N_A_658_369#_c_1617_n 0.00782028f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_723 N_B_c_752_n N_A_658_369#_c_1623_n 0.00104195f $X=4.71 $Y=1.53 $X2=0 $Y2=0
cc_724 N_B_c_754_n N_A_1014_369#_c_1640_n 0.00513411f $X=7.47 $Y=1.53 $X2=0
+ $Y2=0
cc_725 N_B_c_754_n N_A_1014_369#_c_1643_n 0.00484515f $X=7.47 $Y=1.53 $X2=0
+ $Y2=0
cc_726 N_B_M1010_g N_VGND_c_1753_n 0.00121824f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_727 N_B_c_737_n N_VGND_c_1754_n 0.00676915f $X=4.055 $Y=0.73 $X2=0 $Y2=0
cc_728 N_B_c_737_n N_VGND_c_1755_n 0.00208038f $X=4.055 $Y=0.73 $X2=0 $Y2=0
cc_729 N_B_c_738_n N_VGND_c_1755_n 0.0045972f $X=4.92 $Y=0.805 $X2=0 $Y2=0
cc_730 N_B_c_740_n N_VGND_c_1755_n 0.00827538f $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_731 N_B_c_740_n N_VGND_c_1756_n 5.31689e-19 $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_732 N_B_M1030_g N_VGND_c_1757_n 0.00120942f $X=7.18 $Y=0.445 $X2=0 $Y2=0
cc_733 N_B_M1030_g N_VGND_c_1762_n 0.00357877f $X=7.18 $Y=0.445 $X2=0 $Y2=0
cc_734 N_B_M1010_g N_VGND_c_1770_n 0.00357668f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_735 N_B_c_737_n N_VGND_c_1771_n 0.00337001f $X=4.055 $Y=0.73 $X2=0 $Y2=0
cc_736 N_B_c_738_n N_VGND_c_1771_n 0.00469312f $X=4.92 $Y=0.805 $X2=0 $Y2=0
cc_737 N_B_c_740_n N_VGND_c_1772_n 0.0046653f $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_738 N_B_M1010_g N_VGND_c_1774_n 0.00566808f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_739 N_B_c_737_n N_VGND_c_1774_n 0.00512288f $X=4.055 $Y=0.73 $X2=0 $Y2=0
cc_740 N_B_c_738_n N_VGND_c_1774_n 0.00336079f $X=4.92 $Y=0.805 $X2=0 $Y2=0
cc_741 N_B_c_740_n N_VGND_c_1774_n 0.00446764f $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_742 N_B_M1030_g N_VGND_c_1774_n 0.00530375f $X=7.18 $Y=0.445 $X2=0 $Y2=0
cc_743 N_B_c_737_n N_A_658_47#_c_1937_n 0.00758462f $X=4.055 $Y=0.73 $X2=0 $Y2=0
cc_744 N_B_c_738_n N_A_658_47#_c_1937_n 0.00812182f $X=4.92 $Y=0.805 $X2=0 $Y2=0
cc_745 N_B_c_739_n N_A_658_47#_c_1937_n 0.00392189f $X=4.13 $Y=0.805 $X2=0 $Y2=0
cc_746 N_B_c_740_n N_A_658_47#_c_1937_n 0.00310565f $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_747 N_B_c_740_n N_A_658_47#_c_1954_n 0.00158481f $X=4.995 $Y=0.73 $X2=0 $Y2=0
cc_748 N_B_c_740_n N_A_1014_47#_c_1973_n 0.00420459f $X=4.995 $Y=0.73 $X2=0
+ $Y2=0
cc_749 N_CIN_M1009_g N_A_1271_47#_c_1246_n 0.0125611f $X=6.705 $Y=2.165 $X2=0
+ $Y2=0
cc_750 N_CIN_c_988_n N_A_1271_47#_c_1246_n 0.0057196f $X=6.595 $Y=1.6 $X2=0
+ $Y2=0
cc_751 N_CIN_c_993_n N_A_1271_47#_c_1246_n 0.00187747f $X=6.76 $Y=1.52 $X2=0
+ $Y2=0
cc_752 N_CIN_c_994_n N_A_1271_47#_c_1246_n 0.011642f $X=6.76 $Y=1.52 $X2=0 $Y2=0
cc_753 N_CIN_M1037_g N_A_1271_47#_c_1212_n 0.00979993f $X=6.82 $Y=0.445 $X2=0
+ $Y2=0
cc_754 N_CIN_c_994_n N_A_1271_47#_c_1257_n 5.83799e-19 $X=6.76 $Y=1.52 $X2=0
+ $Y2=0
cc_755 N_CIN_M1032_g N_VPWR_c_1376_n 0.00119528f $X=3.215 $Y=2.165 $X2=0 $Y2=0
cc_756 N_CIN_M1013_g N_VPWR_c_1377_n 7.98505e-19 $X=5.415 $Y=2.165 $X2=0 $Y2=0
cc_757 N_CIN_M1013_g N_VPWR_c_1378_n 0.00640108f $X=5.415 $Y=2.165 $X2=0 $Y2=0
cc_758 N_CIN_M1032_g N_VPWR_c_1390_n 0.00541359f $X=3.215 $Y=2.165 $X2=0 $Y2=0
cc_759 N_CIN_M1013_g N_VPWR_c_1392_n 0.00337001f $X=5.415 $Y=2.165 $X2=0 $Y2=0
cc_760 N_CIN_M1009_g N_VPWR_c_1393_n 0.00357877f $X=6.705 $Y=2.165 $X2=0 $Y2=0
cc_761 N_CIN_M1032_g N_VPWR_c_1373_n 0.010123f $X=3.215 $Y=2.165 $X2=0 $Y2=0
cc_762 N_CIN_M1013_g N_VPWR_c_1373_n 0.00397658f $X=5.415 $Y=2.165 $X2=0 $Y2=0
cc_763 N_CIN_M1009_g N_VPWR_c_1373_n 0.00542737f $X=6.705 $Y=2.165 $X2=0 $Y2=0
cc_764 N_CIN_c_984_n N_A_658_369#_c_1617_n 0.0442431f $X=4.17 $Y=1.655 $X2=0
+ $Y2=0
cc_765 N_CIN_c_984_n N_A_658_369#_c_1623_n 0.00577586f $X=4.17 $Y=1.655 $X2=0
+ $Y2=0
cc_766 N_CIN_c_985_n N_A_658_369#_c_1623_n 0.00557804f $X=3.42 $Y=1.655 $X2=0
+ $Y2=0
cc_767 N_CIN_M1013_g N_A_1014_369#_c_1640_n 0.0110354f $X=5.415 $Y=2.165 $X2=0
+ $Y2=0
cc_768 N_CIN_c_988_n N_A_1014_369#_c_1640_n 0.00893804f $X=6.595 $Y=1.6 $X2=0
+ $Y2=0
cc_769 N_CIN_c_990_n N_A_1014_369#_c_1640_n 0.00113985f $X=5.415 $Y=1.52 $X2=0
+ $Y2=0
cc_770 N_CIN_c_991_n N_A_1014_369#_c_1640_n 0.02703f $X=5.58 $Y=1.56 $X2=0 $Y2=0
cc_771 N_CIN_c_991_n N_A_1014_369#_c_1643_n 0.00362847f $X=5.58 $Y=1.56 $X2=0
+ $Y2=0
cc_772 N_CIN_c_994_n A_1356_369# 0.00154519f $X=6.76 $Y=1.52 $X2=-0.19 $Y2=-0.24
cc_773 N_CIN_M1021_g N_VGND_c_1754_n 0.00118455f $X=3.215 $Y=0.445 $X2=0 $Y2=0
cc_774 N_CIN_c_969_n N_VGND_c_1755_n 5.44952e-19 $X=5.417 $Y=0.73 $X2=0 $Y2=0
cc_775 N_CIN_c_973_n N_VGND_c_1755_n 0.00546777f $X=5.22 $Y=1.107 $X2=0 $Y2=0
cc_776 N_CIN_c_969_n N_VGND_c_1756_n 0.00639437f $X=5.417 $Y=0.73 $X2=0 $Y2=0
cc_777 N_CIN_M1037_g N_VGND_c_1762_n 0.00357877f $X=6.82 $Y=0.445 $X2=0 $Y2=0
cc_778 N_CIN_M1021_g N_VGND_c_1770_n 0.00585385f $X=3.215 $Y=0.445 $X2=0 $Y2=0
cc_779 N_CIN_c_969_n N_VGND_c_1772_n 0.00337001f $X=5.417 $Y=0.73 $X2=0 $Y2=0
cc_780 N_CIN_M1021_g N_VGND_c_1774_n 0.00670748f $X=3.215 $Y=0.445 $X2=0 $Y2=0
cc_781 N_CIN_M1037_g N_VGND_c_1774_n 0.00532102f $X=6.82 $Y=0.445 $X2=0 $Y2=0
cc_782 N_CIN_c_969_n N_VGND_c_1774_n 0.00377406f $X=5.417 $Y=0.73 $X2=0 $Y2=0
cc_783 N_CIN_c_973_n N_A_658_47#_c_1937_n 5.77639e-19 $X=5.22 $Y=1.107 $X2=0
+ $Y2=0
cc_784 N_CIN_c_974_n N_A_658_47#_c_1937_n 0.0110711f $X=4.34 $Y=1.107 $X2=0
+ $Y2=0
cc_785 N_CIN_M1021_g N_A_658_47#_c_1938_n 0.00129924f $X=3.215 $Y=0.445 $X2=0
+ $Y2=0
cc_786 N_CIN_c_976_n N_A_658_47#_c_1938_n 2.17239e-19 $X=3.215 $Y=1.19 $X2=0
+ $Y2=0
cc_787 N_CIN_c_977_n N_A_658_47#_c_1938_n 0.00270907f $X=3.335 $Y=1.19 $X2=0
+ $Y2=0
cc_788 N_CIN_c_969_n N_A_1014_47#_c_1972_n 0.00669222f $X=5.417 $Y=0.73 $X2=0
+ $Y2=0
cc_789 N_CIN_c_970_n N_A_1014_47#_c_1972_n 0.00441497f $X=5.417 $Y=0.88 $X2=0
+ $Y2=0
cc_790 N_CIN_c_973_n N_A_1014_47#_c_1972_n 0.00624534f $X=5.22 $Y=1.107 $X2=0
+ $Y2=0
cc_791 N_CIN_c_990_n N_A_1014_47#_c_1972_n 9.85703e-19 $X=5.415 $Y=1.52 $X2=0
+ $Y2=0
cc_792 N_CIN_c_991_n N_A_1014_47#_c_1972_n 0.00195538f $X=5.58 $Y=1.56 $X2=0
+ $Y2=0
cc_793 N_CIN_c_973_n N_A_1014_47#_c_1973_n 0.0111405f $X=5.22 $Y=1.107 $X2=0
+ $Y2=0
cc_794 N_A_1271_47#_c_1230_n N_VPWR_M1026_d 0.00544362f $X=7.935 $Y=2.02 $X2=0
+ $Y2=0
cc_795 N_A_1271_47#_c_1233_n N_VPWR_M1026_d 0.00399486f $X=8.02 $Y=1.935 $X2=0
+ $Y2=0
cc_796 N_A_1271_47#_c_1210_n N_VPWR_M1026_d 0.001562f $X=8.14 $Y=1.555 $X2=0
+ $Y2=0
cc_797 N_A_1271_47#_M1002_g N_VPWR_c_1379_n 0.00671141f $X=8.195 $Y=1.985 $X2=0
+ $Y2=0
cc_798 N_A_1271_47#_M1008_g N_VPWR_c_1379_n 5.32661e-19 $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_799 N_A_1271_47#_c_1230_n N_VPWR_c_1379_n 0.0166961f $X=7.935 $Y=2.02 $X2=0
+ $Y2=0
cc_800 N_A_1271_47#_c_1210_n N_VPWR_c_1379_n 5.96676e-19 $X=8.14 $Y=1.555 $X2=0
+ $Y2=0
cc_801 N_A_1271_47#_M1008_g N_VPWR_c_1380_n 0.00149687f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_802 N_A_1271_47#_M1012_g N_VPWR_c_1380_n 0.00859499f $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_803 N_A_1271_47#_M1025_g N_VPWR_c_1381_n 0.00438629f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_804 N_A_1271_47#_M1002_g N_VPWR_c_1384_n 0.00486043f $X=8.195 $Y=1.985 $X2=0
+ $Y2=0
cc_805 N_A_1271_47#_M1008_g N_VPWR_c_1384_n 0.00557614f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_806 N_A_1271_47#_M1012_g N_VPWR_c_1386_n 0.00542953f $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_807 N_A_1271_47#_M1025_g N_VPWR_c_1386_n 0.00542953f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_808 N_A_1271_47#_c_1246_n N_VPWR_c_1393_n 0.0606537f $X=7.44 $Y=2.295 $X2=0
+ $Y2=0
cc_809 N_A_1271_47#_c_1230_n N_VPWR_c_1393_n 0.00312966f $X=7.935 $Y=2.02 $X2=0
+ $Y2=0
cc_810 N_A_1271_47#_c_1257_n N_VPWR_c_1393_n 0.0108964f $X=7.525 $Y=2.02 $X2=0
+ $Y2=0
cc_811 N_A_1271_47#_M1016_d N_VPWR_c_1373_n 0.00406702f $X=6.355 $Y=1.845 $X2=0
+ $Y2=0
cc_812 N_A_1271_47#_M1002_g N_VPWR_c_1373_n 0.00819893f $X=8.195 $Y=1.985 $X2=0
+ $Y2=0
cc_813 N_A_1271_47#_M1008_g N_VPWR_c_1373_n 0.00986831f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_814 N_A_1271_47#_M1012_g N_VPWR_c_1373_n 0.009908f $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_815 N_A_1271_47#_M1025_g N_VPWR_c_1373_n 0.0105519f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_816 N_A_1271_47#_c_1246_n N_VPWR_c_1373_n 0.0375122f $X=7.44 $Y=2.295 $X2=0
+ $Y2=0
cc_817 N_A_1271_47#_c_1230_n N_VPWR_c_1373_n 0.00650684f $X=7.935 $Y=2.02 $X2=0
+ $Y2=0
cc_818 N_A_1271_47#_c_1257_n N_VPWR_c_1373_n 0.00642843f $X=7.525 $Y=2.02 $X2=0
+ $Y2=0
cc_819 N_A_1271_47#_c_1246_n A_1356_369# 0.00563231f $X=7.44 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_820 N_A_1271_47#_c_1246_n A_1451_371# 0.00398461f $X=7.44 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_821 N_A_1271_47#_c_1257_n A_1451_371# 0.0080653f $X=7.525 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_822 N_A_1271_47#_c_1195_n N_SUM_c_1666_n 0.005977f $X=8.195 $Y=0.995 $X2=0
+ $Y2=0
cc_823 N_A_1271_47#_c_1196_n N_SUM_c_1666_n 0.00485022f $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_824 N_A_1271_47#_c_1199_n N_SUM_c_1666_n 0.0139693f $X=8.055 $Y=0.74 $X2=0
+ $Y2=0
cc_825 N_A_1271_47#_c_1201_n N_SUM_c_1666_n 0.00617628f $X=8.14 $Y=1.075 $X2=0
+ $Y2=0
cc_826 N_A_1271_47#_c_1300_p N_SUM_c_1666_n 0.0199585f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_827 N_A_1271_47#_c_1204_n N_SUM_c_1666_n 0.00367134f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_828 N_A_1271_47#_M1008_g N_SUM_c_1671_n 0.0111746f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_829 N_A_1271_47#_M1012_g N_SUM_c_1671_n 0.0111139f $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_830 N_A_1271_47#_c_1300_p N_SUM_c_1671_n 0.0412347f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_831 N_A_1271_47#_c_1204_n N_SUM_c_1671_n 0.00453387f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_832 N_A_1271_47#_M1002_g N_SUM_c_1672_n 0.0011776f $X=8.195 $Y=1.985 $X2=0
+ $Y2=0
cc_833 N_A_1271_47#_M1008_g N_SUM_c_1672_n 0.00206908f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_834 N_A_1271_47#_c_1202_n N_SUM_c_1672_n 0.00434169f $X=8.14 $Y=1.47 $X2=0
+ $Y2=0
cc_835 N_A_1271_47#_c_1300_p N_SUM_c_1672_n 0.0134703f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_836 N_A_1271_47#_c_1210_n N_SUM_c_1672_n 0.00919212f $X=8.14 $Y=1.555 $X2=0
+ $Y2=0
cc_837 N_A_1271_47#_c_1204_n N_SUM_c_1672_n 0.0012838f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_838 N_A_1271_47#_c_1196_n N_SUM_c_1667_n 0.00850187f $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_839 N_A_1271_47#_c_1197_n N_SUM_c_1667_n 0.00845772f $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_840 N_A_1271_47#_c_1300_p N_SUM_c_1667_n 0.0355133f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_841 N_A_1271_47#_c_1204_n N_SUM_c_1667_n 0.00221825f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_842 N_A_1271_47#_c_1196_n N_SUM_c_1696_n 5.20755e-19 $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_843 N_A_1271_47#_c_1197_n N_SUM_c_1696_n 0.00627667f $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_844 N_A_1271_47#_c_1198_n N_SUM_c_1696_n 0.0108955f $X=9.535 $Y=0.995 $X2=0
+ $Y2=0
cc_845 N_A_1271_47#_M1008_g N_SUM_c_1699_n 7.9249e-19 $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_846 N_A_1271_47#_M1012_g N_SUM_c_1699_n 0.0121185f $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_847 N_A_1271_47#_M1025_g N_SUM_c_1699_n 0.0163599f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_848 N_A_1271_47#_c_1198_n N_SUM_c_1668_n 0.0114727f $X=9.535 $Y=0.995 $X2=0
+ $Y2=0
cc_849 N_A_1271_47#_M1025_g N_SUM_c_1673_n 0.0136897f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_850 N_A_1271_47#_c_1196_n N_SUM_c_1704_n 0.00263861f $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_851 N_A_1271_47#_c_1197_n N_SUM_c_1704_n 5.25981e-19 $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_852 N_A_1271_47#_c_1300_p N_SUM_c_1704_n 0.00205752f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_853 N_A_1271_47#_c_1204_n N_SUM_c_1704_n 7.21164e-19 $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_854 N_A_1271_47#_M1008_g N_SUM_c_1708_n 0.00252508f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_855 N_A_1271_47#_c_1300_p N_SUM_c_1708_n 0.00238329f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_856 N_A_1271_47#_c_1204_n N_SUM_c_1708_n 7.88595e-19 $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_857 N_A_1271_47#_M1002_g N_SUM_c_1711_n 0.00136769f $X=8.195 $Y=1.985 $X2=0
+ $Y2=0
cc_858 N_A_1271_47#_M1008_g N_SUM_c_1711_n 0.00522273f $X=8.615 $Y=1.985 $X2=0
+ $Y2=0
cc_859 N_A_1271_47#_M1012_g N_SUM_c_1711_n 6.90881e-19 $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_860 N_A_1271_47#_c_1210_n N_SUM_c_1711_n 0.00384346f $X=8.14 $Y=1.555 $X2=0
+ $Y2=0
cc_861 N_A_1271_47#_c_1197_n N_SUM_c_1669_n 0.00110513f $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_862 N_A_1271_47#_c_1198_n N_SUM_c_1669_n 0.00138739f $X=9.535 $Y=0.995 $X2=0
+ $Y2=0
cc_863 N_A_1271_47#_c_1300_p N_SUM_c_1669_n 0.0227276f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_864 N_A_1271_47#_c_1204_n N_SUM_c_1669_n 0.00230171f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_865 N_A_1271_47#_M1012_g N_SUM_c_1674_n 0.00170419f $X=9.115 $Y=1.985 $X2=0
+ $Y2=0
cc_866 N_A_1271_47#_M1025_g N_SUM_c_1674_n 0.00199489f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_867 N_A_1271_47#_c_1300_p N_SUM_c_1674_n 0.0228621f $X=9.28 $Y=1.16 $X2=0
+ $Y2=0
cc_868 N_A_1271_47#_c_1204_n N_SUM_c_1674_n 0.00231083f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_869 N_A_1271_47#_c_1198_n SUM 0.0202277f $X=9.535 $Y=0.995 $X2=0 $Y2=0
cc_870 N_A_1271_47#_c_1300_p SUM 0.0104024f $X=9.28 $Y=1.16 $X2=0 $Y2=0
cc_871 N_A_1271_47#_c_1199_n N_VGND_M1003_d 0.00795696f $X=8.055 $Y=0.74 $X2=0
+ $Y2=0
cc_872 N_A_1271_47#_c_1201_n N_VGND_M1003_d 7.72373e-19 $X=8.14 $Y=1.075 $X2=0
+ $Y2=0
cc_873 N_A_1271_47#_c_1195_n N_VGND_c_1757_n 0.00523592f $X=8.195 $Y=0.995 $X2=0
+ $Y2=0
cc_874 N_A_1271_47#_c_1212_n N_VGND_c_1757_n 0.0124309f $X=7.305 $Y=0.38 $X2=0
+ $Y2=0
cc_875 N_A_1271_47#_c_1199_n N_VGND_c_1757_n 0.0186618f $X=8.055 $Y=0.74 $X2=0
+ $Y2=0
cc_876 N_A_1271_47#_c_1196_n N_VGND_c_1758_n 0.00268723f $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_877 N_A_1271_47#_c_1197_n N_VGND_c_1758_n 0.00146448f $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_878 N_A_1271_47#_c_1198_n N_VGND_c_1759_n 0.00316354f $X=9.535 $Y=0.995 $X2=0
+ $Y2=0
cc_879 N_A_1271_47#_c_1212_n N_VGND_c_1762_n 0.0115639f $X=7.305 $Y=0.38 $X2=0
+ $Y2=0
cc_880 N_A_1271_47#_c_1199_n N_VGND_c_1762_n 0.00378546f $X=8.055 $Y=0.74 $X2=0
+ $Y2=0
cc_881 N_A_1271_47#_c_1216_n N_VGND_c_1762_n 0.047666f $X=6.635 $Y=0.425 $X2=0
+ $Y2=0
cc_882 N_A_1271_47#_c_1195_n N_VGND_c_1764_n 0.00475129f $X=8.195 $Y=0.995 $X2=0
+ $Y2=0
cc_883 N_A_1271_47#_c_1196_n N_VGND_c_1764_n 0.00424416f $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_884 N_A_1271_47#_c_1199_n N_VGND_c_1764_n 0.00279992f $X=8.055 $Y=0.74 $X2=0
+ $Y2=0
cc_885 N_A_1271_47#_c_1197_n N_VGND_c_1766_n 0.00425021f $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_886 N_A_1271_47#_c_1198_n N_VGND_c_1766_n 0.00425021f $X=9.535 $Y=0.995 $X2=0
+ $Y2=0
cc_887 N_A_1271_47#_M1017_d N_VGND_c_1774_n 0.00285934f $X=6.355 $Y=0.235 $X2=0
+ $Y2=0
cc_888 N_A_1271_47#_c_1195_n N_VGND_c_1774_n 0.00785437f $X=8.195 $Y=0.995 $X2=0
+ $Y2=0
cc_889 N_A_1271_47#_c_1196_n N_VGND_c_1774_n 0.00593357f $X=8.695 $Y=0.995 $X2=0
+ $Y2=0
cc_890 N_A_1271_47#_c_1197_n N_VGND_c_1774_n 0.00573673f $X=9.115 $Y=0.995 $X2=0
+ $Y2=0
cc_891 N_A_1271_47#_c_1198_n N_VGND_c_1774_n 0.0067844f $X=9.535 $Y=0.995 $X2=0
+ $Y2=0
cc_892 N_A_1271_47#_c_1212_n N_VGND_c_1774_n 0.00651702f $X=7.305 $Y=0.38 $X2=0
+ $Y2=0
cc_893 N_A_1271_47#_c_1199_n N_VGND_c_1774_n 0.012465f $X=8.055 $Y=0.74 $X2=0
+ $Y2=0
cc_894 N_A_1271_47#_c_1216_n N_VGND_c_1774_n 0.0226199f $X=6.635 $Y=0.425 $X2=0
+ $Y2=0
cc_895 N_A_1271_47#_c_1216_n N_A_1014_47#_c_1992_n 0.0162015f $X=6.635 $Y=0.425
+ $X2=0 $Y2=0
cc_896 N_A_1271_47#_c_1212_n A_1379_47# 0.00288105f $X=7.305 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_897 N_A_1271_47#_c_1212_n A_1451_47# 0.00470231f $X=7.305 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_898 N_A_1271_47#_c_1225_n A_1451_47# 0.00165868f $X=7.39 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_899 N_VPWR_c_1373_n N_COUT_M1005_d 0.00216035f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_900 N_VPWR_c_1373_n N_COUT_M1031_d 0.00320325f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_901 N_VPWR_M1011_s N_COUT_c_1542_n 0.00181725f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_902 N_VPWR_c_1374_n N_COUT_c_1542_n 0.0108451f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_903 N_VPWR_M1005_s N_COUT_c_1543_n 0.00388989f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_904 N_VPWR_c_1401_n N_COUT_c_1543_n 0.0112622f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_905 N_VPWR_c_1389_n N_COUT_c_1595_n 0.0128161f $X=1.815 $Y=2.72 $X2=0 $Y2=0
cc_906 N_VPWR_c_1373_n N_COUT_c_1595_n 0.008011f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_907 N_VPWR_c_1373_n N_COUT_c_1585_n 0.0013839f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_908 N_VPWR_c_1382_n N_COUT_c_1586_n 0.0167767f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_909 N_VPWR_c_1373_n N_COUT_c_1586_n 0.0120986f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_910 N_VPWR_c_1373_n A_456_371# 0.0034659f $X=9.89 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_911 N_VPWR_c_1373_n N_A_658_369#_M1032_d 0.00409863f $X=9.89 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_912 N_VPWR_c_1373_n N_A_658_369#_M1038_d 0.00226128f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1390_n N_A_658_369#_c_1629_n 0.0111986f $X=3.68 $Y=2.72 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1373_n N_A_658_369#_c_1629_n 0.00642843f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_915 N_VPWR_M1019_d N_A_658_369#_c_1617_n 0.00319397f $X=3.71 $Y=1.845 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1376_n N_A_658_369#_c_1617_n 0.0158599f $X=3.845 $Y=2.36 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1377_n N_A_658_369#_c_1617_n 0.0131777f $X=4.785 $Y=2 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1390_n N_A_658_369#_c_1617_n 0.00255672f $X=3.68 $Y=2.72 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1391_n N_A_658_369#_c_1617_n 0.00255672f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1373_n N_A_658_369#_c_1617_n 0.0101119f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1377_n N_A_658_369#_c_1618_n 0.0255946f $X=4.785 $Y=2 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1391_n N_A_658_369#_c_1618_n 0.0159201f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1373_n N_A_658_369#_c_1618_n 0.00891562f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1373_n N_A_1014_369#_M1023_d 0.00409863f $X=9.89 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_925 N_VPWR_c_1373_n N_A_1014_369#_M1004_d 0.00516727f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1392_n N_A_1014_369#_c_1651_n 0.0111986f $X=5.46 $Y=2.72 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1373_n N_A_1014_369#_c_1651_n 0.00642843f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_928 N_VPWR_M1013_d N_A_1014_369#_c_1640_n 0.00340913f $X=5.49 $Y=1.845 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1378_n N_A_1014_369#_c_1640_n 0.0158599f $X=5.625 $Y=2.36 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1392_n N_A_1014_369#_c_1640_n 0.00255672f $X=5.46 $Y=2.72 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1393_n N_A_1014_369#_c_1640_n 0.00255672f $X=7.815 $Y=2.72 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1373_n N_A_1014_369#_c_1640_n 0.0101119f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1393_n N_A_1014_369#_c_1658_n 0.0114f $X=7.815 $Y=2.72 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1373_n N_A_1014_369#_c_1658_n 0.00642843f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1373_n A_1356_369# 0.00261003f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_936 N_VPWR_c_1373_n A_1451_371# 0.00323344f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_937 N_VPWR_c_1373_n N_SUM_M1002_s 0.00414458f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_938 N_VPWR_c_1373_n N_SUM_M1012_s 0.00217524f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_939 N_VPWR_M1008_d N_SUM_c_1671_n 0.00471065f $X=8.69 $Y=1.485 $X2=0 $Y2=0
cc_940 N_VPWR_c_1380_n N_SUM_c_1671_n 0.0112622f $X=8.825 $Y=1.96 $X2=0 $Y2=0
cc_941 N_VPWR_c_1380_n N_SUM_c_1699_n 0.0345851f $X=8.825 $Y=1.96 $X2=0 $Y2=0
cc_942 N_VPWR_c_1386_n N_SUM_c_1699_n 0.0150775f $X=9.66 $Y=2.72 $X2=0 $Y2=0
cc_943 N_VPWR_c_1373_n N_SUM_c_1699_n 0.0119688f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_944 N_VPWR_M1025_d N_SUM_c_1673_n 0.00600343f $X=9.61 $Y=1.485 $X2=0 $Y2=0
cc_945 N_VPWR_c_1381_n N_SUM_c_1673_n 0.0121925f $X=9.745 $Y=1.96 $X2=0 $Y2=0
cc_946 N_VPWR_c_1384_n N_SUM_c_1708_n 0.01214f $X=8.74 $Y=2.72 $X2=0 $Y2=0
cc_947 N_VPWR_c_1373_n N_SUM_c_1708_n 0.00842369f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_948 N_COUT_c_1540_n N_VGND_M1020_d 0.00311706f $X=0.845 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_949 N_COUT_c_1539_n N_VGND_M1028_d 0.00162006f $X=1.355 $Y=0.82 $X2=0 $Y2=0
cc_950 N_COUT_c_1539_n N_VGND_c_1752_n 0.0122414f $X=1.355 $Y=0.82 $X2=0 $Y2=0
cc_951 N_COUT_c_1550_n N_VGND_c_1760_n 0.0185358f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_952 N_COUT_c_1540_n N_VGND_c_1760_n 0.00390702f $X=0.845 $Y=0.82 $X2=0 $Y2=0
cc_953 N_COUT_c_1540_n VGND 0.00131872f $X=0.845 $Y=0.82 $X2=0 $Y2=0
cc_954 N_COUT_c_1539_n N_VGND_c_1769_n 0.00193763f $X=1.355 $Y=0.82 $X2=0 $Y2=0
cc_955 N_COUT_c_1578_n N_VGND_c_1769_n 0.0127666f $X=1.52 $Y=0.4 $X2=0 $Y2=0
cc_956 N_COUT_M1020_s N_VGND_c_1774_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_957 N_COUT_M1029_s N_VGND_c_1774_n 0.00219774f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_958 N_COUT_c_1550_n N_VGND_c_1774_n 0.012111f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_959 N_COUT_c_1539_n N_VGND_c_1774_n 0.00444316f $X=1.355 $Y=0.82 $X2=0 $Y2=0
cc_960 N_COUT_c_1540_n N_VGND_c_1774_n 0.0107045f $X=0.845 $Y=0.82 $X2=0 $Y2=0
cc_961 N_COUT_c_1578_n N_VGND_c_1774_n 0.0114218f $X=1.52 $Y=0.4 $X2=0 $Y2=0
cc_962 N_COUT_c_1540_n N_VGND_c_1779_n 0.0127122f $X=0.845 $Y=0.82 $X2=0 $Y2=0
cc_963 N_SUM_c_1667_n N_VGND_M1022_d 0.00162006f $X=9.16 $Y=0.82 $X2=0 $Y2=0
cc_964 N_SUM_c_1668_n N_VGND_M1033_d 0.00406491f $X=9.7 $Y=0.82 $X2=0 $Y2=0
cc_965 N_SUM_c_1667_n N_VGND_c_1758_n 0.0122414f $X=9.16 $Y=0.82 $X2=0 $Y2=0
cc_966 N_SUM_c_1668_n N_VGND_c_1759_n 0.0137399f $X=9.7 $Y=0.82 $X2=0 $Y2=0
cc_967 N_SUM_c_1667_n N_VGND_c_1764_n 0.00193763f $X=9.16 $Y=0.82 $X2=0 $Y2=0
cc_968 N_SUM_c_1704_n N_VGND_c_1764_n 0.0203536f $X=8.485 $Y=0.4 $X2=0 $Y2=0
cc_969 N_SUM_c_1667_n N_VGND_c_1766_n 0.00193763f $X=9.16 $Y=0.82 $X2=0 $Y2=0
cc_970 N_SUM_c_1696_n N_VGND_c_1766_n 0.0171957f $X=9.325 $Y=0.4 $X2=0 $Y2=0
cc_971 N_SUM_c_1668_n N_VGND_c_1766_n 0.00193763f $X=9.7 $Y=0.82 $X2=0 $Y2=0
cc_972 N_SUM_c_1668_n N_VGND_c_1773_n 0.00335113f $X=9.7 $Y=0.82 $X2=0 $Y2=0
cc_973 N_SUM_M1015_s N_VGND_c_1774_n 0.00457293f $X=8.27 $Y=0.235 $X2=0 $Y2=0
cc_974 N_SUM_M1027_s N_VGND_c_1774_n 0.00215764f $X=9.19 $Y=0.235 $X2=0 $Y2=0
cc_975 N_SUM_c_1667_n N_VGND_c_1774_n 0.00825759f $X=9.16 $Y=0.82 $X2=0 $Y2=0
cc_976 N_SUM_c_1696_n N_VGND_c_1774_n 0.0121066f $X=9.325 $Y=0.4 $X2=0 $Y2=0
cc_977 N_SUM_c_1668_n N_VGND_c_1774_n 0.0102792f $X=9.7 $Y=0.82 $X2=0 $Y2=0
cc_978 N_SUM_c_1704_n N_VGND_c_1774_n 0.012337f $X=8.485 $Y=0.4 $X2=0 $Y2=0
cc_979 N_VGND_c_1774_n A_461_47# 0.00286569f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_980 N_VGND_c_1774_n N_A_658_47#_M1021_d 0.00227466f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_981 N_VGND_c_1774_n N_A_658_47#_M1014_d 0.00204709f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_982 N_VGND_c_1770_n N_A_658_47#_c_1962_n 0.0111986f $X=3.68 $Y=0 $X2=0 $Y2=0
cc_983 N_VGND_c_1774_n N_A_658_47#_c_1962_n 0.00304042f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_984 N_VGND_M1018_d N_A_658_47#_c_1937_n 0.00158918f $X=3.71 $Y=0.235 $X2=0
+ $Y2=0
cc_985 N_VGND_c_1754_n N_A_658_47#_c_1937_n 0.0147553f $X=3.845 $Y=0.36 $X2=0
+ $Y2=0
cc_986 N_VGND_c_1770_n N_A_658_47#_c_1937_n 0.00255672f $X=3.68 $Y=0 $X2=0 $Y2=0
cc_987 N_VGND_c_1771_n N_A_658_47#_c_1937_n 0.00255672f $X=4.62 $Y=0 $X2=0 $Y2=0
cc_988 N_VGND_c_1774_n N_A_658_47#_c_1937_n 0.00461038f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_989 N_VGND_c_1755_n N_A_658_47#_c_1954_n 0.0131643f $X=4.785 $Y=0.405 $X2=0
+ $Y2=0
cc_990 N_VGND_c_1771_n N_A_658_47#_c_1954_n 0.0114f $X=4.62 $Y=0 $X2=0 $Y2=0
cc_991 N_VGND_c_1774_n N_A_658_47#_c_1954_n 0.00304042f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_992 N_VGND_c_1774_n N_A_1014_47#_M1000_d 0.00227466f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_993 N_VGND_c_1774_n N_A_1014_47#_M1039_d 0.00263427f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_994 N_VGND_c_1772_n N_A_1014_47#_c_1995_n 0.0111986f $X=5.46 $Y=0 $X2=0 $Y2=0
cc_995 N_VGND_c_1774_n N_A_1014_47#_c_1995_n 0.00304042f $X=9.89 $Y=0 $X2=0
+ $Y2=0
cc_996 N_VGND_M1001_d N_A_1014_47#_c_1972_n 0.00158918f $X=5.49 $Y=0.235 $X2=0
+ $Y2=0
cc_997 N_VGND_c_1756_n N_A_1014_47#_c_1972_n 0.0147553f $X=5.625 $Y=0.36 $X2=0
+ $Y2=0
cc_998 N_VGND_c_1762_n N_A_1014_47#_c_1972_n 0.00255672f $X=7.705 $Y=0 $X2=0
+ $Y2=0
cc_999 N_VGND_c_1772_n N_A_1014_47#_c_1972_n 0.00255672f $X=5.46 $Y=0 $X2=0
+ $Y2=0
cc_1000 N_VGND_c_1774_n N_A_1014_47#_c_1972_n 0.00461038f $X=9.89 $Y=0 $X2=0
+ $Y2=0
cc_1001 N_VGND_c_1762_n N_A_1014_47#_c_1992_n 0.0114f $X=7.705 $Y=0 $X2=0 $Y2=0
cc_1002 N_VGND_c_1774_n N_A_1014_47#_c_1992_n 0.00304042f $X=9.89 $Y=0 $X2=0
+ $Y2=0
cc_1003 N_VGND_c_1774_n A_1379_47# 0.00168648f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1004 N_VGND_c_1774_n A_1451_47# 0.0030831f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__and2_2.spice.SKY130_FD_SC_HD__AND2_2.pxi
* Created: Thu Aug 27 14:06:56 2020
* 
x_PM_SKY130_FD_SC_HD__AND2_2%A N_A_M1002_g N_A_M1001_g A A A N_A_c_56_n
+ N_A_c_57_n PM_SKY130_FD_SC_HD__AND2_2%A
x_PM_SKY130_FD_SC_HD__AND2_2%B N_B_M1000_g N_B_M1006_g B N_B_c_90_n
+ PM_SKY130_FD_SC_HD__AND2_2%B
x_PM_SKY130_FD_SC_HD__AND2_2%A_61_75# N_A_61_75#_M1002_s N_A_61_75#_M1001_d
+ N_A_61_75#_c_124_n N_A_61_75#_M1004_g N_A_61_75#_M1003_g N_A_61_75#_c_125_n
+ N_A_61_75#_M1007_g N_A_61_75#_M1005_g N_A_61_75#_c_126_n N_A_61_75#_c_127_n
+ N_A_61_75#_c_128_n N_A_61_75#_c_129_n N_A_61_75#_c_130_n N_A_61_75#_c_131_n
+ N_A_61_75#_c_138_n N_A_61_75#_c_139_n N_A_61_75#_c_140_n N_A_61_75#_c_132_n
+ N_A_61_75#_c_142_n PM_SKY130_FD_SC_HD__AND2_2%A_61_75#
x_PM_SKY130_FD_SC_HD__AND2_2%VPWR N_VPWR_M1001_s N_VPWR_M1006_d N_VPWR_M1005_s
+ N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n VPWR N_VPWR_c_228_n
+ N_VPWR_c_219_n PM_SKY130_FD_SC_HD__AND2_2%VPWR
x_PM_SKY130_FD_SC_HD__AND2_2%X N_X_M1004_s N_X_M1003_d N_X_c_260_n X X X X X X
+ N_X_c_276_n X PM_SKY130_FD_SC_HD__AND2_2%X
x_PM_SKY130_FD_SC_HD__AND2_2%VGND N_VGND_M1000_d N_VGND_M1007_d N_VGND_c_290_n
+ N_VGND_c_291_n N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n VGND
+ N_VGND_c_295_n N_VGND_c_296_n PM_SKY130_FD_SC_HD__AND2_2%VGND
cc_1 VNB N_A_M1002_g 0.0276839f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.585
cc_2 VNB A 0.0019668f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_3 VNB N_A_c_56_n 0.0362409f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_4 VNB N_A_c_57_n 0.0179007f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.325
cc_5 VNB N_B_M1000_g 0.0214729f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.585
cc_6 VNB N_B_c_90_n 0.0260976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_61_75#_c_124_n 0.0197599f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=2.065
cc_8 VNB N_A_61_75#_c_125_n 0.0225627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_61_75#_c_126_n 0.00808228f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.53
cc_10 VNB N_A_61_75#_c_127_n 0.0188995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_61_75#_c_128_n 0.0219949f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.2
cc_12 VNB N_A_61_75#_c_129_n 0.0162873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_61_75#_c_130_n 0.00748673f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.2
cc_14 VNB N_A_61_75#_c_131_n 0.0100642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_61_75#_c_132_n 0.00335652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_219_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB X 8.36815e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_18 VNB N_VGND_c_290_n 0.00682667f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_VGND_c_291_n 0.0104867f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_20 VNB N_VGND_c_292_n 0.0352669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_293_n 0.0368289f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_22 VNB N_VGND_c_294_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_23 VNB N_VGND_c_295_n 0.0221765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_296_n 0.179269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_A_M1001_g 0.042732f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=2.065
cc_26 VPB A 0.0328541f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_27 VPB A 5.58177e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_28 VPB N_A_c_56_n 0.0111383f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_29 VPB N_A_c_57_n 8.01089e-19 $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.325
cc_30 VPB N_B_M1006_g 0.0392113f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=2.065
cc_31 VPB B 0.00190522f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_B_c_90_n 0.00651062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_61_75#_M1003_g 0.021594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_61_75#_M1005_g 0.0265767f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_35 VPB N_A_61_75#_c_126_n 5.21437e-19 $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.53
cc_36 VPB N_A_61_75#_c_127_n 0.00746182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_61_75#_c_128_n 0.00141902f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.2
cc_38 VPB N_A_61_75#_c_138_n 0.00415653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_61_75#_c_139_n 0.00331457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_61_75#_c_140_n 0.00448261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_61_75#_c_132_n 2.80626e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_61_75#_c_142_n 0.00176402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_220_n 0.0307635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_221_n 0.00720315f $X=-0.19 $Y=1.305 $X2=0.465 $Y2=1.16
cc_45 VPB N_VPWR_c_222_n 0.0104612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_223_n 0.0447066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_224_n 0.0112126f $X=-0.19 $Y=1.305 $X2=0.465 $Y2=1.2
cc_48 VPB N_VPWR_c_225_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.2
cc_49 VPB N_VPWR_c_226_n 0.0195533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_227_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.2
cc_51 VPB N_VPWR_c_228_n 0.0202916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_219_n 0.0621771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB X 0.00121874f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_54 N_A_M1002_g N_B_M1000_g 0.0284572f $X=0.66 $Y=0.585 $X2=0 $Y2=0
cc_55 N_A_M1001_g N_B_M1006_g 0.0284572f $X=0.66 $Y=2.065 $X2=0 $Y2=0
cc_56 A B 0.0167054f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_57 N_A_c_56_n B 2.9595e-19 $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_58 A N_B_c_90_n 0.00173558f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_c_56_n N_B_c_90_n 0.0284572f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_A_61_75#_c_129_n 0.00746013f $X=0.66 $Y=0.585 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_A_61_75#_c_130_n 0.00872515f $X=0.66 $Y=0.585 $X2=0 $Y2=0
cc_62 A N_A_61_75#_c_130_n 0.0115462f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_M1002_g N_A_61_75#_c_131_n 0.00477732f $X=0.66 $Y=0.585 $X2=0 $Y2=0
cc_64 A N_A_61_75#_c_131_n 0.0173113f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_c_56_n N_A_61_75#_c_131_n 0.00725489f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_57_n N_A_61_75#_c_131_n 0.0101632f $X=0.242 $Y=1.325 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_A_61_75#_c_138_n 0.00326606f $X=0.66 $Y=2.065 $X2=0 $Y2=0
cc_68 A N_A_61_75#_c_138_n 0.00100172f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_69 N_A_M1001_g N_A_61_75#_c_140_n 0.00212665f $X=0.66 $Y=2.065 $X2=0 $Y2=0
cc_70 A N_A_61_75#_c_140_n 0.00854343f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_71 A N_A_61_75#_c_140_n 0.00266042f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_72 N_A_M1001_g N_VPWR_c_220_n 0.00517304f $X=0.66 $Y=2.065 $X2=0 $Y2=0
cc_73 A N_VPWR_c_220_n 0.00927177f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_74 A N_VPWR_c_220_n 0.00406435f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_56_n N_VPWR_c_220_n 0.00292944f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VPWR_c_226_n 0.00523993f $X=0.66 $Y=2.065 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_VPWR_c_219_n 0.00519019f $X=0.66 $Y=2.065 $X2=0 $Y2=0
cc_78 N_A_M1002_g N_VGND_c_293_n 0.00441396f $X=0.66 $Y=0.585 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_VGND_c_296_n 0.00541051f $X=0.66 $Y=0.585 $X2=0 $Y2=0
cc_80 N_B_M1000_g N_A_61_75#_c_124_n 0.0169053f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_81 N_B_M1006_g N_A_61_75#_M1003_g 0.0208394f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_82 B N_A_61_75#_c_126_n 2.848e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B_c_90_n N_A_61_75#_c_126_n 0.0207079f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B_M1000_g N_A_61_75#_c_129_n 0.00142377f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_85 N_B_M1000_g N_A_61_75#_c_130_n 0.0132517f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_86 B N_A_61_75#_c_130_n 0.0239051f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B_c_90_n N_A_61_75#_c_130_n 0.00445184f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B_M1006_g N_A_61_75#_c_138_n 0.0101531f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_89 N_B_M1006_g N_A_61_75#_c_139_n 0.011503f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_90 B N_A_61_75#_c_139_n 0.0159296f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_91 N_B_c_90_n N_A_61_75#_c_139_n 0.00116352f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B_M1006_g N_A_61_75#_c_140_n 0.00290243f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_93 B N_A_61_75#_c_140_n 0.00167894f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B_M1000_g N_A_61_75#_c_132_n 0.00157912f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_95 B N_A_61_75#_c_132_n 0.0196812f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B_c_90_n N_A_61_75#_c_132_n 0.0032101f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_M1006_g N_A_61_75#_c_142_n 0.00306f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_98 N_B_M1006_g N_VPWR_c_221_n 0.00636578f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_99 N_B_M1006_g N_VPWR_c_226_n 0.0049636f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_100 N_B_M1006_g N_VPWR_c_219_n 0.00519019f $X=1.08 $Y=2.065 $X2=0 $Y2=0
cc_101 N_B_M1000_g N_VGND_c_290_n 0.00547641f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_102 N_B_M1000_g N_VGND_c_293_n 0.0044865f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_103 N_B_M1000_g N_VGND_c_296_n 0.00541051f $X=1.08 $Y=0.585 $X2=0 $Y2=0
cc_104 N_A_61_75#_c_139_n N_VPWR_M1006_d 0.00735159f $X=1.505 $Y=1.66 $X2=0
+ $Y2=0
cc_105 N_A_61_75#_c_138_n N_VPWR_c_220_n 0.0142628f $X=0.87 $Y=2.13 $X2=0 $Y2=0
cc_106 N_A_61_75#_M1003_g N_VPWR_c_221_n 0.0128908f $X=1.62 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_61_75#_M1005_g N_VPWR_c_221_n 9.31703e-19 $X=2.16 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_61_75#_c_138_n N_VPWR_c_221_n 0.0249299f $X=0.87 $Y=2.13 $X2=0 $Y2=0
cc_109 N_A_61_75#_c_139_n N_VPWR_c_221_n 0.0221013f $X=1.505 $Y=1.66 $X2=0 $Y2=0
cc_110 N_A_61_75#_M1005_g N_VPWR_c_223_n 0.0237337f $X=2.16 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_61_75#_c_138_n N_VPWR_c_226_n 0.0101858f $X=0.87 $Y=2.13 $X2=0 $Y2=0
cc_112 N_A_61_75#_M1003_g N_VPWR_c_228_n 0.0046653f $X=1.62 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_61_75#_M1005_g N_VPWR_c_228_n 0.00389548f $X=2.16 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_61_75#_M1003_g N_VPWR_c_219_n 0.00826408f $X=1.62 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_61_75#_M1005_g N_VPWR_c_219_n 0.00738543f $X=2.16 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_61_75#_c_138_n N_VPWR_c_219_n 0.0103957f $X=0.87 $Y=2.13 $X2=0 $Y2=0
cc_117 N_A_61_75#_c_124_n N_X_c_260_n 0.00391418f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_61_75#_c_127_n N_X_c_260_n 0.00508761f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_61_75#_c_132_n N_X_c_260_n 0.00393781f $X=1.59 $Y=1.325 $X2=0 $Y2=0
cc_120 N_A_61_75#_c_124_n X 0.00532502f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_61_75#_M1003_g X 0.00640518f $X=1.62 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_61_75#_c_125_n X 0.0154728f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_61_75#_M1005_g X 0.0201807f $X=2.16 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_61_75#_c_127_n X 0.00954132f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_61_75#_c_128_n X 0.0166906f $X=2.16 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_61_75#_c_139_n X 0.00909018f $X=1.505 $Y=1.66 $X2=0 $Y2=0
cc_127 N_A_61_75#_c_132_n X 0.0387851f $X=1.59 $Y=1.325 $X2=0 $Y2=0
cc_128 N_A_61_75#_c_142_n X 0.0122272f $X=1.59 $Y=1.575 $X2=0 $Y2=0
cc_129 N_A_61_75#_M1003_g X 0.00503626f $X=1.62 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_61_75#_M1005_g X 0.0107168f $X=2.16 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_61_75#_c_127_n X 0.0047852f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_61_75#_c_132_n X 8.88144e-19 $X=1.59 $Y=1.325 $X2=0 $Y2=0
cc_133 N_A_61_75#_c_125_n N_X_c_276_n 0.01069f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_61_75#_c_130_n A_147_75# 0.00297727f $X=1.505 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_61_75#_c_130_n N_VGND_M1000_d 0.0034258f $X=1.505 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_61_75#_c_124_n N_VGND_c_290_n 0.0044954f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_61_75#_c_129_n N_VGND_c_290_n 0.00513858f $X=0.45 $Y=0.52 $X2=0 $Y2=0
cc_138 N_A_61_75#_c_130_n N_VGND_c_290_n 0.0190303f $X=1.505 $Y=0.81 $X2=0 $Y2=0
cc_139 N_A_61_75#_c_125_n N_VGND_c_292_n 0.0169809f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_61_75#_c_129_n N_VGND_c_293_n 0.0140625f $X=0.45 $Y=0.52 $X2=0 $Y2=0
cc_141 N_A_61_75#_c_130_n N_VGND_c_293_n 0.00788124f $X=1.505 $Y=0.81 $X2=0
+ $Y2=0
cc_142 N_A_61_75#_c_124_n N_VGND_c_295_n 0.00420655f $X=1.62 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_61_75#_c_125_n N_VGND_c_295_n 0.0038803f $X=2.16 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_61_75#_c_132_n N_VGND_c_295_n 0.00212733f $X=1.59 $Y=1.325 $X2=0
+ $Y2=0
cc_145 N_A_61_75#_c_124_n N_VGND_c_296_n 0.0073152f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_61_75#_c_125_n N_VGND_c_296_n 0.00739831f $X=2.16 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_61_75#_c_129_n N_VGND_c_296_n 0.011857f $X=0.45 $Y=0.52 $X2=0 $Y2=0
cc_148 N_A_61_75#_c_130_n N_VGND_c_296_n 0.0178101f $X=1.505 $Y=0.81 $X2=0 $Y2=0
cc_149 N_A_61_75#_c_132_n N_VGND_c_296_n 0.00390104f $X=1.59 $Y=1.325 $X2=0
+ $Y2=0
cc_150 N_VPWR_c_219_n N_X_M1003_d 0.00558844f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_151 N_VPWR_c_223_n X 0.074864f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_152 N_VPWR_c_221_n X 0.0401469f $X=1.41 $Y=2 $X2=0 $Y2=0
cc_153 N_VPWR_c_228_n X 0.0289942f $X=2.385 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_219_n X 0.0165488f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_223_n N_VGND_c_292_n 0.0101475f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_156 X N_VGND_c_292_n 0.0255649f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_157 N_X_c_276_n N_VGND_c_292_n 0.0232886f $X=2.09 $Y=0.545 $X2=0 $Y2=0
cc_158 N_X_c_260_n N_VGND_c_295_n 0.0178654f $X=1.965 $Y=0.4 $X2=0 $Y2=0
cc_159 N_X_c_276_n N_VGND_c_295_n 0.015316f $X=2.09 $Y=0.545 $X2=0 $Y2=0
cc_160 N_X_M1004_s N_VGND_c_296_n 0.00312389f $X=1.695 $Y=0.235 $X2=0 $Y2=0
cc_161 N_X_c_260_n N_VGND_c_296_n 0.011094f $X=1.965 $Y=0.4 $X2=0 $Y2=0
cc_162 N_X_c_276_n N_VGND_c_296_n 0.00903344f $X=2.09 $Y=0.545 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dlclkp_4.spice.SKY130_FD_SC_HD__DLCLKP_4.pxi
* Created: Thu Aug 27 14:16:32 2020
* 
x_PM_SKY130_FD_SC_HD__DLCLKP_4%CLK N_CLK_c_175_n N_CLK_c_164_n N_CLK_M1022_g
+ N_CLK_c_176_n N_CLK_M1010_g N_CLK_M1008_g N_CLK_c_165_n N_CLK_M1018_g
+ N_CLK_c_166_n N_CLK_c_178_n CLK CLK N_CLK_c_168_n N_CLK_c_169_n N_CLK_c_170_n
+ N_CLK_c_171_n N_CLK_c_172_n N_CLK_c_173_n N_CLK_c_174_n
+ PM_SKY130_FD_SC_HD__DLCLKP_4%CLK
x_PM_SKY130_FD_SC_HD__DLCLKP_4%A_27_47# N_A_27_47#_M1022_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1011_g N_A_27_47#_M1000_g N_A_27_47#_M1025_g N_A_27_47#_M1012_g
+ N_A_27_47#_c_296_n N_A_27_47#_c_297_n N_A_27_47#_c_298_n N_A_27_47#_c_308_n
+ N_A_27_47#_c_309_n N_A_27_47#_c_310_n N_A_27_47#_c_299_n N_A_27_47#_c_312_n
+ N_A_27_47#_c_300_n N_A_27_47#_c_301_n N_A_27_47#_c_302_n N_A_27_47#_c_303_n
+ N_A_27_47#_c_314_n N_A_27_47#_c_315_n N_A_27_47#_c_316_n N_A_27_47#_c_317_n
+ N_A_27_47#_c_304_n N_A_27_47#_c_305_n N_A_27_47#_c_319_n N_A_27_47#_c_320_n
+ PM_SKY130_FD_SC_HD__DLCLKP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__DLCLKP_4%GATE N_GATE_c_486_n N_GATE_M1005_g N_GATE_c_487_n
+ N_GATE_M1014_g GATE N_GATE_c_489_n PM_SKY130_FD_SC_HD__DLCLKP_4%GATE
x_PM_SKY130_FD_SC_HD__DLCLKP_4%A_193_47# N_A_193_47#_M1011_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1006_g N_A_193_47#_c_530_n N_A_193_47#_c_531_n
+ N_A_193_47#_M1003_g N_A_193_47#_c_537_n N_A_193_47#_c_533_n
+ N_A_193_47#_c_539_n N_A_193_47#_c_540_n N_A_193_47#_c_541_n
+ N_A_193_47#_c_542_n N_A_193_47#_c_543_n PM_SKY130_FD_SC_HD__DLCLKP_4%A_193_47#
x_PM_SKY130_FD_SC_HD__DLCLKP_4%A_627_153# N_A_627_153#_M1007_s
+ N_A_627_153#_M1017_s N_A_627_153#_c_626_n N_A_627_153#_M1016_g
+ N_A_627_153#_M1009_g N_A_627_153#_c_627_n N_A_627_153#_M1024_g
+ N_A_627_153#_c_628_n N_A_627_153#_c_629_n N_A_627_153#_M1020_g
+ N_A_627_153#_c_630_n N_A_627_153#_c_631_n N_A_627_153#_c_638_n
+ N_A_627_153#_c_639_n N_A_627_153#_c_690_p N_A_627_153#_c_632_n
+ N_A_627_153#_c_640_n N_A_627_153#_c_633_n N_A_627_153#_c_652_n
+ N_A_627_153#_c_653_n N_A_627_153#_c_654_n
+ PM_SKY130_FD_SC_HD__DLCLKP_4%A_627_153#
x_PM_SKY130_FD_SC_HD__DLCLKP_4%A_477_413# N_A_477_413#_M1025_d
+ N_A_477_413#_M1006_d N_A_477_413#_M1017_g N_A_477_413#_c_733_n
+ N_A_477_413#_M1007_g N_A_477_413#_c_734_n N_A_477_413#_c_735_n
+ N_A_477_413#_c_745_n N_A_477_413#_c_751_n N_A_477_413#_c_736_n
+ N_A_477_413#_c_742_n N_A_477_413#_c_737_n N_A_477_413#_c_738_n
+ PM_SKY130_FD_SC_HD__DLCLKP_4%A_477_413#
x_PM_SKY130_FD_SC_HD__DLCLKP_4%A_953_297# N_A_953_297#_M1020_s
+ N_A_953_297#_M1024_d N_A_953_297#_c_825_n N_A_953_297#_M1004_g
+ N_A_953_297#_M1001_g N_A_953_297#_c_826_n N_A_953_297#_M1013_g
+ N_A_953_297#_M1002_g N_A_953_297#_c_827_n N_A_953_297#_M1021_g
+ N_A_953_297#_M1015_g N_A_953_297#_c_828_n N_A_953_297#_M1023_g
+ N_A_953_297#_M1019_g N_A_953_297#_c_829_n N_A_953_297#_c_830_n
+ N_A_953_297#_c_831_n N_A_953_297#_c_832_n N_A_953_297#_c_850_n
+ N_A_953_297#_c_833_n N_A_953_297#_c_855_n N_A_953_297#_c_860_n
+ N_A_953_297#_c_834_n N_A_953_297#_c_845_n N_A_953_297#_c_917_p
+ N_A_953_297#_c_835_n N_A_953_297#_c_870_n N_A_953_297#_c_836_n
+ PM_SKY130_FD_SC_HD__DLCLKP_4%A_953_297#
x_PM_SKY130_FD_SC_HD__DLCLKP_4%VPWR N_VPWR_M1010_d N_VPWR_M1014_s N_VPWR_M1016_d
+ N_VPWR_M1017_d N_VPWR_M1008_d N_VPWR_M1002_s N_VPWR_M1019_s N_VPWR_c_979_n
+ N_VPWR_c_980_n N_VPWR_c_981_n N_VPWR_c_982_n N_VPWR_c_983_n N_VPWR_c_984_n
+ N_VPWR_c_985_n N_VPWR_c_986_n N_VPWR_c_987_n VPWR N_VPWR_c_988_n
+ N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n
+ N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n N_VPWR_c_997_n N_VPWR_c_998_n
+ N_VPWR_c_999_n N_VPWR_c_978_n PM_SKY130_FD_SC_HD__DLCLKP_4%VPWR
x_PM_SKY130_FD_SC_HD__DLCLKP_4%GCLK N_GCLK_M1004_s N_GCLK_M1021_s N_GCLK_M1001_d
+ N_GCLK_M1015_d N_GCLK_c_1115_n N_GCLK_c_1118_n N_GCLK_c_1111_n N_GCLK_c_1125_n
+ N_GCLK_c_1128_n N_GCLK_c_1134_n GCLK GCLK GCLK GCLK GCLK GCLK
+ PM_SKY130_FD_SC_HD__DLCLKP_4%GCLK
x_PM_SKY130_FD_SC_HD__DLCLKP_4%VGND N_VGND_M1022_d N_VGND_M1005_s N_VGND_M1009_d
+ N_VGND_M1007_d N_VGND_M1018_d N_VGND_M1013_d N_VGND_M1023_d N_VGND_c_1188_n
+ N_VGND_c_1189_n N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n
+ N_VGND_c_1193_n N_VGND_c_1194_n N_VGND_c_1195_n N_VGND_c_1196_n
+ N_VGND_c_1197_n VGND N_VGND_c_1198_n N_VGND_c_1199_n N_VGND_c_1200_n
+ N_VGND_c_1201_n N_VGND_c_1202_n N_VGND_c_1203_n N_VGND_c_1204_n
+ N_VGND_c_1205_n N_VGND_c_1206_n N_VGND_c_1207_n N_VGND_c_1208_n
+ N_VGND_c_1209_n PM_SKY130_FD_SC_HD__DLCLKP_4%VGND
cc_1 VNB N_CLK_c_164_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_165_n 0.0159758f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=0.995
cc_3 VNB N_CLK_c_166_n 0.0230896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_4 VNB CLK 0.00750589f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_CLK_c_168_n 0.0420287f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=1.19
cc_6 VNB N_CLK_c_169_n 0.00981446f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_7 VNB N_CLK_c_170_n 3.82824e-19 $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=1.19
cc_8 VNB N_CLK_c_171_n 0.0199736f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_9 VNB N_CLK_c_172_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_10 VNB N_CLK_c_173_n 0.0214554f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=1.16
cc_11 VNB N_CLK_c_174_n 0.0046058f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=1.16
cc_12 VNB N_A_27_47#_M1011_g 0.0411064f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_13 VNB N_A_27_47#_c_296_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_14 VNB N_A_27_47#_c_297_n 0.00193692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_298_n 0.0079398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_299_n 0.00327232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_300_n 7.52483e-19 $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_18 VNB N_A_27_47#_c_301_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=1.16
cc_19 VNB N_A_27_47#_c_302_n 0.0276918f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.19
cc_20 VNB N_A_27_47#_c_303_n 0.00234664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_304_n 0.0233742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_305_n 0.0176244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_GATE_c_486_n 0.0197637f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_24 VNB N_GATE_c_487_n 0.0356574f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.59
cc_25 VNB N_GATE_M1014_g 0.0158452f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_26 VNB N_GATE_c_489_n 0.00594528f $X=-0.19 $Y=-0.24 $X2=5.515 $Y2=1.985
cc_27 VNB N_A_193_47#_c_530_n 0.0118021f $X=-0.19 $Y=-0.24 $X2=5.515 $Y2=1.325
cc_28 VNB N_A_193_47#_c_531_n 0.00846186f $X=-0.19 $Y=-0.24 $X2=5.515 $Y2=1.985
cc_29 VNB N_A_193_47#_M1003_g 0.0443062f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=0.995
cc_30 VNB N_A_193_47#_c_533_n 0.0214412f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_31 VNB N_A_627_153#_c_626_n 0.0179622f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_32 VNB N_A_627_153#_c_627_n 0.0303021f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=0.56
cc_33 VNB N_A_627_153#_c_628_n 0.0305441f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_34 VNB N_A_627_153#_c_629_n 0.0173878f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_35 VNB N_A_627_153#_c_630_n 0.0197988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_627_153#_c_631_n 0.0150294f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_37 VNB N_A_627_153#_c_632_n 0.0025547f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=1.19
cc_38 VNB N_A_627_153#_c_633_n 0.00251059f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_39 VNB N_A_477_413#_c_733_n 0.0229718f $X=-0.19 $Y=-0.24 $X2=5.515 $Y2=1.325
cc_40 VNB N_A_477_413#_c_734_n 0.0438317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_477_413#_c_735_n 0.010276f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=0.995
cc_42 VNB N_A_477_413#_c_736_n 0.00665352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_477_413#_c_737_n 0.00349849f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=1.19
cc_44 VNB N_A_477_413#_c_738_n 0.00582528f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_45 VNB N_A_953_297#_c_825_n 0.0159403f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_46 VNB N_A_953_297#_c_826_n 0.0167443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_953_297#_c_827_n 0.0150503f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_953_297#_c_828_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_953_297#_c_829_n 0.00805142f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=1.19
cc_50 VNB N_A_953_297#_c_830_n 0.0167891f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=1.19
cc_51 VNB N_A_953_297#_c_831_n 0.0544125f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_52 VNB N_A_953_297#_c_832_n 0.00462303f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_53 VNB N_A_953_297#_c_833_n 0.00335865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_953_297#_c_834_n 0.00289461f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=1.19
cc_55 VNB N_A_953_297#_c_835_n 0.00195608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_953_297#_c_836_n 0.00133619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_978_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_GCLK_c_1111_n 5.96696e-19 $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=0.56
cc_59 VNB GCLK 0.00108357f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=1.19
cc_60 VNB N_VGND_c_1188_n 4.11703e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_61 VNB N_VGND_c_1189_n 0.00634462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1190_n 0.00590734f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_63 VNB N_VGND_c_1191_n 0.0189113f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_64 VNB N_VGND_c_1192_n 0.0093552f $X=-0.19 $Y=-0.24 $X2=5.315 $Y2=1.19
cc_65 VNB N_VGND_c_1193_n 0.00231219f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_66 VNB N_VGND_c_1194_n 0.0186688f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_67 VNB N_VGND_c_1195_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=1.325
cc_68 VNB N_VGND_c_1196_n 0.0100062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1197_n 0.0336646f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_70 VNB N_VGND_c_1198_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1199_n 0.0160671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1200_n 0.0410482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1201_n 0.0263071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1202_n 0.0172948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1203_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1204_n 0.00516774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1205_n 0.00514197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1206_n 0.00548191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1207_n 0.00393404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1208_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1209_n 0.395096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VPB N_CLK_c_175_n 0.0127917f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_83 VPB N_CLK_c_176_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_84 VPB N_CLK_M1008_g 0.0228913f $X=-0.19 $Y=1.305 $X2=5.515 $Y2=1.985
cc_85 VPB N_CLK_c_178_n 0.0238508f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_86 VPB CLK 0.0127706f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_87 VPB N_CLK_c_170_n 4.41345e-19 $X=-0.19 $Y=1.305 $X2=5.315 $Y2=1.19
cc_88 VPB N_CLK_c_171_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_89 VPB N_CLK_c_173_n 0.00423052f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=1.16
cc_90 VPB N_CLK_c_174_n 0.00249584f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=1.16
cc_91 VPB N_A_27_47#_M1000_g 0.0384074f $X=-0.19 $Y=1.305 $X2=5.515 $Y2=1.985
cc_92 VPB N_A_27_47#_M1012_g 0.0209898f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_93 VPB N_A_27_47#_c_308_n 0.00104212f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=1.19
cc_94 VPB N_A_27_47#_c_309_n 0.00647333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_c_310_n 0.00379177f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=1.19
cc_96 VPB N_A_27_47#_c_299_n 0.00262797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_47#_c_312_n 0.0299799f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_98 VPB N_A_27_47#_c_300_n 7.331e-19 $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_99 VPB N_A_27_47#_c_314_n 0.00663751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_c_315_n 0.00490944f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=1.19
cc_101 VPB N_A_27_47#_c_316_n 0.00149155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_c_317_n 0.00235505f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_47#_c_304_n 0.0115913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_47#_c_319_n 0.026712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_c_320_n 0.00184933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_GATE_M1014_g 0.0450737f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_107 VPB N_A_193_47#_M1006_g 0.0309903f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_108 VPB N_A_193_47#_c_530_n 0.015594f $X=-0.19 $Y=1.305 $X2=5.515 $Y2=1.325
cc_109 VPB N_A_193_47#_c_531_n 0.00384716f $X=-0.19 $Y=1.305 $X2=5.515 $Y2=1.985
cc_110 VPB N_A_193_47#_c_537_n 0.0108232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_193_47#_c_533_n 0.00140822f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_112 VPB N_A_193_47#_c_539_n 0.0136168f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_113 VPB N_A_193_47#_c_540_n 0.00423565f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=1.19
cc_114 VPB N_A_193_47#_c_541_n 0.00243255f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_115 VPB N_A_193_47#_c_542_n 0.00958545f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_116 VPB N_A_193_47#_c_543_n 0.0143915f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_117 VPB N_A_627_153#_c_626_n 0.0155296f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_118 VPB N_A_627_153#_M1016_g 0.0241492f $X=-0.19 $Y=1.305 $X2=5.515 $Y2=1.325
cc_119 VPB N_A_627_153#_c_627_n 0.0060057f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=0.56
cc_120 VPB N_A_627_153#_M1024_g 0.0231381f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_121 VPB N_A_627_153#_c_638_n 0.00701918f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_122 VPB N_A_627_153#_c_639_n 0.0425139f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=1.19
cc_123 VPB N_A_627_153#_c_640_n 0.0037618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_627_153#_c_633_n 0.0078264f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_125 VPB N_A_477_413#_M1017_g 0.0230236f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_126 VPB N_A_477_413#_c_734_n 0.015757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_477_413#_c_735_n 0.00194612f $X=-0.19 $Y=1.305 $X2=5.575
+ $Y2=0.995
cc_128 VPB N_A_477_413#_c_742_n 0.00863041f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_129 VPB N_A_477_413#_c_737_n 0.00207403f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=1.19
cc_130 VPB N_A_953_297#_M1001_g 0.0188683f $X=-0.19 $Y=1.305 $X2=5.515 $Y2=1.985
cc_131 VPB N_A_953_297#_M1002_g 0.0191667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_953_297#_M1015_g 0.0171325f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_133 VPB N_A_953_297#_M1019_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_134 VPB N_A_953_297#_c_829_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=5.315 $Y2=1.19
cc_135 VPB N_A_953_297#_c_830_n 0.00630337f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=1.19
cc_136 VPB N_A_953_297#_c_831_n 0.00841466f $X=-0.19 $Y=1.305 $X2=0.242
+ $Y2=1.235
cc_137 VPB N_A_953_297#_c_833_n 0.004364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_953_297#_c_845_n 0.00355671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_979_n 0.00106176f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_140 VPB N_VPWR_c_980_n 0.00554306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_981_n 0.0109002f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_142 VPB N_VPWR_c_982_n 0.0170827f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_143 VPB N_VPWR_c_983_n 0.00471272f $X=-0.19 $Y=1.305 $X2=5.315 $Y2=1.19
cc_144 VPB N_VPWR_c_984_n 0.00253902f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_145 VPB N_VPWR_c_985_n 0.00179062f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=1.16
cc_146 VPB N_VPWR_c_986_n 0.00998035f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=1.325
cc_147 VPB N_VPWR_c_987_n 0.0470617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_988_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_989_n 0.0162415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_990_n 0.0385733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_991_n 0.0277693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_992_n 0.017486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_993_n 0.0172948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_994_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_995_n 0.00557046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_996_n 0.00689581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_997_n 0.00545268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_998_n 0.00391734f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_999_n 0.00366786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_978_n 0.0532154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB GCLK 0.00157056f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=1.19
cc_162 N_CLK_c_164_n N_A_27_47#_M1011_g 0.0187834f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_163 N_CLK_c_172_n N_A_27_47#_M1011_g 0.00431651f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_164 N_CLK_c_178_n N_A_27_47#_M1000_g 0.0273371f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_165 N_CLK_c_171_n N_A_27_47#_M1000_g 0.0041981f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_166 N_CLK_c_164_n N_A_27_47#_c_297_n 0.00674622f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_167 N_CLK_c_166_n N_A_27_47#_c_297_n 0.00598065f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_168 N_CLK_c_168_n N_A_27_47#_c_297_n 0.00834405f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_169 N_CLK_c_169_n N_A_27_47#_c_297_n 0.00123352f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_170 N_CLK_c_166_n N_A_27_47#_c_298_n 0.00624006f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_171 CLK N_A_27_47#_c_298_n 0.0182472f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_172 N_CLK_c_169_n N_A_27_47#_c_298_n 0.00215816f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_173 N_CLK_c_171_n N_A_27_47#_c_298_n 7.62625e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_174 N_CLK_c_176_n N_A_27_47#_c_308_n 0.0107434f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_175 N_CLK_c_178_n N_A_27_47#_c_308_n 0.00220936f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_176 N_CLK_c_168_n N_A_27_47#_c_308_n 0.00526871f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_177 N_CLK_c_169_n N_A_27_47#_c_308_n 0.00108512f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_178 N_CLK_c_175_n N_A_27_47#_c_309_n 8.2635e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_179 N_CLK_c_178_n N_A_27_47#_c_309_n 0.00424154f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_180 N_CLK_c_168_n N_A_27_47#_c_310_n 0.00535254f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_181 N_CLK_c_168_n N_A_27_47#_c_299_n 0.0160565f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_182 N_CLK_c_176_n N_A_27_47#_c_312_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_183 N_CLK_c_178_n N_A_27_47#_c_312_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_184 CLK N_A_27_47#_c_312_n 0.0209321f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_185 N_CLK_c_169_n N_A_27_47#_c_312_n 0.00163378f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_186 N_CLK_c_171_n N_A_27_47#_c_312_n 5.90345e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_187 N_CLK_c_168_n N_A_27_47#_c_300_n 0.0233715f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_188 N_CLK_c_169_n N_A_27_47#_c_300_n 0.00217745f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_189 N_CLK_c_171_n N_A_27_47#_c_300_n 0.00320724f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_190 N_CLK_c_166_n N_A_27_47#_c_301_n 0.00179331f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_191 CLK N_A_27_47#_c_301_n 0.0287909f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_192 N_CLK_c_172_n N_A_27_47#_c_301_n 0.00150073f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_193 N_CLK_c_168_n N_A_27_47#_c_302_n 0.00377901f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_194 N_CLK_c_168_n N_A_27_47#_c_303_n 0.0131311f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_195 N_CLK_c_168_n N_A_27_47#_c_314_n 0.0056514f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_196 N_CLK_c_168_n N_A_27_47#_c_315_n 0.0272158f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_197 N_CLK_c_176_n N_A_27_47#_c_316_n 0.00103212f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_198 N_CLK_c_168_n N_A_27_47#_c_316_n 0.0132354f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_199 N_CLK_c_168_n N_A_27_47#_c_317_n 0.0150153f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_200 CLK N_A_27_47#_c_304_n 9.45858e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_201 N_CLK_c_168_n N_A_27_47#_c_304_n 0.0105697f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_202 N_CLK_c_169_n N_A_27_47#_c_304_n 3.75305e-19 $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_203 N_CLK_c_171_n N_A_27_47#_c_304_n 0.0182636f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_204 N_CLK_c_168_n N_A_27_47#_c_319_n 0.00141376f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_205 N_CLK_c_168_n N_GATE_c_487_n 0.00474366f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_206 N_CLK_c_168_n N_GATE_M1014_g 0.00780604f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_207 N_CLK_c_168_n N_GATE_c_489_n 0.0119219f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_208 N_CLK_c_168_n N_A_193_47#_c_530_n 0.00432269f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_209 N_CLK_c_168_n N_A_193_47#_c_531_n 0.00408726f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_210 N_CLK_c_168_n N_A_193_47#_M1003_g 0.00278637f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_211 N_CLK_c_168_n N_A_193_47#_c_533_n 0.0317595f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_212 N_CLK_c_168_n N_A_193_47#_c_543_n 0.0348825f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_213 N_CLK_c_168_n N_A_627_153#_c_627_n 0.00430479f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_214 N_CLK_c_173_n N_A_627_153#_c_627_n 0.0026668f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_215 N_CLK_M1008_g N_A_627_153#_M1024_g 0.00911878f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_CLK_c_168_n N_A_627_153#_c_628_n 0.00602895f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_217 N_CLK_c_170_n N_A_627_153#_c_628_n 0.00156453f $X=5.315 $Y=1.19 $X2=0
+ $Y2=0
cc_218 N_CLK_c_173_n N_A_627_153#_c_628_n 0.00784212f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_219 N_CLK_c_174_n N_A_627_153#_c_628_n 4.69736e-19 $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_CLK_c_165_n N_A_627_153#_c_629_n 0.0414497f $X=5.575 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_CLK_c_168_n N_A_627_153#_c_638_n 0.00757269f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_222 N_CLK_c_168_n N_A_627_153#_c_633_n 0.055142f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_223 N_CLK_c_168_n N_A_627_153#_c_652_n 0.00178106f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_224 N_CLK_c_168_n N_A_627_153#_c_653_n 0.00219349f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_225 N_CLK_c_168_n N_A_627_153#_c_654_n 0.0221464f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_226 N_CLK_c_168_n N_A_477_413#_c_734_n 0.00630685f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_227 N_CLK_c_168_n N_A_477_413#_c_745_n 0.00427749f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_228 N_CLK_c_168_n N_A_477_413#_c_737_n 0.038028f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_229 N_CLK_c_168_n N_A_477_413#_c_738_n 0.0307629f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_230 N_CLK_c_165_n N_A_953_297#_c_825_n 0.026135f $X=5.575 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_CLK_M1008_g N_A_953_297#_M1001_g 0.0230906f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_CLK_c_173_n N_A_953_297#_c_829_n 0.0213193f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_233 N_CLK_c_174_n N_A_953_297#_c_829_n 9.26792e-19 $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_234 N_CLK_M1008_g N_A_953_297#_c_850_n 0.00908082f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_CLK_c_168_n N_A_953_297#_c_833_n 0.0186312f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_236 N_CLK_c_170_n N_A_953_297#_c_833_n 0.00259823f $X=5.315 $Y=1.19 $X2=0
+ $Y2=0
cc_237 N_CLK_c_173_n N_A_953_297#_c_833_n 0.00397818f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_238 N_CLK_c_174_n N_A_953_297#_c_833_n 0.0188569f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_239 N_CLK_c_165_n N_A_953_297#_c_855_n 0.0112703f $X=5.575 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_CLK_c_168_n N_A_953_297#_c_855_n 0.00301679f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_241 N_CLK_c_170_n N_A_953_297#_c_855_n 0.00330575f $X=5.315 $Y=1.19 $X2=0
+ $Y2=0
cc_242 N_CLK_c_173_n N_A_953_297#_c_855_n 0.00285778f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_CLK_c_174_n N_A_953_297#_c_855_n 0.030436f $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_244 N_CLK_M1008_g N_A_953_297#_c_860_n 0.0162803f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_CLK_c_168_n N_A_953_297#_c_860_n 0.0031378f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_246 N_CLK_c_170_n N_A_953_297#_c_860_n 0.00360945f $X=5.315 $Y=1.19 $X2=0
+ $Y2=0
cc_247 N_CLK_c_173_n N_A_953_297#_c_860_n 0.00280181f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_248 N_CLK_c_174_n N_A_953_297#_c_860_n 0.0324026f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_249 N_CLK_c_165_n N_A_953_297#_c_834_n 0.00209837f $X=5.575 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_CLK_c_173_n N_A_953_297#_c_834_n 0.00120633f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_251 N_CLK_M1008_g N_A_953_297#_c_845_n 0.00301185f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_252 N_CLK_c_174_n N_A_953_297#_c_845_n 0.00277809f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_253 N_CLK_c_168_n N_A_953_297#_c_835_n 0.00403531f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_254 N_CLK_c_168_n N_A_953_297#_c_870_n 0.00436956f $X=5.17 $Y=1.19 $X2=0
+ $Y2=0
cc_255 N_CLK_c_170_n N_A_953_297#_c_836_n 9.81534e-19 $X=5.315 $Y=1.19 $X2=0
+ $Y2=0
cc_256 N_CLK_c_173_n N_A_953_297#_c_836_n 8.12038e-19 $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_257 N_CLK_c_174_n N_A_953_297#_c_836_n 0.0206008f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_258 N_CLK_c_176_n N_VPWR_c_979_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_259 N_CLK_M1008_g N_VPWR_c_984_n 0.0172093f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_260 N_CLK_c_176_n N_VPWR_c_988_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_261 N_CLK_M1008_g N_VPWR_c_991_n 0.00525069f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_262 N_CLK_c_176_n N_VPWR_c_978_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_263 N_CLK_M1008_g N_VPWR_c_978_n 0.00965336f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_264 N_CLK_c_164_n N_VGND_c_1188_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_265 N_CLK_c_168_n N_VGND_c_1190_n 0.00215049f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_266 N_CLK_c_168_n N_VGND_c_1192_n 0.00188524f $X=5.17 $Y=1.19 $X2=0 $Y2=0
cc_267 N_CLK_c_165_n N_VGND_c_1193_n 0.0123579f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_268 N_CLK_c_164_n N_VGND_c_1198_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_269 N_CLK_c_166_n N_VGND_c_1198_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_270 N_CLK_c_165_n N_VGND_c_1201_n 0.00261107f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_271 N_CLK_c_164_n N_VGND_c_1209_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_272 N_CLK_c_165_n N_VGND_c_1209_n 0.00330124f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_302_n N_GATE_c_486_n 0.00236006f $X=2.38 $Y=0.87 $X2=-0.19
+ $Y2=-0.24
cc_274 N_A_27_47#_c_303_n N_GATE_c_486_n 3.20776e-19 $X=2.65 $Y=0.87 $X2=-0.19
+ $Y2=-0.24
cc_275 N_A_27_47#_c_305_n N_GATE_c_486_n 0.020383f $X=2.377 $Y=0.705 $X2=-0.19
+ $Y2=-0.24
cc_276 N_A_27_47#_M1011_g N_GATE_c_487_n 0.00345305f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_299_n N_GATE_c_487_n 0.00142118f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_302_n N_GATE_c_487_n 0.0113978f $X=2.38 $Y=0.87 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_303_n N_GATE_c_487_n 4.15796e-19 $X=2.65 $Y=0.87 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_310_n N_GATE_M1014_g 0.0134231f $X=2.505 $Y=1.94 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_299_n N_GATE_M1014_g 0.00229046f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_317_n N_GATE_M1014_g 0.00292531f $X=1.61 $Y=1.87 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_320_n N_GATE_M1014_g 0.00227553f $X=1.695 $Y=1.905 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_302_n N_GATE_c_489_n 9.65794e-19 $X=2.38 $Y=0.87 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_303_n N_GATE_c_489_n 0.0111894f $X=2.65 $Y=0.87 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_315_n N_A_193_47#_M1000_d 6.81311e-19 $X=1.465 $Y=1.87 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1012_g N_A_193_47#_M1006_g 0.0156136f $X=2.85 $Y=2.275 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_310_n N_A_193_47#_M1006_g 0.0130406f $X=2.505 $Y=1.94 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_317_n N_A_193_47#_M1006_g 4.53892e-19 $X=1.61 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_310_n N_A_193_47#_c_530_n 0.00300236f $X=2.505 $Y=1.94 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_299_n N_A_193_47#_c_530_n 0.0116385f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_303_n N_A_193_47#_c_530_n 0.00167722f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_314_n N_A_193_47#_c_530_n 0.00404893f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_319_n N_A_193_47#_c_530_n 0.0188015f $X=2.85 $Y=1.74 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_302_n N_A_193_47#_c_531_n 0.0197699f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_303_n N_A_193_47#_c_531_n 0.0012352f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_299_n N_A_193_47#_M1003_g 0.00536343f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_302_n N_A_193_47#_M1003_g 0.0213151f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_303_n N_A_193_47#_M1003_g 0.0061203f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_305_n N_A_193_47#_M1003_g 0.0123755f $X=2.377 $Y=0.705 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_310_n N_A_193_47#_c_537_n 0.0028551f $X=2.505 $Y=1.94 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_314_n N_A_193_47#_c_537_n 0.00534333f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_319_n N_A_193_47#_c_537_n 0.0161493f $X=2.85 $Y=1.74 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_M1011_g N_A_193_47#_c_533_n 0.0128335f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_297_n N_A_193_47#_c_533_n 0.0103422f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_300_n N_A_193_47#_c_533_n 0.0199464f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_301_n N_A_193_47#_c_533_n 0.0163881f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_M1000_g N_A_193_47#_c_539_n 0.00572366f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_309_n N_A_193_47#_c_539_n 0.0169301f $X=0.695 $Y=1.795 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_315_n N_A_193_47#_c_539_n 0.020099f $X=1.465 $Y=1.87 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_316_n N_A_193_47#_c_539_n 0.00243787f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_317_n N_A_193_47#_c_539_n 0.00316769f $X=1.61 $Y=1.87 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_320_n N_A_193_47#_c_539_n 0.0104976f $X=1.695 $Y=1.905 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_309_n N_A_193_47#_c_540_n 0.0124004f $X=0.695 $Y=1.795 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_300_n N_A_193_47#_c_540_n 0.00358828f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_315_n N_A_193_47#_c_540_n 0.00141747f $X=1.465 $Y=1.87 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_304_n N_A_193_47#_c_540_n 0.00563154f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_310_n N_A_193_47#_c_541_n 0.0210469f $X=2.505 $Y=1.94 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_299_n N_A_193_47#_c_541_n 0.0136802f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_302_n N_A_193_47#_c_541_n 4.30953e-19 $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_303_n N_A_193_47#_c_541_n 0.00114094f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_314_n N_A_193_47#_c_541_n 0.00870241f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_299_n N_A_193_47#_c_542_n 0.00390791f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_310_n N_A_193_47#_c_543_n 0.0142612f $X=2.505 $Y=1.94 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_315_n N_A_193_47#_c_543_n 0.00541768f $X=1.465 $Y=1.87 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_317_n N_A_193_47#_c_543_n 0.00375439f $X=1.61 $Y=1.87 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_320_n N_A_193_47#_c_543_n 0.00969245f $X=1.695 $Y=1.905
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_c_299_n N_A_627_153#_c_626_n 0.00126551f $X=2.65 $Y=1.575
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_M1012_g N_A_627_153#_M1016_g 0.0318529f $X=2.85 $Y=2.275 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_314_n N_A_627_153#_c_639_n 4.25151e-19 $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_319_n N_A_627_153#_c_639_n 0.0318529f $X=2.85 $Y=1.74 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_302_n N_A_477_413#_c_745_n 0.00155649f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_303_n N_A_477_413#_c_745_n 0.0187882f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_305_n N_A_477_413#_c_745_n 0.00406871f $X=2.377 $Y=0.705
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_M1012_g N_A_477_413#_c_751_n 0.00869878f $X=2.85 $Y=2.275
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_310_n N_A_477_413#_c_751_n 0.00214112f $X=2.505 $Y=1.94
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_314_n N_A_477_413#_c_751_n 0.0217886f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_319_n N_A_477_413#_c_751_n 8.02086e-19 $X=2.85 $Y=1.74 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_303_n N_A_477_413#_c_736_n 0.022294f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1012_g N_A_477_413#_c_742_n 0.0074049f $X=2.85 $Y=2.275 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_299_n N_A_477_413#_c_742_n 0.0129827f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_314_n N_A_477_413#_c_742_n 0.0324519f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_319_n N_A_477_413#_c_742_n 0.00260742f $X=2.85 $Y=1.74 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_299_n N_A_477_413#_c_738_n 0.0175246f $X=2.65 $Y=1.575 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_303_n N_A_477_413#_c_738_n 0.00337335f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_319_n N_A_477_413#_c_738_n 5.67091e-19 $X=2.85 $Y=1.74 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_309_n N_VPWR_M1010_d 9.46731e-19 $X=0.695 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_348 N_A_27_47#_c_316_n N_VPWR_M1010_d 0.00195102f $X=0.84 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_349 N_A_27_47#_c_317_n N_VPWR_M1014_s 2.12313e-19 $X=1.61 $Y=1.87 $X2=0 $Y2=0
cc_350 N_A_27_47#_c_320_n N_VPWR_M1014_s 0.00399334f $X=1.695 $Y=1.905 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_M1000_g N_VPWR_c_979_n 0.00836513f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_308_n N_VPWR_c_979_n 0.00355272f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_309_n N_VPWR_c_979_n 0.0110625f $X=0.695 $Y=1.795 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_312_n N_VPWR_c_979_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_316_n N_VPWR_c_979_n 0.004957f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_356 N_A_27_47#_M1000_g N_VPWR_c_980_n 0.00181768f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_315_n N_VPWR_c_980_n 2.23709e-19 $X=1.465 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_317_n N_VPWR_c_980_n 0.00216952f $X=1.61 $Y=1.87 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_320_n N_VPWR_c_980_n 0.0165661f $X=1.695 $Y=1.905 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_308_n N_VPWR_c_988_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_361 N_A_27_47#_c_312_n N_VPWR_c_988_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_362 N_A_27_47#_M1000_g N_VPWR_c_989_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_M1012_g N_VPWR_c_990_n 0.00366098f $X=2.85 $Y=2.275 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_310_n N_VPWR_c_990_n 0.00961689f $X=2.505 $Y=1.94 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_M1000_g N_VPWR_c_978_n 0.00536257f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_M1012_g N_VPWR_c_978_n 0.00544966f $X=2.85 $Y=2.275 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_308_n N_VPWR_c_978_n 0.00396423f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_310_n N_VPWR_c_978_n 0.0167351f $X=2.505 $Y=1.94 $X2=0 $Y2=0
cc_369 N_A_27_47#_c_312_n N_VPWR_c_978_n 0.00993215f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_370 N_A_27_47#_c_315_n N_VPWR_c_978_n 0.0310249f $X=1.465 $Y=1.87 $X2=0 $Y2=0
cc_371 N_A_27_47#_c_316_n N_VPWR_c_978_n 0.0144759f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_372 N_A_27_47#_c_317_n N_VPWR_c_978_n 0.0134286f $X=1.61 $Y=1.87 $X2=0 $Y2=0
cc_373 N_A_27_47#_c_320_n N_VPWR_c_978_n 7.69579e-19 $X=1.695 $Y=1.905 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_310_n A_381_369# 0.00573055f $X=2.505 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_375 N_A_27_47#_c_297_n N_VGND_M1022_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_376 N_A_27_47#_M1011_g N_VGND_c_1188_n 0.00843828f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_297_n N_VGND_c_1188_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_378 N_A_27_47#_c_300_n N_VGND_c_1188_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_304_n N_VGND_c_1188_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_M1011_g N_VGND_c_1189_n 0.00294417f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_305_n N_VGND_c_1189_n 0.00181317f $X=2.377 $Y=0.705 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_296_n N_VGND_c_1198_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_297_n N_VGND_c_1198_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1011_g N_VGND_c_1199_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_302_n N_VGND_c_1200_n 9.43262e-19 $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_303_n N_VGND_c_1200_n 0.00182549f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_305_n N_VGND_c_1200_n 0.00425892f $X=2.377 $Y=0.705 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1022_s N_VGND_c_1209_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1011_g N_VGND_c_1209_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_296_n N_VGND_c_1209_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_297_n N_VGND_c_1209_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_302_n N_VGND_c_1209_n 0.00121904f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_303_n N_VGND_c_1209_n 0.00340834f $X=2.65 $Y=0.87 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_305_n N_VGND_c_1209_n 0.0062921f $X=2.377 $Y=0.705 $X2=0
+ $Y2=0
cc_395 N_GATE_M1014_g N_A_193_47#_M1006_g 0.0355592f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_396 N_GATE_M1014_g N_A_193_47#_c_531_n 0.0286757f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_397 N_GATE_c_486_n N_A_193_47#_c_533_n 0.00636812f $X=1.83 $Y=0.76 $X2=0
+ $Y2=0
cc_398 N_GATE_c_487_n N_A_193_47#_c_533_n 0.00281139f $X=1.83 $Y=1.095 $X2=0
+ $Y2=0
cc_399 N_GATE_M1014_g N_A_193_47#_c_533_n 0.00539787f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_400 N_GATE_c_489_n N_A_193_47#_c_533_n 0.0158678f $X=1.785 $Y=0.93 $X2=0
+ $Y2=0
cc_401 N_GATE_M1014_g N_A_193_47#_c_539_n 0.00918545f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_402 N_GATE_M1014_g N_A_193_47#_c_541_n 0.0022816f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_403 N_GATE_c_487_n N_A_193_47#_c_543_n 0.00397996f $X=1.83 $Y=1.095 $X2=0
+ $Y2=0
cc_404 N_GATE_M1014_g N_A_193_47#_c_543_n 0.0162219f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_405 N_GATE_c_489_n N_A_193_47#_c_543_n 0.0101132f $X=1.785 $Y=0.93 $X2=0
+ $Y2=0
cc_406 N_GATE_c_486_n N_A_477_413#_c_745_n 6.24923e-19 $X=1.83 $Y=0.76 $X2=0
+ $Y2=0
cc_407 N_GATE_M1014_g N_VPWR_c_980_n 0.014031f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_408 N_GATE_M1014_g N_VPWR_c_990_n 0.00259464f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_409 N_GATE_M1014_g N_VPWR_c_978_n 0.00341715f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_410 N_GATE_c_486_n N_VGND_c_1189_n 0.0111586f $X=1.83 $Y=0.76 $X2=0 $Y2=0
cc_411 N_GATE_c_487_n N_VGND_c_1189_n 0.00269535f $X=1.83 $Y=1.095 $X2=0 $Y2=0
cc_412 N_GATE_c_489_n N_VGND_c_1189_n 0.0104173f $X=1.785 $Y=0.93 $X2=0 $Y2=0
cc_413 N_GATE_c_486_n N_VGND_c_1200_n 0.0046653f $X=1.83 $Y=0.76 $X2=0 $Y2=0
cc_414 N_GATE_c_487_n N_VGND_c_1200_n 7.88437e-19 $X=1.83 $Y=1.095 $X2=0 $Y2=0
cc_415 N_GATE_c_486_n N_VGND_c_1209_n 0.00454097f $X=1.83 $Y=0.76 $X2=0 $Y2=0
cc_416 N_GATE_c_487_n N_VGND_c_1209_n 0.0010595f $X=1.83 $Y=1.095 $X2=0 $Y2=0
cc_417 N_GATE_c_489_n N_VGND_c_1209_n 0.00638637f $X=1.785 $Y=0.93 $X2=0 $Y2=0
cc_418 N_A_193_47#_c_530_n N_A_627_153#_c_626_n 0.0142848f $X=2.725 $Y=1.32
+ $X2=0 $Y2=0
cc_419 N_A_193_47#_M1003_g N_A_627_153#_c_630_n 0.0227352f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_420 N_A_193_47#_M1003_g N_A_627_153#_c_631_n 0.0142848f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_421 N_A_193_47#_M1003_g N_A_477_413#_c_745_n 0.0093694f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_422 N_A_193_47#_M1006_g N_A_477_413#_c_751_n 0.00376268f $X=2.31 $Y=2.275
+ $X2=0 $Y2=0
cc_423 N_A_193_47#_M1003_g N_A_477_413#_c_736_n 0.00517821f $X=2.8 $Y=0.415
+ $X2=0 $Y2=0
cc_424 N_A_193_47#_M1006_g N_A_477_413#_c_742_n 9.17726e-19 $X=2.31 $Y=2.275
+ $X2=0 $Y2=0
cc_425 N_A_193_47#_c_530_n N_A_477_413#_c_742_n 5.84404e-19 $X=2.725 $Y=1.32
+ $X2=0 $Y2=0
cc_426 N_A_193_47#_M1003_g N_A_477_413#_c_738_n 0.0025885f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_427 N_A_193_47#_c_539_n N_VPWR_c_979_n 0.0127357f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_428 N_A_193_47#_M1006_g N_VPWR_c_980_n 0.00210053f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_429 N_A_193_47#_c_539_n N_VPWR_c_980_n 0.0189906f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_430 N_A_193_47#_c_543_n N_VPWR_c_980_n 9.77038e-19 $X=2.045 $Y=1.52 $X2=0
+ $Y2=0
cc_431 N_A_193_47#_c_539_n N_VPWR_c_989_n 0.015988f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_432 N_A_193_47#_M1006_g N_VPWR_c_990_n 0.00433717f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_433 N_A_193_47#_M1006_g N_VPWR_c_978_n 0.0065033f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_434 N_A_193_47#_c_539_n N_VPWR_c_978_n 0.00409094f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_435 N_A_193_47#_c_533_n N_VGND_c_1189_n 0.00984039f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_436 N_A_193_47#_M1003_g N_VGND_c_1190_n 0.00174741f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_437 N_A_193_47#_c_533_n N_VGND_c_1199_n 0.0116097f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_438 N_A_193_47#_M1003_g N_VGND_c_1200_n 0.0037981f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_439 N_A_193_47#_M1011_d N_VGND_c_1209_n 0.00394021f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_440 N_A_193_47#_M1003_g N_VGND_c_1209_n 0.00557191f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_441 N_A_193_47#_c_533_n N_VGND_c_1209_n 0.0096527f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_442 N_A_627_153#_M1024_g N_A_477_413#_M1017_g 0.033816f $X=4.69 $Y=1.985
+ $X2=0 $Y2=0
cc_443 N_A_627_153#_c_639_n N_A_477_413#_M1017_g 0.00300925f $X=3.44 $Y=1.7
+ $X2=0 $Y2=0
cc_444 N_A_627_153#_c_640_n N_A_477_413#_M1017_g 0.00755466f $X=4.03 $Y=1.535
+ $X2=0 $Y2=0
cc_445 N_A_627_153#_c_653_n N_A_477_413#_M1017_g 5.32092e-19 $X=3.98 $Y=1.755
+ $X2=0 $Y2=0
cc_446 N_A_627_153#_c_627_n N_A_477_413#_c_733_n 0.00137152f $X=4.69 $Y=1.325
+ $X2=0 $Y2=0
cc_447 N_A_627_153#_c_632_n N_A_477_413#_c_733_n 0.00653044f $X=4.03 $Y=0.995
+ $X2=0 $Y2=0
cc_448 N_A_627_153#_c_626_n N_A_477_413#_c_734_n 0.015703f $X=3.21 $Y=1.535
+ $X2=0 $Y2=0
cc_449 N_A_627_153#_c_638_n N_A_477_413#_c_734_n 0.00914525f $X=3.895 $Y=1.7
+ $X2=0 $Y2=0
cc_450 N_A_627_153#_c_639_n N_A_477_413#_c_734_n 0.00121881f $X=3.44 $Y=1.7
+ $X2=0 $Y2=0
cc_451 N_A_627_153#_c_652_n N_A_477_413#_c_734_n 0.00182108f $X=4.005 $Y=0.58
+ $X2=0 $Y2=0
cc_452 N_A_627_153#_c_653_n N_A_477_413#_c_734_n 0.00212837f $X=3.98 $Y=1.755
+ $X2=0 $Y2=0
cc_453 N_A_627_153#_c_654_n N_A_477_413#_c_734_n 0.0169836f $X=4.03 $Y=1.16
+ $X2=0 $Y2=0
cc_454 N_A_627_153#_c_627_n N_A_477_413#_c_735_n 0.0215424f $X=4.69 $Y=1.325
+ $X2=0 $Y2=0
cc_455 N_A_627_153#_c_633_n N_A_477_413#_c_735_n 0.0245944f $X=4.635 $Y=1.16
+ $X2=0 $Y2=0
cc_456 N_A_627_153#_c_630_n N_A_477_413#_c_745_n 0.0015738f $X=3.242 $Y=0.765
+ $X2=0 $Y2=0
cc_457 N_A_627_153#_c_630_n N_A_477_413#_c_736_n 0.00512255f $X=3.242 $Y=0.765
+ $X2=0 $Y2=0
cc_458 N_A_627_153#_c_631_n N_A_477_413#_c_736_n 0.00542003f $X=3.242 $Y=0.915
+ $X2=0 $Y2=0
cc_459 N_A_627_153#_c_626_n N_A_477_413#_c_742_n 0.0115626f $X=3.21 $Y=1.535
+ $X2=0 $Y2=0
cc_460 N_A_627_153#_M1016_g N_A_477_413#_c_742_n 0.0208289f $X=3.21 $Y=2.275
+ $X2=0 $Y2=0
cc_461 N_A_627_153#_c_638_n N_A_477_413#_c_742_n 0.0249855f $X=3.895 $Y=1.7
+ $X2=0 $Y2=0
cc_462 N_A_627_153#_c_639_n N_A_477_413#_c_742_n 0.00843184f $X=3.44 $Y=1.7
+ $X2=0 $Y2=0
cc_463 N_A_627_153#_c_626_n N_A_477_413#_c_737_n 0.0161482f $X=3.21 $Y=1.535
+ $X2=0 $Y2=0
cc_464 N_A_627_153#_c_631_n N_A_477_413#_c_737_n 0.00165871f $X=3.242 $Y=0.915
+ $X2=0 $Y2=0
cc_465 N_A_627_153#_c_638_n N_A_477_413#_c_737_n 0.0253052f $X=3.895 $Y=1.7
+ $X2=0 $Y2=0
cc_466 N_A_627_153#_c_639_n N_A_477_413#_c_737_n 0.00644091f $X=3.44 $Y=1.7
+ $X2=0 $Y2=0
cc_467 N_A_627_153#_c_654_n N_A_477_413#_c_737_n 0.0252269f $X=4.03 $Y=1.16
+ $X2=0 $Y2=0
cc_468 N_A_627_153#_c_626_n N_A_477_413#_c_738_n 0.00631844f $X=3.21 $Y=1.535
+ $X2=0 $Y2=0
cc_469 N_A_627_153#_M1024_g N_A_953_297#_c_850_n 0.0109082f $X=4.69 $Y=1.985
+ $X2=0 $Y2=0
cc_470 N_A_627_153#_c_690_p N_A_953_297#_c_850_n 0.00306488f $X=3.98 $Y=2.27
+ $X2=0 $Y2=0
cc_471 N_A_627_153#_c_653_n N_A_953_297#_c_850_n 0.00614796f $X=3.98 $Y=1.755
+ $X2=0 $Y2=0
cc_472 N_A_627_153#_c_627_n N_A_953_297#_c_833_n 0.00206342f $X=4.69 $Y=1.325
+ $X2=0 $Y2=0
cc_473 N_A_627_153#_M1024_g N_A_953_297#_c_833_n 0.00427897f $X=4.69 $Y=1.985
+ $X2=0 $Y2=0
cc_474 N_A_627_153#_c_628_n N_A_953_297#_c_833_n 0.0146284f $X=5.08 $Y=1.035
+ $X2=0 $Y2=0
cc_475 N_A_627_153#_c_629_n N_A_953_297#_c_833_n 0.00298516f $X=5.155 $Y=0.96
+ $X2=0 $Y2=0
cc_476 N_A_627_153#_c_633_n N_A_953_297#_c_833_n 0.0238732f $X=4.635 $Y=1.16
+ $X2=0 $Y2=0
cc_477 N_A_627_153#_c_629_n N_A_953_297#_c_855_n 0.0142076f $X=5.155 $Y=0.96
+ $X2=0 $Y2=0
cc_478 N_A_627_153#_c_628_n N_A_953_297#_c_860_n 0.00342326f $X=5.08 $Y=1.035
+ $X2=0 $Y2=0
cc_479 N_A_627_153#_c_627_n N_A_953_297#_c_835_n 0.00395943f $X=4.69 $Y=1.325
+ $X2=0 $Y2=0
cc_480 N_A_627_153#_M1024_g N_A_953_297#_c_870_n 0.0035298f $X=4.69 $Y=1.985
+ $X2=0 $Y2=0
cc_481 N_A_627_153#_c_628_n N_A_953_297#_c_870_n 0.00206525f $X=5.08 $Y=1.035
+ $X2=0 $Y2=0
cc_482 N_A_627_153#_c_653_n N_A_953_297#_c_870_n 0.00412506f $X=3.98 $Y=1.755
+ $X2=0 $Y2=0
cc_483 N_A_627_153#_M1016_g N_VPWR_c_981_n 0.00460314f $X=3.21 $Y=2.275 $X2=0
+ $Y2=0
cc_484 N_A_627_153#_c_638_n N_VPWR_c_981_n 0.0167948f $X=3.895 $Y=1.7 $X2=0
+ $Y2=0
cc_485 N_A_627_153#_c_639_n N_VPWR_c_981_n 0.00529157f $X=3.44 $Y=1.7 $X2=0
+ $Y2=0
cc_486 N_A_627_153#_c_690_p N_VPWR_c_981_n 0.018486f $X=3.98 $Y=2.27 $X2=0 $Y2=0
cc_487 N_A_627_153#_c_690_p N_VPWR_c_982_n 0.0112378f $X=3.98 $Y=2.27 $X2=0
+ $Y2=0
cc_488 N_A_627_153#_c_627_n N_VPWR_c_983_n 0.00176757f $X=4.69 $Y=1.325 $X2=0
+ $Y2=0
cc_489 N_A_627_153#_M1024_g N_VPWR_c_983_n 0.00556318f $X=4.69 $Y=1.985 $X2=0
+ $Y2=0
cc_490 N_A_627_153#_M1016_g N_VPWR_c_990_n 0.00519775f $X=3.21 $Y=2.275 $X2=0
+ $Y2=0
cc_491 N_A_627_153#_M1024_g N_VPWR_c_991_n 0.00564131f $X=4.69 $Y=1.985 $X2=0
+ $Y2=0
cc_492 N_A_627_153#_M1017_s N_VPWR_c_978_n 0.0023739f $X=3.855 $Y=1.485 $X2=0
+ $Y2=0
cc_493 N_A_627_153#_M1016_g N_VPWR_c_978_n 0.0100344f $X=3.21 $Y=2.275 $X2=0
+ $Y2=0
cc_494 N_A_627_153#_M1024_g N_VPWR_c_978_n 0.0110498f $X=4.69 $Y=1.985 $X2=0
+ $Y2=0
cc_495 N_A_627_153#_c_638_n N_VPWR_c_978_n 0.0086096f $X=3.895 $Y=1.7 $X2=0
+ $Y2=0
cc_496 N_A_627_153#_c_639_n N_VPWR_c_978_n 0.00110429f $X=3.44 $Y=1.7 $X2=0
+ $Y2=0
cc_497 N_A_627_153#_c_690_p N_VPWR_c_978_n 0.00827281f $X=3.98 $Y=2.27 $X2=0
+ $Y2=0
cc_498 N_A_627_153#_c_630_n N_VGND_c_1190_n 0.0117279f $X=3.242 $Y=0.765 $X2=0
+ $Y2=0
cc_499 N_A_627_153#_c_652_n N_VGND_c_1190_n 0.00703504f $X=4.005 $Y=0.58 $X2=0
+ $Y2=0
cc_500 N_A_627_153#_c_652_n N_VGND_c_1191_n 0.00690212f $X=4.005 $Y=0.58 $X2=0
+ $Y2=0
cc_501 N_A_627_153#_c_627_n N_VGND_c_1192_n 0.00172952f $X=4.69 $Y=1.325 $X2=0
+ $Y2=0
cc_502 N_A_627_153#_c_629_n N_VGND_c_1192_n 0.00361458f $X=5.155 $Y=0.96 $X2=0
+ $Y2=0
cc_503 N_A_627_153#_c_633_n N_VGND_c_1192_n 0.0135094f $X=4.635 $Y=1.16 $X2=0
+ $Y2=0
cc_504 N_A_627_153#_c_629_n N_VGND_c_1193_n 0.00218204f $X=5.155 $Y=0.96 $X2=0
+ $Y2=0
cc_505 N_A_627_153#_c_630_n N_VGND_c_1200_n 0.00447018f $X=3.242 $Y=0.765 $X2=0
+ $Y2=0
cc_506 N_A_627_153#_c_631_n N_VGND_c_1200_n 0.00129035f $X=3.242 $Y=0.915 $X2=0
+ $Y2=0
cc_507 N_A_627_153#_c_629_n N_VGND_c_1201_n 0.00436487f $X=5.155 $Y=0.96 $X2=0
+ $Y2=0
cc_508 N_A_627_153#_M1007_s N_VGND_c_1209_n 0.00375142f $X=3.88 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_627_153#_c_629_n N_VGND_c_1209_n 0.00747881f $X=5.155 $Y=0.96 $X2=0
+ $Y2=0
cc_510 N_A_627_153#_c_630_n N_VGND_c_1209_n 0.00782321f $X=3.242 $Y=0.765 $X2=0
+ $Y2=0
cc_511 N_A_627_153#_c_631_n N_VGND_c_1209_n 0.0017268f $X=3.242 $Y=0.915 $X2=0
+ $Y2=0
cc_512 N_A_627_153#_c_652_n N_VGND_c_1209_n 0.00761394f $X=4.005 $Y=0.58 $X2=0
+ $Y2=0
cc_513 N_A_477_413#_M1017_g N_A_953_297#_c_850_n 0.00115681f $X=4.19 $Y=1.985
+ $X2=0 $Y2=0
cc_514 N_A_477_413#_c_733_n N_A_953_297#_c_833_n 0.001765f $X=4.215 $Y=0.995
+ $X2=0 $Y2=0
cc_515 N_A_477_413#_c_733_n N_A_953_297#_c_835_n 0.00358276f $X=4.215 $Y=0.995
+ $X2=0 $Y2=0
cc_516 N_A_477_413#_M1017_g N_A_953_297#_c_870_n 5.16476e-19 $X=4.19 $Y=1.985
+ $X2=0 $Y2=0
cc_517 N_A_477_413#_c_751_n N_VPWR_c_980_n 0.00644392f $X=2.915 $Y=2.31 $X2=0
+ $Y2=0
cc_518 N_A_477_413#_M1017_g N_VPWR_c_981_n 0.00249422f $X=4.19 $Y=1.985 $X2=0
+ $Y2=0
cc_519 N_A_477_413#_M1017_g N_VPWR_c_982_n 0.00585385f $X=4.19 $Y=1.985 $X2=0
+ $Y2=0
cc_520 N_A_477_413#_M1017_g N_VPWR_c_983_n 0.00210243f $X=4.19 $Y=1.985 $X2=0
+ $Y2=0
cc_521 N_A_477_413#_c_751_n N_VPWR_c_990_n 0.0210957f $X=2.915 $Y=2.31 $X2=0
+ $Y2=0
cc_522 N_A_477_413#_c_742_n N_VPWR_c_990_n 0.011081f $X=3.1 $Y=2.015 $X2=0 $Y2=0
cc_523 N_A_477_413#_M1006_d N_VPWR_c_978_n 0.00356601f $X=2.385 $Y=2.065 $X2=0
+ $Y2=0
cc_524 N_A_477_413#_M1017_g N_VPWR_c_978_n 0.012235f $X=4.19 $Y=1.985 $X2=0
+ $Y2=0
cc_525 N_A_477_413#_c_751_n N_VPWR_c_978_n 0.0154439f $X=2.915 $Y=2.31 $X2=0
+ $Y2=0
cc_526 N_A_477_413#_c_742_n N_VPWR_c_978_n 0.0096884f $X=3.1 $Y=2.015 $X2=0
+ $Y2=0
cc_527 N_A_477_413#_c_742_n A_585_413# 0.00101795f $X=3.1 $Y=2.015 $X2=-0.19
+ $Y2=-0.24
cc_528 N_A_477_413#_c_745_n N_VGND_c_1189_n 0.00264829f $X=2.905 $Y=0.45 $X2=0
+ $Y2=0
cc_529 N_A_477_413#_c_733_n N_VGND_c_1190_n 0.00419493f $X=4.215 $Y=0.995 $X2=0
+ $Y2=0
cc_530 N_A_477_413#_c_734_n N_VGND_c_1190_n 0.00179389f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_531 N_A_477_413#_c_745_n N_VGND_c_1190_n 0.0104349f $X=2.905 $Y=0.45 $X2=0
+ $Y2=0
cc_532 N_A_477_413#_c_737_n N_VGND_c_1190_n 0.0103619f $X=3.69 $Y=1.16 $X2=0
+ $Y2=0
cc_533 N_A_477_413#_c_733_n N_VGND_c_1191_n 0.00585385f $X=4.215 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_A_477_413#_c_733_n N_VGND_c_1192_n 0.0053182f $X=4.215 $Y=0.995 $X2=0
+ $Y2=0
cc_535 N_A_477_413#_c_745_n N_VGND_c_1200_n 0.0221422f $X=2.905 $Y=0.45 $X2=0
+ $Y2=0
cc_536 N_A_477_413#_M1025_d N_VGND_c_1209_n 0.00242229f $X=2.44 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_A_477_413#_c_733_n N_VGND_c_1209_n 0.0133299f $X=4.215 $Y=0.995 $X2=0
+ $Y2=0
cc_538 N_A_477_413#_c_745_n N_VGND_c_1209_n 0.0222941f $X=2.905 $Y=0.45 $X2=0
+ $Y2=0
cc_539 N_A_477_413#_c_745_n A_575_47# 0.00355017f $X=2.905 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_540 N_A_477_413#_c_736_n A_575_47# 0.00146881f $X=2.99 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_541 N_A_953_297#_c_860_n N_VPWR_M1008_d 0.00612881f $X=5.91 $Y=1.58 $X2=0
+ $Y2=0
cc_542 N_A_953_297#_M1001_g N_VPWR_c_984_n 0.00541497f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_543 N_A_953_297#_c_850_n N_VPWR_c_984_n 0.0193231f $X=4.95 $Y=2.3 $X2=0 $Y2=0
cc_544 N_A_953_297#_c_860_n N_VPWR_c_984_n 0.0166452f $X=5.91 $Y=1.58 $X2=0
+ $Y2=0
cc_545 N_A_953_297#_M1001_g N_VPWR_c_985_n 9.98731e-19 $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_546 N_A_953_297#_M1002_g N_VPWR_c_985_n 0.00909783f $X=6.505 $Y=1.985 $X2=0
+ $Y2=0
cc_547 N_A_953_297#_M1015_g N_VPWR_c_985_n 0.00151876f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_548 N_A_953_297#_M1019_g N_VPWR_c_987_n 0.00322031f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_549 N_A_953_297#_c_850_n N_VPWR_c_991_n 0.0178522f $X=4.95 $Y=2.3 $X2=0 $Y2=0
cc_550 N_A_953_297#_M1001_g N_VPWR_c_992_n 0.00541763f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_551 N_A_953_297#_M1002_g N_VPWR_c_992_n 0.00319306f $X=6.505 $Y=1.985 $X2=0
+ $Y2=0
cc_552 N_A_953_297#_M1015_g N_VPWR_c_993_n 0.00422131f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_553 N_A_953_297#_M1019_g N_VPWR_c_993_n 0.00541359f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_554 N_A_953_297#_M1024_d N_VPWR_c_978_n 0.0195597f $X=4.765 $Y=1.485 $X2=0
+ $Y2=0
cc_555 N_A_953_297#_M1001_g N_VPWR_c_978_n 0.00996513f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_556 N_A_953_297#_M1002_g N_VPWR_c_978_n 0.00407575f $X=6.505 $Y=1.985 $X2=0
+ $Y2=0
cc_557 N_A_953_297#_M1015_g N_VPWR_c_978_n 0.00569458f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_558 N_A_953_297#_M1019_g N_VPWR_c_978_n 0.0104605f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_559 N_A_953_297#_c_850_n N_VPWR_c_978_n 0.0107624f $X=4.95 $Y=2.3 $X2=0 $Y2=0
cc_560 N_A_953_297#_c_860_n N_GCLK_M1001_d 0.00281912f $X=5.91 $Y=1.58 $X2=0
+ $Y2=0
cc_561 N_A_953_297#_c_825_n N_GCLK_c_1115_n 0.00315572f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_A_953_297#_c_826_n N_GCLK_c_1115_n 0.00462854f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_563 N_A_953_297#_c_827_n N_GCLK_c_1115_n 4.36062e-19 $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_564 N_A_953_297#_c_826_n N_GCLK_c_1118_n 0.00844123f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_565 N_A_953_297#_c_831_n N_GCLK_c_1118_n 0.00318912f $X=7.345 $Y=1.16 $X2=0
+ $Y2=0
cc_566 N_A_953_297#_c_917_p N_GCLK_c_1118_n 0.00830729f $X=6.415 $Y=1.16 $X2=0
+ $Y2=0
cc_567 N_A_953_297#_c_825_n N_GCLK_c_1111_n 6.38332e-19 $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_568 N_A_953_297#_c_826_n N_GCLK_c_1111_n 0.0024004f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_569 N_A_953_297#_c_830_n N_GCLK_c_1111_n 0.00122612f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_570 N_A_953_297#_c_917_p N_GCLK_c_1111_n 0.0105553f $X=6.415 $Y=1.16 $X2=0
+ $Y2=0
cc_571 N_A_953_297#_c_826_n N_GCLK_c_1125_n 5.19281e-19 $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_572 N_A_953_297#_c_827_n N_GCLK_c_1125_n 0.00618985f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_573 N_A_953_297#_c_828_n N_GCLK_c_1125_n 0.00528656f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_574 N_A_953_297#_c_825_n N_GCLK_c_1128_n 0.00367156f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_575 N_A_953_297#_c_826_n N_GCLK_c_1128_n 0.00759403f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_576 N_A_953_297#_c_830_n N_GCLK_c_1128_n 0.0024765f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_577 N_A_953_297#_c_855_n N_GCLK_c_1128_n 0.00223888f $X=5.91 $Y=0.8 $X2=0
+ $Y2=0
cc_578 N_A_953_297#_c_917_p N_GCLK_c_1128_n 0.00480939f $X=6.415 $Y=1.16 $X2=0
+ $Y2=0
cc_579 N_A_953_297#_c_836_n N_GCLK_c_1128_n 5.63789e-19 $X=6.025 $Y=1.172 $X2=0
+ $Y2=0
cc_580 N_A_953_297#_M1001_g N_GCLK_c_1134_n 0.004721f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_581 N_A_953_297#_c_830_n N_GCLK_c_1134_n 0.00336509f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_582 N_A_953_297#_c_860_n N_GCLK_c_1134_n 0.00363279f $X=5.91 $Y=1.58 $X2=0
+ $Y2=0
cc_583 N_A_953_297#_c_917_p N_GCLK_c_1134_n 0.00741015f $X=6.415 $Y=1.16 $X2=0
+ $Y2=0
cc_584 N_A_953_297#_M1001_g GCLK 0.00638255f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_585 N_A_953_297#_M1002_g GCLK 0.00481144f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_586 N_A_953_297#_M1002_g GCLK 0.0124661f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_587 N_A_953_297#_M1015_g GCLK 0.00818783f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_588 N_A_953_297#_M1019_g GCLK 0.00241889f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_589 N_A_953_297#_c_831_n GCLK 0.00228188f $X=7.345 $Y=1.16 $X2=0 $Y2=0
cc_590 N_A_953_297#_c_917_p GCLK 0.00481708f $X=6.415 $Y=1.16 $X2=0 $Y2=0
cc_591 N_A_953_297#_c_826_n GCLK 0.00132182f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_592 N_A_953_297#_M1002_g GCLK 0.00713368f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_593 N_A_953_297#_c_827_n GCLK 0.0107211f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_594 N_A_953_297#_M1015_g GCLK 0.0109427f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_595 N_A_953_297#_c_828_n GCLK 0.0081063f $X=7.345 $Y=0.995 $X2=0 $Y2=0
cc_596 N_A_953_297#_M1019_g GCLK 0.012448f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_597 N_A_953_297#_c_831_n GCLK 0.0423903f $X=7.345 $Y=1.16 $X2=0 $Y2=0
cc_598 N_A_953_297#_c_860_n GCLK 0.00572583f $X=5.91 $Y=1.58 $X2=0 $Y2=0
cc_599 N_A_953_297#_c_834_n GCLK 0.00514489f $X=6.015 $Y=1.055 $X2=0 $Y2=0
cc_600 N_A_953_297#_c_845_n GCLK 0.00670136f $X=6.025 $Y=1.495 $X2=0 $Y2=0
cc_601 N_A_953_297#_c_917_p GCLK 0.0192907f $X=6.415 $Y=1.16 $X2=0 $Y2=0
cc_602 N_A_953_297#_M1002_g GCLK 4.53016e-19 $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_603 N_A_953_297#_M1015_g GCLK 0.0064464f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_604 N_A_953_297#_M1019_g GCLK 0.00528656f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_605 N_A_953_297#_c_855_n N_VGND_M1018_d 0.00426075f $X=5.91 $Y=0.8 $X2=0
+ $Y2=0
cc_606 N_A_953_297#_c_832_n N_VGND_c_1192_n 0.0347929f $X=4.945 $Y=0.455 $X2=0
+ $Y2=0
cc_607 N_A_953_297#_c_825_n N_VGND_c_1193_n 0.00282934f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_608 N_A_953_297#_c_855_n N_VGND_c_1193_n 0.0164498f $X=5.91 $Y=0.8 $X2=0
+ $Y2=0
cc_609 N_A_953_297#_c_825_n N_VGND_c_1194_n 0.00420655f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_610 N_A_953_297#_c_826_n N_VGND_c_1194_n 0.00420765f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_611 N_A_953_297#_c_855_n N_VGND_c_1194_n 0.00188806f $X=5.91 $Y=0.8 $X2=0
+ $Y2=0
cc_612 N_A_953_297#_c_826_n N_VGND_c_1195_n 0.00268723f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_613 N_A_953_297#_c_827_n N_VGND_c_1195_n 0.00146448f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_614 N_A_953_297#_c_828_n N_VGND_c_1197_n 0.00322031f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_615 N_A_953_297#_c_832_n N_VGND_c_1201_n 0.0166184f $X=4.945 $Y=0.455 $X2=0
+ $Y2=0
cc_616 N_A_953_297#_c_855_n N_VGND_c_1201_n 0.00664634f $X=5.91 $Y=0.8 $X2=0
+ $Y2=0
cc_617 N_A_953_297#_c_827_n N_VGND_c_1202_n 0.00422131f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_618 N_A_953_297#_c_828_n N_VGND_c_1202_n 0.00541359f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_619 N_A_953_297#_M1020_s N_VGND_c_1209_n 0.00220649f $X=4.82 $Y=0.235 $X2=0
+ $Y2=0
cc_620 N_A_953_297#_c_825_n N_VGND_c_1209_n 0.00595102f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_621 N_A_953_297#_c_826_n N_VGND_c_1209_n 0.00596406f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_622 N_A_953_297#_c_827_n N_VGND_c_1209_n 0.00569458f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_623 N_A_953_297#_c_828_n N_VGND_c_1209_n 0.0104605f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_624 N_A_953_297#_c_832_n N_VGND_c_1209_n 0.0116214f $X=4.945 $Y=0.455 $X2=0
+ $Y2=0
cc_625 N_A_953_297#_c_855_n N_VGND_c_1209_n 0.0182519f $X=5.91 $Y=0.8 $X2=0
+ $Y2=0
cc_626 N_A_953_297#_c_855_n A_1046_47# 0.0044541f $X=5.91 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_627 N_VPWR_c_978_n A_381_369# 0.00416708f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_628 N_VPWR_c_978_n A_585_413# 0.00170448f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_629 N_VPWR_c_978_n N_GCLK_M1001_d 0.00316777f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_630 N_VPWR_c_978_n N_GCLK_M1015_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_631 N_VPWR_c_984_n N_GCLK_c_1134_n 0.0119478f $X=5.755 $Y=2 $X2=0 $Y2=0
cc_632 N_VPWR_c_984_n GCLK 0.0302744f $X=5.755 $Y=2 $X2=0 $Y2=0
cc_633 N_VPWR_c_985_n GCLK 0.021358f $X=6.715 $Y=2.34 $X2=0 $Y2=0
cc_634 N_VPWR_c_992_n GCLK 0.0196063f $X=6.54 $Y=2.72 $X2=0 $Y2=0
cc_635 N_VPWR_c_978_n GCLK 0.0123353f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_636 N_VPWR_M1002_s GCLK 0.00415786f $X=6.58 $Y=1.485 $X2=0 $Y2=0
cc_637 N_VPWR_c_985_n GCLK 0.0155388f $X=6.715 $Y=2.34 $X2=0 $Y2=0
cc_638 N_VPWR_c_992_n GCLK 0.00197418f $X=6.54 $Y=2.72 $X2=0 $Y2=0
cc_639 N_VPWR_c_993_n GCLK 0.00219911f $X=7.47 $Y=2.72 $X2=0 $Y2=0
cc_640 N_VPWR_c_978_n GCLK 0.00918168f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_641 N_VPWR_M1002_s GCLK 0.00426184f $X=6.58 $Y=1.485 $X2=0 $Y2=0
cc_642 N_VPWR_c_993_n GCLK 0.0189039f $X=7.47 $Y=2.72 $X2=0 $Y2=0
cc_643 N_VPWR_c_978_n GCLK 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_644 N_VPWR_c_987_n N_VGND_c_1197_n 0.00917978f $X=7.555 $Y=1.66 $X2=0 $Y2=0
cc_645 N_GCLK_c_1118_n N_VGND_M1013_d 0.00330466f $X=6.75 $Y=0.8 $X2=0 $Y2=0
cc_646 GCLK N_VGND_M1013_d 4.63659e-19 $X=7.045 $Y=0.765 $X2=0 $Y2=0
cc_647 N_GCLK_c_1118_n N_VGND_c_1194_n 0.0020257f $X=6.75 $Y=0.8 $X2=0 $Y2=0
cc_648 N_GCLK_c_1128_n N_VGND_c_1194_n 0.0239883f $X=6.375 $Y=0.4 $X2=0 $Y2=0
cc_649 N_GCLK_c_1118_n N_VGND_c_1195_n 0.0087883f $X=6.75 $Y=0.8 $X2=0 $Y2=0
cc_650 GCLK N_VGND_c_1195_n 0.00370896f $X=7.045 $Y=0.765 $X2=0 $Y2=0
cc_651 N_GCLK_c_1125_n N_VGND_c_1202_n 0.0189039f $X=7.135 $Y=0.38 $X2=0 $Y2=0
cc_652 GCLK N_VGND_c_1202_n 0.00219911f $X=7.045 $Y=0.765 $X2=0 $Y2=0
cc_653 N_GCLK_M1004_s N_VGND_c_1209_n 0.00288308f $X=6.07 $Y=0.235 $X2=0 $Y2=0
cc_654 N_GCLK_M1021_s N_VGND_c_1209_n 0.00215201f $X=7 $Y=0.235 $X2=0 $Y2=0
cc_655 N_GCLK_c_1118_n N_VGND_c_1209_n 0.00434076f $X=6.75 $Y=0.8 $X2=0 $Y2=0
cc_656 N_GCLK_c_1125_n N_VGND_c_1209_n 0.0122217f $X=7.135 $Y=0.38 $X2=0 $Y2=0
cc_657 N_GCLK_c_1128_n N_VGND_c_1209_n 0.015484f $X=6.375 $Y=0.4 $X2=0 $Y2=0
cc_658 GCLK N_VGND_c_1209_n 0.00438298f $X=7.045 $Y=0.765 $X2=0 $Y2=0
cc_659 N_VGND_c_1209_n A_381_47# 0.0139761f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_660 N_VGND_c_1209_n A_575_47# 0.00554895f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_661 N_VGND_c_1209_n A_1046_47# 0.00348377f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24

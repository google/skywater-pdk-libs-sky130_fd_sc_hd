# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.790000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 0.305000 9.575000 0.820000 ;
        RECT 9.230000 1.505000 9.575000 2.395000 ;
        RECT 9.405000 0.820000 9.575000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.530000 1.055000 3.990000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.635000 3.250000 0.785000 ;
        RECT 1.760000 0.785000 1.990000 0.835000 ;
        RECT 1.760000 0.835000 1.930000 1.685000 ;
        RECT 1.870000 0.615000 3.250000 0.635000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.065000 0.785000 3.250000 1.095000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.810000 0.805000 ;
      RECT 0.180000  1.795000 0.845000 1.965000 ;
      RECT 0.180000  1.965000 0.350000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.520000  2.135000 0.850000 2.635000 ;
      RECT 0.615000  0.805000 0.810000 0.970000 ;
      RECT 0.615000  0.970000 0.845000 1.795000 ;
      RECT 1.015000  0.345000 1.230000 0.715000 ;
      RECT 1.020000  0.715000 1.230000 2.465000 ;
      RECT 1.420000  0.260000 1.790000 0.465000 ;
      RECT 1.420000  0.465000 1.590000 1.860000 ;
      RECT 1.420000  1.860000 3.220000 2.075000 ;
      RECT 1.420000  2.075000 1.710000 2.445000 ;
      RECT 1.880000  2.245000 2.210000 2.635000 ;
      RECT 1.960000  0.085000 2.305000 0.445000 ;
      RECT 2.115000  0.960000 2.460000 1.130000 ;
      RECT 2.115000  1.130000 2.290000 1.860000 ;
      RECT 2.690000  2.245000 3.560000 2.415000 ;
      RECT 2.820000  0.275000 3.590000 0.445000 ;
      RECT 3.050000  1.305000 3.270000 1.635000 ;
      RECT 3.050000  1.635000 3.220000 1.860000 ;
      RECT 3.390000  1.825000 4.350000 1.995000 ;
      RECT 3.390000  1.995000 3.560000 2.245000 ;
      RECT 3.420000  0.445000 3.590000 0.715000 ;
      RECT 3.420000  0.715000 4.350000 0.885000 ;
      RECT 3.730000  2.165000 3.925000 2.635000 ;
      RECT 3.760000  0.085000 3.960000 0.545000 ;
      RECT 4.180000  0.285000 4.460000 0.615000 ;
      RECT 4.180000  0.615000 4.350000 0.715000 ;
      RECT 4.180000  0.885000 4.350000 1.825000 ;
      RECT 4.180000  1.995000 4.350000 2.065000 ;
      RECT 4.180000  2.065000 4.420000 2.440000 ;
      RECT 4.520000  0.780000 5.100000 1.035000 ;
      RECT 4.520000  1.035000 4.760000 1.905000 ;
      RECT 4.630000  0.705000 5.100000 0.780000 ;
      RECT 4.660000  2.190000 5.730000 2.360000 ;
      RECT 4.700000  0.365000 5.440000 0.535000 ;
      RECT 4.950000  1.655000 5.390000 2.010000 ;
      RECT 5.270000  0.535000 5.440000 1.315000 ;
      RECT 5.270000  1.315000 6.070000 1.485000 ;
      RECT 5.560000  1.485000 6.070000 1.575000 ;
      RECT 5.560000  1.575000 5.730000 2.190000 ;
      RECT 5.610000  0.765000 6.410000 1.065000 ;
      RECT 5.610000  1.065000 5.780000 1.095000 ;
      RECT 5.690000  0.085000 6.060000 0.585000 ;
      RECT 5.900000  1.245000 6.070000 1.315000 ;
      RECT 5.900000  1.835000 6.070000 2.635000 ;
      RECT 6.240000  0.365000 6.700000 0.535000 ;
      RECT 6.240000  0.535000 6.410000 0.765000 ;
      RECT 6.240000  1.065000 6.410000 2.135000 ;
      RECT 6.240000  2.135000 6.490000 2.465000 ;
      RECT 6.580000  0.705000 7.130000 1.035000 ;
      RECT 6.580000  1.245000 6.770000 1.965000 ;
      RECT 6.715000  2.165000 7.600000 2.335000 ;
      RECT 6.930000  0.365000 7.470000 0.535000 ;
      RECT 6.940000  1.035000 7.130000 1.575000 ;
      RECT 6.940000  1.575000 7.260000 1.905000 ;
      RECT 7.300000  0.535000 7.470000 0.995000 ;
      RECT 7.300000  0.995000 8.365000 1.325000 ;
      RECT 7.300000  1.325000 7.600000 1.405000 ;
      RECT 7.430000  1.405000 7.600000 2.165000 ;
      RECT 7.715000  0.085000 8.085000 0.615000 ;
      RECT 7.770000  1.575000 8.705000 1.905000 ;
      RECT 7.790000  2.135000 8.095000 2.635000 ;
      RECT 8.355000  0.300000 8.705000 0.825000 ;
      RECT 8.435000  1.905000 8.705000 2.455000 ;
      RECT 8.535000  0.825000 8.705000 0.995000 ;
      RECT 8.535000  0.995000 9.235000 1.325000 ;
      RECT 8.535000  1.325000 8.705000 1.575000 ;
      RECT 8.875000  0.085000 9.045000 0.695000 ;
      RECT 8.875000  1.625000 9.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.640000  1.785000 0.810000 1.955000 ;
      RECT 1.040000  0.765000 1.210000 0.935000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.590000  1.785000 6.760000 1.955000 ;
      RECT 6.630000  0.765000 6.800000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.580000 1.755000 0.870000 1.800000 ;
      RECT 0.580000 1.800000 6.820000 1.940000 ;
      RECT 0.580000 1.940000 0.870000 1.985000 ;
      RECT 0.980000 0.735000 1.270000 0.780000 ;
      RECT 0.980000 0.780000 6.860000 0.920000 ;
      RECT 0.980000 0.920000 1.270000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.530000 1.755000 6.820000 1.800000 ;
      RECT 6.530000 1.940000 6.820000 1.985000 ;
      RECT 6.570000 0.735000 6.860000 0.780000 ;
      RECT 6.570000 0.920000 6.860000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxtp_1
END LIBRARY

* File: sky130_fd_sc_hd__o41ai_1.pex.spice
* Created: Thu Aug 27 14:42:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O41AI_1%B1 3 7 9 15
r26 12 15 40.336 $w=2.9e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r27 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r28 5 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r29 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r30 1 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r31 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%A4 3 7 9 10 11 12 23 37
c37 9 0 2.46038e-19 $X=1.07 $Y=1.105
r38 37 38 2.0058 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=1.155 $Y2=1.245
r39 21 23 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.155 $Y=1.16
+ $X2=1.245 $Y2=1.16
r40 18 21 58.876 $w=2.7e-07 $l=2.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.155 $Y2=1.16
r41 11 12 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=1.87
+ $X2=1.167 $Y2=2.21
r42 10 11 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=1.53
+ $X2=1.167 $Y2=1.87
r43 9 37 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.155 $Y=1.16 $X2=1.155
+ $Y2=1.19
r44 9 10 10.202 $w=3.03e-07 $l=2.7e-07 $layer=LI1_cond $X=1.167 $Y=1.26
+ $X2=1.167 $Y2=1.53
r45 9 38 0.566775 $w=3.03e-07 $l=1.5e-08 $layer=LI1_cond $X=1.167 $Y=1.26
+ $X2=1.167 $Y2=1.245
r46 9 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.16 $X2=1.155 $Y2=1.16
r47 5 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.245 $Y=1.025
+ $X2=1.245 $Y2=1.16
r48 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.245 $Y=1.025
+ $X2=1.245 $Y2=0.56
r49 1 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r50 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295 $X2=0.89
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%A3 1 3 6 8 9 10 11 18 32
c39 18 0 1.18336e-19 $X=1.665 $Y=1.16
r40 32 33 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.665 $Y=1.19
+ $X2=1.665 $Y2=1.245
r41 10 11 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.66 $Y=1.87
+ $X2=1.66 $Y2=2.21
r42 9 10 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.66 $Y=1.53 $X2=1.66
+ $Y2=1.87
r43 8 32 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.665 $Y=1.16 $X2=1.665
+ $Y2=1.19
r44 8 9 9.72374 $w=3.18e-07 $l=2.7e-07 $layer=LI1_cond $X=1.66 $Y=1.26 $X2=1.66
+ $Y2=1.53
r45 8 33 0.540208 $w=3.18e-07 $l=1.5e-08 $layer=LI1_cond $X=1.66 $Y=1.26
+ $X2=1.66 $Y2=1.245
r46 8 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.16 $X2=1.665 $Y2=1.16
r47 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.325
+ $X2=1.665 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.665 $Y=1.325
+ $X2=1.665 $Y2=1.985
r49 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=0.995
+ $X2=1.665 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.665 $Y=0.995
+ $X2=1.665 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%A2 3 6 10 11 13 14 15 21 33
r41 23 33 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.16 $Y=1.585
+ $X2=2.16 $Y2=1.53
r42 14 15 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=1.87
+ $X2=2.16 $Y2=2.21
r43 13 33 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.16 $Y=1.515
+ $X2=2.16 $Y2=1.53
r44 13 31 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.515 $X2=2.16
+ $Y2=1.415
r45 13 14 9.15175 $w=3.38e-07 $l=2.7e-07 $layer=LI1_cond $X=2.16 $Y=1.6 $X2=2.16
+ $Y2=1.87
r46 13 23 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.16 $Y=1.6
+ $X2=2.16 $Y2=1.585
r47 11 22 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.16
+ $X2=2.155 $Y2=1.325
r48 11 21 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.16
+ $X2=2.155 $Y2=0.995
r49 10 31 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.165 $Y=1.16
+ $X2=2.165 $Y2=1.415
r50 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.16 $X2=2.165 $Y2=1.16
r51 6 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.085 $Y=1.985
+ $X2=2.085 $Y2=1.325
r52 3 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.085 $Y=0.56
+ $X2=2.085 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%A1 3 6 8 11 13
r26 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.16
+ $X2=2.655 $Y2=1.325
r27 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.16
+ $X2=2.655 $Y2=0.995
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.16 $X2=2.665 $Y2=1.16
r29 8 12 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=2.995 $Y=1.2
+ $X2=2.665 $Y2=1.2
r30 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.585 $Y=1.985
+ $X2=2.585 $Y2=1.325
r31 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.585 $Y=0.56
+ $X2=2.585 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%VPWR 1 2 7 9 13 15 19 21 34
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r40 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r42 25 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 24 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 22 30 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r46 22 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 21 33 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=2.72
+ $X2=2.925 $Y2=2.72
r48 21 27 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.63 $Y=2.72 $X2=2.53
+ $Y2=2.72
r49 19 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 19 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.795 $Y=1.66
+ $X2=2.795 $Y2=2.34
r52 13 33 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.795 $Y=2.635
+ $X2=2.925 $Y2=2.72
r53 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.795 $Y=2.635
+ $X2=2.795 $Y2=2.34
r54 9 12 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r55 7 30 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r56 7 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r57 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.485 $X2=2.795 $Y2=2.34
r58 2 15 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.485 $X2=2.795 $Y2=1.66
r59 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r60 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%Y 1 2 7 9 13 17 18 19 26 30
c34 30 0 1.71822e-19 $X=0.695 $Y=0.905
c35 18 0 1.35704e-19 $X=0.695 $Y=0.85
c36 7 0 1.10786e-19 $X=0.68 $Y=1.65
r37 18 30 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.82
+ $X2=0.695 $Y2=0.905
r38 18 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.695 $Y=0.92
+ $X2=0.695 $Y2=1.19
r39 18 30 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.695 $Y=0.92
+ $X2=0.695 $Y2=0.905
r40 17 26 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=0.51
+ $X2=0.255 $Y2=0.38
r41 16 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=1.485
+ $X2=0.695 $Y2=1.19
r42 14 17 7.62646 $w=3.38e-07 $l=2.25e-07 $layer=LI1_cond $X=0.255 $Y=0.735
+ $X2=0.255 $Y2=0.51
r43 13 18 8.18414 $w=3.08e-07 $l=1.85e-07 $layer=LI1_cond $X=0.425 $Y=0.82
+ $X2=0.61 $Y2=0.82
r44 13 14 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.425 $Y=0.82
+ $X2=0.255 $Y2=0.735
r45 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.66 $X2=0.68
+ $Y2=2.34
r46 7 16 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.65
+ $X2=0.68 $Y2=1.485
r47 7 9 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.68 $Y=1.65 $X2=0.68
+ $Y2=1.66
r48 2 11 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r49 2 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r50 1 26 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%A_109_47# 1 2 3 13 14 15 18 20 24 27 30
c58 1 0 1.35704e-19 $X=0.545 $Y=0.235
r59 27 29 9.16063 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.955 $Y=0.38
+ $X2=0.955 $Y2=0.565
r60 22 24 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.795 $Y=0.735
+ $X2=2.795 $Y2=0.38
r61 21 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.82
+ $X2=1.875 $Y2=0.82
r62 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.63 $Y=0.82
+ $X2=2.795 $Y2=0.735
r63 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.63 $Y=0.82 $X2=2.04
+ $Y2=0.82
r64 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.735
+ $X2=1.875 $Y2=0.82
r65 16 18 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.875 $Y=0.735
+ $X2=1.875 $Y2=0.38
r66 14 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0.82
+ $X2=1.875 $Y2=0.82
r67 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.71 $Y=0.82 $X2=1.12
+ $Y2=0.82
r68 13 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.035 $Y=0.72
+ $X2=1.035 $Y2=0.565
r69 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=0.735
+ $X2=1.12 $Y2=0.82
r70 11 13 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.035 $Y=0.735
+ $X2=1.035 $Y2=0.72
r71 3 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.66
+ $Y=0.235 $X2=2.795 $Y2=0.38
r72 2 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.74
+ $Y=0.235 $X2=1.875 $Y2=0.38
r73 1 27 182 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.955 $Y2=0.38
r74 1 13 182 $w=1.7e-07 $l=6.91195e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=1.035 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r48 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r50 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r51 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r52 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 24 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r54 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r55 21 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r56 19 31 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.07
+ $Y2=0
r57 19 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.335
+ $Y2=0
r58 18 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.99
+ $Y2=0
r59 18 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.335
+ $Y2=0
r60 16 28 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.15
+ $Y2=0
r61 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.415
+ $Y2=0
r62 15 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=2.07
+ $Y2=0
r63 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.415
+ $Y2=0
r64 11 20 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0
r65 11 13 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0.38
r66 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=0.085
+ $X2=1.415 $Y2=0
r67 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.415 $Y=0.085
+ $X2=1.415 $Y2=0.38
r68 2 13 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=2.16
+ $Y=0.235 $X2=2.375 $Y2=0.38
r69 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.32
+ $Y=0.235 $X2=1.455 $Y2=0.38
.ends


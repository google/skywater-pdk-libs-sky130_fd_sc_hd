* File: sky130_fd_sc_hd__dlxtn_4.pex.spice
* Created: Thu Aug 27 14:18:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLXTN_4%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%A_27_47# 1 2 9 13 17 20 24 28 29 30 38 42 45
+ 47 52 54 56 57 60 63 64 68 71 75 79
c167 20 0 1.41946e-19 $X=3.335 $Y=2.275
c168 13 0 2.6965e-20 $X=0.89 $Y=2.135
c169 9 0 2.6965e-20 $X=0.89 $Y=0.445
r170 64 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.095 $Y=1.53
+ $X2=3.095 $Y2=1.415
r171 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.53
+ $X2=3.015 $Y2=1.53
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r173 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=3.015 $Y2=1.53
r175 56 57 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=0.84 $Y2=1.53
r176 52 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.87
+ $X2=2.8 $Y2=0.705
r177 51 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0.87
+ $X2=3.01 $Y2=0.87
r178 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=0.87 $X2=2.8 $Y2=0.87
r179 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r180 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r181 46 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r182 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r183 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r184 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r185 39 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.335 $Y2=1.74
r186 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r187 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.53
r188 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.74
r189 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=0.87
r190 34 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.415
r191 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r192 31 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r193 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r194 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r195 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r196 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r197 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r198 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r199 18 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=1.74
r200 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=2.275
r201 17 71 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.79 $Y=0.415
+ $X2=2.79 $Y2=0.705
r202 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r203 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r204 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r206 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 32 0 1.12109e-19 $X=2.255 $Y=0.93
c84 18 0 7.13094e-20 $X=1.97 $Y=0.7
r85 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r86 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r87 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r88 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r89 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r90 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r92 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r93 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r94 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r95 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r96 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r97 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r98 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r99 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r101 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c112 38 0 1.41946e-19 $X=2.67 $Y=1.52
r113 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r114 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.612 $Y=1.87
+ $X2=2.612 $Y2=1.52
r115 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.87
+ $X2=2.555 $Y2=1.87
r116 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r117 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=2.555 $Y2=1.87
r119 26 27 1.37376 $w=1.4e-07 $l=1.11e-06 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=1.3 $Y2=1.87
r120 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r121 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r122 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r123 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r124 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r125 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r126 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.22 $Y=1.245
+ $X2=3.22 $Y2=0.415
r127 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r128 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=3.22 $Y2=1.245
r129 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=2.805 $Y2=1.32
r130 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r131 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r132 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%A_724_21# 1 2 9 13 15 17 20 22 24 27 29 31
+ 34 36 38 41 43 46 50 53 55 58 62 66 67 77
c124 29 0 1.62185e-19 $X=5.99 $Y=0.995
r125 76 77 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=5.99 $Y=1.16
+ $X2=6.43 $Y2=1.16
r126 75 76 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=5.535 $Y=1.16
+ $X2=5.99 $Y2=1.16
r127 74 75 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.115 $Y=1.16
+ $X2=5.535 $Y2=1.16
r128 62 64 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.58
+ $X2=4.495 $Y2=0.745
r129 59 74 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.1 $Y=1.16
+ $X2=5.115 $Y2=1.16
r130 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=1.16 $X2=5.1 $Y2=1.16
r131 56 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.605 $Y=1.16
+ $X2=4.52 $Y2=1.16
r132 56 58 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.605 $Y=1.16
+ $X2=5.1 $Y2=1.16
r133 55 66 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.52 $Y=1.535
+ $X2=4.495 $Y2=1.7
r134 54 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=1.325
+ $X2=4.52 $Y2=1.16
r135 54 55 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.52 $Y=1.325
+ $X2=4.52 $Y2=1.535
r136 53 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=0.995
+ $X2=4.52 $Y2=1.16
r137 53 64 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.52 $Y=0.995
+ $X2=4.52 $Y2=0.745
r138 48 66 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=1.865
+ $X2=4.495 $Y2=1.7
r139 48 50 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.495 $Y=1.865
+ $X2=4.495 $Y2=2.27
r140 46 68 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.695 $Y2=1.7
r141 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r142 43 66 0.463323 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.385 $Y=1.7
+ $X2=4.495 $Y2=1.7
r143 43 45 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.385 $Y=1.7
+ $X2=3.925 $Y2=1.7
r144 39 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.16
r145 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.985
r146 36 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=1.16
r147 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=0.56
r148 32 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.99 $Y=1.325
+ $X2=5.99 $Y2=1.16
r149 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.99 $Y=1.325
+ $X2=5.99 $Y2=1.985
r150 29 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.99 $Y=0.995
+ $X2=5.99 $Y2=1.16
r151 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.99 $Y=0.995
+ $X2=5.99 $Y2=0.56
r152 25 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.325
+ $X2=5.535 $Y2=1.16
r153 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.535 $Y=1.325
+ $X2=5.535 $Y2=1.985
r154 22 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=0.995
+ $X2=5.535 $Y2=1.16
r155 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.535 $Y=0.995
+ $X2=5.535 $Y2=0.56
r156 18 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.325
+ $X2=5.115 $Y2=1.16
r157 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.115 $Y=1.325
+ $X2=5.115 $Y2=1.985
r158 15 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=0.995
+ $X2=5.115 $Y2=1.16
r159 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.115 $Y=0.995
+ $X2=5.115 $Y2=0.56
r160 11 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=1.7
r161 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=2.275
r162 7 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=1.7
r163 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=0.445
r164 2 66 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.47 $Y2=1.755
r165 2 50 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.47 $Y2=2.27
r166 1 62 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.345
+ $Y=0.235 $X2=4.47 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%A_561_413# 1 2 7 9 12 14 15 16 20 25 26 27
+ 30
c82 26 0 1.57048e-19 $X=3.565 $Y=1.325
c83 15 0 1.24075e-19 $X=4.68 $Y=1.16
r84 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r85 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.65 $Y=1.16
+ $X2=4.115 $Y2=1.16
r86 26 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.49 $Y2=1.16
r87 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=2.255
r88 25 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.415 $Y=0.995
+ $X2=3.49 $Y2=1.16
r89 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=0.995
r90 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.565 $Y2=2.255
r91 20 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.065 $Y2=2.34
r92 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r93 16 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.005 $Y2=0.45
r94 14 31 85.682 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=4.605 $Y=1.16
+ $X2=4.115 $Y2=1.16
r95 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.605 $Y=1.16
+ $X2=4.68 $Y2=1.16
r96 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.68 $Y=1.325
+ $X2=4.68 $Y2=1.16
r97 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.68 $Y=1.325
+ $X2=4.68 $Y2=1.985
r98 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.68 $Y=0.995
+ $X2=4.68 $Y2=1.16
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.68 $Y=0.995 $X2=4.68
+ $Y2=0.56
r100 2 22 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=3.065 $Y2=2.34
r101 1 18 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3.005 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 37 41 43 45
+ 47 49 54 59 67 73 76 79 82 85 89
r110 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r111 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r112 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r113 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r114 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r115 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r116 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r117 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 71 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r119 71 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r121 68 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.82 $Y2=2.72
r122 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=6.21 $Y2=2.72
r123 67 88 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.727 $Y2=2.72
r124 67 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 66 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r126 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r127 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 63 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r129 62 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r130 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r131 60 76 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r132 60 62 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r133 59 79 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=3.97 $Y2=2.72
r134 59 65 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=3.45 $Y2=2.72
r135 58 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 58 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r138 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r139 55 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 54 76 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r141 54 57 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r142 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r143 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r144 47 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r145 47 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r146 43 88 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.685 $Y=2.635
+ $X2=6.727 $Y2=2.72
r147 43 45 35.4598 $w=2.58e-07 $l=8e-07 $layer=LI1_cond $X=6.685 $Y=2.635
+ $X2=6.685 $Y2=1.835
r148 39 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r149 39 41 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=1.835
r150 38 82 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.07 $Y=2.72
+ $X2=4.927 $Y2=2.72
r151 37 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.82 $Y2=2.72
r152 37 38 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.07 $Y2=2.72
r153 33 82 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.927 $Y=2.635
+ $X2=4.927 $Y2=2.72
r154 33 35 36.3929 $w=2.83e-07 $l=9e-07 $layer=LI1_cond $X=4.927 $Y=2.635
+ $X2=4.927 $Y2=1.735
r155 32 79 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.12 $Y=2.72
+ $X2=3.97 $Y2=2.72
r156 31 82 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=4.927 $Y2=2.72
r157 31 32 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=4.12 $Y2=2.72
r158 27 79 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.72
r159 27 29 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.3
r160 23 76 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r161 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r162 19 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r163 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r164 6 45 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=6.505
+ $Y=1.485 $X2=6.64 $Y2=1.835
r165 5 41 300 $w=1.7e-07 $l=4.26615e-07 $layer=licon1_PDIFF $count=2 $X=5.61
+ $Y=1.485 $X2=5.78 $Y2=1.835
r166 4 35 300 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=2 $X=4.755
+ $Y=1.485 $X2=4.905 $Y2=1.735
r167 3 29 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=2.065 $X2=3.905 $Y2=2.3
r168 2 25 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r169 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%Q 1 2 3 4 14 17 18 20 21 22 23 24 25 26 27
+ 28 29 30 47 60
c45 21 0 1.62185e-19 $X=5.38 $Y=0.51
c46 20 0 1.24075e-19 $X=5.44 $Y=1.16
r47 58 60 21.7684 $w=2.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.25 $Y=1.325
+ $X2=6.25 $Y2=1.835
r48 30 66 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.705 $Y=1.16
+ $X2=6.385 $Y2=1.16
r49 28 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.25 $Y=1.87
+ $X2=6.25 $Y2=2.21
r50 28 60 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.25 $Y=1.87
+ $X2=6.25 $Y2=1.835
r51 27 50 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.25 $Y=0.85
+ $X2=6.25 $Y2=0.995
r52 27 55 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=6.25 $Y=0.85 $X2=6.25
+ $Y2=0.55
r53 26 55 1.70732 $w=2.68e-07 $l=4e-08 $layer=LI1_cond $X=6.25 $Y=0.51 $X2=6.25
+ $Y2=0.55
r54 25 50 7.45556 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=1.16
+ $X2=6.25 $Y2=0.995
r55 25 58 7.45556 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=1.16
+ $X2=6.25 $Y2=1.325
r56 25 47 4.99091 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=6.25 $Y=1.16
+ $X2=6.115 $Y2=1.16
r57 25 66 4.99091 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=6.25 $Y=1.16
+ $X2=6.385 $Y2=1.16
r58 24 47 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.785 $Y=1.16
+ $X2=6.115 $Y2=1.16
r59 22 23 15.1637 $w=2.83e-07 $l=3.75e-07 $layer=LI1_cond $X=5.382 $Y=1.835
+ $X2=5.382 $Y2=2.21
r60 21 74 11.3641 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=5.382 $Y=0.51
+ $X2=5.382 $Y2=0.745
r61 19 24 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.525 $Y=1.16
+ $X2=5.785 $Y2=1.16
r62 19 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.525 $Y=1.16
+ $X2=5.44 $Y2=1.16
r63 17 22 8.00645 $w=2.83e-07 $l=1.98e-07 $layer=LI1_cond $X=5.382 $Y=1.637
+ $X2=5.382 $Y2=1.835
r64 17 18 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=5.382 $Y=1.637
+ $X2=5.382 $Y2=1.495
r65 15 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.44 $Y=1.325
+ $X2=5.44 $Y2=1.16
r66 15 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.44 $Y=1.325
+ $X2=5.44 $Y2=1.495
r67 14 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.44 $Y=0.995
+ $X2=5.44 $Y2=1.16
r68 14 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.44 $Y=0.995
+ $X2=5.44 $Y2=0.745
r69 4 60 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=6.065
+ $Y=1.485 $X2=6.2 $Y2=1.835
r70 3 22 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=1.485 $X2=5.325 $Y2=1.835
r71 2 55 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=6.065
+ $Y=0.235 $X2=6.2 $Y2=0.55
r72 1 21 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.19
+ $Y=0.235 $X2=5.325 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_4%VGND 1 2 3 4 5 6 21 25 29 31 35 37 41 43 45
+ 47 49 54 59 67 73 76 79 82 85 89
c112 89 0 2.71124e-20 $X=6.67 $Y=0
c113 2 0 7.13094e-20 $X=1.905 $Y=0.235
r114 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r115 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r116 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r117 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r118 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r119 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r120 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r121 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r122 71 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r123 71 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r124 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r125 68 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=0 $X2=5.82
+ $Y2=0
r126 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=6.21 $Y2=0
r127 67 88 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.727 $Y2=0
r128 67 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.21
+ $Y2=0
r129 66 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r130 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r131 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r132 63 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r133 62 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r134 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r135 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r136 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r137 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.905
+ $Y2=0
r138 59 65 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.45
+ $Y2=0
r139 58 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r140 58 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r141 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r142 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r143 55 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r144 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r145 54 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r146 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r147 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r148 47 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r149 47 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r150 43 88 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.685 $Y=0.085
+ $X2=6.727 $Y2=0
r151 43 45 20.611 $w=2.58e-07 $l=4.65e-07 $layer=LI1_cond $X=6.685 $Y=0.085
+ $X2=6.685 $Y2=0.55
r152 39 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r153 39 41 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.55
r154 38 82 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.07 $Y=0 $X2=4.927
+ $Y2=0
r155 37 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=0 $X2=5.82
+ $Y2=0
r156 37 38 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.07 $Y2=0
r157 33 82 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.927 $Y=0.085
+ $X2=4.927 $Y2=0
r158 33 35 18.803 $w=2.83e-07 $l=4.65e-07 $layer=LI1_cond $X=4.927 $Y=0.085
+ $X2=4.927 $Y2=0.55
r159 32 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.905
+ $Y2=0
r160 31 82 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.785 $Y=0
+ $X2=4.927 $Y2=0
r161 31 32 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=4.785 $Y=0
+ $X2=4.07 $Y2=0
r162 27 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r163 27 29 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0.445
r164 23 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r165 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r166 19 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r167 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r168 6 45 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.64 $Y2=0.55
r169 5 41 182 $w=1.7e-07 $l=3.90864e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.235 $X2=5.78 $Y2=0.55
r170 4 35 182 $w=1.7e-07 $l=3.82721e-07 $layer=licon1_NDIFF $count=1 $X=4.755
+ $Y=0.235 $X2=4.905 $Y2=0.55
r171 3 29 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.235 $X2=3.905 $Y2=0.445
r172 2 25 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r173 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o2111ai_1.pex.spice
* Created: Thu Aug 27 14:34:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2111AI_1%D1 3 7 9 10 14
c31 14 0 7.45289e-20 $X=0.65 $Y=1.16
c32 9 0 1.59109e-19 $X=0.69 $Y=1.19
r33 14 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.65 $Y=1.16
+ $X2=0.65 $Y2=1.295
r34 14 16 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.65 $Y=1.16
+ $X2=0.65 $Y2=1.025
r35 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.65 $Y=1.16 $X2=0.65
+ $Y2=1.53
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.65
+ $Y=1.16 $X2=0.65 $Y2=1.16
r37 7 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.74 $Y=0.56
+ $X2=0.74 $Y2=1.025
r38 3 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.67 $Y=1.985
+ $X2=0.67 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%C1 3 7 9 10 14
c38 3 0 7.34074e-20 $X=1.1 $Y=0.56
r39 14 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.19 $Y=1.16
+ $X2=1.19 $Y2=1.295
r40 14 16 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.19 $Y=1.16
+ $X2=1.19 $Y2=1.025
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.16 $X2=1.19 $Y2=1.16
r42 10 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=1.53
+ $X2=1.19 $Y2=1.16
r43 9 15 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=1.19 $Y=0.51 $X2=1.19
+ $Y2=1.16
r44 7 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.1 $Y=1.985 $X2=1.1
+ $Y2=1.295
r45 3 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.1 $Y=0.56 $X2=1.1
+ $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%B1 3 7 9 10 14 15
c35 15 0 1.52049e-19 $X=1.73 $Y=1.16
c36 3 0 9.68735e-20 $X=1.64 $Y=0.56
r37 14 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.73 $Y2=1.295
r38 14 16 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.73 $Y2=1.025
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r40 9 10 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=1.19 $X2=1.67
+ $Y2=1.53
r41 9 15 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=1.67 $Y=1.19 $X2=1.67
+ $Y2=1.16
r42 7 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.64 $Y=1.985
+ $X2=1.64 $Y2=1.295
r43 3 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.64 $Y=0.56
+ $X2=1.64 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%A2 3 7 9 11 16 27
c38 27 0 9.68735e-20 $X=2.442 $Y=1.305
c39 3 0 9.08294e-20 $X=2.195 $Y=0.56
r40 20 27 4.17786 $w=3.45e-07 $l=3.1e-07 $layer=LI1_cond $X=2.442 $Y=1.615
+ $X2=2.442 $Y2=1.305
r41 17 27 3.02878 $w=6.18e-07 $l=1.57e-07 $layer=LI1_cond $X=2.285 $Y=1.305
+ $X2=2.442 $Y2=1.305
r42 16 19 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.285 $Y=1.16
+ $X2=2.285 $Y2=1.295
r43 16 18 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.285 $Y=1.16
+ $X2=2.285 $Y2=1.025
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=1.16 $X2=2.285 $Y2=1.16
r45 11 20 19.8755 $w=3.43e-07 $l=5.95e-07 $layer=LI1_cond $X=2.442 $Y=2.21
+ $X2=2.442 $Y2=1.615
r46 9 17 4.14769 $w=6.18e-07 $l=2.15e-07 $layer=LI1_cond $X=2.07 $Y=1.305
+ $X2=2.285 $Y2=1.305
r47 7 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.195 $Y=1.985
+ $X2=2.195 $Y2=1.295
r48 3 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.195 $Y=0.56
+ $X2=2.195 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%A1 3 7 9 14
c26 9 0 1.21874e-20 $X=2.99 $Y=1.19
r27 11 14 44.473 $w=2.9e-07 $l=2.15e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=2.95 $Y2=1.16
r28 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r29 5 11 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.735 $Y=1.305
+ $X2=2.735 $Y2=1.16
r30 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.735 $Y=1.305
+ $X2=2.735 $Y2=1.985
r31 1 11 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.735 $Y=1.015
+ $X2=2.735 $Y2=1.16
r32 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.735 $Y=1.015
+ $X2=2.735 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%VPWR 1 2 3 12 16 18 20 23 24 26 27 28 37
+ 46
r53 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 39 42 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 37 45 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=3.002 $Y2=2.72
r60 37 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 36 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 28 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 26 35 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.21 $Y=2.72 $X2=1.15
+ $Y2=2.72
r66 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=2.72
+ $X2=1.375 $Y2=2.72
r67 25 39 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.54 $Y=2.72 $X2=1.61
+ $Y2=2.72
r68 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=2.72
+ $X2=1.375 $Y2=2.72
r69 23 31 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.29 $Y=2.72 $X2=0.23
+ $Y2=2.72
r70 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.29 $Y=2.72
+ $X2=0.455 $Y2=2.72
r71 22 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.62 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=2.72
+ $X2=0.455 $Y2=2.72
r73 18 45 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.95 $Y=2.635
+ $X2=3.002 $Y2=2.72
r74 18 20 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=2.95 $Y=2.635
+ $X2=2.95 $Y2=1.88
r75 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=2.635
+ $X2=1.375 $Y2=2.72
r76 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.375 $Y=2.635
+ $X2=1.375 $Y2=2.34
r77 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=2.635
+ $X2=0.455 $Y2=2.72
r78 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.455 $Y=2.635
+ $X2=0.455 $Y2=2.34
r79 3 20 300 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.485 $X2=2.95 $Y2=1.88
r80 2 16 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.485 $X2=1.375 $Y2=2.34
r81 1 12 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.485 $X2=0.455 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%Y 1 2 3 12 14 16 18 20 22 25 26 37
c49 22 0 7.45289e-20 $X=0.885 $Y=1.885
r50 26 41 27.1832 $w=3.98e-07 $l=9e-07 $layer=LI1_cond $X=0.2 $Y=1.785 $X2=0.2
+ $Y2=0.885
r51 25 41 12.209 $w=6.03e-07 $l=3.75e-07 $layer=LI1_cond $X=0.387 $Y=0.51
+ $X2=0.387 $Y2=0.885
r52 25 37 2.17469 $w=6.03e-07 $l=1.1e-07 $layer=LI1_cond $X=0.387 $Y=0.51
+ $X2=0.387 $Y2=0.4
r53 20 26 14.5886 $w=4.08e-07 $l=4.75e-07 $layer=LI1_cond $X=0.79 $Y=1.905
+ $X2=0.315 $Y2=1.905
r54 20 22 5.07612 $w=2.4e-07 $l=1.17e-07 $layer=LI1_cond $X=0.79 $Y=1.905
+ $X2=0.907 $Y2=1.905
r55 16 24 2.92029 $w=3.45e-07 $l=1.2e-07 $layer=LI1_cond $X=1.922 $Y=2.025
+ $X2=1.922 $Y2=1.905
r56 16 18 10.5223 $w=3.43e-07 $l=3.15e-07 $layer=LI1_cond $X=1.922 $Y=2.025
+ $X2=1.922 $Y2=2.34
r57 15 22 5.07612 $w=2.4e-07 $l=1.18e-07 $layer=LI1_cond $X=1.025 $Y=1.905
+ $X2=0.907 $Y2=1.905
r58 14 24 4.18576 $w=2.4e-07 $l=1.72e-07 $layer=LI1_cond $X=1.75 $Y=1.905
+ $X2=1.922 $Y2=1.905
r59 14 15 34.8134 $w=2.38e-07 $l=7.25e-07 $layer=LI1_cond $X=1.75 $Y=1.905
+ $X2=1.025 $Y2=1.905
r60 10 22 1.41848 $w=2.35e-07 $l=1.2e-07 $layer=LI1_cond $X=0.907 $Y=2.025
+ $X2=0.907 $Y2=1.905
r61 10 12 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=0.907 $Y=2.025
+ $X2=0.907 $Y2=2.3
r62 3 24 600 $w=1.7e-07 $l=4.95984e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.485 $X2=1.93 $Y2=1.885
r63 3 18 600 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.485 $X2=1.93 $Y2=2.34
r64 2 22 600 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=1.485 $X2=0.885 $Y2=1.885
r65 2 12 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=1.485 $X2=0.885 $Y2=2.3
r66 1 37 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.4
+ $Y=0.235 $X2=0.525 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%A_343_47# 1 2 7 9 11 15
r24 13 15 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.95 $Y=0.625
+ $X2=2.95 $Y2=0.4
r25 12 18 4.72967 $w=2e-07 $l=1.73e-07 $layer=LI1_cond $X=2.095 $Y=0.725
+ $X2=1.922 $Y2=0.725
r26 11 13 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.785 $Y=0.725
+ $X2=2.95 $Y2=0.625
r27 11 12 38.2636 $w=1.98e-07 $l=6.9e-07 $layer=LI1_cond $X=2.785 $Y=0.725
+ $X2=2.095 $Y2=0.725
r28 7 18 2.73391 $w=3.45e-07 $l=1e-07 $layer=LI1_cond $X=1.922 $Y=0.625
+ $X2=1.922 $Y2=0.725
r29 7 9 7.51593 $w=3.43e-07 $l=2.25e-07 $layer=LI1_cond $X=1.922 $Y=0.625
+ $X2=1.922 $Y2=0.4
r30 2 15 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.81
+ $Y=0.235 $X2=2.95 $Y2=0.4
r31 1 18 182 $w=1.7e-07 $l=6.02993e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.235 $X2=1.93 $Y2=0.74
r32 1 9 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.235 $X2=1.93 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_1%VGND 1 6 8 10 20 21 24
r35 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r36 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r37 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r38 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.45
+ $Y2=0
r39 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.99
+ $Y2=0
r40 17 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r41 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r42 12 16 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r43 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.45
+ $Y2=0
r44 10 16 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.07
+ $Y2=0
r45 8 17 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r46 8 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r47 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085 $X2=2.45
+ $Y2=0
r48 4 6 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.37
r49 1 6 182 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.45 $Y2=0.37
.ends


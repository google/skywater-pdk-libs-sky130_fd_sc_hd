* File: sky130_fd_sc_hd__decap_12.spice.SKY130_FD_SC_HD__DECAP_12.pxi
* Created: Thu Aug 27 14:13:22 2020
* 
x_PM_SKY130_FD_SC_HD__DECAP_12%VGND N_VGND_M1001_s N_VGND_M1000_g N_VGND_c_18_n
+ N_VGND_c_19_n VGND N_VGND_c_20_n N_VGND_c_21_n N_VGND_c_22_n N_VGND_c_23_n
+ PM_SKY130_FD_SC_HD__DECAP_12%VGND
x_PM_SKY130_FD_SC_HD__DECAP_12%VPWR N_VPWR_M1000_s N_VPWR_M1001_g N_VPWR_c_48_n
+ N_VPWR_c_49_n VPWR N_VPWR_c_44_n N_VPWR_c_45_n N_VPWR_c_46_n N_VPWR_c_47_n
+ PM_SKY130_FD_SC_HD__DECAP_12%VPWR
cc_1 VNB N_VGND_c_18_n 0.0304509f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=0.385
cc_2 VNB N_VGND_c_19_n 0.0927556f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=0.385
cc_3 VNB N_VGND_c_20_n 0.0491357f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.87
cc_4 VNB N_VGND_c_21_n 0.0241734f $X=-0.19 $Y=-0.24 $X2=2.645 $Y2=1.87
cc_5 VNB N_VGND_c_22_n 0.0439157f $X=-0.19 $Y=-0.24 $X2=5.26 $Y2=0.475
cc_6 VNB N_VGND_c_23_n 0.274429f $X=-0.19 $Y=-0.24 $X2=5.29 $Y2=0
cc_7 VNB N_VPWR_c_44_n 0.173698f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.29
cc_8 VNB N_VPWR_c_45_n 0.266152f $X=-0.19 $Y=-0.24 $X2=2.48 $Y2=1.87
cc_9 VNB N_VPWR_c_46_n 0.0177273f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0
cc_10 VNB N_VPWR_c_47_n 0.231782f $X=-0.19 $Y=-0.24 $X2=5.26 $Y2=0.385
cc_11 VPB N_VGND_c_19_n 0.0068688f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=0.385
cc_12 VPB N_VGND_c_20_n 0.129851f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.87
cc_13 VPB N_VGND_c_21_n 0.235821f $X=-0.19 $Y=1.305 $X2=2.645 $Y2=1.87
cc_14 VPB N_VPWR_c_48_n 0.0281269f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=0.385
cc_15 VPB N_VPWR_c_49_n 0.0597303f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=0.385
cc_16 VPB N_VPWR_c_46_n 0.0955067f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=0
cc_17 VPB N_VPWR_c_47_n 0.0426425f $X=-0.19 $Y=1.305 $X2=5.26 $Y2=0.385
cc_18 N_VGND_c_19_n N_VPWR_c_48_n 0.164206f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_19 N_VGND_c_20_n N_VPWR_c_48_n 0.157227f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_20 N_VGND_c_21_n N_VPWR_c_48_n 0.124986f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_21 N_VGND_c_19_n N_VPWR_c_49_n 0.0561345f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_22 N_VGND_c_20_n N_VPWR_c_49_n 0.0493583f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_23 N_VGND_c_18_n N_VPWR_c_44_n 0.0203068f $X=4.96 $Y=0.385 $X2=0 $Y2=0
cc_24 N_VGND_c_19_n N_VPWR_c_44_n 0.247023f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_25 N_VGND_c_20_n N_VPWR_c_44_n 0.147138f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_26 N_VGND_c_21_n N_VPWR_c_44_n 0.00421128f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_27 N_VGND_c_18_n N_VPWR_c_45_n 0.216233f $X=4.96 $Y=0.385 $X2=0 $Y2=0
cc_28 N_VGND_c_19_n N_VPWR_c_45_n 0.00648593f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_29 N_VGND_c_21_n N_VPWR_c_45_n 0.15829f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_30 N_VGND_c_22_n N_VPWR_c_45_n 0.0242057f $X=5.26 $Y=0.475 $X2=0 $Y2=0
cc_31 N_VGND_c_18_n N_VPWR_c_46_n 0.179033f $X=4.96 $Y=0.385 $X2=0 $Y2=0
cc_32 N_VGND_c_19_n N_VPWR_c_46_n 0.0327855f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_33 N_VGND_c_21_n N_VPWR_c_46_n 0.324097f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_34 N_VGND_c_22_n N_VPWR_c_46_n 0.0425452f $X=5.26 $Y=0.475 $X2=0 $Y2=0

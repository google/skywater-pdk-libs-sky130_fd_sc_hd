* File: sky130_fd_sc_hd__or3b_1.pex.spice
* Created: Thu Aug 27 14:43:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR3B_1%C_N 1 3 6 8 14 17
c22 8 0 1.57334e-19 $X=0.15 $Y=1.105
r23 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r24 8 17 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r25 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r26 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r27 4 6 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r28 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r29 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%A_109_93# 1 2 9 13 15 16 17 19 23
c43 15 0 1.57334e-19 $X=1.335 $Y=1.16
r44 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.16 $X2=1.135 $Y2=1.16
r45 21 27 17.669 $w=2.9e-07 $l=4.2e-07 $layer=LI1_cond $X=0.68 $Y=1.16 $X2=0.68
+ $Y2=0.74
r46 21 23 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=1.135 $Y2=1.16
r47 17 21 9.01297 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=1.16
r48 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=1.63
r49 15 24 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.135 $Y2=1.16
r50 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.41 $Y2=1.16
r51 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r52 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.695
r53 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r54 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.475
r55 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.63
r56 1 27 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%B 2 4 7 8 9 10 11 12 18
r42 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=2.28 $X2=1.825 $Y2=2.28
r43 12 18 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.61 $Y=2.29
+ $X2=1.825 $Y2=2.29
r44 11 12 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=2.29
+ $X2=1.61 $Y2=2.29
r45 10 11 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=2.29
+ $X2=1.15 $Y2=2.29
r46 8 9 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.8 $Y=0.76 $X2=1.8
+ $Y2=0.91
r47 7 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.475 $X2=1.83
+ $Y2=0.76
r48 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.77 $Y=1.695
+ $X2=1.77 $Y2=0.91
r49 2 17 34.1986 $w=3.29e-07 $l=1.60156e-07 $layer=POLY_cond $X=1.77 $Y=2.145
+ $X2=1.825 $Y2=2.28
r50 2 4 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.77 $Y=2.145 $X2=1.77
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%A 1 3 7 9 10 11 17 18
c52 18 0 1.20602e-19 $X=1.647 $Y=1.325
r53 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.16 $X2=2.23 $Y2=1.16
r54 11 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.07 $Y=1.16 $X2=2.23
+ $Y2=1.16
r55 11 22 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.07 $Y=1.16 $X2=1.77
+ $Y2=1.16
r56 10 18 9.64289 $w=2.43e-07 $l=2.05e-07 $layer=LI1_cond $X=1.647 $Y=1.53
+ $X2=1.647 $Y2=1.325
r57 9 18 4.01731 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=1.647 $Y=1.16
+ $X2=1.647 $Y2=1.325
r58 9 22 2.99472 $w=3.3e-07 $l=1.23e-07 $layer=LI1_cond $X=1.647 $Y=1.16
+ $X2=1.77 $Y2=1.16
r59 5 16 38.9235 $w=2.69e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.25 $Y=0.995
+ $X2=2.23 $Y2=1.16
r60 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.25 $Y=0.995 $X2=2.25
+ $Y2=0.475
r61 1 16 38.9235 $w=2.69e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.245 $Y=1.325
+ $X2=2.23 $Y2=1.16
r62 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.245 $Y=1.325
+ $X2=2.245 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%A_215_53# 1 2 3 12 15 19 21 22 23 27 29 31 36
+ 38 42 43 48 49 50 53
c100 48 0 1.14153e-19 $X=2.71 $Y=1.16
c101 36 0 1.06604e-19 $X=2.605 $Y=1.495
r102 49 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=1.325
r103 49 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=0.995
r104 48 51 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.657 $Y=1.16
+ $X2=2.657 $Y2=1.325
r105 48 50 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.657 $Y=1.16
+ $X2=2.657 $Y2=0.995
r106 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.16 $X2=2.71 $Y2=1.16
r107 43 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.115 $Y=1.58
+ $X2=2.115 $Y2=1.87
r108 38 40 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.19 $Y=1.685
+ $X2=1.19 $Y2=1.87
r109 36 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.605 $Y=1.495
+ $X2=2.605 $Y2=1.325
r110 33 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.605 $Y=0.825
+ $X2=2.605 $Y2=0.995
r111 32 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=1.58
+ $X2=2.115 $Y2=1.58
r112 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.52 $Y=1.58
+ $X2=2.605 $Y2=1.495
r113 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.52 $Y=1.58 $X2=2.2
+ $Y2=1.58
r114 30 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=0.74
+ $X2=2.04 $Y2=0.74
r115 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.52 $Y=0.74
+ $X2=2.605 $Y2=0.825
r116 29 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.52 $Y=0.74
+ $X2=2.125 $Y2=0.74
r117 25 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.655
+ $X2=2.04 $Y2=0.74
r118 25 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.04 $Y=0.655
+ $X2=2.04 $Y2=0.47
r119 24 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.87
+ $X2=1.19 $Y2=1.87
r120 23 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.87
+ $X2=2.115 $Y2=1.87
r121 23 24 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.03 $Y=1.87
+ $X2=1.355 $Y2=1.87
r122 21 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=2.04 $Y2=0.74
r123 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=1.285 $Y2=0.74
r124 17 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.155 $Y=0.655
+ $X2=1.285 $Y2=0.74
r125 17 19 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.155 $Y=0.655
+ $X2=1.155 $Y2=0.42
r126 15 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.735 $Y=1.985
+ $X2=2.735 $Y2=1.325
r127 12 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.735 $Y=0.56
+ $X2=2.735 $Y2=0.995
r128 3 38 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.685
r129 2 27 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.265 $X2=2.04 $Y2=0.47
r130 1 19 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.265 $X2=1.2 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%VPWR 1 2 7 9 13 15 17 27 28 34
c33 9 0 1.56946e-19 $X=0.26 $Y=1.66
c34 2 0 1.06604e-19 $X=2.32 $Y=1.485
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r37 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r38 25 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.65 $Y=2.72 $X2=2.51
+ $Y2=2.72
r39 25 27 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.65 $Y=2.72
+ $X2=2.99 $Y2=2.72
r40 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 21 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 20 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 18 31 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r46 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 17 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.37 $Y=2.72 $X2=2.51
+ $Y2=2.72
r48 17 23 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.37 $Y=2.72 $X2=2.07
+ $Y2=2.72
r49 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 11 34 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.635
+ $X2=2.51 $Y2=2.72
r52 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.51 $Y=2.635
+ $X2=2.51 $Y2=2
r53 7 31 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r54 7 9 43.2166 $w=2.58e-07 $l=9.75e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=1.66
r55 2 13 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.485 $X2=2.52 $Y2=2
r56 1 9 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%X 1 2 12 14 15 16
r18 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=2.997 $Y=1.632
+ $X2=2.997 $Y2=1.845
r19 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.997 $Y=1.632
+ $X2=2.997 $Y2=1.495
r20 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=2.945 $Y=0.587
+ $X2=3.05 $Y2=0.587
r21 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.05 $Y=0.76 $X2=3.05
+ $Y2=0.587
r22 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.05 $Y=0.76
+ $X2=3.05 $Y2=1.495
r23 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.485 $X2=2.945 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.945 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_1%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
c53 12 0 1.56946e-19 $X=0.26 $Y=0.73
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r55 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r56 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r57 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 34 46 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.482
+ $Y2=0
r59 34 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.99
+ $Y2=0
r60 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r61 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r64 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.07
+ $Y2=0
r65 29 46 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.482
+ $Y2=0
r66 29 32 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.07
+ $Y2=0
r67 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r68 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 25 40 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r70 25 27 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=1.15
+ $Y2=0
r71 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r72 24 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.15
+ $Y2=0
r73 22 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r74 22 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 18 46 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.482 $Y=0.085
+ $X2=2.482 $Y2=0
r76 18 20 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.482 $Y=0.085
+ $X2=2.482 $Y2=0.4
r77 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r78 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.4
r79 10 40 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r80 10 12 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.73
r81 3 20 182 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.265 $X2=2.505 $Y2=0.4
r82 2 16 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.265 $X2=1.62 $Y2=0.4
r83 1 12 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.73
.ends


* File: sky130_fd_sc_hd__or4_1.spice
* Created: Thu Aug 27 14:43:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4_1.pex.spice"
.subckt sky130_fd_sc_hd__or4_1  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1005 N_A_27_297#_M1005_d N_D_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.1092 PD=0.75 PS=1.36 NRD=7.14 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g N_A_27_297#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0693 PD=0.69 PS=0.75 NRD=0 NRS=7.14 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_27_297#_M1004_d N_B_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_297#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_27_297#_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.123773 PD=1.84 PS=1.2028 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 A_109_297# N_D_M1008_g N_A_27_297#_M1008_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0693 AS=0.1092 PD=0.75 PS=1.36 NRD=51.5943 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1000 A_205_297# N_C_M1000_g A_109_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0693 PD=0.63 PS=0.75 NRD=23.443 NRS=51.5943 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 A_277_297# N_B_M1002_g A_205_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=51.5943 NRS=23.443 M=1 R=2.8 SA=75001 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_277_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.0693 PD=0.792676 PS=0.75 NRD=72.1217 NRS=51.5943 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_297#_M1001_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.208803 PD=2.54 PS=1.88732 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_59 VPB 0 1.1436e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__or4_1.pxi.spice"
*
.ends
*
*

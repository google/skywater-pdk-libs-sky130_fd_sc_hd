* File: sky130_fd_sc_hd__o41a_1.pxi.spice
* Created: Tue Sep  1 19:26:20 2020
* 
x_PM_SKY130_FD_SC_HD__O41A_1%A_103_21# N_A_103_21#_M1004_s N_A_103_21#_M1000_d
+ N_A_103_21#_c_66_n N_A_103_21#_M1011_g N_A_103_21#_M1002_g N_A_103_21#_c_71_n
+ N_A_103_21#_c_67_n N_A_103_21#_c_84_p N_A_103_21#_c_68_n N_A_103_21#_c_69_n
+ N_A_103_21#_c_73_n PM_SKY130_FD_SC_HD__O41A_1%A_103_21#
x_PM_SKY130_FD_SC_HD__O41A_1%B1 N_B1_M1000_g N_B1_c_119_n N_B1_M1004_g B1
+ N_B1_c_121_n PM_SKY130_FD_SC_HD__O41A_1%B1
x_PM_SKY130_FD_SC_HD__O41A_1%A4 N_A4_c_149_n N_A4_M1008_g N_A4_c_150_n
+ N_A4_M1007_g A4 A4 A4 N_A4_c_153_n PM_SKY130_FD_SC_HD__O41A_1%A4
x_PM_SKY130_FD_SC_HD__O41A_1%A3 N_A3_M1005_g N_A3_M1001_g A3 A3 A3 N_A3_c_187_n
+ N_A3_c_191_n N_A3_c_188_n PM_SKY130_FD_SC_HD__O41A_1%A3
x_PM_SKY130_FD_SC_HD__O41A_1%A2 N_A2_M1010_g N_A2_M1006_g A2 A2 A2 N_A2_c_221_n
+ N_A2_c_222_n N_A2_c_223_n PM_SKY130_FD_SC_HD__O41A_1%A2
x_PM_SKY130_FD_SC_HD__O41A_1%A1 N_A1_M1003_g N_A1_M1009_g A1 N_A1_c_257_n
+ N_A1_c_258_n PM_SKY130_FD_SC_HD__O41A_1%A1
x_PM_SKY130_FD_SC_HD__O41A_1%X N_X_M1011_s N_X_M1002_s X X X X X X N_X_c_282_n X
+ X PM_SKY130_FD_SC_HD__O41A_1%X
x_PM_SKY130_FD_SC_HD__O41A_1%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_c_303_n
+ N_VPWR_c_304_n N_VPWR_c_305_n VPWR N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_308_n N_VPWR_c_302_n PM_SKY130_FD_SC_HD__O41A_1%VPWR
x_PM_SKY130_FD_SC_HD__O41A_1%VGND N_VGND_M1011_d N_VGND_M1007_d N_VGND_M1010_d
+ N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n
+ N_VGND_c_359_n N_VGND_c_360_n VGND N_VGND_c_361_n N_VGND_c_362_n
+ N_VGND_c_363_n N_VGND_c_364_n PM_SKY130_FD_SC_HD__O41A_1%VGND
x_PM_SKY130_FD_SC_HD__O41A_1%A_321_47# N_A_321_47#_M1004_d N_A_321_47#_M1005_d
+ N_A_321_47#_M1003_d N_A_321_47#_c_442_n N_A_321_47#_c_414_n
+ N_A_321_47#_c_415_n N_A_321_47#_c_449_n N_A_321_47#_c_416_n
+ N_A_321_47#_c_417_n N_A_321_47#_c_418_n PM_SKY130_FD_SC_HD__O41A_1%A_321_47#
cc_1 VNB N_A_103_21#_c_66_n 0.0224361f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_2 VNB N_A_103_21#_c_67_n 0.00558415f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=0.38
cc_3 VNB N_A_103_21#_c_68_n 0.0309014f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_4 VNB N_A_103_21#_c_69_n 0.0121363f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1
cc_5 VNB N_B1_c_119_n 0.0198752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB B1 0.00682009f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.56
cc_7 VNB N_B1_c_121_n 0.0315249f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.985
cc_8 VNB N_A4_c_149_n 0.0280081f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=0.235
cc_9 VNB N_A4_c_150_n 0.0171835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A3_c_187_n 0.0253555f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.455
cc_11 VNB N_A3_c_188_n 0.0182152f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=0.38
cc_12 VNB N_A2_c_221_n 0.0238843f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.455
cc_13 VNB N_A2_c_222_n 0.00172914f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=0.715
cc_14 VNB N_A2_c_223_n 0.0182931f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=0.38
cc_15 VNB A1 0.013263f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.56
cc_16 VNB N_A1_c_257_n 0.0294134f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.985
cc_17 VNB N_A1_c_258_n 0.0227197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0298109f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.56
cc_19 VNB N_X_c_282_n 0.0183576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_302_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_354_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.985
cc_22 VNB N_VGND_c_355_n 0.00561552f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=0.715
cc_23 VNB N_VGND_c_356_n 0.0055721f $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=1.745
cc_24 VNB N_VGND_c_357_n 0.0217162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_358_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_26 VNB N_VGND_c_359_n 0.0190293f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_27 VNB N_VGND_c_360_n 0.00631567f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1
cc_28 VNB N_VGND_c_361_n 0.0309953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_362_n 0.0201086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_363_n 0.225904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_364_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_321_47#_c_414_n 0.00877451f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.285
cc_33 VNB N_A_321_47#_c_415_n 0.00528521f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.455
cc_34 VNB N_A_321_47#_c_416_n 0.0180479f $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=1.745
cc_35 VNB N_A_321_47#_c_417_n 0.0183265f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_36 VNB N_A_321_47#_c_418_n 0.0079689f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_37 VPB N_A_103_21#_M1002_g 0.0215593f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.985
cc_38 VPB N_A_103_21#_c_71_n 0.00208437f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.455
cc_39 VPB N_A_103_21#_c_68_n 0.0100731f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_40 VPB N_A_103_21#_c_73_n 0.00328457f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.62
cc_41 VPB N_B1_M1000_g 0.0207711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B1_c_121_n 0.0095959f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.985
cc_43 VPB N_A4_c_149_n 0.00801975f $X=-0.19 $Y=1.305 $X2=1.195 $Y2=0.235
cc_44 VPB N_A4_M1008_g 0.0222316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A4_c_153_n 0.00105896f $X=-0.19 $Y=1.305 $X2=1.32 $Y2=0.715
cc_46 VPB N_A3_M1001_g 0.0210481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A3_c_187_n 0.0064814f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.455
cc_48 VPB N_A3_c_191_n 9.91125e-19 $X=-0.19 $Y=1.305 $X2=1.32 $Y2=0.715
cc_49 VPB N_A2_M1006_g 0.0197733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A2_c_221_n 0.00633674f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.455
cc_51 VPB N_A2_c_222_n 0.00292695f $X=-0.19 $Y=1.305 $X2=1.32 $Y2=0.715
cc_52 VPB N_A1_M1009_g 0.026598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB A1 0.00421218f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=0.56
cc_54 VPB N_A1_c_257_n 0.00583605f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.985
cc_55 VPB X 0.00830535f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=0.56
cc_56 VPB X 0.0369374f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.985
cc_57 VPB X 0.018114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_303_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.59 $Y2=0.56
cc_59 VPB N_VPWR_c_304_n 0.013819f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.985
cc_60 VPB N_VPWR_c_305_n 0.039714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_306_n 0.0230659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_307_n 0.0645052f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_63 VPB N_VPWR_c_308_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_302_n 0.049963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 N_A_103_21#_M1002_g N_B1_M1000_g 0.0187154f $X=0.8 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_103_21#_c_73_n N_B1_M1000_g 0.0207999f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_67 N_A_103_21#_c_67_n N_B1_c_119_n 0.00603017f $X=1.32 $Y=0.38 $X2=0 $Y2=0
cc_68 N_A_103_21#_c_69_n N_B1_c_119_n 0.00563732f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_69 N_A_103_21#_c_69_n B1 0.0346336f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_70 N_A_103_21#_c_73_n B1 0.0241809f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_71 N_A_103_21#_c_71_n N_B1_c_121_n 0.0044842f $X=0.975 $Y=1.455 $X2=0 $Y2=0
cc_72 N_A_103_21#_c_68_n N_B1_c_121_n 0.0217072f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_103_21#_c_69_n N_B1_c_121_n 0.0125846f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_74 N_A_103_21#_c_73_n N_B1_c_121_n 0.00771966f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_75 N_A_103_21#_c_84_p N_A4_M1008_g 0.0072064f $X=1.51 $Y=1.96 $X2=0 $Y2=0
cc_76 N_A_103_21#_c_73_n N_A4_M1008_g 0.00270688f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_77 N_A_103_21#_c_67_n N_A4_c_150_n 4.59528e-19 $X=1.32 $Y=0.38 $X2=0 $Y2=0
cc_78 N_A_103_21#_c_84_p N_A4_c_153_n 0.0343747f $X=1.51 $Y=1.96 $X2=0 $Y2=0
cc_79 N_A_103_21#_c_73_n N_A4_c_153_n 0.0167217f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_80 N_A_103_21#_c_66_n X 0.0104506f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_103_21#_M1002_g X 0.00231917f $X=0.8 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_103_21#_c_71_n X 0.00583732f $X=0.975 $Y=1.455 $X2=0 $Y2=0
cc_83 N_A_103_21#_c_69_n X 0.0351395f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_84 N_A_103_21#_c_66_n N_X_c_282_n 0.0176602f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_103_21#_M1002_g X 0.0257823f $X=0.8 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_103_21#_c_68_n X 0.0029035f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_103_21#_c_69_n X 0.00690646f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_88 N_A_103_21#_c_73_n X 0.0191457f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_89 N_A_103_21#_c_73_n N_VPWR_M1002_d 0.00168581f $X=1.51 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_103_21#_M1002_g N_VPWR_c_303_n 0.0129874f $X=0.8 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_103_21#_c_73_n N_VPWR_c_303_n 0.0176682f $X=1.51 $Y=1.62 $X2=0 $Y2=0
cc_92 N_A_103_21#_M1002_g N_VPWR_c_306_n 0.0046653f $X=0.8 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_103_21#_c_84_p N_VPWR_c_307_n 0.0173023f $X=1.51 $Y=1.96 $X2=0 $Y2=0
cc_94 N_A_103_21#_M1000_d N_VPWR_c_302_n 0.0136451f $X=1.295 $Y=1.485 $X2=0
+ $Y2=0
cc_95 N_A_103_21#_M1002_g N_VPWR_c_302_n 0.00934473f $X=0.8 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_103_21#_c_84_p N_VPWR_c_302_n 0.0095654f $X=1.51 $Y=1.96 $X2=0 $Y2=0
cc_97 N_A_103_21#_c_69_n N_VGND_M1011_d 0.00529577f $X=0.975 $Y=1 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_103_21#_c_66_n N_VGND_c_354_n 0.00438629f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_103_21#_c_67_n N_VGND_c_354_n 0.0154051f $X=1.32 $Y=0.38 $X2=0 $Y2=0
cc_100 N_A_103_21#_c_68_n N_VGND_c_354_n 9.52068e-19 $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_103_21#_c_69_n N_VGND_c_354_n 0.0132445f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_102 N_A_103_21#_c_66_n N_VGND_c_357_n 0.00585385f $X=0.59 $Y=0.995 $X2=0
+ $Y2=0
cc_103 N_A_103_21#_c_67_n N_VGND_c_361_n 0.0191165f $X=1.32 $Y=0.38 $X2=0 $Y2=0
cc_104 N_A_103_21#_c_69_n N_VGND_c_361_n 0.00455475f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_105 N_A_103_21#_M1004_s N_VGND_c_363_n 0.00209863f $X=1.195 $Y=0.235 $X2=0
+ $Y2=0
cc_106 N_A_103_21#_c_66_n N_VGND_c_363_n 0.0130305f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_103_21#_c_67_n N_VGND_c_363_n 0.0123122f $X=1.32 $Y=0.38 $X2=0 $Y2=0
cc_108 N_A_103_21#_c_69_n N_VGND_c_363_n 0.00826911f $X=0.975 $Y=1 $X2=0 $Y2=0
cc_109 N_A_103_21#_c_69_n N_A_321_47#_c_415_n 0.00808484f $X=0.975 $Y=1 $X2=0
+ $Y2=0
cc_110 B1 N_A4_c_149_n 0.00135064f $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_111 N_B1_c_121_n N_A4_c_149_n 0.0203981f $X=1.44 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_112 N_B1_M1000_g N_A4_M1008_g 0.0214206f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B1_c_119_n N_A4_c_150_n 0.023537f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B1_M1000_g N_A4_c_153_n 0.00105744f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_115 B1 N_A4_c_153_n 0.0168625f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B1_c_121_n N_A4_c_153_n 4.70936e-19 $X=1.44 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B1_M1000_g N_VPWR_c_303_n 0.0116043f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B1_M1000_g N_VPWR_c_307_n 0.0046653f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_VPWR_c_302_n 0.00851192f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_c_119_n N_VGND_c_354_n 0.00211786f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_119_n N_VGND_c_361_n 0.00541964f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B1_c_119_n N_VGND_c_363_n 0.0110552f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B1_c_119_n N_A_321_47#_c_415_n 6.10199e-19 $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_124 B1 N_A_321_47#_c_415_n 0.0033403f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_125 N_A4_M1008_g N_A3_M1001_g 0.0297627f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A4_c_153_n N_A3_M1001_g 0.00793238f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A4_c_149_n N_A3_c_187_n 0.0213209f $X=1.89 $Y=1.325 $X2=0 $Y2=0
cc_128 N_A4_c_153_n N_A3_c_187_n 8.70727e-19 $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A4_c_149_n N_A3_c_191_n 8.90747e-19 $X=1.89 $Y=1.325 $X2=0 $Y2=0
cc_130 N_A4_M1008_g N_A3_c_191_n 9.94192e-19 $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A4_c_153_n N_A3_c_191_n 0.086339f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A4_c_150_n N_A3_c_188_n 0.0178111f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A4_M1008_g N_VPWR_c_303_n 9.06371e-19 $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A4_M1008_g N_VPWR_c_307_n 0.00445128f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A4_c_153_n N_VPWR_c_307_n 0.0140494f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A4_M1008_g N_VPWR_c_302_n 0.00812503f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A4_c_153_n N_VPWR_c_302_n 0.0116719f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A4_c_153_n A_393_297# 0.0128822f $X=2.03 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_139 N_A4_c_150_n N_VGND_c_355_n 0.00318876f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A4_c_150_n N_VGND_c_361_n 0.00439206f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A4_c_150_n N_VGND_c_363_n 0.00619524f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A4_c_149_n N_A_321_47#_c_414_n 0.00609178f $X=1.89 $Y=1.325 $X2=0 $Y2=0
cc_143 N_A4_c_150_n N_A_321_47#_c_414_n 0.0118392f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A4_c_153_n N_A_321_47#_c_414_n 0.02565f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A4_c_149_n N_A_321_47#_c_415_n 4.48324e-19 $X=1.89 $Y=1.325 $X2=0 $Y2=0
cc_146 N_A3_M1001_g N_A2_M1006_g 0.0386094f $X=2.48 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A3_c_191_n N_A2_M1006_g 0.00370451f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A3_c_187_n N_A2_c_221_n 0.0215729f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A3_c_191_n N_A2_c_221_n 2.88395e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A3_M1001_g N_A2_c_222_n 0.00105245f $X=2.48 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A3_c_187_n N_A2_c_222_n 0.00142573f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A3_c_191_n N_A2_c_222_n 0.0696548f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A3_c_188_n N_A2_c_223_n 0.0159796f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A3_M1001_g N_VPWR_c_307_n 0.00374292f $X=2.48 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A3_c_191_n N_VPWR_c_307_n 0.0139564f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A3_M1001_g N_VPWR_c_302_n 0.00600416f $X=2.48 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A3_c_191_n N_VPWR_c_302_n 0.0114332f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A3_c_191_n A_511_297# 0.00923629f $X=2.57 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_159 N_A3_c_188_n N_VGND_c_355_n 0.00318876f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A3_c_188_n N_VGND_c_359_n 0.00439206f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A3_c_188_n N_VGND_c_363_n 0.00641625f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A3_c_187_n N_A_321_47#_c_414_n 6.13264e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A3_c_191_n N_A_321_47#_c_414_n 0.01331f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A3_c_188_n N_A_321_47#_c_414_n 0.0109589f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A3_c_187_n N_A_321_47#_c_418_n 0.00398638f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A3_c_191_n N_A_321_47#_c_418_n 0.0136799f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A2_M1006_g N_A1_M1009_g 0.0349353f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A2_c_222_n N_A1_M1009_g 0.012037f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A2_c_221_n A1 8.63316e-19 $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A2_c_222_n A1 0.016464f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A2_c_221_n N_A1_c_257_n 0.021693f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_c_222_n N_A1_c_257_n 3.12795e-19 $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A2_c_223_n N_A1_c_258_n 0.017202f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_M1006_g N_VPWR_c_305_n 0.00208619f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A2_c_222_n N_VPWR_c_305_n 0.0412132f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A2_M1006_g N_VPWR_c_307_n 0.00372875f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_c_222_n N_VPWR_c_307_n 0.0149675f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A2_M1006_g N_VPWR_c_302_n 0.00591481f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_c_222_n N_VPWR_c_302_n 0.0129095f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A2_c_222_n A_619_297# 0.0117991f $X=3.11 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_181 N_A2_c_223_n N_VGND_c_356_n 0.00317203f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_223_n N_VGND_c_359_n 0.00439206f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_223_n N_VGND_c_363_n 0.00650478f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_221_n N_A_321_47#_c_416_n 0.00445034f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A2_c_222_n N_A_321_47#_c_416_n 0.0286482f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_c_223_n N_A_321_47#_c_416_n 0.0133132f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A2_c_223_n N_A_321_47#_c_417_n 8.45515e-19 $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_M1009_g N_VPWR_c_305_n 0.0208805f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_189 A1 N_VPWR_c_305_n 0.0224218f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A1_c_257_n N_VPWR_c_305_n 0.00396625f $X=3.65 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A1_M1009_g N_VPWR_c_307_n 0.0046653f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A1_M1009_g N_VPWR_c_302_n 0.00827284f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A1_c_258_n N_VGND_c_356_n 0.00317203f $X=3.65 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_258_n N_VGND_c_362_n 0.00435288f $X=3.65 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_258_n N_VGND_c_363_n 0.0071386f $X=3.65 $Y=0.995 $X2=0 $Y2=0
cc_196 A1 N_A_321_47#_c_416_n 0.0374637f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A1_c_257_n N_A_321_47#_c_416_n 0.00460678f $X=3.65 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A1_c_258_n N_A_321_47#_c_416_n 0.0108508f $X=3.65 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_258_n N_A_321_47#_c_417_n 0.00630239f $X=3.65 $Y=0.995 $X2=0 $Y2=0
cc_200 X N_VPWR_c_303_n 0.0345427f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_201 X N_VPWR_c_306_n 0.0370719f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_202 N_X_M1002_s N_VPWR_c_302_n 0.00748091f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_203 X N_VPWR_c_302_n 0.0201416f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_204 N_X_c_282_n N_VGND_c_357_n 0.0238087f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_205 N_X_M1011_s N_VGND_c_363_n 0.00624411f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_206 N_X_c_282_n N_VGND_c_363_n 0.0130117f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_207 N_VPWR_c_302_n A_393_297# 0.0109267f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_208 N_VPWR_c_302_n A_511_297# 0.00915523f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_209 N_VPWR_c_302_n A_619_297# 0.0104998f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_210 N_VGND_c_363_n N_A_321_47#_M1004_d 0.00433464f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_211 N_VGND_c_363_n N_A_321_47#_M1005_d 0.00340968f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_363_n N_A_321_47#_M1003_d 0.00242111f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_361_n N_A_321_47#_c_442_n 0.00545209f $X=2.05 $Y=0 $X2=0 $Y2=0
cc_214 N_VGND_c_363_n N_A_321_47#_c_442_n 0.00583023f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_M1007_d N_A_321_47#_c_414_n 0.00305665f $X=2.025 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_VGND_c_355_n N_A_321_47#_c_414_n 0.0189571f $X=2.215 $Y=0.38 $X2=0
+ $Y2=0
cc_217 N_VGND_c_359_n N_A_321_47#_c_414_n 0.00233081f $X=3.125 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_361_n N_A_321_47#_c_414_n 0.00251982f $X=2.05 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_363_n N_A_321_47#_c_414_n 0.0107865f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_359_n N_A_321_47#_c_449_n 0.0211894f $X=3.125 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_363_n N_A_321_47#_c_449_n 0.0126169f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_M1010_d N_A_321_47#_c_416_n 0.00324783f $X=3.095 $Y=0.235 $X2=0
+ $Y2=0
cc_223 N_VGND_c_356_n N_A_321_47#_c_416_n 0.0196698f $X=3.29 $Y=0.38 $X2=0 $Y2=0
cc_224 N_VGND_c_359_n N_A_321_47#_c_416_n 0.00244976f $X=3.125 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_362_n N_A_321_47#_c_416_n 0.00204854f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_363_n N_A_321_47#_c_416_n 0.00984583f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_362_n N_A_321_47#_c_417_n 0.0209906f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_363_n N_A_321_47#_c_417_n 0.0125034f $X=3.91 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o21a_2.spice.SKY130_FD_SC_HD__O21A_2.pxi
* Created: Thu Aug 27 14:35:16 2020
* 
x_PM_SKY130_FD_SC_HD__O21A_2%A_79_21# N_A_79_21#_M1004_s N_A_79_21#_M1006_d
+ N_A_79_21#_c_53_n N_A_79_21#_M1003_g N_A_79_21#_M1001_g N_A_79_21#_c_54_n
+ N_A_79_21#_M1009_g N_A_79_21#_M1008_g N_A_79_21#_c_55_n N_A_79_21#_c_61_n
+ N_A_79_21#_c_65_p N_A_79_21#_c_86_p N_A_79_21#_c_56_n N_A_79_21#_c_57_n
+ N_A_79_21#_c_78_p N_A_79_21#_c_79_p N_A_79_21#_c_62_n N_A_79_21#_c_58_n
+ PM_SKY130_FD_SC_HD__O21A_2%A_79_21#
x_PM_SKY130_FD_SC_HD__O21A_2%B1 N_B1_M1004_g N_B1_M1006_g B1 N_B1_c_128_n
+ N_B1_c_129_n N_B1_c_130_n PM_SKY130_FD_SC_HD__O21A_2%B1
x_PM_SKY130_FD_SC_HD__O21A_2%A2 N_A2_M1007_g N_A2_M1002_g N_A2_c_164_n
+ N_A2_c_165_n A2 N_A2_c_166_n PM_SKY130_FD_SC_HD__O21A_2%A2
x_PM_SKY130_FD_SC_HD__O21A_2%A1 N_A1_c_208_n N_A1_M1005_g N_A1_M1000_g A1
+ N_A1_c_210_n PM_SKY130_FD_SC_HD__O21A_2%A1
x_PM_SKY130_FD_SC_HD__O21A_2%VPWR N_VPWR_M1001_d N_VPWR_M1008_d N_VPWR_M1000_d
+ N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n VPWR
+ N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_234_n
+ PM_SKY130_FD_SC_HD__O21A_2%VPWR
x_PM_SKY130_FD_SC_HD__O21A_2%X N_X_M1003_s N_X_M1001_s X N_X_c_283_n
+ PM_SKY130_FD_SC_HD__O21A_2%X
x_PM_SKY130_FD_SC_HD__O21A_2%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1007_d
+ N_VGND_c_300_n N_VGND_c_301_n N_VGND_c_302_n N_VGND_c_303_n VGND
+ N_VGND_c_304_n N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n
+ N_VGND_c_309_n PM_SKY130_FD_SC_HD__O21A_2%VGND
x_PM_SKY130_FD_SC_HD__O21A_2%A_384_47# N_A_384_47#_M1004_d N_A_384_47#_M1005_d
+ N_A_384_47#_c_352_n N_A_384_47#_c_355_n N_A_384_47#_c_351_n
+ PM_SKY130_FD_SC_HD__O21A_2%A_384_47#
cc_1 VNB N_A_79_21#_c_53_n 0.0215607f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_54_n 0.0190895f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_3 VNB N_A_79_21#_c_55_n 0.00225496f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.16
cc_4 VNB N_A_79_21#_c_56_n 0.0113762f $X=-0.19 $Y=-0.24 $X2=1.63 $Y2=0.635
cc_5 VNB N_A_79_21#_c_57_n 0.00486842f $X=-0.19 $Y=-0.24 $X2=1.63 $Y2=0.385
cc_6 VNB N_A_79_21#_c_58_n 0.063262f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.165
cc_7 VNB N_B1_c_128_n 0.0278553f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_8 VNB N_B1_c_129_n 0.0025398f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_9 VNB N_B1_c_130_n 0.0202542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A2_c_164_n 0.00607245f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_11 VNB N_A2_c_165_n 0.0218879f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_12 VNB N_A2_c_166_n 0.0168009f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.335
cc_13 VNB N_A1_c_208_n 0.0224385f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.235
cc_14 VNB A1 0.0137693f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB N_A1_c_210_n 0.0365663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_234_n 0.136896f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.33
cc_17 VNB N_X_c_283_n 6.33903e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.335
cc_18 VNB N_VGND_c_300_n 0.0101667f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.335
cc_19 VNB N_VGND_c_301_n 0.0378482f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_20 VNB N_VGND_c_302_n 0.00523275f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.56
cc_21 VNB N_VGND_c_303_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_304_n 0.0155725f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.16
cc_23 VNB N_VGND_c_305_n 0.026809f $X=-0.19 $Y=-0.24 $X2=1.275 $Y2=1.895
cc_24 VNB N_VGND_c_306_n 0.0160722f $X=-0.19 $Y=-0.24 $X2=2.06 $Y2=2.3
cc_25 VNB N_VGND_c_307_n 0.183653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_308_n 0.00510127f $X=-0.19 $Y=-0.24 $X2=2.095 $Y2=1.895
cc_27 VNB N_VGND_c_309_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.165
cc_28 VNB N_A_384_47#_c_351_n 0.0130293f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.56
cc_29 VPB N_A_79_21#_M1001_g 0.024604f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_30 VPB N_A_79_21#_M1008_g 0.0206041f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_31 VPB N_A_79_21#_c_61_n 0.00221288f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=1.785
cc_32 VPB N_A_79_21#_c_62_n 0.00531935f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.33
cc_33 VPB N_A_79_21#_c_58_n 0.0161708f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.165
cc_34 VPB N_B1_M1006_g 0.0225734f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_B1_c_128_n 0.00841604f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB N_B1_c_129_n 0.00127164f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A2_M1002_g 0.01892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A2_c_164_n 0.0055088f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_39 VPB N_A2_c_165_n 0.00619625f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_40 VPB A2 0.00138521f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.995
cc_41 VPB N_A1_M1000_g 0.0227219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB A1 0.00875776f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_43 VPB N_A1_c_210_n 0.0100499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_235_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.335
cc_45 VPB N_VPWR_c_236_n 0.0383544f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_46 VPB N_VPWR_c_237_n 0.0103006f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.995
cc_47 VPB N_VPWR_c_238_n 0.035072f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.56
cc_48 VPB N_VPWR_c_239_n 0.0256981f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.16
cc_49 VPB N_VPWR_c_240_n 0.0155667f $X=-0.19 $Y=1.305 $X2=2.06 $Y2=2.3
cc_50 VPB N_VPWR_c_241_n 0.0167584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_234_n 0.043034f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.33
cc_52 VPB N_X_c_283_n 0.00108493f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.335
cc_53 N_A_79_21#_c_61_n N_B1_M1006_g 0.00412643f $X=1.19 $Y=1.785 $X2=0 $Y2=0
cc_54 N_A_79_21#_c_65_p N_B1_M1006_g 0.015797f $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_55 N_A_79_21#_c_62_n N_B1_M1006_g 0.00102633f $X=1.11 $Y=1.33 $X2=0 $Y2=0
cc_56 N_A_79_21#_c_55_n N_B1_c_128_n 4.48662e-19 $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_79_21#_c_65_p N_B1_c_128_n 8.5331e-19 $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_58 N_A_79_21#_c_56_n N_B1_c_128_n 0.00547797f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_58_n N_B1_c_128_n 0.0176117f $X=0.895 $Y=1.165 $X2=0 $Y2=0
cc_60 N_A_79_21#_c_55_n N_B1_c_129_n 0.048325f $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_65_p N_B1_c_129_n 0.0283525f $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_56_n N_B1_c_129_n 0.0257333f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_58_n N_B1_c_129_n 0.00222428f $X=0.895 $Y=1.165 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_55_n N_B1_c_130_n 0.00353599f $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_56_n N_B1_c_130_n 0.00265201f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_57_n N_B1_c_130_n 0.00571981f $X=1.63 $Y=0.385 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_78_p N_A2_M1002_g 0.00298068f $X=2.095 $Y=2.005 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_79_p N_A2_M1002_g 0.00859804f $X=2.06 $Y=2.3 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_78_p N_A2_c_164_n 0.00814514f $X=2.095 $Y=2.005 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_78_p N_A2_c_165_n 2.1987e-19 $X=2.095 $Y=2.005 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_57_n N_A2_c_166_n 6.71456e-19 $X=1.63 $Y=0.385 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_79_p N_A1_M1000_g 0.00139349f $X=2.06 $Y=2.3 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_61_n N_VPWR_M1008_d 0.00964918f $X=1.19 $Y=1.785 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_65_p N_VPWR_M1008_d 0.0177752f $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_86_p N_VPWR_M1008_d 0.00642291f $X=1.275 $Y=1.895 $X2=0 $Y2=0
cc_76 N_A_79_21#_M1001_g N_VPWR_c_236_n 0.00573151f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_78_p N_VPWR_c_238_n 5.86816e-19 $X=2.095 $Y=2.005 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_79_p N_VPWR_c_238_n 0.0124858f $X=2.06 $Y=2.3 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_65_p N_VPWR_c_239_n 0.00208303f $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_79_p N_VPWR_c_239_n 0.0156896f $X=2.06 $Y=2.3 $X2=0 $Y2=0
cc_81 N_A_79_21#_M1001_g N_VPWR_c_240_n 0.00564131f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_79_21#_M1008_g N_VPWR_c_240_n 0.00486043f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_83 N_A_79_21#_M1001_g N_VPWR_c_241_n 4.96225e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_79_21#_M1008_g N_VPWR_c_241_n 0.00981811f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_85 N_A_79_21#_c_65_p N_VPWR_c_241_n 0.0346085f $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_86_p N_VPWR_c_241_n 0.0137948f $X=1.275 $Y=1.895 $X2=0 $Y2=0
cc_87 N_A_79_21#_M1006_d N_VPWR_c_234_n 0.00243647f $X=1.92 $Y=1.485 $X2=0 $Y2=0
cc_88 N_A_79_21#_M1001_g N_VPWR_c_234_n 0.0110238f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_79_21#_M1008_g N_VPWR_c_234_n 0.00816366f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_90 N_A_79_21#_c_65_p N_VPWR_c_234_n 0.00599596f $X=1.965 $Y=1.895 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_86_p N_VPWR_c_234_n 7.64972e-19 $X=1.275 $Y=1.895 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_79_p N_VPWR_c_234_n 0.00975383f $X=2.06 $Y=2.3 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_53_n N_X_c_283_n 0.0145651f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_79_21#_M1001_g N_X_c_283_n 0.0244565f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_54_n N_X_c_283_n 0.00193944f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_79_21#_M1008_g N_X_c_283_n 0.00243172f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_55_n N_X_c_283_n 0.034655f $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_61_n N_X_c_283_n 0.0141566f $X=1.19 $Y=1.785 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_58_n N_X_c_283_n 0.0307534f $X=0.895 $Y=1.165 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_55_n N_VGND_M1009_d 6.10963e-19 $X=1.11 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_56_n N_VGND_M1009_d 0.00348222f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_53_n N_VGND_c_301_n 0.00312525f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_53_n N_VGND_c_302_n 4.75139e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_54_n N_VGND_c_302_n 0.00767711f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_105 N_A_79_21#_c_56_n N_VGND_c_302_n 0.0208852f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_57_n N_VGND_c_302_n 0.0161705f $X=1.63 $Y=0.385 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_57_n N_VGND_c_303_n 0.00600743f $X=1.63 $Y=0.385 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_53_n N_VGND_c_304_n 0.00564131f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_54_n N_VGND_c_304_n 0.00486043f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_110 N_A_79_21#_c_56_n N_VGND_c_305_n 0.00354429f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_57_n N_VGND_c_305_n 0.0202676f $X=1.63 $Y=0.385 $X2=0 $Y2=0
cc_112 N_A_79_21#_M1004_s N_VGND_c_307_n 0.00213418f $X=1.505 $Y=0.235 $X2=0
+ $Y2=0
cc_113 N_A_79_21#_c_53_n N_VGND_c_307_n 0.0110238f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_54_n N_VGND_c_307_n 0.00821218f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_79_21#_c_56_n N_VGND_c_307_n 0.0069915f $X=1.63 $Y=0.635 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_57_n N_VGND_c_307_n 0.0122675f $X=1.63 $Y=0.385 $X2=0 $Y2=0
cc_117 N_B1_M1006_g N_A2_M1002_g 0.0233461f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B1_c_129_n N_A2_M1002_g 7.89099e-19 $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_c_128_n N_A2_c_164_n 0.00261027f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_c_129_n N_A2_c_164_n 0.0315002f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B1_c_128_n N_A2_c_165_n 0.0210165f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B1_c_129_n N_A2_c_165_n 3.70396e-19 $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_123 N_B1_c_129_n A2 0.00458368f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_124 N_B1_c_130_n N_A2_c_166_n 0.023072f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B1_c_129_n N_VPWR_M1008_d 0.00508292f $X=1.69 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B1_M1006_g N_VPWR_c_239_n 0.00362954f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B1_M1006_g N_VPWR_c_241_n 0.00996925f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B1_M1006_g N_VPWR_c_234_n 0.00428526f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B1_c_130_n N_VGND_c_302_n 0.00233012f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_130_n N_VGND_c_303_n 0.00167142f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_130_n N_VGND_c_305_n 0.00547881f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_130_n N_VGND_c_307_n 0.0112188f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_166_n N_A1_c_208_n 0.0218582f $X=2.295 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A2_M1002_g N_A1_M1000_g 0.0423381f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_135 A2 N_A1_M1000_g 0.00806207f $X=2.44 $Y=1.785 $X2=0 $Y2=0
cc_136 N_A2_c_164_n A1 0.0230042f $X=2.405 $Y=1.212 $X2=0 $Y2=0
cc_137 N_A2_c_165_n A1 3.67608e-19 $X=2.295 $Y=1.16 $X2=0 $Y2=0
cc_138 A2 A1 0.00293999f $X=2.44 $Y=1.785 $X2=0 $Y2=0
cc_139 N_A2_c_164_n N_A1_c_210_n 0.00355634f $X=2.405 $Y=1.212 $X2=0 $Y2=0
cc_140 N_A2_c_165_n N_A1_c_210_n 0.0210605f $X=2.295 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_M1002_g N_VPWR_c_238_n 0.00260307f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_142 A2 N_VPWR_c_238_n 0.0234683f $X=2.44 $Y=1.785 $X2=0 $Y2=0
cc_143 N_A2_M1002_g N_VPWR_c_239_n 0.0054895f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_144 A2 N_VPWR_c_239_n 0.00318925f $X=2.44 $Y=1.785 $X2=0 $Y2=0
cc_145 N_A2_M1002_g N_VPWR_c_241_n 0.00113943f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A2_M1002_g N_VPWR_c_234_n 0.0100878f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_147 A2 N_VPWR_c_234_n 0.00566607f $X=2.44 $Y=1.785 $X2=0 $Y2=0
cc_148 A2 A_470_297# 0.0136633f $X=2.44 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_149 N_A2_c_166_n N_VGND_c_303_n 0.00807531f $X=2.295 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A2_c_166_n N_VGND_c_305_n 0.00410216f $X=2.295 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A2_c_166_n N_VGND_c_307_n 0.00475398f $X=2.295 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_164_n N_A_384_47#_c_352_n 0.027146f $X=2.405 $Y=1.212 $X2=0 $Y2=0
cc_153 N_A2_c_165_n N_A_384_47#_c_352_n 0.0023628f $X=2.295 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_c_166_n N_A_384_47#_c_352_n 0.0105491f $X=2.295 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A2_c_164_n N_A_384_47#_c_355_n 0.00974409f $X=2.405 $Y=1.212 $X2=0
+ $Y2=0
cc_156 N_A2_c_165_n N_A_384_47#_c_355_n 9.30233e-19 $X=2.295 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_M1000_g N_VPWR_c_238_n 0.0219476f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_158 A1 N_VPWR_c_238_n 0.0196616f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A1_c_210_n N_VPWR_c_238_n 0.00139451f $X=2.975 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_M1000_g N_VPWR_c_239_n 0.00486043f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A1_M1000_g N_VPWR_c_234_n 0.00842581f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A1_c_208_n N_VGND_c_303_n 0.0137629f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_208_n N_VGND_c_306_n 0.00410216f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_208_n N_VGND_c_307_n 0.00569615f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_208_n N_A_384_47#_c_352_n 0.0148746f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_166 A1 N_A_384_47#_c_351_n 0.0199632f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A1_c_210_n N_A_384_47#_c_351_n 0.00178274f $X=2.975 $Y=1.16 $X2=0 $Y2=0
cc_168 N_VPWR_c_234_n N_X_M1001_s 0.00375437f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_240_n N_X_c_283_n 0.0146562f $X=0.945 $Y=2.495 $X2=0 $Y2=0
cc_170 N_VPWR_c_234_n N_X_c_283_n 0.00922188f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_171 N_VPWR_c_234_n A_470_297# 0.00766774f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_172 N_X_c_283_n N_VGND_c_304_n 0.0146562f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_173 N_X_M1003_s N_VGND_c_307_n 0.00375437f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_174 N_X_c_283_n N_VGND_c_307_n 0.00922188f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_175 N_VGND_c_307_n N_A_384_47#_M1004_d 0.00421987f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_176 N_VGND_c_307_n N_A_384_47#_M1005_d 0.00264396f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_177 N_VGND_M1007_d N_A_384_47#_c_352_n 0.00430242f $X=2.35 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_VGND_c_303_n N_A_384_47#_c_352_n 0.0163248f $X=2.51 $Y=0.38 $X2=0 $Y2=0
cc_179 N_VGND_c_305_n N_A_384_47#_c_352_n 0.00261733f $X=2.345 $Y=0 $X2=0 $Y2=0
cc_180 N_VGND_c_306_n N_A_384_47#_c_352_n 0.00261733f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_181 N_VGND_c_307_n N_A_384_47#_c_352_n 0.0097386f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_182 N_VGND_c_305_n N_A_384_47#_c_355_n 0.00533689f $X=2.345 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_c_307_n N_A_384_47#_c_355_n 0.00689411f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_184 N_VGND_c_306_n N_A_384_47#_c_351_n 0.00671053f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_185 N_VGND_c_307_n N_A_384_47#_c_351_n 0.0088263f $X=2.99 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nor2b_2.spice.SKY130_FD_SC_HD__NOR2B_2.pxi
* Created: Thu Aug 27 14:31:45 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2B_2%A N_A_c_63_n N_A_M1003_g N_A_M1001_g N_A_c_64_n
+ N_A_M1005_g N_A_M1008_g A N_A_c_65_n PM_SKY130_FD_SC_HD__NOR2B_2%A
x_PM_SKY130_FD_SC_HD__NOR2B_2%A_251_21# N_A_251_21#_M1000_s N_A_251_21#_M1009_s
+ N_A_251_21#_c_100_n N_A_251_21#_M1002_g N_A_251_21#_M1006_g
+ N_A_251_21#_c_101_n N_A_251_21#_M1004_g N_A_251_21#_M1007_g
+ N_A_251_21#_c_102_n N_A_251_21#_c_103_n N_A_251_21#_c_104_n
+ N_A_251_21#_c_105_n N_A_251_21#_c_106_n N_A_251_21#_c_107_n
+ N_A_251_21#_c_115_n N_A_251_21#_c_108_n N_A_251_21#_c_109_n
+ N_A_251_21#_c_116_n PM_SKY130_FD_SC_HD__NOR2B_2%A_251_21#
x_PM_SKY130_FD_SC_HD__NOR2B_2%B_N N_B_N_M1000_g N_B_N_M1009_g B_N B_N B_N
+ N_B_N_c_186_n N_B_N_c_187_n PM_SKY130_FD_SC_HD__NOR2B_2%B_N
x_PM_SKY130_FD_SC_HD__NOR2B_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1008_s
+ N_A_27_297#_M1007_d N_A_27_297#_c_219_n N_A_27_297#_c_220_n
+ N_A_27_297#_c_221_n N_A_27_297#_c_222_n N_A_27_297#_c_246_p
+ N_A_27_297#_c_231_n N_A_27_297#_c_223_n N_A_27_297#_c_224_n
+ N_A_27_297#_c_225_n PM_SKY130_FD_SC_HD__NOR2B_2%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR2B_2%VPWR N_VPWR_M1001_d N_VPWR_M1009_d N_VPWR_c_264_n
+ N_VPWR_c_265_n N_VPWR_c_266_n VPWR N_VPWR_c_267_n N_VPWR_c_268_n
+ N_VPWR_c_269_n N_VPWR_c_263_n PM_SKY130_FD_SC_HD__NOR2B_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR2B_2%Y N_Y_M1003_s N_Y_M1002_d N_Y_M1006_s N_Y_c_309_n
+ N_Y_c_304_n N_Y_c_305_n N_Y_c_306_n N_Y_c_307_n Y N_Y_c_319_n
+ PM_SKY130_FD_SC_HD__NOR2B_2%Y
x_PM_SKY130_FD_SC_HD__NOR2B_2%VGND N_VGND_M1003_d N_VGND_M1005_d N_VGND_M1004_s
+ N_VGND_M1000_d N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n
+ N_VGND_c_363_n VGND N_VGND_c_364_n N_VGND_c_365_n
+ PM_SKY130_FD_SC_HD__NOR2B_2%VGND
cc_1 VNB N_A_c_63_n 0.0216649f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_64_n 0.0160882f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A_c_65_n 0.0436153f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_4 VNB N_A_251_21#_c_100_n 0.0160831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_251_21#_c_101_n 0.0195312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_251_21#_c_102_n 0.0273917f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_7 VNB N_A_251_21#_c_103_n 6.18364e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_251_21#_c_104_n 0.0335288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_251_21#_c_105_n 0.00440548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_251_21#_c_106_n 0.00106425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_251_21#_c_107_n 0.00209644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_251_21#_c_108_n 0.00656081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_251_21#_c_109_n 0.00296896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB B_N 0.0165774f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_15 VNB B_N 0.00131519f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_16 VNB N_B_N_c_186_n 0.029221f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_17 VNB N_B_N_c_187_n 0.0404958f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_18 VNB N_VPWR_c_263_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_304_n 0.00429176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_305_n 0.00222618f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_21 VNB N_Y_c_306_n 0.00181222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_307_n 8.0856e-19 $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_23 VNB N_VGND_c_354_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_24 VNB N_VGND_c_355_n 0.0345494f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_25 VNB N_VGND_c_356_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_26 VNB N_VGND_c_357_n 0.00536469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_358_n 0.0131666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_359_n 0.0314647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_360_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_361_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_362_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_363_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_364_n 0.0213925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_365_n 0.194897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_M1001_g 0.025044f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_36 VPB N_A_M1008_g 0.0183967f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_37 VPB N_A_c_65_n 0.0047988f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_38 VPB N_A_251_21#_M1006_g 0.0187755f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_39 VPB N_A_251_21#_M1007_g 0.0224801f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_40 VPB N_A_251_21#_c_102_n 0.00417579f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_41 VPB N_A_251_21#_c_104_n 0.0129763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_251_21#_c_106_n 0.0035431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_251_21#_c_115_n 0.0107634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_251_21#_c_116_n 0.0116985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B_N_M1009_g 0.0622965f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_46 VPB B_N 0.0352637f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_47 VPB N_B_N_c_186_n 0.00841919f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_48 VPB N_A_27_297#_c_219_n 0.0151088f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_49 VPB N_A_27_297#_c_220_n 0.0318598f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_50 VPB N_A_27_297#_c_221_n 0.00264631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_297#_c_222_n 0.00424874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_223_n 0.00610479f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_53 VPB N_A_27_297#_c_224_n 0.00186102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_297#_c_225_n 0.00454996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_264_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_56 VPB N_VPWR_c_265_n 0.0128556f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.325
cc_57 VPB N_VPWR_c_266_n 0.00517963f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_58 VPB N_VPWR_c_267_n 0.0174493f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_59 VPB N_VPWR_c_268_n 0.0495297f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_60 VPB N_VPWR_c_269_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_263_n 0.0546744f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_Y_c_306_n 0.00266976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 N_A_c_64_n N_A_251_21#_c_100_n 0.0192417f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A_M1008_g N_A_251_21#_M1006_g 0.0192417f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_65 A N_A_251_21#_c_102_n 8.91259e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_66 N_A_c_65_n N_A_251_21#_c_102_n 0.0192417f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_A_27_297#_c_221_n 0.0169301f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_M1008_g N_A_27_297#_c_221_n 0.0153285f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_69 A N_A_27_297#_c_221_n 0.0318513f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_65_n N_A_27_297#_c_221_n 0.00215121f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_M1001_g N_VPWR_c_264_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_M1008_g N_VPWR_c_264_n 0.00302074f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_M1001_g N_VPWR_c_267_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_M1008_g N_VPWR_c_268_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1001_g N_VPWR_c_263_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1008_g N_VPWR_c_263_n 0.010464f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_c_63_n N_Y_c_309_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_c_64_n N_Y_c_309_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_c_64_n N_Y_c_304_n 0.0092324f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_80 A N_Y_c_304_n 0.0037556f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_c_63_n N_Y_c_305_n 0.00240075f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_c_64_n N_Y_c_305_n 9.88607e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_83 A N_Y_c_305_n 0.0265925f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A_c_65_n N_Y_c_305_n 0.00227419f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_85 A N_Y_c_306_n 0.00655643f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_65_n N_Y_c_306_n 0.001358f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_c_64_n N_Y_c_319_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_c_63_n N_VGND_c_355_n 0.00344836f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_c_64_n N_VGND_c_356_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_c_63_n N_VGND_c_360_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_c_64_n N_VGND_c_360_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A_c_63_n N_VGND_c_365_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_64_n N_VGND_c_365_n 0.0057435f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_251_21#_c_115_n N_B_N_M1009_g 0.012849f $X=2.48 $Y=2.28 $X2=0 $Y2=0
cc_95 N_A_251_21#_c_116_n N_B_N_M1009_g 0.0042507f $X=2.48 $Y=1.53 $X2=0 $Y2=0
cc_96 N_A_251_21#_c_104_n B_N 4.9878e-19 $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_251_21#_c_105_n B_N 7.17163e-19 $X=2.322 $Y=1.075 $X2=0 $Y2=0
cc_98 N_A_251_21#_c_106_n B_N 0.00235945f $X=2.345 $Y=1.445 $X2=0 $Y2=0
cc_99 N_A_251_21#_c_109_n B_N 0.0153846f $X=2.322 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_251_21#_c_106_n B_N 0.00629384f $X=2.345 $Y=1.445 $X2=0 $Y2=0
cc_101 N_A_251_21#_c_115_n B_N 0.0163902f $X=2.48 $Y=2.28 $X2=0 $Y2=0
cc_102 N_A_251_21#_c_116_n B_N 0.00824612f $X=2.48 $Y=1.53 $X2=0 $Y2=0
cc_103 N_A_251_21#_c_104_n N_B_N_c_186_n 0.00848254f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_251_21#_c_106_n N_B_N_c_186_n 0.00326297f $X=2.345 $Y=1.445 $X2=0
+ $Y2=0
cc_105 N_A_251_21#_c_109_n N_B_N_c_186_n 6.87544e-19 $X=2.322 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_A_251_21#_c_105_n N_B_N_c_187_n 0.00509776f $X=2.322 $Y=1.075 $X2=0
+ $Y2=0
cc_107 N_A_251_21#_c_107_n N_B_N_c_187_n 8.35068e-19 $X=2.48 $Y=0.725 $X2=0
+ $Y2=0
cc_108 N_A_251_21#_c_108_n N_B_N_c_187_n 5.53506e-19 $X=2.48 $Y=0.81 $X2=0 $Y2=0
cc_109 N_A_251_21#_M1006_g N_A_27_297#_c_222_n 3.45391e-19 $X=1.33 $Y=1.985
+ $X2=0 $Y2=0
cc_110 N_A_251_21#_M1006_g N_A_27_297#_c_231_n 0.0121747f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_251_21#_M1007_g N_A_27_297#_c_231_n 0.0121306f $X=1.75 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_251_21#_M1007_g N_A_27_297#_c_223_n 9.36283e-19 $X=1.75 $Y=1.985
+ $X2=0 $Y2=0
cc_113 N_A_251_21#_c_103_n N_A_27_297#_c_223_n 0.0152874f $X=2.215 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_A_251_21#_c_104_n N_A_27_297#_c_223_n 0.00724241f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_A_251_21#_c_115_n N_A_27_297#_c_223_n 0.0142206f $X=2.48 $Y=2.28 $X2=0
+ $Y2=0
cc_116 N_A_251_21#_c_116_n N_A_27_297#_c_223_n 0.0137022f $X=2.48 $Y=1.53 $X2=0
+ $Y2=0
cc_117 N_A_251_21#_c_103_n N_A_27_297#_c_224_n 9.87727e-19 $X=2.215 $Y=1.16
+ $X2=0 $Y2=0
cc_118 N_A_251_21#_c_104_n N_A_27_297#_c_224_n 6.15165e-19 $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_119 N_A_251_21#_c_115_n N_A_27_297#_c_224_n 0.0226471f $X=2.48 $Y=2.28 $X2=0
+ $Y2=0
cc_120 N_A_251_21#_c_115_n N_A_27_297#_c_225_n 0.00984577f $X=2.48 $Y=2.28 $X2=0
+ $Y2=0
cc_121 N_A_251_21#_M1006_g N_VPWR_c_268_n 0.00357877f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_251_21#_M1007_g N_VPWR_c_268_n 0.00357877f $X=1.75 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_251_21#_c_115_n N_VPWR_c_268_n 0.0112447f $X=2.48 $Y=2.28 $X2=0 $Y2=0
cc_124 N_A_251_21#_M1009_s N_VPWR_c_263_n 0.00529598f $X=2.355 $Y=2.065 $X2=0
+ $Y2=0
cc_125 N_A_251_21#_M1006_g N_VPWR_c_263_n 0.00525237f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_251_21#_M1007_g N_VPWR_c_263_n 0.00655123f $X=1.75 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_251_21#_c_115_n N_VPWR_c_263_n 0.00645481f $X=2.48 $Y=2.28 $X2=0
+ $Y2=0
cc_128 N_A_251_21#_c_100_n N_Y_c_309_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_251_21#_c_100_n N_Y_c_304_n 0.0120621f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_251_21#_c_100_n N_Y_c_306_n 0.00267866f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_251_21#_M1006_g N_Y_c_306_n 0.00355132f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_251_21#_c_101_n N_Y_c_306_n 0.0013426f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_251_21#_M1007_g N_Y_c_306_n 0.00199909f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_251_21#_c_102_n N_Y_c_306_n 0.0238478f $X=1.825 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_251_21#_c_103_n N_Y_c_306_n 0.0109102f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_251_21#_c_105_n N_Y_c_306_n 0.00589498f $X=2.322 $Y=1.075 $X2=0 $Y2=0
cc_137 N_A_251_21#_c_106_n N_Y_c_306_n 0.00610516f $X=2.345 $Y=1.445 $X2=0 $Y2=0
cc_138 N_A_251_21#_c_100_n N_Y_c_307_n 0.00206444f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_251_21#_c_101_n N_Y_c_307_n 0.00345997f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_251_21#_c_100_n N_Y_c_319_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_251_21#_c_101_n N_Y_c_319_n 0.00539651f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_251_21#_c_100_n N_VGND_c_356_n 0.00146448f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_251_21#_c_101_n N_VGND_c_357_n 0.00338128f $X=1.75 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A_251_21#_c_103_n N_VGND_c_357_n 0.0129839f $X=2.215 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_251_21#_c_104_n N_VGND_c_357_n 0.00429275f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_251_21#_c_107_n N_VGND_c_357_n 0.0119909f $X=2.48 $Y=0.725 $X2=0
+ $Y2=0
cc_147 N_A_251_21#_c_108_n N_VGND_c_357_n 0.0132324f $X=2.48 $Y=0.81 $X2=0 $Y2=0
cc_148 N_A_251_21#_c_107_n N_VGND_c_359_n 0.00127149f $X=2.48 $Y=0.725 $X2=0
+ $Y2=0
cc_149 N_A_251_21#_c_100_n N_VGND_c_362_n 0.00423334f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A_251_21#_c_101_n N_VGND_c_362_n 0.00541359f $X=1.75 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A_251_21#_c_107_n N_VGND_c_364_n 0.00509579f $X=2.48 $Y=0.725 $X2=0
+ $Y2=0
cc_152 N_A_251_21#_c_108_n N_VGND_c_364_n 0.00273515f $X=2.48 $Y=0.81 $X2=0
+ $Y2=0
cc_153 N_A_251_21#_c_100_n N_VGND_c_365_n 0.0057435f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A_251_21#_c_101_n N_VGND_c_365_n 0.0108276f $X=1.75 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_A_251_21#_c_107_n N_VGND_c_365_n 0.0055979f $X=2.48 $Y=0.725 $X2=0
+ $Y2=0
cc_156 N_A_251_21#_c_108_n N_VGND_c_365_n 0.00480544f $X=2.48 $Y=0.81 $X2=0
+ $Y2=0
cc_157 N_B_N_M1009_g N_A_27_297#_c_223_n 8.49741e-19 $X=2.69 $Y=2.275 $X2=0
+ $Y2=0
cc_158 B_N N_VPWR_c_265_n 0.00159942f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_159 N_B_N_M1009_g N_VPWR_c_266_n 0.00482366f $X=2.69 $Y=2.275 $X2=0 $Y2=0
cc_160 B_N N_VPWR_c_266_n 0.00955496f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_161 N_B_N_M1009_g N_VPWR_c_268_n 0.00585385f $X=2.69 $Y=2.275 $X2=0 $Y2=0
cc_162 N_B_N_M1009_g N_VPWR_c_263_n 0.0128967f $X=2.69 $Y=2.275 $X2=0 $Y2=0
cc_163 B_N N_VPWR_c_263_n 0.00322535f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_164 N_B_N_c_187_n N_VGND_c_357_n 0.00722462f $X=2.757 $Y=0.995 $X2=0 $Y2=0
cc_165 B_N N_VGND_c_359_n 0.0161764f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_166 N_B_N_c_186_n N_VGND_c_359_n 0.00287932f $X=2.765 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B_N_c_187_n N_VGND_c_359_n 0.0146349f $X=2.757 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B_N_c_187_n N_VGND_c_364_n 0.00585385f $X=2.757 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B_N_c_187_n N_VGND_c_365_n 0.0130111f $X=2.757 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_27_297#_c_221_n N_VPWR_M1001_d 0.00166915f $X=0.995 $Y=1.55 $X2=-0.19
+ $Y2=1.305
cc_171 N_A_27_297#_c_221_n N_VPWR_c_264_n 0.0128751f $X=0.995 $Y=1.55 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_c_220_n N_VPWR_c_267_n 0.0208267f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_173 N_A_27_297#_c_246_p N_VPWR_c_268_n 0.0143053f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_c_231_n N_VPWR_c_268_n 0.0330174f $X=1.835 $Y=2.38 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_c_225_n N_VPWR_c_268_n 0.0187799f $X=1.98 $Y=2.295 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_M1001_s N_VPWR_c_263_n 0.00260431f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_M1008_s N_VPWR_c_263_n 0.00246446f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_M1007_d N_VPWR_c_263_n 0.0020932f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_179 N_A_27_297#_c_220_n N_VPWR_c_263_n 0.0122467f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_246_p N_VPWR_c_263_n 0.00962794f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_181 N_A_27_297#_c_231_n N_VPWR_c_263_n 0.0204627f $X=1.835 $Y=2.38 $X2=0
+ $Y2=0
cc_182 N_A_27_297#_c_225_n N_VPWR_c_263_n 0.0111575f $X=1.98 $Y=2.295 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_231_n N_Y_M1006_s 0.00312348f $X=1.835 $Y=2.38 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_221_n N_Y_c_304_n 0.00202983f $X=0.995 $Y=1.55 $X2=0 $Y2=0
cc_185 N_A_27_297#_c_222_n N_Y_c_304_n 0.00932875f $X=1.12 $Y=1.655 $X2=0 $Y2=0
cc_186 N_A_27_297#_c_222_n N_Y_c_306_n 0.0033804f $X=1.12 $Y=1.655 $X2=0 $Y2=0
cc_187 N_A_27_297#_c_231_n N_Y_c_306_n 0.0118865f $X=1.835 $Y=2.38 $X2=0 $Y2=0
cc_188 N_A_27_297#_c_223_n N_Y_c_306_n 0.0031162f $X=1.96 $Y=1.63 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_219_n N_VGND_c_355_n 0.0114749f $X=0.245 $Y=1.655 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_263_n N_Y_M1006_s 0.00216833f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_191 N_Y_c_304_n N_VGND_M1005_d 0.00161804f $X=1.375 $Y=0.81 $X2=0 $Y2=0
cc_192 N_Y_c_305_n N_VGND_c_355_n 0.00752789f $X=0.865 $Y=0.81 $X2=0 $Y2=0
cc_193 N_Y_c_304_n N_VGND_c_356_n 0.0122105f $X=1.375 $Y=0.81 $X2=0 $Y2=0
cc_194 N_Y_c_307_n N_VGND_c_357_n 0.00750114f $X=1.54 $Y=0.81 $X2=0 $Y2=0
cc_195 N_Y_c_309_n N_VGND_c_360_n 0.0188385f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_196 N_Y_c_304_n N_VGND_c_360_n 0.00198102f $X=1.375 $Y=0.81 $X2=0 $Y2=0
cc_197 N_Y_c_304_n N_VGND_c_362_n 0.00198102f $X=1.375 $Y=0.81 $X2=0 $Y2=0
cc_198 N_Y_c_319_n N_VGND_c_362_n 0.0188871f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_199 N_Y_M1003_s N_VGND_c_365_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_200 N_Y_M1002_d N_VGND_c_365_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_201 N_Y_c_309_n N_VGND_c_365_n 0.0122019f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_202 N_Y_c_304_n N_VGND_c_365_n 0.00833546f $X=1.375 $Y=0.81 $X2=0 $Y2=0
cc_203 N_Y_c_319_n N_VGND_c_365_n 0.0122172f $X=1.54 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__ebufn_4.pex.spice
* Created: Tue Sep  1 19:07:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EBUFN_4%A 3 6 8 9 13 15
c33 6 0 8.64755e-20 $X=0.47 $Y=1.985
r34 13 16 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.552 $Y=1.16
+ $X2=0.552 $Y2=1.325
r35 13 15 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.552 $Y=1.16
+ $X2=0.552 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.16 $X2=0.575 $Y2=1.16
r37 9 14 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.635 $Y=1.53
+ $X2=0.635 $Y2=1.16
r38 8 14 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=0.635 $Y=0.85
+ $X2=0.635 $Y2=1.16
r39 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r40 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%TE_B 3 5 7 8 9 10 12 13 15 17 18 20 22 23 25
+ 27 28 29 30 31
c84 31 0 8.64755e-20 $X=1.155 $Y=0.85
r85 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.16 $X2=1.115 $Y2=1.16
r86 33 35 19.4094 $w=2.98e-07 $l=1.2e-07 $layer=POLY_cond $X=0.995 $Y=1.247
+ $X2=1.115 $Y2=1.247
r87 31 36 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.115 $Y=0.85
+ $X2=1.115 $Y2=1.16
r88 25 27 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.195 $Y=1.47
+ $X2=3.195 $Y2=2.015
r89 24 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.85 $Y=1.395
+ $X2=2.775 $Y2=1.395
r90 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.12 $Y=1.395
+ $X2=3.195 $Y2=1.47
r91 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.12 $Y=1.395
+ $X2=2.85 $Y2=1.395
r92 20 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.775 $Y=1.47
+ $X2=2.775 $Y2=1.395
r93 20 22 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.775 $Y=1.47
+ $X2=2.775 $Y2=2.015
r94 19 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.43 $Y=1.395
+ $X2=2.355 $Y2=1.395
r95 18 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.395
+ $X2=2.775 $Y2=1.395
r96 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.7 $Y=1.395
+ $X2=2.43 $Y2=1.395
r97 15 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=1.47
+ $X2=2.355 $Y2=1.395
r98 15 17 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.355 $Y=1.47
+ $X2=2.355 $Y2=2.015
r99 14 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=1.395
+ $X2=1.935 $Y2=1.395
r100 13 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=1.395
+ $X2=2.355 $Y2=1.395
r101 13 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.28 $Y=1.395
+ $X2=2.01 $Y2=1.395
r102 10 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.47
+ $X2=1.935 $Y2=1.395
r103 10 12 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.935 $Y=1.47
+ $X2=1.935 $Y2=2.015
r104 9 35 89.5107 $w=2.98e-07 $l=5.49036e-07 $layer=POLY_cond $X=1.595 $Y=1.395
+ $X2=1.115 $Y2=1.247
r105 8 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.86 $Y=1.395
+ $X2=1.935 $Y2=1.395
r106 8 9 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.86 $Y=1.395
+ $X2=1.595 $Y2=1.395
r107 5 33 18.8112 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.247
r108 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.985
r109 1 33 18.8112 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.995 $Y=1.025
+ $X2=0.995 $Y2=1.247
r110 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.995 $Y=1.025
+ $X2=0.995 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%A_214_47# 1 2 7 9 10 11 12 14 15 17 19 20 24
+ 25 26 27 33 36 38 41 48 49 50
c94 50 0 8.82398e-20 $X=3.645 $Y=0.96
c95 49 0 9.17735e-20 $X=3.645 $Y=1.035
r96 49 50 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.645 $Y=1.035
+ $X2=3.645 $Y2=0.96
r97 42 49 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.645 $Y=1.16
+ $X2=3.645 $Y2=1.035
r98 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.645
+ $Y=1.16 $X2=3.645 $Y2=1.16
r99 39 48 1.68792 $w=2.5e-07 $l=1.38e-07 $layer=LI1_cond $X=1.725 $Y=1.15
+ $X2=1.587 $Y2=1.15
r100 39 41 88.5076 $w=2.48e-07 $l=1.92e-06 $layer=LI1_cond $X=1.725 $Y=1.15
+ $X2=3.645 $Y2=1.15
r101 37 48 4.76867 $w=2.75e-07 $l=1.25e-07 $layer=LI1_cond $X=1.587 $Y=1.275
+ $X2=1.587 $Y2=1.15
r102 37 38 13.4102 $w=2.73e-07 $l=3.2e-07 $layer=LI1_cond $X=1.587 $Y=1.275
+ $X2=1.587 $Y2=1.595
r103 36 48 4.76867 $w=2.75e-07 $l=1.25e-07 $layer=LI1_cond $X=1.587 $Y=1.025
+ $X2=1.587 $Y2=1.15
r104 35 36 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=1.587 $Y=0.595
+ $X2=1.587 $Y2=1.025
r105 31 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.227 $Y=1.68
+ $X2=1.587 $Y2=1.68
r106 31 33 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=1.227 $Y=1.765
+ $X2=1.227 $Y2=1.96
r107 27 35 6.916 $w=3.4e-07 $l=2.28451e-07 $layer=LI1_cond $X=1.45 $Y=0.425
+ $X2=1.587 $Y2=0.595
r108 27 29 8.30437 $w=3.38e-07 $l=2.45e-07 $layer=LI1_cond $X=1.45 $Y=0.425
+ $X2=1.205 $Y2=0.425
r109 24 50 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.56 $Y=0.56 $X2=3.56
+ $Y2=0.96
r110 21 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.215 $Y=1.035
+ $X2=3.14 $Y2=1.035
r111 20 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.035
+ $X2=3.645 $Y2=1.035
r112 20 21 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.48 $Y=1.035
+ $X2=3.215 $Y2=1.035
r113 17 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.14 $Y=0.96
+ $X2=3.14 $Y2=1.035
r114 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.14 $Y=0.96 $X2=3.14
+ $Y2=0.56
r115 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.795 $Y=1.035
+ $X2=2.72 $Y2=1.035
r116 15 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.065 $Y=1.035
+ $X2=3.14 $Y2=1.035
r117 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.065 $Y=1.035
+ $X2=2.795 $Y2=1.035
r118 12 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.72 $Y=0.96
+ $X2=2.72 $Y2=1.035
r119 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.72 $Y=0.96 $X2=2.72
+ $Y2=0.56
r120 10 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.645 $Y=1.035
+ $X2=2.72 $Y2=1.035
r121 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.645 $Y=1.035
+ $X2=2.375 $Y2=1.035
r122 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.3 $Y=0.96
+ $X2=2.375 $Y2=1.035
r123 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.3 $Y=0.96 $X2=2.3
+ $Y2=0.56
r124 2 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.205 $Y2=1.96
r125 1 29 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.205 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 39 41 45
+ 50 51 54 57 69 70
c99 57 0 2.39919e-19 $X=4.395 $Y=1.19
r100 68 70 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.27 $Y=1.16 $X2=5.36
+ $Y2=1.16
r101 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.27
+ $Y=1.16 $X2=5.27 $Y2=1.16
r102 66 68 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=4.94 $Y=1.16
+ $X2=5.27 $Y2=1.16
r103 65 66 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.52 $Y=1.16
+ $X2=4.94 $Y2=1.16
r104 64 69 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=4.25 $Y=1.15
+ $X2=5.27 $Y2=1.15
r105 63 65 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.52 $Y2=1.16
r106 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.25
+ $Y=1.16 $X2=4.25 $Y2=1.16
r107 60 63 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=4.1 $Y=1.16
+ $X2=4.25 $Y2=1.16
r108 57 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.395 $Y=1.19
+ $X2=4.395 $Y2=1.19
r109 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.19
+ $X2=0.235 $Y2=1.19
r110 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.38 $Y=1.19
+ $X2=0.235 $Y2=1.19
r111 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.25 $Y=1.19
+ $X2=4.395 $Y2=1.19
r112 50 51 4.7896 $w=1.4e-07 $l=3.87e-06 $layer=MET1_cond $X=4.25 $Y=1.19
+ $X2=0.38 $Y2=1.19
r113 49 54 28.1981 $w=2.33e-07 $l=5.75e-07 $layer=LI1_cond $X=0.202 $Y=1.765
+ $X2=0.202 $Y2=1.19
r114 47 54 25.7461 $w=2.33e-07 $l=5.25e-07 $layer=LI1_cond $X=0.202 $Y=0.665
+ $X2=0.202 $Y2=1.19
r115 45 47 9.88221 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.215 $Y=0.445
+ $X2=0.215 $Y2=0.665
r116 39 49 5.89299 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.895
+ $X2=0.215 $Y2=1.765
r117 39 41 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.215 $Y=1.895
+ $X2=0.215 $Y2=1.96
r118 35 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.36 $Y=1.295
+ $X2=5.36 $Y2=1.16
r119 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.36 $Y=1.295
+ $X2=5.36 $Y2=1.985
r120 31 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.36 $Y=1.025
+ $X2=5.36 $Y2=1.16
r121 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.36 $Y=1.025
+ $X2=5.36 $Y2=0.56
r122 27 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.94 $Y=1.295
+ $X2=4.94 $Y2=1.16
r123 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.94 $Y=1.295
+ $X2=4.94 $Y2=1.985
r124 23 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.94 $Y=1.025
+ $X2=4.94 $Y2=1.16
r125 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.94 $Y=1.025
+ $X2=4.94 $Y2=0.56
r126 19 65 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.52 $Y=1.295
+ $X2=4.52 $Y2=1.16
r127 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.52 $Y=1.295
+ $X2=4.52 $Y2=1.985
r128 15 65 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.52 $Y=1.025
+ $X2=4.52 $Y2=1.16
r129 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.52 $Y=1.025
+ $X2=4.52 $Y2=0.56
r130 11 60 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.1 $Y=1.295
+ $X2=4.1 $Y2=1.16
r131 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.1 $Y=1.295
+ $X2=4.1 $Y2=1.985
r132 7 60 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.1 $Y=1.025
+ $X2=4.1 $Y2=1.16
r133 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.1 $Y=1.025 $X2=4.1
+ $Y2=0.56
r134 2 41 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r135 1 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%VPWR 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r75 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r76 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r77 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r79 42 45 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=5.75 $Y2=2.72
r80 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 41 44 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=5.75 $Y2=2.72
r82 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=2.72
+ $X2=2.985 $Y2=2.72
r84 39 41 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.15 $Y=2.72 $X2=3.45
+ $Y2=2.72
r85 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r88 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.145 $Y2=2.72
r89 35 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.53 $Y2=2.72
r90 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=2.72
+ $X2=2.985 $Y2=2.72
r91 34 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.82 $Y=2.72
+ $X2=2.53 $Y2=2.72
r92 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r93 33 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r95 30 48 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.722 $Y2=2.72
r96 30 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.61 $Y2=2.72
r97 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=2.145 $Y2=2.72
r98 29 32 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=2.72 $X2=1.61
+ $Y2=2.72
r99 24 48 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.722 $Y2=2.72
r100 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r101 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r102 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r103 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=2.635
+ $X2=2.985 $Y2=2.72
r104 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.985 $Y=2.635
+ $X2=2.985 $Y2=2.36
r105 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.635
+ $X2=2.145 $Y2=2.72
r106 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.145 $Y=2.635
+ $X2=2.145 $Y2=2.36
r107 10 48 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.722 $Y=2.635
+ $X2=0.722 $Y2=2.72
r108 10 12 17.0784 $w=4.13e-07 $l=6.15e-07 $layer=LI1_cond $X=0.722 $Y=2.635
+ $X2=0.722 $Y2=2.02
r109 3 20 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.545 $X2=2.985 $Y2=2.36
r110 2 16 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.545 $X2=2.145 $Y2=2.36
r111 1 12 300 $w=1.7e-07 $l=6.1632e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.72 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%A_320_309# 1 2 3 4 5 18 22 25 26 30 36
r51 35 36 15.8179 $w=5.68e-07 $l=5.15e-07 $layer=LI1_cond $X=3.835 $Y=2.18
+ $X2=3.32 $Y2=2.18
r52 28 30 17.6264 $w=5.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.73 $Y=2.18
+ $X2=5.57 $Y2=2.18
r53 26 35 1.15411 $w=5.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.89 $Y=2.18
+ $X2=3.835 $Y2=2.18
r54 26 28 17.6264 $w=5.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.89 $Y=2.18
+ $X2=4.73 $Y2=2.18
r55 25 33 5.00066 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=2 $X2=2.565
+ $Y2=2
r56 25 36 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=2.65 $Y=2 $X2=3.32
+ $Y2=2
r57 20 33 1.60063 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.565 $Y=2.105
+ $X2=2.565 $Y2=2
r58 20 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.565 $Y=2.105
+ $X2=2.565 $Y2=2.3
r59 16 33 54.3736 $w=1.97e-07 $l=8.78e-07 $layer=LI1_cond $X=1.687 $Y=2
+ $X2=2.565 $Y2=2
r60 16 18 9.17251 $w=2.43e-07 $l=1.95e-07 $layer=LI1_cond $X=1.687 $Y=2.105
+ $X2=1.687 $Y2=2.3
r61 5 30 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.435
+ $Y=1.485 $X2=5.57 $Y2=2.02
r62 4 28 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=4.595
+ $Y=1.485 $X2=4.73 $Y2=2.02
r63 3 35 150 $w=1.7e-07 $l=7.66551e-07 $layer=licon1_PDIFF $count=4 $X=3.27
+ $Y=1.545 $X2=3.835 $Y2=2.02
r64 2 22 600 $w=1.7e-07 $l=8.19726e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.545 $X2=2.565 $Y2=2.3
r65 1 18 600 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.545 $X2=1.725 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%Z 1 2 3 4 13 19 20 21 22 23 24 25 26 27 28
+ 41 61
c66 13 0 8.82398e-20 $X=5.675 $Y=0.735
r67 28 41 3.05577 $w=2.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.785 $Y=1.585
+ $X2=5.675 $Y2=1.585
r68 27 28 9.70706 $w=3.88e-07 $l=2.55e-07 $layer=LI1_cond $X=5.785 $Y=1.19
+ $X2=5.785 $Y2=1.445
r69 26 61 3.56518 $w=2.2e-07 $l=1.2e-07 $layer=LI1_cond $X=5.785 $Y=0.735
+ $X2=5.785 $Y2=0.855
r70 26 27 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=5.785 $Y=0.895
+ $X2=5.785 $Y2=1.19
r71 26 61 2.09535 $w=2.18e-07 $l=4e-08 $layer=LI1_cond $X=5.785 $Y=0.895
+ $X2=5.785 $Y2=0.855
r72 25 41 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.315 $Y=1.585
+ $X2=5.675 $Y2=1.585
r73 25 58 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=1.585
+ $X2=5.15 $Y2=1.585
r74 24 58 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=1.585
+ $X2=5.15 $Y2=1.585
r75 24 54 22.4315 $w=2.78e-07 $l=5.45e-07 $layer=LI1_cond $X=4.855 $Y=1.585
+ $X2=4.31 $Y2=1.585
r76 23 54 15.4345 $w=2.78e-07 $l=3.75e-07 $layer=LI1_cond $X=3.935 $Y=1.585
+ $X2=4.31 $Y2=1.585
r77 22 23 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=3.475 $Y=1.585
+ $X2=3.935 $Y2=1.585
r78 21 22 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=3.015 $Y=1.585
+ $X2=3.475 $Y2=1.585
r79 20 21 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=2.555 $Y=1.585
+ $X2=3.015 $Y2=1.585
r80 19 20 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=2.095 $Y=1.585
+ $X2=2.555 $Y2=1.585
r81 15 18 40.3355 $w=2.38e-07 $l=8.4e-07 $layer=LI1_cond $X=4.31 $Y=0.735
+ $X2=5.15 $Y2=0.735
r82 13 26 3.26808 $w=2.4e-07 $l=1.1e-07 $layer=LI1_cond $X=5.675 $Y=0.735
+ $X2=5.785 $Y2=0.735
r83 13 18 25.2097 $w=2.38e-07 $l=5.25e-07 $layer=LI1_cond $X=5.675 $Y=0.735
+ $X2=5.15 $Y2=0.735
r84 4 58 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.485 $X2=5.15 $Y2=1.64
r85 3 54 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=1.485 $X2=4.31 $Y2=1.64
r86 2 18 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.15 $Y2=0.76
r87 1 15 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.235 $X2=4.31 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48 51
+ 54
r79 54 55 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r80 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r81 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r82 45 55 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=3.45
+ $Y2=0
r83 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r84 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.35
+ $Y2=0
r85 42 44 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=5.75 $Y2=0
r86 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r87 41 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r88 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r89 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.51
+ $Y2=0
r90 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.99
+ $Y2=0
r91 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.35
+ $Y2=0
r92 37 40 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=2.99
+ $Y2=0
r93 36 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r94 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r95 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r96 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r97 32 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r98 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r99 30 48 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.722
+ $Y2=0
r100 30 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.15
+ $Y2=0
r101 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.51
+ $Y2=0
r102 29 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.07 $Y2=0
r103 24 48 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.722 $Y2=0
r104 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r105 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r106 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r107 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r108 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.36
r109 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0
r110 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0.36
r111 10 48 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.722 $Y=0.085
+ $X2=0.722 $Y2=0
r112 10 12 7.63667 $w=4.13e-07 $l=2.75e-07 $layer=LI1_cond $X=0.722 $Y=0.085
+ $X2=0.722 $Y2=0.36
r113 3 20 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.235 $X2=3.35 $Y2=0.36
r114 2 16 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.235 $X2=2.51 $Y2=0.36
r115 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_4%A_393_47# 1 2 3 4 5 16 19 20 21 24 30 34 36
r59 32 34 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=4.73 $Y=0.35
+ $X2=5.57 $Y2=0.35
r60 30 32 44.0718 $w=1.88e-07 $l=7.55e-07 $layer=LI1_cond $X=3.975 $Y=0.35
+ $X2=4.73 $Y2=0.35
r61 27 29 3.77524 $w=2.88e-07 $l=9.5e-08 $layer=LI1_cond $X=3.83 $Y=0.655
+ $X2=3.83 $Y2=0.56
r62 26 30 7.20849 $w=1.9e-07 $l=1.86548e-07 $layer=LI1_cond $X=3.83 $Y=0.445
+ $X2=3.975 $Y2=0.35
r63 26 29 4.57003 $w=2.88e-07 $l=1.15e-07 $layer=LI1_cond $X=3.83 $Y=0.445
+ $X2=3.83 $Y2=0.56
r64 25 36 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.755 $X2=2.93
+ $Y2=0.755
r65 24 27 7.11991 $w=2e-07 $l=1.88481e-07 $layer=LI1_cond $X=3.685 $Y=0.755
+ $X2=3.83 $Y2=0.655
r66 24 25 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=3.685 $Y=0.755
+ $X2=3.015 $Y2=0.755
r67 21 36 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.93 $Y=0.655 $X2=2.93
+ $Y2=0.755
r68 21 23 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.93 $Y=0.655
+ $X2=2.93 $Y2=0.56
r69 19 36 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.755 $X2=2.93
+ $Y2=0.755
r70 19 20 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=2.845 $Y=0.755
+ $X2=2.175 $Y2=0.755
r71 16 20 7.06569 $w=2e-07 $l=1.83303e-07 $layer=LI1_cond $X=2.035 $Y=0.655
+ $X2=2.175 $Y2=0.755
r72 16 18 4.13929 $w=2.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.035 $Y=0.655
+ $X2=2.035 $Y2=0.56
r73 5 34 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.235 $X2=5.57 $Y2=0.36
r74 4 32 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.595
+ $Y=0.235 $X2=4.73 $Y2=0.36
r75 3 29 182 $w=1.7e-07 $l=4.11096e-07 $layer=licon1_NDIFF $count=1 $X=3.635
+ $Y=0.235 $X2=3.83 $Y2=0.56
r76 2 23 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.93 $Y2=0.56
r77 1 18 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.235 $X2=2.09 $Y2=0.56
.ends


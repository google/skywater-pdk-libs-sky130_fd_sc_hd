* File: sky130_fd_sc_hd__or3_2.spice
* Created: Tue Sep  1 19:27:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or3_2.pex.spice"
.subckt sky130_fd_sc_hd__or3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_30_53#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_30_53#_M1009_d N_B_M1009_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_30_53#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1008_d N_A_30_53#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.123773 AS=0.08775 PD=1.2028 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_30_53#_M1006_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.08775 PD=1.87 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 A_112_297# N_C_M1005_g N_A_30_53#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_184_297# N_B_M1002_g A_112_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=51.5943 NRS=23.443 M=1 R=2.8 SA=75000.5
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_184_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.0693 PD=0.792676 PS=0.75 NRD=72.1217 NRS=51.5943 M=1 R=2.8
+ SA=75001 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1007_d N_A_30_53#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.208803 AS=0.135 PD=1.88732 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_30_53#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.315 AS=0.135 PD=2.63 PS=1.27 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_58 VPB 0 2.32308e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__or3_2.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.810000 1.495000 9.575000 1.615000 ;
        RECT 8.810000 1.615000 9.140000 2.460000 ;
        RECT 8.890000 0.265000 9.135000 0.765000 ;
        RECT 8.890000 0.765000 9.575000 0.825000 ;
        RECT 8.975000 0.825000 9.575000 0.855000 ;
        RECT 8.975000 1.445000 9.575000 1.495000 ;
        RECT 8.990000 0.855000 9.575000 0.895000 ;
        RECT 9.020000 0.895000 9.575000 1.445000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.340000 1.005000 ;
        RECT 6.660000 1.005000 7.010000 1.065000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.455000  0.085000 1.785000 0.465000 ;
        RECT 3.610000  0.085000 4.020000 0.525000 ;
        RECT 4.760000  0.085000 5.080000 0.545000 ;
        RECT 6.690000  0.085000 7.330000 0.565000 ;
        RECT 8.390000  0.085000 8.720000 0.825000 ;
        RECT 9.305000  0.085000 9.575000 0.595000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.455000 2.135000 1.785000 2.635000 ;
        RECT 3.430000 2.255000 3.810000 2.635000 ;
        RECT 4.330000 2.255000 4.660000 2.635000 ;
        RECT 5.920000 2.255000 6.340000 2.635000 ;
        RECT 7.010000 1.945000 7.340000 2.635000 ;
        RECT 8.470000 1.495000 8.640000 2.635000 ;
        RECT 9.310000 1.785000 9.575000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.345000 0.345000 0.635000 ;
      RECT 0.085000 0.635000 0.835000 0.805000 ;
      RECT 0.085000 1.795000 0.835000 1.965000 ;
      RECT 0.085000 1.965000 0.345000 2.465000 ;
      RECT 0.605000 0.805000 0.835000 1.795000 ;
      RECT 1.005000 0.565000 1.235000 2.045000 ;
      RECT 1.015000 0.345000 1.235000 0.565000 ;
      RECT 1.015000 2.045000 1.235000 2.465000 ;
      RECT 1.430000 0.635000 2.125000 0.825000 ;
      RECT 1.430000 0.825000 1.600000 1.795000 ;
      RECT 1.430000 1.795000 2.125000 1.965000 ;
      RECT 1.955000 0.305000 2.125000 0.635000 ;
      RECT 1.955000 1.965000 2.125000 2.465000 ;
      RECT 2.350000 0.705000 2.570000 1.575000 ;
      RECT 2.350000 1.575000 2.850000 1.955000 ;
      RECT 2.360000 2.250000 3.190000 2.420000 ;
      RECT 2.425000 0.265000 3.440000 0.465000 ;
      RECT 2.750000 0.645000 3.100000 1.015000 ;
      RECT 3.020000 1.195000 3.440000 1.235000 ;
      RECT 3.020000 1.235000 4.370000 1.405000 ;
      RECT 3.020000 1.405000 3.190000 2.250000 ;
      RECT 3.270000 0.465000 3.440000 1.195000 ;
      RECT 3.360000 1.575000 3.610000 1.835000 ;
      RECT 3.360000 1.835000 4.710000 2.085000 ;
      RECT 3.990000 2.085000 4.160000 2.375000 ;
      RECT 4.120000 1.405000 4.370000 1.565000 ;
      RECT 4.310000 0.295000 4.560000 0.725000 ;
      RECT 4.310000 0.725000 4.710000 1.065000 ;
      RECT 4.540000 1.065000 4.710000 1.835000 ;
      RECT 4.880000 0.725000 6.150000 0.895000 ;
      RECT 4.880000 0.895000 5.050000 1.655000 ;
      RECT 4.880000 1.655000 5.400000 1.965000 ;
      RECT 5.110000 2.165000 5.740000 2.415000 ;
      RECT 5.220000 1.065000 5.400000 1.475000 ;
      RECT 5.570000 1.235000 7.490000 1.405000 ;
      RECT 5.570000 1.405000 5.740000 1.915000 ;
      RECT 5.570000 1.915000 6.780000 2.085000 ;
      RECT 5.570000 2.085000 5.740000 2.165000 ;
      RECT 5.640000 0.305000 6.490000 0.475000 ;
      RECT 5.800000 0.895000 6.150000 1.015000 ;
      RECT 5.910000 1.575000 7.880000 1.745000 ;
      RECT 6.320000 0.475000 6.490000 1.235000 ;
      RECT 6.540000 2.085000 6.780000 2.375000 ;
      RECT 7.140000 1.175000 7.490000 1.235000 ;
      RECT 7.510000 1.745000 7.880000 1.765000 ;
      RECT 7.510000 1.765000 7.680000 2.375000 ;
      RECT 7.530000 0.350000 7.880000 0.680000 ;
      RECT 7.690000 0.680000 7.880000 1.575000 ;
      RECT 7.970000 1.915000 8.300000 2.425000 ;
      RECT 8.050000 0.345000 8.220000 0.995000 ;
      RECT 8.050000 0.995000 8.850000 1.325000 ;
      RECT 8.050000 1.325000 8.300000 1.915000 ;
    LAYER mcon ;
      RECT 0.605000 1.785000 0.775000 1.955000 ;
      RECT 1.065000 0.765000 1.235000 0.935000 ;
      RECT 2.445000 1.785000 2.615000 1.955000 ;
      RECT 2.905000 0.765000 3.075000 0.935000 ;
      RECT 5.205000 1.785000 5.375000 1.955000 ;
      RECT 5.225000 1.105000 5.395000 1.275000 ;
    LAYER met1 ;
      RECT 0.545000 1.755000 0.835000 1.800000 ;
      RECT 0.545000 1.800000 5.435000 1.940000 ;
      RECT 0.545000 1.940000 0.835000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.455000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.165000 1.075000 5.455000 1.120000 ;
      RECT 5.165000 1.260000 5.455000 1.305000 ;
  END
END sky130_fd_sc_hd__dfstp_2
END LIBRARY

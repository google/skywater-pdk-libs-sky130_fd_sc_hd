# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__mux2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.995000 1.750000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.435000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.740000 1.325000 ;
        RECT 0.570000 0.635000 2.850000 0.805000 ;
        RECT 0.570000 0.805000 0.740000 0.995000 ;
        RECT 2.680000 0.805000 2.850000 0.995000 ;
        RECT 2.680000 0.995000 3.395000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.915000 0.255000 4.085000 0.635000 ;
        RECT 3.915000 0.635000 5.430000 0.805000 ;
        RECT 3.915000 1.575000 5.430000 1.745000 ;
        RECT 3.915000 1.745000 4.085000 2.465000 ;
        RECT 4.755000 0.255000 4.925000 0.635000 ;
        RECT 4.755000 1.745000 4.925000 2.465000 ;
        RECT 5.200000 0.805000 5.430000 1.575000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.295000 0.345000 0.625000 ;
      RECT 0.090000  0.625000 0.260000 1.495000 ;
      RECT 0.090000  1.495000 1.080000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  1.835000 0.820000 2.635000 ;
      RECT 0.910000  0.995000 1.080000 1.495000 ;
      RECT 0.990000  1.935000 1.340000 2.275000 ;
      RECT 0.990000  2.275000 2.770000 2.445000 ;
      RECT 1.530000  1.935000 3.245000 2.105000 ;
      RECT 1.975000  0.295000 3.230000 0.465000 ;
      RECT 1.980000  1.595000 3.735000 1.765000 ;
      RECT 3.060000  0.465000 3.230000 0.655000 ;
      RECT 3.060000  0.655000 3.735000 0.825000 ;
      RECT 3.075000  2.105000 3.245000 2.465000 ;
      RECT 3.415000  0.085000 3.745000 0.465000 ;
      RECT 3.415000  2.255000 3.745000 2.635000 ;
      RECT 3.565000  0.825000 3.735000 1.075000 ;
      RECT 3.565000  1.075000 5.030000 1.245000 ;
      RECT 3.565000  1.245000 3.735000 1.595000 ;
      RECT 3.565000  1.765000 3.735000 1.785000 ;
      RECT 4.255000  0.085000 4.585000 0.465000 ;
      RECT 4.255000  1.915000 4.585000 2.635000 ;
      RECT 5.095000  0.085000 5.425000 0.465000 ;
      RECT 5.095000  1.915000 5.425000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_4

* File: sky130_fd_sc_hd__nor4bb_1.spice.SKY130_FD_SC_HD__NOR4BB_1.pxi
* Created: Thu Aug 27 14:33:24 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4BB_1%C_N N_C_N_M1010_g N_C_N_M1002_g C_N C_N
+ N_C_N_c_77_n N_C_N_c_78_n N_C_N_c_79_n PM_SKY130_FD_SC_HD__NOR4BB_1%C_N
x_PM_SKY130_FD_SC_HD__NOR4BB_1%D_N N_D_N_M1008_g N_D_N_M1011_g D_N N_D_N_c_111_n
+ N_D_N_c_112_n PM_SKY130_FD_SC_HD__NOR4BB_1%D_N
x_PM_SKY130_FD_SC_HD__NOR4BB_1%A_205_93# N_A_205_93#_M1008_d N_A_205_93#_M1011_d
+ N_A_205_93#_c_143_n N_A_205_93#_M1003_g N_A_205_93#_M1007_g
+ N_A_205_93#_c_144_n N_A_205_93#_c_145_n N_A_205_93#_c_152_n
+ N_A_205_93#_c_153_n N_A_205_93#_c_146_n N_A_205_93#_c_147_n
+ N_A_205_93#_c_148_n PM_SKY130_FD_SC_HD__NOR4BB_1%A_205_93#
x_PM_SKY130_FD_SC_HD__NOR4BB_1%A_27_410# N_A_27_410#_M1002_s N_A_27_410#_M1010_s
+ N_A_27_410#_c_208_n N_A_27_410#_M1005_g N_A_27_410#_M1004_g
+ N_A_27_410#_c_209_n N_A_27_410#_c_214_n N_A_27_410#_c_215_n
+ N_A_27_410#_c_216_n N_A_27_410#_c_217_n N_A_27_410#_c_218_n
+ N_A_27_410#_c_219_n N_A_27_410#_c_210_n N_A_27_410#_c_211_n
+ N_A_27_410#_c_221_n PM_SKY130_FD_SC_HD__NOR4BB_1%A_27_410#
x_PM_SKY130_FD_SC_HD__NOR4BB_1%B N_B_c_289_n N_B_M1006_g N_B_M1001_g B
+ N_B_c_290_n N_B_c_291_n PM_SKY130_FD_SC_HD__NOR4BB_1%B
x_PM_SKY130_FD_SC_HD__NOR4BB_1%A N_A_M1009_g N_A_M1000_g A N_A_c_330_n
+ N_A_c_331_n N_A_c_332_n PM_SKY130_FD_SC_HD__NOR4BB_1%A
x_PM_SKY130_FD_SC_HD__NOR4BB_1%VPWR N_VPWR_M1010_d N_VPWR_M1000_d N_VPWR_c_358_n
+ N_VPWR_c_359_n N_VPWR_c_360_n VPWR N_VPWR_c_361_n N_VPWR_c_362_n
+ N_VPWR_c_363_n N_VPWR_c_357_n PM_SKY130_FD_SC_HD__NOR4BB_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR4BB_1%Y N_Y_M1003_d N_Y_M1006_d N_Y_M1007_s N_Y_c_404_n
+ N_Y_c_403_n N_Y_c_445_p N_Y_c_432_n N_Y_c_420_n Y
+ PM_SKY130_FD_SC_HD__NOR4BB_1%Y
x_PM_SKY130_FD_SC_HD__NOR4BB_1%VGND N_VGND_M1002_d N_VGND_M1003_s N_VGND_M1005_d
+ N_VGND_M1009_d N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n
+ N_VGND_c_467_n VGND N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n
+ N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n VGND
+ PM_SKY130_FD_SC_HD__NOR4BB_1%VGND
cc_1 VNB N_C_N_c_77_n 0.023255f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_2 VNB N_C_N_c_78_n 0.00587728f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_3 VNB N_C_N_c_79_n 0.020759f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_4 VNB D_N 0.00229145f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_5 VNB N_D_N_c_111_n 0.0258825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_D_N_c_112_n 0.0189315f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_7 VNB N_A_205_93#_c_143_n 0.0180526f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.675
cc_8 VNB N_A_205_93#_c_144_n 0.0256525f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_9 VNB N_A_205_93#_c_145_n 0.0080853f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_10 VNB N_A_205_93#_c_146_n 0.0113249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_205_93#_c_147_n 0.00330492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_205_93#_c_148_n 0.00273059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_c_208_n 0.0169951f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.675
cc_14 VNB N_A_27_410#_c_209_n 0.0224435f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_15 VNB N_A_27_410#_c_210_n 0.0220289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_410#_c_211_n 0.0187759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B_c_289_n 0.0170187f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_18 VNB N_B_c_290_n 0.0185667f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_19 VNB N_B_c_291_n 0.00563386f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_20 VNB A 0.0158416f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_21 VNB N_A_c_330_n 0.0276092f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_22 VNB N_A_c_331_n 0.0213312f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_23 VNB N_A_c_332_n 0.00142889f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.19
cc_24 VNB N_VPWR_c_357_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_403_n 0.00291513f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_26 VNB N_VGND_c_463_n 0.0151102f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_27 VNB N_VGND_c_464_n 0.00881627f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.53
cc_28 VNB N_VGND_c_465_n 0.00423911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_466_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_467_n 0.0258009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_468_n 0.0196515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_469_n 0.0129543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_470_n 0.0136663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_471_n 0.0242066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_472_n 0.00507259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_473_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_474_n 0.219556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_C_N_M1010_g 0.056069f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.26
cc_39 VPB N_C_N_c_77_n 0.00471554f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_40 VPB N_C_N_c_78_n 0.00237324f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_41 VPB N_D_N_M1011_g 0.0219639f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_42 VPB D_N 5.1145e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_43 VPB N_D_N_c_111_n 0.00579592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_205_93#_M1007_g 0.0215438f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_45 VPB N_A_205_93#_c_144_n 0.0115474f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_46 VPB N_A_205_93#_c_145_n 5.21632e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_47 VPB N_A_205_93#_c_152_n 0.00988601f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.325
cc_48 VPB N_A_205_93#_c_153_n 0.00341854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_205_93#_c_147_n 0.00167012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_410#_M1004_g 0.0179385f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_51 VPB N_A_27_410#_c_209_n 0.0273492f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_52 VPB N_A_27_410#_c_214_n 0.0149581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_410#_c_215_n 0.0064407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_410#_c_216_n 0.00590134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_410#_c_217_n 0.00953976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_410#_c_218_n 0.00358648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_410#_c_219_n 0.00212219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_410#_c_210_n 0.00695225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_410#_c_221_n 0.0117133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_B_M1001_g 0.0179103f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_61 VPB B 0.00283213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_B_c_290_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_63 VPB N_B_c_291_n 0.00203325f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_64 VPB N_A_M1000_g 0.0212562f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_65 VPB N_A_c_330_n 0.00693428f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_66 VPB N_A_c_332_n 0.0169994f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.19
cc_67 VPB N_VPWR_c_358_n 0.00656694f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_68 VPB N_VPWR_c_359_n 0.0103102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_360_n 0.0266763f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_70 VPB N_VPWR_c_361_n 0.0144618f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_71 VPB N_VPWR_c_362_n 0.0595127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_363_n 0.00518909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_357_n 0.0519452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_Y_c_404_n 0.00357658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_Y_c_403_n 0.00108648f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_76 N_C_N_M1010_g N_D_N_M1011_g 0.0242889f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_77 N_C_N_c_78_n N_D_N_M1011_g 0.00412866f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C_N_c_77_n D_N 2.85663e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C_N_c_78_n D_N 0.0259635f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_80 N_C_N_c_77_n N_D_N_c_111_n 0.019221f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_81 N_C_N_c_78_n N_D_N_c_111_n 0.00225922f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C_N_c_79_n N_D_N_c_112_n 0.0106782f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_83 N_C_N_M1010_g N_A_205_93#_c_152_n 2.23982e-19 $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_84 N_C_N_c_78_n N_A_205_93#_c_152_n 0.0115417f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_85 N_C_N_c_78_n N_A_205_93#_c_147_n 0.0063226f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_86 N_C_N_M1010_g N_A_27_410#_c_209_n 0.0141141f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_87 N_C_N_c_77_n N_A_27_410#_c_209_n 0.00753785f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_88 N_C_N_c_78_n N_A_27_410#_c_209_n 0.0529229f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_89 N_C_N_c_79_n N_A_27_410#_c_209_n 0.00528758f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C_N_M1010_g N_A_27_410#_c_215_n 0.0155459f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_91 N_C_N_c_77_n N_A_27_410#_c_215_n 7.20588e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_92 N_C_N_c_78_n N_A_27_410#_c_215_n 0.0259102f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_93 N_C_N_M1010_g N_A_27_410#_c_216_n 0.00281901f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_94 N_C_N_c_79_n N_A_27_410#_c_211_n 3.38304e-19 $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_95 N_C_N_c_78_n N_VPWR_M1010_d 0.00454723f $X=0.515 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_96 N_C_N_M1010_g N_VPWR_c_358_n 0.00962285f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_97 N_C_N_M1010_g N_VPWR_c_361_n 0.00331133f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_98 N_C_N_M1010_g N_VPWR_c_357_n 0.00482357f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_99 N_C_N_c_78_n N_VGND_c_463_n 0.0113325f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C_N_c_79_n N_VGND_c_463_n 0.00422655f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_101 N_C_N_c_79_n N_VGND_c_471_n 0.00510437f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_102 N_C_N_c_79_n N_VGND_c_474_n 0.00512902f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_103 D_N N_A_205_93#_c_144_n 9.69012e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_104 N_D_N_c_111_n N_A_205_93#_c_144_n 0.0160964f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_105 N_D_N_M1011_g N_A_205_93#_c_152_n 0.00334116f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_106 D_N N_A_205_93#_c_152_n 0.0142775f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_107 N_D_N_c_111_n N_A_205_93#_c_152_n 0.0036075f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_108 N_D_N_M1011_g N_A_205_93#_c_153_n 0.0030911f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_109 D_N N_A_205_93#_c_146_n 0.0128769f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_110 N_D_N_c_111_n N_A_205_93#_c_146_n 0.00284091f $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_D_N_c_112_n N_A_205_93#_c_146_n 3.44947e-19 $X=1.035 $Y=0.995 $X2=0
+ $Y2=0
cc_112 D_N N_A_205_93#_c_147_n 0.0267936f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_113 N_D_N_c_111_n N_A_205_93#_c_147_n 9.94404e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_D_N_c_112_n N_A_205_93#_c_148_n 0.00422007f $X=1.035 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_D_N_M1011_g N_A_27_410#_c_215_n 0.0137665f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_116 D_N N_A_27_410#_c_215_n 0.00121337f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_117 N_D_N_M1011_g N_VPWR_c_362_n 5.42132e-19 $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_118 N_D_N_M1011_g N_Y_c_404_n 4.13604e-19 $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_119 N_D_N_c_112_n N_VGND_c_463_n 0.00289858f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_120 N_D_N_c_112_n N_VGND_c_464_n 0.00311391f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_121 N_D_N_c_112_n N_VGND_c_468_n 0.00510437f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_122 N_D_N_c_112_n N_VGND_c_474_n 0.00512902f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_205_93#_c_143_n N_A_27_410#_c_208_n 0.0231911f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_205_93#_M1007_g N_A_27_410#_M1004_g 0.0608997f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_205_93#_M1011_d N_A_27_410#_c_215_n 0.00155839f $X=1.03 $Y=1.485
+ $X2=0 $Y2=0
cc_126 N_A_205_93#_c_152_n N_A_27_410#_c_215_n 0.0119231f $X=1.41 $Y=1.62 $X2=0
+ $Y2=0
cc_127 N_A_205_93#_M1007_g N_A_27_410#_c_216_n 0.00251023f $X=1.89 $Y=1.985
+ $X2=0 $Y2=0
cc_128 N_A_205_93#_M1007_g N_A_27_410#_c_217_n 0.011647f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_205_93#_c_152_n N_A_27_410#_c_217_n 0.00861067f $X=1.41 $Y=1.62 $X2=0
+ $Y2=0
cc_130 N_A_205_93#_M1007_g N_A_27_410#_c_219_n 8.35144e-19 $X=1.89 $Y=1.985
+ $X2=0 $Y2=0
cc_131 N_A_205_93#_c_145_n N_A_27_410#_c_219_n 3.18783e-19 $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_205_93#_c_145_n N_A_27_410#_c_210_n 0.0202445f $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_205_93#_M1007_g N_VPWR_c_362_n 0.00357877f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_205_93#_M1007_g N_VPWR_c_357_n 0.00666937f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_205_93#_c_152_n N_Y_M1007_s 0.00256692f $X=1.41 $Y=1.62 $X2=0 $Y2=0
cc_136 N_A_205_93#_c_153_n N_Y_M1007_s 4.24137e-19 $X=1.5 $Y=1.525 $X2=0 $Y2=0
cc_137 N_A_205_93#_M1007_g N_Y_c_404_n 0.00706004f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_205_93#_c_144_n N_Y_c_404_n 0.00327613f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_205_93#_c_152_n N_Y_c_404_n 0.00782608f $X=1.41 $Y=1.62 $X2=0 $Y2=0
cc_140 N_A_205_93#_c_147_n N_Y_c_404_n 0.00247032f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_205_93#_c_143_n N_Y_c_403_n 0.00446329f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_205_93#_M1007_g N_Y_c_403_n 0.0208794f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_205_93#_c_145_n N_Y_c_403_n 0.00911914f $X=1.89 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_205_93#_c_152_n N_Y_c_403_n 0.0106646f $X=1.41 $Y=1.62 $X2=0 $Y2=0
cc_145 N_A_205_93#_c_153_n N_Y_c_403_n 0.0103106f $X=1.5 $Y=1.525 $X2=0 $Y2=0
cc_146 N_A_205_93#_c_147_n N_Y_c_403_n 0.0235082f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_205_93#_c_148_n N_Y_c_403_n 0.00871448f $X=1.547 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_205_93#_c_143_n N_Y_c_420_n 0.00757831f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_205_93#_c_146_n N_Y_c_420_n 0.0101936f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_150 N_A_205_93#_c_146_n N_VGND_M1003_s 0.00245866f $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_151 N_A_205_93#_c_148_n N_VGND_M1003_s 6.03459e-19 $X=1.547 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_205_93#_c_146_n N_VGND_c_463_n 8.07382e-19 $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_153 N_A_205_93#_c_143_n N_VGND_c_464_n 0.00933051f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A_205_93#_c_144_n N_VGND_c_464_n 0.00389571f $X=1.815 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_205_93#_c_146_n N_VGND_c_464_n 0.00795191f $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_156 N_A_205_93#_c_147_n N_VGND_c_464_n 0.00323367f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_205_93#_c_146_n N_VGND_c_468_n 0.0100902f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_158 N_A_205_93#_c_143_n N_VGND_c_469_n 0.00351131f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_205_93#_c_143_n N_VGND_c_474_n 0.00439928f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_205_93#_c_146_n N_VGND_c_474_n 0.013836f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_161 N_A_27_410#_c_208_n N_B_c_289_n 0.0208152f $X=2.31 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_27_410#_M1004_g N_B_M1001_g 0.0454356f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_27_410#_c_219_n N_B_M1001_g 5.37697e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_27_410#_M1004_g B 8.46082e-19 $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_27_410#_c_219_n N_B_c_290_n 3.60807e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_27_410#_c_210_n N_B_c_290_n 0.0203108f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_27_410#_M1004_g N_B_c_291_n 0.0011933f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_27_410#_c_219_n N_B_c_291_n 0.0362271f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_27_410#_c_210_n N_B_c_291_n 0.00203858f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_27_410#_c_215_n N_VPWR_M1010_d 0.00552714f $X=1.035 $Y=1.977
+ $X2=-0.19 $Y2=-0.24
cc_171 N_A_27_410#_c_215_n N_VPWR_c_358_n 0.0208172f $X=1.035 $Y=1.977 $X2=0
+ $Y2=0
cc_172 N_A_27_410#_c_216_n N_VPWR_c_358_n 0.00399771f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_173 N_A_27_410#_c_218_n N_VPWR_c_358_n 0.0139001f $X=1.205 $Y=2.38 $X2=0
+ $Y2=0
cc_174 N_A_27_410#_c_214_n N_VPWR_c_361_n 0.0168539f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_175 N_A_27_410#_c_215_n N_VPWR_c_361_n 0.00236787f $X=1.035 $Y=1.977 $X2=0
+ $Y2=0
cc_176 N_A_27_410#_M1004_g N_VPWR_c_362_n 0.00357668f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_410#_c_215_n N_VPWR_c_362_n 0.00336708f $X=1.035 $Y=1.977 $X2=0
+ $Y2=0
cc_178 N_A_27_410#_c_217_n N_VPWR_c_362_n 0.0711203f $X=2.225 $Y=2.38 $X2=0
+ $Y2=0
cc_179 N_A_27_410#_c_218_n N_VPWR_c_362_n 0.0120427f $X=1.205 $Y=2.38 $X2=0
+ $Y2=0
cc_180 N_A_27_410#_M1004_g N_VPWR_c_357_n 0.00546639f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_27_410#_c_214_n N_VPWR_c_357_n 0.00987378f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_182 N_A_27_410#_c_215_n N_VPWR_c_357_n 0.0109951f $X=1.035 $Y=1.977 $X2=0
+ $Y2=0
cc_183 N_A_27_410#_c_217_n N_VPWR_c_357_n 0.0431508f $X=2.225 $Y=2.38 $X2=0
+ $Y2=0
cc_184 N_A_27_410#_c_218_n N_VPWR_c_357_n 0.00651993f $X=1.205 $Y=2.38 $X2=0
+ $Y2=0
cc_185 N_A_27_410#_c_217_n N_Y_M1007_s 0.00480304f $X=2.225 $Y=2.38 $X2=0 $Y2=0
cc_186 N_A_27_410#_M1004_g N_Y_c_404_n 6.40012e-19 $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_27_410#_c_215_n N_Y_c_404_n 0.00773156f $X=1.035 $Y=1.977 $X2=0 $Y2=0
cc_188 N_A_27_410#_c_216_n N_Y_c_404_n 0.00327505f $X=1.12 $Y=2.295 $X2=0 $Y2=0
cc_189 N_A_27_410#_c_217_n N_Y_c_404_n 0.032695f $X=2.225 $Y=2.38 $X2=0 $Y2=0
cc_190 N_A_27_410#_c_208_n N_Y_c_403_n 0.00356321f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_27_410#_M1004_g N_Y_c_403_n 0.00197712f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_27_410#_c_215_n N_Y_c_403_n 0.00202317f $X=1.035 $Y=1.977 $X2=0 $Y2=0
cc_193 N_A_27_410#_c_219_n N_Y_c_403_n 0.0535214f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_27_410#_c_210_n N_Y_c_403_n 0.00190451f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_27_410#_c_208_n N_Y_c_432_n 0.0116657f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_27_410#_c_219_n N_Y_c_432_n 0.0121845f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_27_410#_c_210_n N_Y_c_432_n 0.00108358f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_27_410#_c_210_n N_Y_c_420_n 0.00108358f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_410#_c_217_n A_393_297# 0.00649847f $X=2.225 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_200 N_A_27_410#_c_211_n N_VGND_c_463_n 0.0106535f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_201 N_A_27_410#_c_208_n N_VGND_c_464_n 6.85849e-19 $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_27_410#_c_208_n N_VGND_c_465_n 0.0016712f $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_27_410#_c_208_n N_VGND_c_469_n 0.00427293f $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_27_410#_c_211_n N_VGND_c_471_n 0.00972557f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_205 N_A_27_410#_c_208_n N_VGND_c_474_n 0.00582284f $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_27_410#_c_211_n N_VGND_c_474_n 0.0107261f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_207 N_B_M1001_g N_A_M1000_g 0.0559517f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_208 B N_A_M1000_g 0.00414093f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_209 N_B_c_290_n A 9.33416e-19 $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B_c_291_n A 0.0239216f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B_c_290_n N_A_c_330_n 0.021289f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B_c_291_n N_A_c_330_n 0.00221729f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B_c_289_n N_A_c_331_n 0.0241532f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_214 B N_A_c_332_n 0.00286498f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_215 N_B_c_291_n N_A_c_332_n 0.00824651f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B_M1001_g N_VPWR_c_360_n 0.00181357f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B_M1001_g N_VPWR_c_362_n 0.00529104f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_218 B N_VPWR_c_362_n 0.0117355f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_219 N_B_M1001_g N_VPWR_c_357_n 0.00957803f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_220 B N_VPWR_c_357_n 0.00947667f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_221 N_B_c_289_n N_Y_c_432_n 0.0113209f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_222 B N_Y_c_432_n 0.00479918f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_223 N_B_c_290_n N_Y_c_432_n 5.02391e-19 $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B_c_291_n N_Y_c_432_n 0.0215897f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_225 B A_477_297# 0.003296f $X=2.905 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_226 B A_573_297# 0.00328672f $X=2.905 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_227 N_B_c_289_n N_VGND_c_465_n 0.0016712f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B_c_289_n N_VGND_c_467_n 8.53588e-19 $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B_c_289_n N_VGND_c_470_n 0.00427293f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B_c_289_n N_VGND_c_474_n 0.00582284f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_332_n N_VPWR_M1000_d 0.0043956f $X=3.45 $Y=1.49 $X2=0 $Y2=0
cc_232 N_A_M1000_g N_VPWR_c_360_n 0.0137706f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_233 A N_VPWR_c_360_n 9.17937e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_234 N_A_c_330_n N_VPWR_c_360_n 5.61471e-19 $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_c_332_n N_VPWR_c_360_n 0.021134f $X=3.45 $Y=1.49 $X2=0 $Y2=0
cc_236 N_A_M1000_g N_VPWR_c_362_n 0.0046653f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_M1000_g N_VPWR_c_357_n 0.00799591f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_238 A N_VGND_c_467_n 0.0246263f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A_c_330_n N_VGND_c_467_n 0.00413601f $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_c_331_n N_VGND_c_467_n 0.0119667f $X=3.302 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_c_331_n N_VGND_c_470_n 0.0046653f $X=3.302 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_331_n N_VGND_c_474_n 0.00799591f $X=3.302 $Y=0.995 $X2=0 $Y2=0
cc_243 N_VPWR_c_357_n N_Y_M1007_s 0.00210147f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_357_n A_393_297# 0.00216832f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_245 N_VPWR_c_357_n A_477_297# 0.0137589f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_246 N_VPWR_c_357_n A_573_297# 0.00397011f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_247 N_Y_c_404_n A_393_297# 0.00180053f $X=1.855 $Y=2.04 $X2=-0.19 $Y2=-0.24
cc_248 N_Y_c_403_n A_393_297# 0.00395835f $X=1.955 $Y=1.955 $X2=-0.19 $Y2=-0.24
cc_249 N_Y_c_432_n N_VGND_M1005_d 0.00915616f $X=2.885 $Y=0.74 $X2=0 $Y2=0
cc_250 N_Y_c_432_n N_VGND_c_465_n 0.0165818f $X=2.885 $Y=0.74 $X2=0 $Y2=0
cc_251 N_Y_c_445_p N_VGND_c_469_n 0.00930397f $X=2.1 $Y=0.495 $X2=0 $Y2=0
cc_252 N_Y_c_420_n N_VGND_c_469_n 0.00470974f $X=2.215 $Y=0.74 $X2=0 $Y2=0
cc_253 N_Y_c_432_n N_VGND_c_470_n 0.00251419f $X=2.885 $Y=0.74 $X2=0 $Y2=0
cc_254 Y N_VGND_c_470_n 0.00906533f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_255 N_Y_M1003_d N_VGND_c_474_n 0.00247227f $X=1.965 $Y=0.235 $X2=0 $Y2=0
cc_256 N_Y_M1006_d N_VGND_c_474_n 0.00403782f $X=2.865 $Y=0.235 $X2=0 $Y2=0
cc_257 N_Y_c_445_p N_VGND_c_474_n 0.00731608f $X=2.1 $Y=0.495 $X2=0 $Y2=0
cc_258 N_Y_c_432_n N_VGND_c_474_n 0.00538285f $X=2.885 $Y=0.74 $X2=0 $Y2=0
cc_259 N_Y_c_420_n N_VGND_c_474_n 0.00793983f $X=2.215 $Y=0.74 $X2=0 $Y2=0
cc_260 Y N_VGND_c_474_n 0.00735151f $X=2.905 $Y=0.425 $X2=0 $Y2=0

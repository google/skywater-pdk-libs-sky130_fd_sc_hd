* File: sky130_fd_sc_hd__and3_2.pxi.spice
* Created: Thu Aug 27 14:07:41 2020
* 
x_PM_SKY130_FD_SC_HD__AND3_2%A N_A_M1000_g N_A_M1001_g A N_A_c_58_n
+ PM_SKY130_FD_SC_HD__AND3_2%A
x_PM_SKY130_FD_SC_HD__AND3_2%B N_B_c_83_n N_B_M1007_g N_B_M1006_g B N_B_c_88_n
+ PM_SKY130_FD_SC_HD__AND3_2%B
x_PM_SKY130_FD_SC_HD__AND3_2%C N_C_M1008_g N_C_M1005_g C C N_C_c_128_n
+ PM_SKY130_FD_SC_HD__AND3_2%C
x_PM_SKY130_FD_SC_HD__AND3_2%A_29_311# N_A_29_311#_M1001_s N_A_29_311#_M1000_s
+ N_A_29_311#_M1006_d N_A_29_311#_c_174_n N_A_29_311#_M1003_g
+ N_A_29_311#_M1002_g N_A_29_311#_c_175_n N_A_29_311#_M1004_g
+ N_A_29_311#_M1009_g N_A_29_311#_c_182_n N_A_29_311#_c_176_n
+ N_A_29_311#_c_183_n N_A_29_311#_c_184_n N_A_29_311#_c_177_n
+ N_A_29_311#_c_186_n N_A_29_311#_c_210_n N_A_29_311#_c_187_n
+ N_A_29_311#_c_178_n N_A_29_311#_c_213_n N_A_29_311#_c_189_n
+ N_A_29_311#_c_179_n PM_SKY130_FD_SC_HD__AND3_2%A_29_311#
x_PM_SKY130_FD_SC_HD__AND3_2%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_M1009_s
+ N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n
+ N_VPWR_c_300_n VPWR N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n
+ N_VPWR_c_289_n PM_SKY130_FD_SC_HD__AND3_2%VPWR
x_PM_SKY130_FD_SC_HD__AND3_2%X N_X_M1003_s N_X_M1002_d N_X_c_339_n N_X_c_348_n
+ N_X_c_341_n X X X N_X_c_363_n X N_X_c_364_n PM_SKY130_FD_SC_HD__AND3_2%X
x_PM_SKY130_FD_SC_HD__AND3_2%VGND N_VGND_M1008_d N_VGND_M1004_d N_VGND_c_376_n
+ N_VGND_c_377_n N_VGND_c_378_n VGND N_VGND_c_379_n N_VGND_c_380_n
+ N_VGND_c_381_n N_VGND_c_382_n PM_SKY130_FD_SC_HD__AND3_2%VGND
cc_1 VNB N_A_M1001_g 0.0336848f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.475
cc_2 VNB A 0.022558f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A_c_58_n 0.0369784f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_4 VNB N_B_c_83_n 0.00432773f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_5 VNB N_B_M1007_g 0.0357978f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.765
cc_6 VNB N_C_M1008_g 0.0266361f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.765
cc_7 VNB C 3.82421e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_8 VNB C 0.0105161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_c_128_n 0.0208659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_29_311#_c_174_n 0.0176896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_29_311#_c_175_n 0.0202412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_29_311#_c_176_n 0.011913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_29_311#_c_177_n 0.00415939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_29_311#_c_178_n 0.00379462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_29_311#_c_179_n 0.0412129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_289_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_339_n 7.18219e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0226639f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_19 VNB N_VGND_c_376_n 0.00310376f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_20 VNB N_VGND_c_377_n 0.0101986f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_21 VNB N_VGND_c_378_n 0.0245278f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_22 VNB N_VGND_c_379_n 0.0397582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_380_n 0.0153644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_381_n 0.00510766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_382_n 0.172646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_M1000_g 0.0303289f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.765
cc_27 VPB N_A_c_58_n 0.00858848f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_28 VPB N_B_c_83_n 0.0111753f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.325
cc_29 VPB N_B_M1006_g 0.012812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB B 0.00962821f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_31 VPB N_B_c_88_n 0.0424452f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_32 VPB N_C_M1005_g 0.0205767f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.475
cc_33 VPB N_C_c_128_n 0.00466733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_29_311#_M1002_g 0.020779f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_35 VPB N_A_29_311#_M1009_g 0.0231123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_29_311#_c_182_n 0.0141199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_29_311#_c_183_n 0.00305118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_29_311#_c_184_n 0.00925693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_29_311#_c_177_n 0.00114652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_29_311#_c_186_n 0.00324769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_29_311#_c_187_n 0.00654569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_29_311#_c_178_n 0.00121877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_29_311#_c_189_n 0.0016468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_29_311#_c_179_n 0.00855278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_290_n 0.00144702f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_46 VPB N_VPWR_c_291_n 0.0220356f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_47 VPB N_VPWR_c_292_n 0.00443251f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_48 VPB N_VPWR_c_293_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=0.85
cc_49 VPB N_VPWR_c_294_n 0.0376795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_295_n 0.0177674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_296_n 0.0516155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_297_n 0.00410958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_289_n 0.0497826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_X_c_341_n 5.92182e-19 $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_55 VPB X 0.0119579f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_56 N_A_M1000_g N_B_c_83_n 0.00908734f $X=0.48 $Y=1.765 $X2=-0.19 $Y2=-0.24
cc_57 N_A_c_58_n N_B_c_83_n 0.0370039f $X=0.485 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_58 N_A_M1001_g N_B_M1007_g 0.0370039f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_59 A N_B_M1007_g 4.09557e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_B_M1006_g 0.0143746f $X=0.48 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_A_29_311#_c_176_n 0.012673f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_62 A N_A_29_311#_c_176_n 0.023752f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_58_n N_A_29_311#_c_176_n 0.00106793f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_A_29_311#_c_183_n 0.0148709f $X=0.48 $Y=1.765 $X2=0 $Y2=0
cc_65 A N_A_29_311#_c_183_n 0.00820785f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_66 N_A_c_58_n N_A_29_311#_c_183_n 0.00144512f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_67 A N_A_29_311#_c_184_n 0.0210059f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_68 N_A_c_58_n N_A_29_311#_c_184_n 0.00543798f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_A_29_311#_c_177_n 0.0023763f $X=0.48 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_M1001_g N_A_29_311#_c_177_n 0.00973945f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_71 A N_A_29_311#_c_177_n 0.0376093f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_VPWR_c_290_n 0.00874185f $X=0.48 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_VPWR_c_300_n 0.00256209f $X=0.48 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_M1000_g N_VPWR_c_296_n 0.00483317f $X=0.48 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_M1001_g N_VGND_c_379_n 0.00347765f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VGND_c_382_n 0.00564484f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_77 A N_VGND_c_382_n 0.00154089f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_78 N_B_M1007_g N_C_M1008_g 0.0529454f $X=0.845 $Y=0.475 $X2=0 $Y2=0
cc_79 N_B_c_83_n N_C_M1005_g 0.0122963f $X=0.845 $Y=1.26 $X2=0 $Y2=0
cc_80 B N_C_M1005_g 0.00230876f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_81 N_B_M1007_g C 0.0055249f $X=0.845 $Y=0.475 $X2=0 $Y2=0
cc_82 N_B_c_83_n N_C_c_128_n 0.00410295f $X=0.845 $Y=1.26 $X2=0 $Y2=0
cc_83 N_B_c_88_n N_A_29_311#_M1002_g 0.00208277f $X=0.98 $Y=2.3 $X2=0 $Y2=0
cc_84 N_B_M1007_g N_A_29_311#_c_176_n 0.00808008f $X=0.845 $Y=0.475 $X2=0 $Y2=0
cc_85 N_B_c_83_n N_A_29_311#_c_177_n 0.0051802f $X=0.845 $Y=1.26 $X2=0 $Y2=0
cc_86 N_B_M1007_g N_A_29_311#_c_177_n 0.0151777f $X=0.845 $Y=0.475 $X2=0 $Y2=0
cc_87 N_B_c_83_n N_A_29_311#_c_186_n 0.00427695f $X=0.845 $Y=1.26 $X2=0 $Y2=0
cc_88 N_B_M1006_g N_A_29_311#_c_186_n 0.00379139f $X=0.9 $Y=1.765 $X2=0 $Y2=0
cc_89 B N_A_29_311#_c_186_n 0.00496204f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_90 N_B_c_88_n N_A_29_311#_c_186_n 3.69348e-19 $X=0.98 $Y=2.3 $X2=0 $Y2=0
cc_91 B N_A_29_311#_c_210_n 0.0138456f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_92 N_B_c_88_n N_A_29_311#_c_210_n 2.414e-19 $X=0.98 $Y=2.3 $X2=0 $Y2=0
cc_93 B N_A_29_311#_c_187_n 0.00127347f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_94 N_B_c_83_n N_A_29_311#_c_213_n 0.00206648f $X=0.845 $Y=1.26 $X2=0 $Y2=0
cc_95 N_B_M1006_g N_A_29_311#_c_213_n 0.0045522f $X=0.9 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B_M1006_g N_VPWR_c_290_n 0.00394037f $X=0.9 $Y=1.765 $X2=0 $Y2=0
cc_97 B N_VPWR_c_291_n 0.0314336f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_98 N_B_c_88_n N_VPWR_c_291_n 0.00627151f $X=0.98 $Y=2.3 $X2=0 $Y2=0
cc_99 N_B_M1006_g N_VPWR_c_292_n 0.00232967f $X=0.9 $Y=1.765 $X2=0 $Y2=0
cc_100 B N_VPWR_c_292_n 0.02606f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_101 N_B_c_88_n N_VPWR_c_292_n 0.00132334f $X=0.98 $Y=2.3 $X2=0 $Y2=0
cc_102 N_B_M1006_g N_VPWR_c_300_n 0.00373989f $X=0.9 $Y=1.765 $X2=0 $Y2=0
cc_103 N_B_M1006_g N_VPWR_c_296_n 0.00956409f $X=0.9 $Y=1.765 $X2=0 $Y2=0
cc_104 B N_VPWR_c_296_n 0.0275814f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_105 B N_VPWR_c_289_n 0.0169635f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_106 N_B_c_88_n N_VPWR_c_289_n 0.00893764f $X=0.98 $Y=2.3 $X2=0 $Y2=0
cc_107 N_B_M1007_g N_VGND_c_379_n 0.00382191f $X=0.845 $Y=0.475 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_VGND_c_382_n 0.00577482f $X=0.845 $Y=0.475 $X2=0 $Y2=0
cc_109 N_C_M1008_g N_A_29_311#_c_174_n 0.0141959f $X=1.25 $Y=0.475 $X2=0 $Y2=0
cc_110 C N_A_29_311#_c_174_n 5.7347e-19 $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_111 C N_A_29_311#_c_174_n 0.00248723f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_112 N_C_M1005_g N_A_29_311#_M1002_g 0.0179714f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_113 N_C_M1008_g N_A_29_311#_c_176_n 2.65899e-19 $X=1.25 $Y=0.475 $X2=0 $Y2=0
cc_114 C N_A_29_311#_c_176_n 0.0212766f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_115 N_C_M1008_g N_A_29_311#_c_177_n 6.82237e-19 $X=1.25 $Y=0.475 $X2=0 $Y2=0
cc_116 N_C_M1005_g N_A_29_311#_c_177_n 5.2097e-19 $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_117 C N_A_29_311#_c_177_n 0.0524879f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_118 N_C_c_128_n N_A_29_311#_c_177_n 4.86221e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_119 C N_A_29_311#_c_186_n 0.00109917f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_120 N_C_M1005_g N_A_29_311#_c_210_n 0.00517698f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_121 N_C_M1005_g N_A_29_311#_c_187_n 0.0100433f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_122 C N_A_29_311#_c_187_n 0.0103212f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_123 N_C_c_128_n N_A_29_311#_c_187_n 2.44767e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C_M1005_g N_A_29_311#_c_178_n 0.00213111f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_125 C N_A_29_311#_c_178_n 0.0194111f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_126 N_C_c_128_n N_A_29_311#_c_178_n 0.002428f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_127 N_C_M1005_g N_A_29_311#_c_189_n 0.00228114f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_128 C N_A_29_311#_c_189_n 0.0209596f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_129 N_C_c_128_n N_A_29_311#_c_189_n 0.00367993f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_130 C N_A_29_311#_c_179_n 8.54806e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_131 N_C_c_128_n N_A_29_311#_c_179_n 0.021264f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_132 N_C_M1005_g N_VPWR_c_291_n 0.00178962f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_133 N_C_M1005_g N_VPWR_c_292_n 0.00430676f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_134 N_C_M1005_g N_VPWR_c_300_n 2.74587e-19 $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_135 N_C_M1005_g N_VPWR_c_289_n 0.00222661f $X=1.375 $Y=1.695 $X2=0 $Y2=0
cc_136 C N_X_c_339_n 0.00573711f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_137 C X 0.00257428f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_138 C A_184_53# 0.00372867f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_139 N_C_M1008_g N_VGND_c_376_n 0.00596669f $X=1.25 $Y=0.475 $X2=0 $Y2=0
cc_140 C N_VGND_c_376_n 0.0198952f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_141 N_C_M1008_g N_VGND_c_379_n 0.00362558f $X=1.25 $Y=0.475 $X2=0 $Y2=0
cc_142 C N_VGND_c_379_n 0.0104247f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_143 C N_VGND_c_379_n 0.00277151f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_144 N_C_M1008_g N_VGND_c_382_n 0.00545964f $X=1.25 $Y=0.475 $X2=0 $Y2=0
cc_145 C N_VGND_c_382_n 0.00800021f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_146 C N_VGND_c_382_n 0.00471768f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_147 N_A_29_311#_c_183_n N_VPWR_M1000_d 2.87715e-19 $X=0.64 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_29_311#_c_213_n N_VPWR_M1000_d 0.00141996f $X=0.767 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A_29_311#_c_187_n N_VPWR_M1005_d 0.00393107f $X=1.66 $Y=1.51 $X2=0
+ $Y2=0
cc_150 N_A_29_311#_M1002_g N_VPWR_c_292_n 0.00318952f $X=1.87 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_29_311#_c_210_n N_VPWR_c_292_n 0.00593175f $X=1.165 $Y=1.725 $X2=0
+ $Y2=0
cc_152 N_A_29_311#_c_187_n N_VPWR_c_292_n 0.0138923f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A_29_311#_c_179_n N_VPWR_c_292_n 3.76018e-19 $X=2.29 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_29_311#_M1009_g N_VPWR_c_294_n 0.00588529f $X=2.29 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_29_311#_c_183_n N_VPWR_c_300_n 0.00403101f $X=0.64 $Y=1.51 $X2=0
+ $Y2=0
cc_156 N_A_29_311#_c_210_n N_VPWR_c_300_n 0.00762619f $X=1.165 $Y=1.725 $X2=0
+ $Y2=0
cc_157 N_A_29_311#_c_213_n N_VPWR_c_300_n 0.0127607f $X=0.767 $Y=1.51 $X2=0
+ $Y2=0
cc_158 N_A_29_311#_M1002_g N_VPWR_c_295_n 0.00585385f $X=1.87 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_29_311#_M1009_g N_VPWR_c_295_n 0.00541359f $X=2.29 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_29_311#_c_182_n N_VPWR_c_296_n 0.0219674f $X=0.27 $Y=1.76 $X2=0 $Y2=0
cc_161 N_A_29_311#_c_183_n N_VPWR_c_296_n 0.00511706f $X=0.64 $Y=1.51 $X2=0
+ $Y2=0
cc_162 N_A_29_311#_M1002_g N_VPWR_c_289_n 0.011733f $X=1.87 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_29_311#_M1009_g N_VPWR_c_289_n 0.0104557f $X=2.29 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_29_311#_c_182_n N_VPWR_c_289_n 0.00100952f $X=0.27 $Y=1.76 $X2=0
+ $Y2=0
cc_165 N_A_29_311#_c_174_n N_X_c_339_n 0.00252432f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_29_311#_c_175_n N_X_c_339_n 0.00913332f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_29_311#_c_179_n N_X_c_339_n 3.85946e-19 $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_29_311#_M1009_g N_X_c_348_n 0.00150631f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_29_311#_c_179_n N_X_c_348_n 8.89396e-19 $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_29_311#_M1002_g N_X_c_341_n 0.00505032f $X=1.87 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_29_311#_M1009_g N_X_c_341_n 0.0115133f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_29_311#_c_187_n N_X_c_341_n 0.0110921f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A_29_311#_c_179_n N_X_c_341_n 2.90425e-19 $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_29_311#_c_175_n X 0.00137437f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_29_311#_c_179_n X 0.00154919f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_29_311#_c_174_n X 8.79604e-19 $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_29_311#_M1002_g X 8.16932e-19 $X=1.87 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_29_311#_c_175_n X 0.0090066f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_29_311#_M1009_g X 0.0111022f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_29_311#_c_187_n X 0.00168047f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A_29_311#_c_178_n X 0.0335499f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_29_311#_c_179_n X 0.0231283f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_29_311#_c_175_n N_X_c_363_n 0.00462562f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_29_311#_M1009_g N_X_c_364_n 0.00608919f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_29_311#_c_176_n A_112_53# 0.00191292f $X=0.64 $Y=0.437 $X2=-0.19
+ $Y2=-0.24
cc_186 N_A_29_311#_c_177_n A_112_53# 0.00132529f $X=0.767 $Y=1.425 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_29_311#_c_174_n N_VGND_c_376_n 0.00937747f $X=1.855 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_29_311#_c_175_n N_VGND_c_376_n 6.48221e-19 $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_29_311#_c_178_n N_VGND_c_376_n 0.00482106f $X=1.805 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_29_311#_c_179_n N_VGND_c_376_n 5.18654e-19 $X=2.29 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_29_311#_c_175_n N_VGND_c_378_n 0.00543359f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_29_311#_c_176_n N_VGND_c_379_n 0.0355665f $X=0.64 $Y=0.437 $X2=0
+ $Y2=0
cc_193 N_A_29_311#_c_174_n N_VGND_c_380_n 0.00486043f $X=1.855 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_29_311#_c_175_n N_VGND_c_380_n 0.00541359f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_29_311#_c_174_n N_VGND_c_382_n 0.0082748f $X=1.855 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_29_311#_c_175_n N_VGND_c_382_n 0.0106216f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_29_311#_c_176_n N_VGND_c_382_n 0.0278067f $X=0.64 $Y=0.437 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_289_n N_X_M1002_d 0.0030199f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_294_n X 0.0220198f $X=2.5 $Y=1.96 $X2=0 $Y2=0
cc_200 N_VPWR_c_295_n N_X_c_364_n 0.0160313f $X=2.415 $Y=2.72 $X2=0 $Y2=0
cc_201 N_VPWR_c_289_n N_X_c_364_n 0.0103071f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_202 X N_VGND_c_378_n 0.0233099f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_203 N_X_c_363_n N_VGND_c_380_n 0.0150309f $X=2.105 $Y=0.59 $X2=0 $Y2=0
cc_204 N_X_M1003_s N_VGND_c_382_n 0.00393857f $X=1.93 $Y=0.235 $X2=0 $Y2=0
cc_205 N_X_c_363_n N_VGND_c_382_n 0.00938555f $X=2.105 $Y=0.59 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkinv_4.spice
* Created: Tue Sep  1 19:01:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkinv_4.pex.spice"
.subckt sky130_fd_sc_hd__clkinv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.1386
+ AS=0.0588 PD=1.5 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.3 SB=75001.6 A=0.063
+ P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75001.2 A=0.063
+ P=1.14 MULT=1
MM1008 N_VGND_M1003_d N_A_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.7 A=0.063
+ P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.1659
+ AS=0.0588 PD=1.63 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.3 A=0.063
+ P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.305 PD=1.28 PS=2.61 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.4
+ A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7 SB=75002 A=0.15
+ P=2.3 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1 SB=75001.6 A=0.15
+ P=2.3 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75001.1 A=0.15
+ P=2.3 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75000.7 A=0.15
+ P=2.3 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.345 PD=1.28 PS=2.69 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4 SB=75000.3
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__clkinv_4.pxi.spice"
*
.ends
*
*

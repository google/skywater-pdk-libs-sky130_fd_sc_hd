* File: sky130_fd_sc_hd__maj3_2.spice
* Created: Tue Sep  1 19:14:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__maj3_2.pex.spice"
.subckt sky130_fd_sc_hd__maj3_2  VNB VPB C A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C	C
* VPB	VPB
* VNB	VNB
MM1008 A_129_47# N_C_M1008_g N_A_47_47#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g A_129_47# VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5 SB=75002.9
+ A=0.063 P=1.14 MULT=1
MM1001 A_285_47# N_A_M1001_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_47_47#_M1002_d N_B_M1002_g A_285_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1000 A_441_47# N_B_M1000_g N_A_47_47#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_C_M1011_g A_441_47# VNB NSHORT L=0.15 W=0.42 AD=0.127354
+ AS=0.0441 PD=0.981308 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_X_M1012_d N_A_47_47#_M1012_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.197096 PD=0.92 PS=1.51869 NRD=0 NRS=41.532 M=1 R=4.33333
+ SA=75001.9 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1012_d N_A_47_47#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1755 PD=0.92 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 A_129_369# N_C_M1009_g N_A_47_47#_M1009_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1664 PD=0.85 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.3 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_129_369# VPB PHIGHVT L=0.15 W=0.64 AD=0.0864
+ AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.5
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1003 A_285_369# N_A_M1003_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001 SB=75002.5
+ A=0.096 P=1.58 MULT=1
MM1005 N_A_47_47#_M1005_d N_B_M1005_g A_285_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.3
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1014 A_441_369# N_B_M1014_g N_A_47_47#_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g A_441_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.184976 AS=0.0672 PD=1.24878 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75002.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1010_d N_A_47_47#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.289024 AS=0.135 PD=1.95122 PS=1.27 NRD=64.025 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_47_47#_M1007_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.135 PD=2.54 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__maj3_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__xnor3_1.spice.pex
* Created: Thu Aug 27 14:49:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_78_199# 1 2 9 12 14 15 16 18 19 21 23 25
+ 26 28 33 35 36 39
c97 12 0 1.74668e-19 $X=0.49 $Y=1.985
r98 35 36 15.2541 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=2.34 $Y=0.355
+ $X2=2.07 $Y2=0.355
r99 33 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.16
+ $X2=0.555 $Y2=1.325
r100 33 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.16
+ $X2=0.555 $Y2=0.995
r101 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.16 $X2=0.585 $Y2=1.16
r102 30 32 24.4 $w=1.9e-07 $l=3.8e-07 $layer=LI1_cond $X=0.602 $Y=0.78 $X2=0.602
+ $Y2=1.16
r103 26 28 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=1.22 $Y=2.32
+ $X2=2.265 $Y2=2.32
r104 25 36 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.105 $Y=0.34
+ $X2=2.07 $Y2=0.34
r105 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=2.235
+ $X2=1.22 $Y2=2.32
r106 22 23 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.135 $Y=2.045
+ $X2=1.135 $Y2=2.235
r107 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.02 $Y=0.425
+ $X2=1.105 $Y2=0.34
r108 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.02 $Y=0.425
+ $X2=1.02 $Y2=0.695
r109 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=1.96
+ $X2=1.135 $Y2=2.045
r110 18 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.05 $Y=1.96
+ $X2=0.705 $Y2=1.96
r111 17 30 1.386 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.705 $Y=0.78
+ $X2=0.602 $Y2=0.78
r112 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.935 $Y=0.78
+ $X2=1.02 $Y2=0.695
r113 16 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.935 $Y=0.78
+ $X2=0.705 $Y2=0.78
r114 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=1.875
+ $X2=0.705 $Y2=1.96
r115 14 32 10.7577 $w=1.9e-07 $l=1.73767e-07 $layer=LI1_cond $X=0.62 $Y=1.325
+ $X2=0.602 $Y2=1.16
r116 14 15 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.62 $Y=1.325
+ $X2=0.62 $Y2=1.875
r117 12 40 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.985
+ $X2=0.49 $Y2=1.325
r118 9 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
r119 2 28 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.625 $X2=2.265 $Y2=2.32
r120 1 35 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.195
+ $Y=0.245 $X2=2.34 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%C 1 3 4 6 9 11 13 15 16 17 18
c64 1 0 1.70967e-19 $X=1.005 $Y=0.995
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.16 $X2=1.915 $Y2=1.16
r66 18 22 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.07 $Y=1.2
+ $X2=1.915 $Y2=1.2
r67 16 21 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.98 $Y=1.16
+ $X2=1.915 $Y2=1.16
r68 16 17 5.03009 $w=3.3e-07 $l=1.14254e-07 $layer=POLY_cond $X=1.98 $Y=1.16
+ $X2=2.087 $Y2=1.175
r69 14 21 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=1.08 $Y=1.16
+ $X2=1.915 $Y2=1.16
r70 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.08 $Y=1.16
+ $X2=1.005 $Y2=1.16
r71 11 17 37.0704 $w=1.5e-07 $l=1.95806e-07 $layer=POLY_cond $X=2.12 $Y=0.995
+ $X2=2.087 $Y2=1.175
r72 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.12 $Y=0.995
+ $X2=2.12 $Y2=0.565
r73 7 17 37.0704 $w=1.5e-07 $l=1.95346e-07 $layer=POLY_cond $X=2.055 $Y=1.355
+ $X2=2.087 $Y2=1.175
r74 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.055 $Y=1.355
+ $X2=2.055 $Y2=2.045
r75 4 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.325
+ $X2=1.005 $Y2=1.16
r76 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.005 $Y=1.325
+ $X2=1.005 $Y2=1.805
r77 1 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.16
r78 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_216_93# 1 2 7 9 12 13 18 20 23 24 28 29 32
c75 13 0 1.74668e-19 $X=1.275 $Y=1.62
r76 29 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.54 $Y=1.16
+ $X2=2.54 $Y2=0.995
r77 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.16 $X2=2.54 $Y2=1.16
r78 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.435 $Y=1.16
+ $X2=2.54 $Y2=1.16
r79 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=1.325
+ $X2=2.435 $Y2=1.16
r80 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.435 $Y=1.325
+ $X2=2.435 $Y2=1.535
r81 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=1.62
+ $X2=1.36 $Y2=1.62
r82 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.35 $Y=1.62
+ $X2=2.435 $Y2=1.535
r83 20 21 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.35 $Y=1.62
+ $X2=1.445 $Y2=1.62
r84 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=1.535
+ $X2=1.36 $Y2=1.62
r85 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.36 $Y=1.535
+ $X2=1.36 $Y2=0.76
r86 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.62
+ $X2=1.36 $Y2=1.62
r87 13 15 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=1.275 $Y=1.62 $X2=1.215
+ $Y2=1.62
r88 12 32 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.56 $Y=0.565
+ $X2=2.56 $Y2=0.995
r89 7 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.54 $Y=1.325
+ $X2=2.54 $Y2=1.16
r90 7 9 186.373 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.54 $Y=1.325 $X2=2.54
+ $Y2=1.905
r91 2 15 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.485 $X2=1.215 $Y2=1.62
r92 1 18 182 $w=1.7e-07 $l=4.11856e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.465 $X2=1.36 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_735_297# 1 2 9 13 15 17 19 21 22 23 27 35
+ 37 38 39 40 47 49 50 58
c169 49 0 1.83334e-19 $X=6.67 $Y=0.85
c170 27 0 1.36535e-19 $X=3.945 $Y=1.58
c171 15 0 1.24749e-19 $X=6.845 $Y=1.28
r172 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=1.11 $X2=6.79 $Y2=1.11
r173 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.72 $Y=0.85
+ $X2=6.72 $Y2=1.11
r174 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0.85
+ $X2=6.67 $Y2=0.85
r175 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.85
r176 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0.85
+ $X2=3.91 $Y2=0.85
r177 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=0.85
+ $X2=5.29 $Y2=0.85
r178 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.525 $Y=0.85
+ $X2=6.67 $Y2=0.85
r179 39 40 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=6.525 $Y=0.85
+ $X2=5.435 $Y2=0.85
r180 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=0.85
+ $X2=3.91 $Y2=0.85
r181 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=0.85
+ $X2=5.29 $Y2=0.85
r182 37 38 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=5.145 $Y=0.85
+ $X2=4.055 $Y2=0.85
r183 35 47 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.85
r184 31 35 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=5.12 $Y=1.132
+ $X2=5.27 $Y2=1.132
r185 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.16 $X2=5.12 $Y2=1.16
r186 28 58 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=3.945 $Y=1.445
+ $X2=3.945 $Y2=0.74
r187 27 28 1.42499 $w=2.4e-07 $l=1.35e-07 $layer=LI1_cond $X=3.945 $Y=1.58
+ $X2=3.945 $Y2=1.445
r188 25 27 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.81 $Y=1.58
+ $X2=3.945 $Y2=1.58
r189 22 32 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=5.38 $Y=1.16
+ $X2=5.12 $Y2=1.16
r190 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.38 $Y=1.16
+ $X2=5.455 $Y2=1.16
r191 19 55 38.945 $w=2.68e-07 $l=1.92678e-07 $layer=POLY_cond $X=6.85 $Y=0.945
+ $X2=6.79 $Y2=1.11
r192 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=6.85 $Y=0.945
+ $X2=6.85 $Y2=0.535
r193 15 55 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=6.845 $Y=1.28
+ $X2=6.79 $Y2=1.11
r194 15 17 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.845 $Y=1.28
+ $X2=6.845 $Y2=2.065
r195 11 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.325
+ $X2=5.455 $Y2=1.16
r196 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.455 $Y=1.325
+ $X2=5.455 $Y2=1.805
r197 7 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=0.995
+ $X2=5.455 $Y2=1.16
r198 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.455 $Y=0.995
+ $X2=5.455 $Y2=0.455
r199 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.81 $Y2=1.63
r200 1 58 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.235 $X2=3.98 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%B 3 7 9 10 13 18 19 20 23 27 31 34 35 37 38
+ 41
r121 37 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.395 $Y=1.53
+ $X2=6.67 $Y2=1.53
r122 35 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.16
+ $X2=6.31 $Y2=1.325
r123 35 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.16
+ $X2=6.31 $Y2=0.995
r124 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.16 $X2=6.31 $Y2=1.16
r125 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.31 $Y=1.445
+ $X2=6.395 $Y2=1.53
r126 32 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.31 $Y=1.445
+ $X2=6.31 $Y2=1.16
r127 28 30 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.6 $Y=1.16
+ $X2=3.77 $Y2=1.16
r128 27 42 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.33 $Y=1.965
+ $X2=6.33 $Y2=1.325
r129 25 27 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.33 $Y=2.465
+ $X2=6.33 $Y2=1.965
r130 23 41 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.25 $Y=0.565
+ $X2=6.25 $Y2=0.995
r131 19 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.255 $Y=2.54
+ $X2=6.33 $Y2=2.465
r132 19 20 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=6.255 $Y=2.54
+ $X2=4.775 $Y2=2.54
r133 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.7 $Y=2.465
+ $X2=4.775 $Y2=2.54
r134 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.7 $Y=2.465
+ $X2=4.7 $Y2=1.905
r135 15 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.7 $Y=1.235
+ $X2=4.7 $Y2=1.16
r136 15 18 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.7 $Y=1.235
+ $X2=4.7 $Y2=1.905
r137 11 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.7 $Y=1.085
+ $X2=4.7 $Y2=1.16
r138 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=4.7 $Y=1.085
+ $X2=4.7 $Y2=0.565
r139 10 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=1.16
+ $X2=3.77 $Y2=1.16
r140 9 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.625 $Y=1.16
+ $X2=4.7 $Y2=1.16
r141 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.625 $Y=1.16
+ $X2=3.845 $Y2=1.16
r142 5 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=1.085
+ $X2=3.77 $Y2=1.16
r143 5 7 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.77 $Y=1.085
+ $X2=3.77 $Y2=0.56
r144 1 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.6 $Y=1.235 $X2=3.6
+ $Y2=1.16
r145 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.6 $Y=1.235 $X2=3.6
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A 3 6 8 11 12 13
c44 13 0 1.83334e-19 $X=7.28 $Y=0.995
r45 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.28 $Y=1.16
+ $X2=7.28 $Y2=1.325
r46 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.28 $Y=1.16
+ $X2=7.28 $Y2=0.995
r47 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.16 $X2=7.27 $Y2=1.16
r48 8 12 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=7.13 $Y=1.2 $X2=7.27
+ $Y2=1.2
r49 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.35 $Y=1.985
+ $X2=7.35 $Y2=1.325
r50 3 13 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.35 $Y=0.555
+ $X2=7.35 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_841_297# 1 2 3 4 13 15 18 22 24 28 29 30
+ 31 36 37 38 41 44 45
c135 36 0 1.4656e-19 $X=7.77 $Y=1.16
c136 31 0 1.06604e-19 $X=7.71 $Y=1.495
c137 30 0 1.40536e-19 $X=7.71 $Y=1.325
r138 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.51
+ $X2=7.13 $Y2=0.51
r139 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0.51
+ $X2=4.37 $Y2=0.51
r140 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=0.51
+ $X2=4.37 $Y2=0.51
r141 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.51
+ $X2=7.13 $Y2=0.51
r142 37 38 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=6.985 $Y=0.51
+ $X2=4.515 $Y2=0.51
r143 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.77
+ $Y=1.16 $X2=7.77 $Y2=1.16
r144 33 35 20.4335 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=7.74 $Y=0.82
+ $X2=7.74 $Y2=1.16
r145 32 45 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=7.16 $Y=0.735
+ $X2=7.16 $Y2=0.51
r146 30 35 10.2745 $w=2.03e-07 $l=1.79374e-07 $layer=LI1_cond $X=7.71 $Y=1.325
+ $X2=7.74 $Y2=1.16
r147 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.71 $Y=1.325
+ $X2=7.71 $Y2=1.495
r148 29 32 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.305 $Y=0.82
+ $X2=7.16 $Y2=0.735
r149 28 33 1.77774 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.625 $Y=0.82
+ $X2=7.74 $Y2=0.82
r150 28 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.625 $Y=0.82
+ $X2=7.305 $Y2=0.82
r151 24 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.625 $Y=1.6
+ $X2=7.71 $Y2=1.495
r152 24 26 25.6147 $w=2.08e-07 $l=4.85e-07 $layer=LI1_cond $X=7.625 $Y=1.6
+ $X2=7.14 $Y2=1.6
r153 20 41 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=0.595
+ $X2=4.33 $Y2=0.43
r154 20 22 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.33 $Y=0.595
+ $X2=4.33 $Y2=1.94
r155 16 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.77 $Y=1.325
+ $X2=7.77 $Y2=1.16
r156 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.77 $Y=1.325
+ $X2=7.77 $Y2=1.985
r157 13 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.77 $Y=0.995
+ $X2=7.77 $Y2=1.16
r158 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.77 $Y=0.995
+ $X2=7.77 $Y2=0.555
r159 4 26 600 $w=1.7e-07 $l=2.32164e-07 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.645 $X2=7.14 $Y2=1.62
r160 3 22 600 $w=1.7e-07 $l=5.13712e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.485 $X2=4.33 $Y2=1.94
r161 2 45 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=6.925
+ $Y=0.235 $X2=7.14 $Y2=0.625
r162 1 41 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.365
+ $Y=0.245 $X2=4.49 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%X 1 2 9 13 14 15 16 19
r21 16 23 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=2.3
r22 16 19 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.62
r23 14 19 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=0.225 $Y=1.58
+ $X2=0.225 $Y2=1.62
r24 14 15 5.97229 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=1.58
+ $X2=0.225 $Y2=1.44
r25 13 15 24.2248 $w=2.43e-07 $l=5.15e-07 $layer=LI1_cond $X=0.207 $Y=0.925
+ $X2=0.207 $Y2=1.44
r26 7 13 5.81426 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=0.795
+ $X2=0.215 $Y2=0.925
r27 7 9 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=0.215 $Y=0.795
+ $X2=0.215 $Y2=0.56
r28 2 23 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r29 2 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r30 1 9 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%VPWR 1 2 3 12 16 20 22 24 29 37 47 48 51 54
+ 57
c91 3 0 1.06604e-19 $X=7.425 $Y=1.485
r92 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r93 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r94 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 48 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r96 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r97 45 57 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.73 $Y=2.72
+ $X2=7.562 $Y2=2.72
r98 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.73 $Y=2.72 $X2=8.05
+ $Y2=2.72
r99 44 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r100 43 44 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r101 41 44 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=7.13 $Y2=2.72
r102 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r103 40 43 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=7.13 $Y2=2.72
r104 40 41 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r105 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=2.72
+ $X2=3.39 $Y2=2.72
r106 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.555 $Y=2.72
+ $X2=3.91 $Y2=2.72
r107 37 57 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.395 $Y=2.72
+ $X2=7.562 $Y2=2.72
r108 37 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.395 $Y=2.72
+ $X2=7.13 $Y2=2.72
r109 36 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r110 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r111 33 36 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r112 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 32 35 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r114 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r115 30 51 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.702 $Y2=2.72
r116 30 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=2.72
+ $X2=3.39 $Y2=2.72
r118 29 35 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r119 24 51 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.702 $Y2=2.72
r120 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r121 22 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r123 18 57 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.562 $Y=2.635
+ $X2=7.562 $Y2=2.72
r124 18 20 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=7.562 $Y=2.635
+ $X2=7.562 $Y2=2.36
r125 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.39 $Y=2.635
+ $X2=3.39 $Y2=2.72
r126 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.39 $Y=2.635
+ $X2=3.39 $Y2=2.32
r127 10 51 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.702 $Y=2.635
+ $X2=0.702 $Y2=2.72
r128 10 12 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.702 $Y=2.635
+ $X2=0.702 $Y2=2.3
r129 3 20 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=2.36
r130 2 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=2.175 $X2=3.39 $Y2=2.32
r131 1 12 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.705 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_331_325# 1 2 3 4 13 17 22 24 25 28 29 30
+ 32 35 39 43 45 46 48
c149 29 0 1.36535e-19 $X=4.585 $Y=2.36
r150 46 47 14.9388 $w=1.96e-07 $l=2.4e-07 $layer=LI1_cond $X=4.67 $Y=0.772
+ $X2=4.91 $Y2=0.772
r151 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.22 $Y=1.12
+ $X2=3.33 $Y2=1.12
r152 37 47 1.57051 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.91 $Y=0.655
+ $X2=4.91 $Y2=0.772
r153 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.91 $Y=0.655
+ $X2=4.91 $Y2=0.545
r154 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=2.36
+ $X2=4.67 $Y2=2.36
r155 33 35 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=4.755 $Y=2.36
+ $X2=6.625 $Y2=2.36
r156 32 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=2.275
+ $X2=4.67 $Y2=2.36
r157 31 46 1.57051 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.67 $Y=0.89
+ $X2=4.67 $Y2=0.772
r158 31 32 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.67 $Y=0.89
+ $X2=4.67 $Y2=2.275
r159 29 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=2.36
+ $X2=4.67 $Y2=2.36
r160 29 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.585 $Y=2.36
+ $X2=4.06 $Y2=2.36
r161 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=2.275
+ $X2=4.06 $Y2=2.36
r162 27 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.975 $Y=2.065
+ $X2=3.975 $Y2=2.275
r163 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.98
+ $X2=3.33 $Y2=1.98
r164 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=1.98
+ $X2=3.975 $Y2=2.065
r165 25 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.89 $Y=1.98
+ $X2=3.415 $Y2=1.98
r166 24 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.895
+ $X2=3.33 $Y2=1.98
r167 23 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.205
+ $X2=3.33 $Y2=1.12
r168 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.33 $Y=1.205
+ $X2=3.33 $Y2=1.895
r169 22 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.035
+ $X2=3.22 $Y2=1.12
r170 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.22 $Y=0.455
+ $X2=3.22 $Y2=1.035
r171 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.135 $Y=0.37
+ $X2=3.22 $Y2=0.455
r172 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.135 $Y=0.37
+ $X2=2.84 $Y2=0.37
r173 13 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=1.98
+ $X2=3.33 $Y2=1.98
r174 13 15 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.245 $Y=1.98
+ $X2=1.845 $Y2=1.98
r175 4 35 600 $w=1.7e-07 $l=8.17634e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=1.645 $X2=6.625 $Y2=2.36
r176 3 15 600 $w=1.7e-07 $l=4.39858e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.625 $X2=1.845 $Y2=1.98
r177 2 39 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.245 $X2=4.91 $Y2=0.545
r178 1 19 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.245 $X2=2.84 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_355_49# 1 2 3 4 13 16 17 19 21 24 26 30 32
+ 33 35 36 39 42
c129 32 0 1.24749e-19 $X=6.47 $Y=0.38
r130 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.53
+ $X2=5.29 $Y2=1.53
r131 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.53
+ $X2=2.99 $Y2=1.53
r132 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.53
+ $X2=2.99 $Y2=1.53
r133 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.53
+ $X2=5.29 $Y2=1.53
r134 35 36 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=5.145 $Y=1.53
+ $X2=3.135 $Y2=1.53
r135 32 33 13.3743 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=6.47 $Y=0.36
+ $X2=6.225 $Y2=0.36
r136 28 30 10.6148 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.91 $Y=0.765
+ $X2=2.125 $Y2=0.765
r137 26 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.715 $Y=0.34
+ $X2=6.225 $Y2=0.34
r138 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.63 $Y=0.425
+ $X2=5.715 $Y2=0.34
r139 23 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=5.63 $Y=0.425
+ $X2=5.63 $Y2=1.445
r140 22 43 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=5.35 $Y=1.53
+ $X2=5.142 $Y2=1.53
r141 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.545 $Y=1.53
+ $X2=5.63 $Y2=1.445
r142 21 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.545 $Y=1.53
+ $X2=5.35 $Y2=1.53
r143 17 43 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.142 $Y=1.615
+ $X2=5.142 $Y2=1.53
r144 17 19 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=5.142 $Y=1.615
+ $X2=5.142 $Y2=1.62
r145 16 39 8.59825 $w=3.35e-07 $l=1.55997e-07 $layer=LI1_cond $X=2.88 $Y=1.375
+ $X2=2.882 $Y2=1.53
r146 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.88 $Y=0.795
+ $X2=2.88 $Y2=1.375
r147 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.795 $Y=0.71
+ $X2=2.88 $Y2=0.795
r148 13 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.795 $Y=0.71
+ $X2=2.125 $Y2=0.71
r149 4 19 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=4.775
+ $Y=1.485 $X2=5.11 $Y2=1.62
r150 3 39 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=1.485 $X2=2.855 $Y2=1.61
r151 2 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.325
+ $Y=0.245 $X2=6.47 $Y2=0.38
r152 1 28 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.245 $X2=1.91 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%A_1106_49# 1 2 3 4 15 18 23 26 29 31 36
c67 29 0 1.17772e-19 $X=7.71 $Y=1.99
r68 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.98 $Y=0.42
+ $X2=8.11 $Y2=0.42
r69 28 29 14.5869 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.985 $Y=1.99
+ $X2=7.71 $Y2=1.99
r70 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.11 $Y=1.875
+ $X2=8.11 $Y2=1.99
r71 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.11 $Y=0.585
+ $X2=8.11 $Y2=0.42
r72 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=8.11 $Y=0.585
+ $X2=8.11 $Y2=1.875
r73 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=8.047 $Y=1.99
+ $X2=8.11 $Y2=1.99
r74 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=8.047 $Y=1.99
+ $X2=7.985 $Y2=1.99
r75 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=8.047 $Y=2.105
+ $X2=8.047 $Y2=2.3
r76 20 29 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=6.12 $Y=2.02
+ $X2=7.71 $Y2=2.02
r77 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.055 $Y=2.02
+ $X2=6.12 $Y2=2.02
r78 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.97 $Y=1.935
+ $X2=6.055 $Y2=2.02
r79 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=5.97 $Y=1.935
+ $X2=5.97 $Y2=0.76
r80 4 28 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=7.845
+ $Y=1.485 $X2=7.985 $Y2=1.96
r81 4 23 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=7.845
+ $Y=1.485 $X2=7.985 $Y2=2.3
r82 3 20 600 $w=1.7e-07 $l=8.14709e-07 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=1.485 $X2=6.12 $Y2=2.02
r83 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.845
+ $Y=0.235 $X2=7.98 $Y2=0.42
r84 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=5.53
+ $Y=0.245 $X2=5.97 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_1%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
c101 47 0 1.70967e-19 $X=8.05 $Y=0
c102 20 0 2.87884e-20 $X=7.56 $Y=0.4
c103 3 0 1.40536e-19 $X=7.425 $Y=0.235
r104 50 51 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r105 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r106 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r107 43 44 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r108 41 44 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=7.13 $Y2=0
r109 40 43 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=7.13
+ $Y2=0
r110 40 41 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r111 38 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r112 38 51 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=0.69 $Y2=0
r113 37 38 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r114 35 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.64
+ $Y2=0
r115 35 37 175.171 $w=1.68e-07 $l=2.685e-06 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=3.45 $Y2=0
r116 30 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.64
+ $Y2=0
r117 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r118 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 26 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.475 $Y=0 $X2=7.13
+ $Y2=0
r121 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.475 $Y=0 $X2=7.56
+ $Y2=0
r122 25 46 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.645 $Y=0
+ $X2=8.05 $Y2=0
r123 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.645 $Y=0 $X2=7.56
+ $Y2=0
r124 23 37 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.45
+ $Y2=0
r125 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.56
+ $Y2=0
r126 22 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.645 $Y=0
+ $X2=3.91 $Y2=0
r127 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.56
+ $Y2=0
r128 18 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=0.085
+ $X2=7.56 $Y2=0
r129 18 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.56 $Y=0.085
+ $X2=7.56 $Y2=0.4
r130 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0
r131 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0.36
r132 10 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=0.085
+ $X2=0.64 $Y2=0
r133 10 12 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.64 $Y=0.085
+ $X2=0.64 $Y2=0.36
r134 3 20 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.56 $Y2=0.4
r135 2 16 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.235 $X2=3.56 $Y2=0.36
r136 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
M1000 a_316_47# B a_232_47# VNB nshort w=650000u l=150000u
+  ad=2.5025e+11p pd=2.07e+06u as=1.755e+11p ps=1.84e+06u
M1001 VPWR B Y VPB phighvt w=1e+06u l=150000u
+  ad=6.765e+11p pd=5.44e+06u as=5.5e+11p ps=5.1e+06u
M1002 a_232_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.005e+11p ps=1.97e+06u
M1003 VPWR A_N a_53_93# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1004 VGND A_N a_53_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 Y a_53_93# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_53_93# a_316_47# VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1007 Y C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

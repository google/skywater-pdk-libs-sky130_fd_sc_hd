# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_3
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 1.295000 2.465000 ;
        RECT 0.775000 1.005000 1.295000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.085000 2.080000 1.295000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 1.380000 0.085000 ;
        RECT 0.085000  0.085000 1.295000 0.835000 ;
        RECT 0.085000  0.835000 0.605000 1.375000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 1.380000 2.805000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
END sky130_fd_sc_hd__lpflow_decapkapwr_3

* File: sky130_fd_sc_hd__a21oi_4.spice
* Created: Thu Aug 27 14:01:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a21oi_4  VNB VPB B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_Y_M1008_d N_B1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75005
+ A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1008_d N_B1_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75004.5
+ A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1014_d N_B1_M1014_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1 SB=75004.1
+ A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1014_d N_B1_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.104 PD=0.93 PS=0.97 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75001.5 SB=75003.7
+ A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1023_s N_A2_M1000_g N_A_462_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.091 PD=0.97 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_462_47#_M1000_s N_A1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1004 N_A_462_47#_M1004_d N_A1_M1004_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1018 N_A_462_47#_M1004_d N_A1_M1018_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1019 N_A_462_47#_M1019_d N_A1_M1019_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_462_47#_M1019_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1005_d N_A2_M1017_g N_A_462_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A2_M1021_g N_A_462_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_28_297#_M1006_d N_B1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75005
+ A=0.15 P=2.3 MULT=1
MM1011 N_A_28_297#_M1011_d N_B1_M1011_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1012 N_A_28_297#_M1011_d N_B1_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75004.1
+ A=0.15 P=2.3 MULT=1
MM1022 N_A_28_297#_M1022_d N_B1_M1022_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.14 PD=1.31 PS=1.28 NRD=5.8903 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_28_297#_M1022_d VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.155 PD=1.29 PS=1.31 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1001_d N_A1_M1002_g N_A_28_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.14 PD=1.29 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_28_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1007_d N_A1_M1009_g N_A_28_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A1_M1015_g N_A_28_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.7
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1015_d N_A2_M1010_g N_A_28_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_A2_M1016_g N_A_28_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1016_d N_A2_M1020_g N_A_28_297#_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75005 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_48 VNB 0 1.1531e-19 $X=0.15 $Y=-0.085
c_88 VPB 0 3.12905e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__a21oi_4.pxi.spice"
*
.ends
*
*

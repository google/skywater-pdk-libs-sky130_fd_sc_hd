* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR B2 a_397_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.3e+11p pd=5.06e+06u as=5.3e+11p ps=5.06e+06u
M1001 a_481_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=1.755e+11p ps=1.84e+06u
M1002 Y a_109_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=9.035e+11p ps=6.68e+06u
M1003 a_397_297# a_109_47# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.4e+11p ps=2.68e+06u
M1004 VGND B1 a_481_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_109_47# A2_N a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1006 VGND A2_N a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1007 a_109_297# A1_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_109_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_397_297# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__o21ai_4.spice
* Created: Thu Aug 27 14:35:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21ai_4.pex.spice"
.subckt sky130_fd_sc_hd__o21ai_4  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A1_M1012_g N_A_32_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1012_d N_A1_M1017_g N_A_32_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A1_M1021_g N_A_32_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1021_d N_A2_M1005_g N_A_32_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_32_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1009_d N_A2_M1018_g N_A_32_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A2_M1019_g N_A_32_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.091 PD=0.97 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1019_d N_A1_M1022_g N_A_32_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.091 PD=0.97 PS=0.93 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_32_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1001_d N_B1_M1003_g N_A_32_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1010_d N_B1_M1010_g N_A_32_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1010_d N_B1_M1015_g N_A_32_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.18525 PD=0.93 PS=1.87 NRD=0 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_115_297#_M1002_d N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75005
+ A=0.15 P=2.3 MULT=1
MM1004 N_A_115_297#_M1002_d N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1007 N_A_115_297#_M1007_d N_A1_M1007_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75004.1
+ A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g N_A_115_297#_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1000_d N_A2_M1008_g N_A_115_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1013 N_Y_M1013_d N_A2_M1013_g N_A_115_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1016 N_Y_M1013_d N_A2_M1016_g N_A_115_297#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1020 N_A_115_297#_M1016_s N_A1_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.16 PD=1.28 PS=1.32 NRD=0 NRS=3.9203 M=1 R=6.66667 SA=75003.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1020_s N_B1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75003.7 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_B1_M1011_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1014 N_VPWR_M1011_d N_B1_M1014_g N_Y_M1014_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_B1_M1023_g N_Y_M1014_s VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75005 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__o21ai_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__dfstp_2.pxi.spice
* Created: Thu Aug 27 14:15:22 2020
* 
x_PM_SKY130_FD_SC_HD__DFSTP_2%CLK N_CLK_c_227_n N_CLK_c_222_n N_CLK_M1029_g
+ N_CLK_c_228_n N_CLK_M1017_g N_CLK_c_223_n N_CLK_c_229_n CLK CLK N_CLK_c_225_n
+ N_CLK_c_226_n PM_SKY130_FD_SC_HD__DFSTP_2%CLK
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_27_47# N_A_27_47#_M1029_s N_A_27_47#_M1017_s
+ N_A_27_47#_M1019_g N_A_27_47#_M1000_g N_A_27_47#_c_267_n N_A_27_47#_M1028_g
+ N_A_27_47#_M1031_g N_A_27_47#_M1005_g N_A_27_47#_M1012_g N_A_27_47#_c_268_n
+ N_A_27_47#_c_269_n N_A_27_47#_c_270_n N_A_27_47#_c_284_n N_A_27_47#_c_386_p
+ N_A_27_47#_c_271_n N_A_27_47#_c_272_n N_A_27_47#_c_273_n N_A_27_47#_c_274_n
+ N_A_27_47#_c_275_n N_A_27_47#_c_276_n N_A_27_47#_c_288_n N_A_27_47#_c_277_n
+ N_A_27_47#_c_278_n N_A_27_47#_c_289_n N_A_27_47#_c_290_n N_A_27_47#_c_291_n
+ N_A_27_47#_c_292_n N_A_27_47#_c_293_n N_A_27_47#_c_279_n N_A_27_47#_c_295_n
+ N_A_27_47#_c_296_n N_A_27_47#_c_297_n N_A_27_47#_c_298_n N_A_27_47#_c_280_n
+ PM_SKY130_FD_SC_HD__DFSTP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DFSTP_2%D N_D_M1010_g N_D_M1023_g D D N_D_c_548_n
+ N_D_c_549_n PM_SKY130_FD_SC_HD__DFSTP_2%D
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_193_47# N_A_193_47#_M1019_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1011_g N_A_193_47#_c_589_n N_A_193_47#_c_590_n
+ N_A_193_47#_M1018_g N_A_193_47#_c_592_n N_A_193_47#_M1014_g
+ N_A_193_47#_c_594_n N_A_193_47#_M1024_g N_A_193_47#_c_595_n
+ N_A_193_47#_c_614_n N_A_193_47#_c_596_n N_A_193_47#_c_615_n
+ N_A_193_47#_c_597_n N_A_193_47#_c_598_n N_A_193_47#_c_599_n
+ N_A_193_47#_c_600_n N_A_193_47#_c_601_n N_A_193_47#_c_602_n
+ N_A_193_47#_c_603_n N_A_193_47#_c_604_n N_A_193_47#_c_605_n
+ N_A_193_47#_c_606_n N_A_193_47#_c_607_n PM_SKY130_FD_SC_HD__DFSTP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_652_21# N_A_652_21#_M1007_d N_A_652_21#_M1026_d
+ N_A_652_21#_M1022_g N_A_652_21#_M1009_g N_A_652_21#_c_803_n
+ N_A_652_21#_c_887_p N_A_652_21#_c_804_n N_A_652_21#_c_798_n
+ N_A_652_21#_c_799_n N_A_652_21#_c_806_n N_A_652_21#_c_807_n
+ N_A_652_21#_c_808_n N_A_652_21#_c_800_n PM_SKY130_FD_SC_HD__DFSTP_2%A_652_21#
x_PM_SKY130_FD_SC_HD__DFSTP_2%SET_B N_SET_B_c_912_n N_SET_B_M1026_g
+ N_SET_B_M1004_g N_SET_B_M1002_g N_SET_B_c_916_n N_SET_B_M1001_g
+ N_SET_B_c_927_n N_SET_B_c_917_n N_SET_B_c_918_n SET_B N_SET_B_c_920_n
+ N_SET_B_c_921_n N_SET_B_c_922_n N_SET_B_c_923_n
+ PM_SKY130_FD_SC_HD__DFSTP_2%SET_B
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_476_47# N_A_476_47#_M1028_d N_A_476_47#_M1011_d
+ N_A_476_47#_c_1047_n N_A_476_47#_M1007_g N_A_476_47#_c_1048_n
+ N_A_476_47#_M1020_g N_A_476_47#_c_1049_n N_A_476_47#_M1016_g
+ N_A_476_47#_c_1050_n N_A_476_47#_M1021_g N_A_476_47#_c_1051_n
+ N_A_476_47#_c_1074_n N_A_476_47#_c_1079_n N_A_476_47#_c_1059_n
+ N_A_476_47#_c_1052_n N_A_476_47#_c_1053_n N_A_476_47#_c_1054_n
+ N_A_476_47#_c_1055_n N_A_476_47#_c_1056_n
+ PM_SKY130_FD_SC_HD__DFSTP_2%A_476_47#
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_1178_261# N_A_1178_261#_M1013_d
+ N_A_1178_261#_M1027_d N_A_1178_261#_M1015_g N_A_1178_261#_M1033_g
+ N_A_1178_261#_c_1205_n N_A_1178_261#_c_1210_n N_A_1178_261#_c_1211_n
+ N_A_1178_261#_c_1264_p N_A_1178_261#_c_1206_n N_A_1178_261#_c_1213_n
+ N_A_1178_261#_c_1214_n N_A_1178_261#_c_1207_n
+ PM_SKY130_FD_SC_HD__DFSTP_2%A_1178_261#
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_1028_413# N_A_1028_413#_M1014_d
+ N_A_1028_413#_M1005_d N_A_1028_413#_M1001_s N_A_1028_413#_M1027_g
+ N_A_1028_413#_M1013_g N_A_1028_413#_c_1284_n N_A_1028_413#_c_1285_n
+ N_A_1028_413#_M1030_g N_A_1028_413#_c_1296_n N_A_1028_413#_M1006_g
+ N_A_1028_413#_c_1287_n N_A_1028_413#_c_1305_n N_A_1028_413#_c_1298_n
+ N_A_1028_413#_c_1313_n N_A_1028_413#_c_1288_n N_A_1028_413#_c_1289_n
+ N_A_1028_413#_c_1300_n N_A_1028_413#_c_1290_n N_A_1028_413#_c_1301_n
+ N_A_1028_413#_c_1302_n N_A_1028_413#_c_1384_n N_A_1028_413#_c_1291_n
+ N_A_1028_413#_c_1292_n PM_SKY130_FD_SC_HD__DFSTP_2%A_1028_413#
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_1602_47# N_A_1602_47#_M1030_s
+ N_A_1602_47#_M1006_s N_A_1602_47#_c_1442_n N_A_1602_47#_M1003_g
+ N_A_1602_47#_M1025_g N_A_1602_47#_c_1443_n N_A_1602_47#_M1008_g
+ N_A_1602_47#_M1032_g N_A_1602_47#_c_1444_n N_A_1602_47#_c_1450_n
+ N_A_1602_47#_c_1445_n N_A_1602_47#_c_1452_n N_A_1602_47#_c_1446_n
+ N_A_1602_47#_c_1447_n PM_SKY130_FD_SC_HD__DFSTP_2%A_1602_47#
x_PM_SKY130_FD_SC_HD__DFSTP_2%VPWR N_VPWR_M1017_d N_VPWR_M1023_s N_VPWR_M1009_d
+ N_VPWR_M1020_d N_VPWR_M1015_d N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_M1032_d
+ N_VPWR_c_1518_n N_VPWR_c_1519_n N_VPWR_c_1520_n N_VPWR_c_1521_n
+ N_VPWR_c_1522_n N_VPWR_c_1523_n N_VPWR_c_1524_n N_VPWR_c_1525_n VPWR VPWR
+ N_VPWR_c_1526_n N_VPWR_c_1527_n N_VPWR_c_1528_n N_VPWR_c_1529_n
+ N_VPWR_c_1530_n N_VPWR_c_1531_n N_VPWR_c_1532_n N_VPWR_c_1533_n
+ N_VPWR_c_1534_n N_VPWR_c_1535_n N_VPWR_c_1536_n N_VPWR_c_1537_n
+ N_VPWR_c_1538_n N_VPWR_c_1539_n N_VPWR_c_1517_n
+ PM_SKY130_FD_SC_HD__DFSTP_2%VPWR
x_PM_SKY130_FD_SC_HD__DFSTP_2%A_381_47# N_A_381_47#_M1010_d N_A_381_47#_M1023_d
+ N_A_381_47#_c_1688_n N_A_381_47#_c_1693_n N_A_381_47#_c_1689_n
+ N_A_381_47#_c_1695_n N_A_381_47#_c_1691_n N_A_381_47#_c_1697_n
+ N_A_381_47#_c_1698_n PM_SKY130_FD_SC_HD__DFSTP_2%A_381_47#
x_PM_SKY130_FD_SC_HD__DFSTP_2%Q N_Q_M1003_s N_Q_M1025_s Q Q Q Q Q Q N_Q_c_1758_n
+ N_Q_c_1771_n N_Q_c_1756_n Q PM_SKY130_FD_SC_HD__DFSTP_2%Q
x_PM_SKY130_FD_SC_HD__DFSTP_2%VGND N_VGND_M1029_d N_VGND_M1010_s N_VGND_M1022_d
+ N_VGND_M1021_s N_VGND_M1002_d N_VGND_M1030_d N_VGND_M1008_d N_VGND_c_1787_n
+ N_VGND_c_1788_n N_VGND_c_1789_n N_VGND_c_1790_n N_VGND_c_1791_n
+ N_VGND_c_1792_n N_VGND_c_1793_n N_VGND_c_1794_n VGND VGND N_VGND_c_1795_n
+ N_VGND_c_1796_n N_VGND_c_1797_n N_VGND_c_1798_n N_VGND_c_1799_n
+ N_VGND_c_1800_n N_VGND_c_1801_n N_VGND_c_1802_n N_VGND_c_1803_n
+ N_VGND_c_1804_n N_VGND_c_1805_n N_VGND_c_1806_n N_VGND_c_1807_n
+ PM_SKY130_FD_SC_HD__DFSTP_2%VGND
cc_1 VNB N_CLK_c_222_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_223_n 0.0233701f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK 0.016129f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_c_225_n 0.0195341f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_CLK_c_226_n 0.0141401f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1019_g 0.0365111f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_267_n 0.0180457f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_8 VNB N_A_27_47#_c_268_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_9 VNB N_A_27_47#_c_269_n 0.00157584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_270_n 0.00786724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_271_n 0.00246572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_272_n 0.00445416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_273_n 0.0327378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_274_n 0.00637933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_275_n 0.00815721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_276_n 0.00156937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_277_n 0.00533129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_278_n 0.0270495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_279_n 0.0229519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_280_n 0.0161153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_D_M1010_g 0.0205663f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_22 VNB N_D_c_548_n 0.0258802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_D_c_549_n 0.00442451f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_24 VNB N_A_193_47#_c_589_n 0.0132632f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_25 VNB N_A_193_47#_c_590_n 0.00435992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_M1018_g 0.0199482f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_27 VNB N_A_193_47#_c_592_n 0.00803437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_M1014_g 0.034159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_c_594_n 0.0101649f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_30 VNB N_A_193_47#_c_595_n 0.018279f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_31 VNB N_A_193_47#_c_596_n 0.00411907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_597_n 0.0194566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_598_n 0.0054023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_599_n 0.00105673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_600_n 0.016384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_601_n 0.00113053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_602_n 0.011972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_603_n 0.00189817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_604_n 0.00500582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_605_n 0.00145914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_193_47#_c_606_n 0.00217053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_193_47#_c_607_n 0.0246637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_652_21#_M1022_g 0.0422386f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_44 VNB N_A_652_21#_c_798_n 0.00136482f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_45 VNB N_A_652_21#_c_799_n 0.00314488f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_46 VNB N_A_652_21#_c_800_n 0.00513705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_SET_B_c_912_n 0.0308821f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_48 VNB N_SET_B_M1026_g 0.00706345f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_49 VNB N_SET_B_M1004_g 0.0179723f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_50 VNB N_SET_B_M1002_g 0.0183771f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_51 VNB N_SET_B_c_916_n 0.00782548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_SET_B_c_917_n 0.0247676f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_53 VNB N_SET_B_c_918_n 0.00482639f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_54 VNB SET_B 0.00646661f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_55 VNB N_SET_B_c_920_n 0.013319f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_56 VNB N_SET_B_c_921_n 0.00185354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_SET_B_c_922_n 4.87659e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_923_n 0.00285341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_476_47#_c_1047_n 0.017726f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_60 VNB N_A_476_47#_c_1048_n 0.0138425f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_61 VNB N_A_476_47#_c_1049_n 0.0550461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_476_47#_c_1050_n 0.0177765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_476_47#_c_1051_n 0.00507008f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_64 VNB N_A_476_47#_c_1052_n 0.00430167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_476_47#_c_1053_n 0.00446117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_476_47#_c_1054_n 0.00393532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_476_47#_c_1055_n 0.00107462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_476_47#_c_1056_n 0.0145441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1178_261#_M1033_g 0.0397645f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_70 VNB N_A_1178_261#_c_1205_n 0.00851883f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1178_261#_c_1206_n 0.00717892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1178_261#_c_1207_n 0.00543457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1028_413#_M1013_g 0.0322348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1028_413#_c_1284_n 0.0388051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1028_413#_c_1285_n 0.0124415f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_76 VNB N_A_1028_413#_M1030_g 0.0246021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1028_413#_c_1287_n 0.00547482f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_78 VNB N_A_1028_413#_c_1288_n 0.00490305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1028_413#_c_1289_n 0.0010444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1028_413#_c_1290_n 0.00489285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1028_413#_c_1291_n 8.99453e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1028_413#_c_1292_n 0.00431952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1602_47#_c_1442_n 0.0159483f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_84 VNB N_A_1602_47#_c_1443_n 0.019415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1602_47#_c_1444_n 0.00182991f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_86 VNB N_A_1602_47#_c_1445_n 0.00194757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1602_47#_c_1446_n 0.00279295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1602_47#_c_1447_n 0.0363082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VPWR_c_1517_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_381_47#_c_1688_n 0.00886009f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_91 VNB N_A_381_47#_c_1689_n 0.00231118f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_92 VNB Q 0.0193767f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_93 VNB N_Q_c_1756_n 0.00636192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1787_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_95 VNB N_VGND_c_1788_n 0.00493513f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_96 VNB N_VGND_c_1789_n 0.00404464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1790_n 0.0199361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1791_n 0.00985311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1792_n 4.08532e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1793_n 0.0100799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1794_n 0.0188231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1795_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1796_n 0.0164074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1797_n 0.0451324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1798_n 0.0408311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1799_n 0.0285572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1800_n 0.0152636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1801_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1802_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1803_n 0.0056662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1804_n 0.00612673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1805_n 0.0156869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1806_n 0.00439458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1807_n 0.457663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VPB N_CLK_c_227_n 0.0118979f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_116 VPB N_CLK_c_228_n 0.0184083f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_117 VPB N_CLK_c_229_n 0.0238007f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_118 VPB CLK 0.0152043f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_119 VPB N_CLK_c_225_n 0.0100928f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_120 VPB N_A_27_47#_M1000_g 0.0364881f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_121 VPB N_A_27_47#_M1031_g 0.021588f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_122 VPB N_A_27_47#_M1005_g 0.0202797f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_123 VPB N_A_27_47#_c_284_n 0.00103857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_271_n 0.00335104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_47#_c_272_n 0.00245013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_27_47#_c_274_n 0.00546282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_288_n 0.0299306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_289_n 0.0140517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_290_n 0.00181346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_291_n 0.0108096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_292_n 0.0015212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_293_n 0.00372072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_279_n 0.0117644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_295_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_296_n 0.00564526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_297_n 0.0279259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_298_n 0.00620409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_D_M1023_g 0.0293669f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_139 VPB N_D_c_548_n 0.00538482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_D_c_549_n 0.00459652f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_141 VPB N_A_193_47#_M1011_g 0.0465266f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_142 VPB N_A_193_47#_c_589_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_143 VPB N_A_193_47#_c_590_n 0.00328709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_193_47#_c_594_n 0.0110035f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_145 VPB N_A_193_47#_M1024_g 0.0394871f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_146 VPB N_A_193_47#_c_595_n 0.0125421f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_147 VPB N_A_193_47#_c_614_n 0.00566154f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_148 VPB N_A_193_47#_c_615_n 0.00134324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_193_47#_c_602_n 0.0112434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_193_47#_c_606_n 0.00217264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_652_21#_M1022_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_152 VPB N_A_652_21#_M1009_g 0.0208799f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_153 VPB N_A_652_21#_c_803_n 0.00189033f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_154 VPB N_A_652_21#_c_804_n 0.00247793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_652_21#_c_799_n 0.00270641f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_156 VPB N_A_652_21#_c_806_n 0.00460198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_652_21#_c_807_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_158 VPB N_A_652_21#_c_808_n 0.00112185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_SET_B_M1026_g 0.0474843f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_160 VPB N_SET_B_c_916_n 0.0166983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_SET_B_M1001_g 0.0382157f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_162 VPB N_SET_B_c_927_n 0.00527828f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_163 VPB N_A_476_47#_M1020_g 0.0334449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_476_47#_M1016_g 0.0319093f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_165 VPB N_A_476_47#_c_1059_n 0.0121124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_476_47#_c_1053_n 0.00542515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_476_47#_c_1054_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_476_47#_c_1055_n 0.00262972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_476_47#_c_1056_n 0.0306997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1178_261#_M1015_g 0.0268094f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_171 VPB N_A_1178_261#_c_1205_n 0.0294612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1178_261#_c_1210_n 0.0164657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_1178_261#_c_1211_n 0.0160465f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_174 VPB N_A_1178_261#_c_1206_n 0.00334108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1178_261#_c_1213_n 0.0176565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1178_261#_c_1214_n 0.0110714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1028_413#_M1027_g 0.026322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1028_413#_c_1284_n 0.0284854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1028_413#_c_1285_n 0.00812887f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_180 VPB N_A_1028_413#_c_1296_n 0.0179641f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_181 VPB N_A_1028_413#_c_1287_n 0.00353272f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_182 VPB N_A_1028_413#_c_1298_n 0.00422026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1028_413#_c_1288_n 0.00190145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1028_413#_c_1300_n 0.0149543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1028_413#_c_1301_n 0.0037282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1028_413#_c_1302_n 2.86428e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1028_413#_c_1291_n 4.61735e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1028_413#_c_1292_n 0.00430849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1602_47#_M1025_g 0.0187885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1602_47#_M1032_g 0.022286f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_191 VPB N_A_1602_47#_c_1450_n 5.65061e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1602_47#_c_1445_n 0.00337528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1602_47#_c_1452_n 0.00624721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1602_47#_c_1447_n 0.00706808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1518_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_196 VPB N_VPWR_c_1519_n 0.00580969f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_197 VPB N_VPWR_c_1520_n 0.0114969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1521_n 3.97306e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1522_n 0.00364239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1523_n 0.00411693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1524_n 0.00998201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1525_n 0.0318786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1526_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1527_n 0.0163044f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1528_n 0.0416374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1529_n 0.0307572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1530_n 0.01851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1531_n 0.0306694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1532_n 0.0181025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1533_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1534_n 0.00507833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1535_n 0.0091704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1536_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1537_n 0.011387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1538_n 0.00504924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1539_n 0.00324235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1517_n 0.0641099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_381_47#_c_1688_n 0.00802497f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_219 VPB N_A_381_47#_c_1691_n 0.00187115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB Q 0.00753886f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_221 VPB N_Q_c_1758_n 0.00862547f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_222 N_CLK_c_222_n N_A_27_47#_M1019_g 0.020058f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_223 CLK N_A_27_47#_M1019_g 3.07529e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_224 N_CLK_c_226_n N_A_27_47#_M1019_g 0.00498861f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_225 N_CLK_c_229_n N_A_27_47#_M1000_g 0.028055f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_226 CLK N_A_27_47#_M1000_g 5.68848e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_227 N_CLK_c_225_n N_A_27_47#_M1000_g 0.00521293f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_228 N_CLK_c_222_n N_A_27_47#_c_269_n 0.00695828f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_229 N_CLK_c_223_n N_A_27_47#_c_269_n 0.00799602f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_230 CLK N_A_27_47#_c_269_n 0.00698378f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_231 N_CLK_c_223_n N_A_27_47#_c_270_n 0.00636033f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_232 CLK N_A_27_47#_c_270_n 0.0224397f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_233 N_CLK_c_225_n N_A_27_47#_c_270_n 7.17088e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_234 N_CLK_c_228_n N_A_27_47#_c_284_n 0.0129687f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_235 N_CLK_c_229_n N_A_27_47#_c_284_n 0.0013404f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_236 CLK N_A_27_47#_c_284_n 0.00690269f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_237 N_CLK_c_223_n N_A_27_47#_c_271_n 0.00191059f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_238 N_CLK_c_229_n N_A_27_47#_c_271_n 0.00441254f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_239 CLK N_A_27_47#_c_271_n 0.0517134f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_240 N_CLK_c_225_n N_A_27_47#_c_271_n 0.00100166f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_241 N_CLK_c_226_n N_A_27_47#_c_271_n 0.00247465f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_242 N_CLK_c_228_n N_A_27_47#_c_288_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_243 N_CLK_c_229_n N_A_27_47#_c_288_n 0.00374438f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_244 CLK N_A_27_47#_c_288_n 0.0236151f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_245 N_CLK_c_225_n N_A_27_47#_c_288_n 5.66731e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_246 N_CLK_c_228_n N_A_27_47#_c_290_n 0.00106507f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_247 CLK N_A_27_47#_c_279_n 0.00162145f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_248 N_CLK_c_225_n N_A_27_47#_c_279_n 0.0169859f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_249 N_CLK_c_228_n N_VPWR_c_1518_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_250 N_CLK_c_228_n N_VPWR_c_1526_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_251 N_CLK_c_228_n N_VPWR_c_1517_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_252 N_CLK_c_222_n N_VGND_c_1787_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_253 N_CLK_c_222_n N_VGND_c_1795_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_254 N_CLK_c_223_n N_VGND_c_1795_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_255 N_CLK_c_222_n N_VGND_c_1807_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_267_n N_D_M1010_g 0.0210908f $X=2.305 $Y=0.705 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_272_n N_D_M1010_g 0.00120175f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_296_n N_D_M1023_g 7.92917e-19 $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_272_n N_D_c_548_n 0.00106119f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_273_n N_D_c_548_n 0.00155965f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_272_n N_D_c_549_n 0.0453933f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_273_n N_D_c_549_n 2.37218e-19 $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_289_n N_D_c_549_n 0.00575757f $X=2.385 $Y=1.87 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_296_n N_D_c_549_n 0.00408526f $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_289_n N_A_193_47#_M1000_d 5.39371e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1031_g N_A_193_47#_M1011_g 0.0191849f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_272_n N_A_193_47#_M1011_g 0.0053439f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_289_n N_A_193_47#_M1011_g 0.00702647f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_292_n N_A_193_47#_M1011_g 5.22576e-19 $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_295_n N_A_193_47#_M1011_g 0.0174486f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_296_n N_A_193_47#_M1011_g 0.010416f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_272_n N_A_193_47#_c_589_n 0.0101526f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_291_n N_A_193_47#_c_589_n 3.63007e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_295_n N_A_193_47#_c_589_n 0.0212215f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_296_n N_A_193_47#_c_589_n 0.00655916f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_272_n N_A_193_47#_c_590_n 0.00204176f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_273_n N_A_193_47#_c_590_n 0.0232669f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_267_n N_A_193_47#_M1018_g 0.0128045f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_272_n N_A_193_47#_M1018_g 4.48322e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_273_n N_A_193_47#_M1018_g 0.0214244f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_274_n N_A_193_47#_M1014_g 0.00402103f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_282 N_A_27_47#_c_275_n N_A_193_47#_M1014_g 0.0116603f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_277_n N_A_193_47#_M1014_g 0.00281779f $X=5.975 $Y=0.81 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_278_n N_A_193_47#_M1014_g 0.0209674f $X=5.985 $Y=0.93 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_280_n N_A_193_47#_M1014_g 0.0117187f $X=5.995 $Y=0.765 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1005_g N_A_193_47#_M1024_g 0.0175645f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_274_n N_A_193_47#_M1024_g 0.00215568f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_288 N_A_27_47#_c_293_n N_A_193_47#_M1024_g 0.00434444f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_297_n N_A_193_47#_M1024_g 0.0159766f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_298_n N_A_193_47#_M1024_g 0.00180554f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_274_n N_A_193_47#_c_595_n 0.00355331f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_275_n N_A_193_47#_c_595_n 0.00394592f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_293_n N_A_193_47#_c_595_n 5.11972e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_297_n N_A_193_47#_c_595_n 0.0106615f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_298_n N_A_193_47#_c_595_n 0.00101144f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1000_g N_A_193_47#_c_614_n 2.1943e-19 $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1019_g N_A_193_47#_c_596_n 5.60719e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_269_n N_A_193_47#_c_596_n 0.00285924f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_289_n N_A_193_47#_c_615_n 0.00680899f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_290_n N_A_193_47#_c_615_n 8.29293e-19 $X=0.835 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_279_n N_A_193_47#_c_615_n 0.0133915f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_272_n N_A_193_47#_c_597_n 0.0173405f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_273_n N_A_193_47#_c_597_n 0.0059767f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_M1019_g N_A_193_47#_c_598_n 0.00656242f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_269_n N_A_193_47#_c_598_n 0.00214831f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_271_n N_A_193_47#_c_598_n 0.00506081f $X=0.75 $Y=1.235 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_272_n N_A_193_47#_c_599_n 0.00886175f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_274_n N_A_193_47#_c_600_n 0.0118781f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_275_n N_A_193_47#_c_600_n 0.00159218f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_293_n N_A_193_47#_c_600_n 9.05104e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_297_n N_A_193_47#_c_600_n 8.971e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_298_n N_A_193_47#_c_600_n 0.00270751f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_291_n N_A_193_47#_c_601_n 0.0945834f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1019_g N_A_193_47#_c_602_n 0.0133915f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_269_n N_A_193_47#_c_602_n 0.00935521f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_386_p N_A_193_47#_c_602_n 0.0085177f $X=0.72 $Y=1.795 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_271_n N_A_193_47#_c_602_n 0.0719147f $X=0.75 $Y=1.235 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_289_n N_A_193_47#_c_602_n 0.0182528f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_290_n N_A_193_47#_c_602_n 0.0010354f $X=0.835 $Y=1.87 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_272_n N_A_193_47#_c_603_n 5.02791e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_267_n N_A_193_47#_c_604_n 5.21885e-19 $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_272_n N_A_193_47#_c_604_n 0.0209059f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_273_n N_A_193_47#_c_604_n 0.00155193f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_295_n N_A_193_47#_c_604_n 3.45191e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_296_n N_A_193_47#_c_604_n 0.00332918f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_274_n N_A_193_47#_c_605_n 0.00256294f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_275_n N_A_193_47#_c_605_n 0.0014885f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_293_n N_A_193_47#_c_605_n 0.0132733f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_298_n N_A_193_47#_c_605_n 0.00178603f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_274_n N_A_193_47#_c_606_n 0.0285015f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_275_n N_A_193_47#_c_606_n 0.0123304f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_293_n N_A_193_47#_c_606_n 6.9568e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_297_n N_A_193_47#_c_606_n 6.19272e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_298_n N_A_193_47#_c_606_n 0.0119993f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_272_n N_A_193_47#_c_607_n 0.00673428f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_272_n N_A_652_21#_M1022_g 5.35023e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_291_n N_A_652_21#_M1009_g 0.00197541f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_291_n N_A_652_21#_c_803_n 0.0147195f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_M1005_g N_A_652_21#_c_804_n 6.75516e-19 $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_291_n N_A_652_21#_c_804_n 0.021867f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_293_n N_A_652_21#_c_804_n 9.32161e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_298_n N_A_652_21#_c_804_n 0.0093814f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_274_n N_A_652_21#_c_799_n 0.041895f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_291_n N_A_652_21#_c_799_n 0.00686718f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_297_n N_A_652_21#_c_799_n 2.22171e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_298_n N_A_652_21#_c_799_n 0.0136142f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_291_n N_A_652_21#_c_806_n 0.0157473f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_M1031_g N_A_652_21#_c_807_n 0.0161874f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_291_n N_A_652_21#_c_807_n 0.00193898f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_295_n N_A_652_21#_c_807_n 0.00927772f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_291_n N_A_652_21#_c_808_n 0.00782494f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_274_n N_A_652_21#_c_800_n 0.0132853f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_276_n N_A_652_21#_c_800_n 0.0121054f $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_291_n N_SET_B_M1026_g 0.00205491f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_274_n N_SET_B_c_920_n 0.00399047f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_275_n N_SET_B_c_920_n 0.0294013f $X=5.8 $Y=0.81 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_276_n N_SET_B_c_920_n 0.00574094f $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_277_n N_SET_B_c_920_n 0.0175891f $X=5.975 $Y=0.81 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_274_n N_A_476_47#_c_1048_n 2.94773e-19 $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_291_n N_A_476_47#_M1020_g 0.00187886f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_274_n N_A_476_47#_c_1049_n 0.00469727f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_275_n N_A_476_47#_c_1049_n 0.0078216f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_276_n N_A_476_47#_c_1049_n 0.00630303f $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_297_n N_A_476_47#_c_1049_n 0.00228498f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_291_n N_A_476_47#_M1016_g 0.00301713f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_297_n N_A_476_47#_M1016_g 0.0626672f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_298_n N_A_476_47#_M1016_g 0.00172662f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_275_n N_A_476_47#_c_1050_n 0.00414107f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_M1031_g N_A_476_47#_c_1074_n 0.0090453f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_291_n N_A_476_47#_c_1074_n 0.00517144f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_292_n N_A_476_47#_c_1074_n 0.00306479f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_295_n N_A_476_47#_c_1074_n 0.00186639f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_296_n N_A_476_47#_c_1074_n 0.015267f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_272_n N_A_476_47#_c_1079_n 0.00676006f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_273_n N_A_476_47#_c_1079_n 9.25786e-19 $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_M1031_g N_A_476_47#_c_1059_n 0.00650943f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_272_n N_A_476_47#_c_1059_n 0.00666284f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_291_n N_A_476_47#_c_1059_n 0.013911f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_292_n N_A_476_47#_c_1059_n 0.00145075f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_295_n N_A_476_47#_c_1059_n 0.00203066f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_296_n N_A_476_47#_c_1059_n 0.0283088f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_291_n N_A_476_47#_c_1053_n 0.00472657f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_272_n N_A_476_47#_c_1054_n 0.007273f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_291_n N_A_476_47#_c_1054_n 0.00456576f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_c_291_n N_A_476_47#_c_1055_n 0.00248872f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_274_n N_A_476_47#_c_1056_n 0.00640057f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_291_n N_A_476_47#_c_1056_n 0.00148193f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_277_n N_A_1178_261#_M1033_g 8.03923e-19 $X=5.975 $Y=0.81
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_280_n N_A_1178_261#_M1033_g 0.0627625f $X=5.995 $Y=0.765
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_277_n N_A_1178_261#_c_1205_n 2.97133e-19 $X=5.975 $Y=0.81
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_278_n N_A_1178_261#_c_1205_n 0.0161765f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_M1005_g N_A_1028_413#_c_1305_n 0.00493733f $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_293_n N_A_1028_413#_c_1305_n 0.00403604f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_297_n N_A_1028_413#_c_1305_n 9.00165e-19 $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_298_n N_A_1028_413#_c_1305_n 0.0148431f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_274_n N_A_1028_413#_c_1298_n 0.00537793f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_293_n N_A_1028_413#_c_1298_n 0.00776519f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_297_n N_A_1028_413#_c_1298_n 4.1977e-19 $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_298_n N_A_1028_413#_c_1298_n 0.0211547f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_275_n N_A_1028_413#_c_1313_n 0.0059175f $X=5.8 $Y=0.81 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_277_n N_A_1028_413#_c_1313_n 0.0140112f $X=5.975 $Y=0.81
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_278_n N_A_1028_413#_c_1313_n 6.91335e-19 $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_280_n N_A_1028_413#_c_1313_n 0.00790984f $X=5.995 $Y=0.765
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_275_n N_A_1028_413#_c_1288_n 0.00194166f $X=5.8 $Y=0.81
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_277_n N_A_1028_413#_c_1288_n 0.0194146f $X=5.975 $Y=0.81
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_278_n N_A_1028_413#_c_1288_n 0.00260024f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_275_n N_A_1028_413#_c_1289_n 0.00570635f $X=5.8 $Y=0.81
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_277_n N_A_1028_413#_c_1290_n 0.0219337f $X=5.975 $Y=0.81
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_278_n N_A_1028_413#_c_1290_n 0.00160679f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_280_n N_A_1028_413#_c_1290_n 0.00257842f $X=5.995 $Y=0.765
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_M1005_g N_A_1028_413#_c_1302_n 0.0010081f $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_386_p N_VPWR_M1017_d 7.14517e-19 $X=0.72 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_413 N_A_27_47#_c_290_n N_VPWR_M1017_d 0.00181761f $X=0.835 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_414 N_A_27_47#_M1000_g N_VPWR_c_1518_n 0.00837918f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_284_n N_VPWR_c_1518_n 0.00328949f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_386_p N_VPWR_c_1518_n 0.0133733f $X=0.72 $Y=1.795 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_288_n N_VPWR_c_1518_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_418 N_A_27_47#_c_289_n N_VPWR_c_1518_n 2.78216e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_290_n N_VPWR_c_1518_n 0.00348405f $X=0.835 $Y=1.87 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1000_g N_VPWR_c_1519_n 0.00191658f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_289_n N_VPWR_c_1519_n 0.00166908f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1005_g N_VPWR_c_1521_n 0.0019199f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_291_n N_VPWR_c_1521_n 0.001212f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_424 N_A_27_47#_c_284_n N_VPWR_c_1526_n 0.0018545f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_288_n N_VPWR_c_1526_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_426 N_A_27_47#_M1000_g N_VPWR_c_1527_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_M1031_g N_VPWR_c_1528_n 0.00367119f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_M1005_g N_VPWR_c_1529_n 0.00427125f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_298_n N_VPWR_c_1529_n 0.0032218f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_291_n N_VPWR_c_1535_n 0.0014214f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_M1000_g N_VPWR_c_1517_n 0.00536257f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1031_g N_VPWR_c_1517_n 0.00563088f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_M1005_g N_VPWR_c_1517_n 0.00577339f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_284_n N_VPWR_c_1517_n 0.00394611f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_288_n N_VPWR_c_1517_n 0.00993215f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_289_n N_VPWR_c_1517_n 0.0726622f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_290_n N_VPWR_c_1517_n 0.01448f $X=0.835 $Y=1.87 $X2=0 $Y2=0
cc_438 N_A_27_47#_c_291_n N_VPWR_c_1517_n 0.111929f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_439 N_A_27_47#_c_292_n N_VPWR_c_1517_n 0.0160044f $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_c_293_n N_VPWR_c_1517_n 0.016077f $X=5.29 $Y=1.87 $X2=0 $Y2=0
cc_441 N_A_27_47#_c_296_n N_VPWR_c_1517_n 2.46058e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_298_n N_VPWR_c_1517_n 0.00246615f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_289_n N_A_381_47#_M1023_d 8.84929e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_267_n N_A_381_47#_c_1693_n 0.00223782f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_272_n N_A_381_47#_c_1693_n 0.00713576f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_289_n N_A_381_47#_c_1695_n 0.019313f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_289_n N_A_381_47#_c_1691_n 0.015767f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_267_n N_A_381_47#_c_1697_n 0.00399753f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_449 N_A_27_47#_c_289_n N_A_381_47#_c_1698_n 0.0109514f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_292_n N_A_381_47#_c_1698_n 0.00146426f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_451 N_A_27_47#_c_296_n N_A_381_47#_c_1698_n 0.00827001f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_269_n N_VGND_M1029_d 0.00162876f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_453 N_A_27_47#_M1019_g N_VGND_c_1787_n 0.00826572f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_269_n N_VGND_c_1787_n 0.0165953f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_279_n N_VGND_c_1787_n 5.88506e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_M1019_g N_VGND_c_1788_n 0.00296886f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_267_n N_VGND_c_1788_n 0.00120909f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_275_n N_VGND_c_1791_n 0.0017326f $X=5.8 $Y=0.81 $X2=0 $Y2=0
cc_459 N_A_27_47#_c_276_n N_VGND_c_1791_n 0.0129707f $X=5.05 $Y=0.81 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_268_n N_VGND_c_1795_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_269_n N_VGND_c_1795_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_M1019_g N_VGND_c_1796_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_267_n N_VGND_c_1797_n 0.00556304f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_272_n N_VGND_c_1797_n 0.00113905f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_273_n N_VGND_c_1797_n 2.48118e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_275_n N_VGND_c_1798_n 0.00797153f $X=5.8 $Y=0.81 $X2=0 $Y2=0
cc_467 N_A_27_47#_c_280_n N_VGND_c_1798_n 0.00368123f $X=5.995 $Y=0.765 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_M1029_s N_VGND_c_1807_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1019_g N_VGND_c_1807_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_267_n N_VGND_c_1807_n 0.00678262f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_268_n N_VGND_c_1807_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_269_n N_VGND_c_1807_n 0.0057651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_272_n N_VGND_c_1807_n 0.00122477f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_275_n N_VGND_c_1807_n 0.00610816f $X=5.8 $Y=0.81 $X2=0 $Y2=0
cc_475 N_A_27_47#_c_276_n N_VGND_c_1807_n 4.92512e-19 $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_280_n N_VGND_c_1807_n 0.00526484f $X=5.995 $Y=0.765 $X2=0
+ $Y2=0
cc_477 N_D_M1023_g N_A_193_47#_c_590_n 0.0303627f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_478 N_D_c_548_n N_A_193_47#_c_590_n 0.00467503f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_479 N_D_c_549_n N_A_193_47#_c_590_n 0.00330794f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_480 N_D_M1023_g N_A_193_47#_c_614_n 6.25863e-19 $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_481 N_D_M1010_g N_A_193_47#_c_596_n 0.00306188f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_482 N_D_M1023_g N_A_193_47#_c_615_n 0.00288262f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_483 N_D_M1010_g N_A_193_47#_c_597_n 0.00395556f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_484 N_D_c_548_n N_A_193_47#_c_597_n 8.88354e-19 $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_485 N_D_c_549_n N_A_193_47#_c_597_n 0.0127149f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_486 N_D_M1010_g N_A_193_47#_c_602_n 6.53696e-19 $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_487 N_D_M1023_g N_A_193_47#_c_602_n 0.00119126f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_488 N_D_M1023_g N_VPWR_c_1519_n 0.0116766f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_489 N_D_M1023_g N_VPWR_c_1528_n 0.0035268f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_490 N_D_M1023_g N_VPWR_c_1517_n 0.00402871f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_491 N_D_M1010_g N_A_381_47#_c_1688_n 0.00557005f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_492 N_D_M1023_g N_A_381_47#_c_1688_n 0.0115166f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_493 N_D_c_548_n N_A_381_47#_c_1688_n 0.00753248f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_494 N_D_c_549_n N_A_381_47#_c_1688_n 0.0473419f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_495 N_D_M1010_g N_A_381_47#_c_1693_n 0.0126635f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_496 N_D_c_548_n N_A_381_47#_c_1693_n 0.0014463f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_497 N_D_c_549_n N_A_381_47#_c_1693_n 0.0217898f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_498 N_D_M1023_g N_A_381_47#_c_1695_n 0.011823f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_499 N_D_c_549_n N_A_381_47#_c_1695_n 0.0109323f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_500 N_D_c_549_n N_A_381_47#_c_1698_n 0.0137404f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_501 N_D_M1010_g N_VGND_c_1788_n 0.00942273f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_502 N_D_M1010_g N_VGND_c_1797_n 0.00339367f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_503 N_D_M1010_g N_VGND_c_1807_n 0.00393034f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_504 N_A_193_47#_M1018_g N_A_652_21#_M1022_g 0.024565f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_505 N_A_193_47#_c_592_n N_A_652_21#_M1022_g 0.0114519f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_506 N_A_193_47#_c_600_n N_A_652_21#_M1022_g 9.99732e-19 $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_507 N_A_193_47#_c_603_n N_A_652_21#_M1022_g 0.00631121f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_508 N_A_193_47#_c_604_n N_A_652_21#_M1022_g 0.00191013f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_509 N_A_193_47#_c_607_n N_A_652_21#_M1022_g 0.0200607f $X=2.915 $Y=0.93 $X2=0
+ $Y2=0
cc_510 N_A_193_47#_c_600_n N_A_652_21#_c_803_n 5.47854e-19 $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_511 N_A_193_47#_c_600_n N_A_652_21#_c_804_n 0.00115455f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_512 N_A_193_47#_c_600_n N_A_652_21#_c_799_n 0.0140676f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_513 N_A_193_47#_c_600_n N_A_652_21#_c_806_n 8.37667e-19 $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_514 N_A_193_47#_c_600_n N_A_652_21#_c_800_n 0.00655125f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_515 N_A_193_47#_c_600_n N_SET_B_c_912_n 0.00381498f $X=5.165 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_516 N_A_193_47#_c_600_n N_SET_B_M1026_g 0.00121673f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_517 N_A_193_47#_c_600_n SET_B 0.00570533f $X=5.165 $Y=1.19 $X2=0 $Y2=0
cc_518 N_A_193_47#_M1014_g N_SET_B_c_920_n 0.00419104f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_519 N_A_193_47#_c_595_n N_SET_B_c_920_n 0.00120258f $X=5.47 $Y=1.26 $X2=0
+ $Y2=0
cc_520 N_A_193_47#_c_600_n N_SET_B_c_920_n 0.0878381f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_521 N_A_193_47#_c_605_n N_SET_B_c_920_n 0.02693f $X=5.31 $Y=1.19 $X2=0 $Y2=0
cc_522 N_A_193_47#_c_606_n N_SET_B_c_920_n 0.00112669f $X=5.31 $Y=1.19 $X2=0
+ $Y2=0
cc_523 N_A_193_47#_c_600_n N_SET_B_c_921_n 0.0263312f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_524 N_A_193_47#_c_600_n N_A_476_47#_c_1048_n 0.00253485f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_525 N_A_193_47#_c_595_n N_A_476_47#_c_1049_n 0.00912806f $X=5.47 $Y=1.26
+ $X2=0 $Y2=0
cc_526 N_A_193_47#_c_600_n N_A_476_47#_c_1049_n 0.00101093f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_527 N_A_193_47#_c_606_n N_A_476_47#_c_1049_n 3.19592e-19 $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_528 N_A_193_47#_M1014_g N_A_476_47#_c_1050_n 0.0518139f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_529 N_A_193_47#_M1011_g N_A_476_47#_c_1074_n 0.00278769f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_530 N_A_193_47#_M1018_g N_A_476_47#_c_1079_n 0.008828f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_531 N_A_193_47#_c_597_n N_A_476_47#_c_1079_n 0.00573977f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_532 N_A_193_47#_c_603_n N_A_476_47#_c_1079_n 0.00194059f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_533 N_A_193_47#_c_604_n N_A_476_47#_c_1079_n 0.0194974f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_534 N_A_193_47#_c_607_n N_A_476_47#_c_1079_n 5.24271e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_535 N_A_193_47#_M1011_g N_A_476_47#_c_1059_n 8.73767e-19 $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_536 N_A_193_47#_c_601_n N_A_476_47#_c_1059_n 3.07745e-19 $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_M1018_g N_A_476_47#_c_1052_n 0.00118778f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_538 N_A_193_47#_c_592_n N_A_476_47#_c_1052_n 7.74259e-19 $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_539 N_A_193_47#_c_600_n N_A_476_47#_c_1052_n 0.0146154f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_540 N_A_193_47#_c_603_n N_A_476_47#_c_1052_n 0.0134967f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_541 N_A_193_47#_c_604_n N_A_476_47#_c_1052_n 0.0244992f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_542 N_A_193_47#_c_607_n N_A_476_47#_c_1052_n 7.73887e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_c_600_n N_A_476_47#_c_1053_n 0.0232188f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_544 N_A_193_47#_c_592_n N_A_476_47#_c_1054_n 0.00262762f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_600_n N_A_476_47#_c_1054_n 0.0121342f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_601_n N_A_476_47#_c_1054_n 0.00535278f $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_c_604_n N_A_476_47#_c_1054_n 0.00527199f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_c_607_n N_A_476_47#_c_1054_n 5.70501e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_600_n N_A_476_47#_c_1055_n 0.00996075f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_550 N_A_193_47#_c_594_n N_A_476_47#_c_1056_n 5.76045e-19 $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_551 N_A_193_47#_c_595_n N_A_476_47#_c_1056_n 0.00482213f $X=5.47 $Y=1.26
+ $X2=0 $Y2=0
cc_552 N_A_193_47#_c_600_n N_A_476_47#_c_1056_n 0.00412912f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_553 N_A_193_47#_M1014_g N_A_1178_261#_M1033_g 0.00229504f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_554 N_A_193_47#_c_594_n N_A_1178_261#_c_1205_n 0.0407174f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_555 N_A_193_47#_M1024_g N_A_1178_261#_c_1210_n 0.0407174f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_556 N_A_193_47#_M1024_g N_A_1028_413#_c_1305_n 0.00768489f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_557 N_A_193_47#_c_594_n N_A_1028_413#_c_1298_n 0.00103911f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_558 N_A_193_47#_M1024_g N_A_1028_413#_c_1298_n 0.0101662f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_559 N_A_193_47#_c_606_n N_A_1028_413#_c_1298_n 0.00496139f $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_560 N_A_193_47#_c_594_n N_A_1028_413#_c_1289_n 0.00829662f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_561 N_A_193_47#_c_605_n N_A_1028_413#_c_1289_n 0.00200974f $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_562 N_A_193_47#_c_606_n N_A_1028_413#_c_1289_n 0.0123133f $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_563 N_A_193_47#_M1024_g N_A_1028_413#_c_1300_n 2.49577e-19 $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_564 N_A_193_47#_M1014_g N_A_1028_413#_c_1290_n 0.00204758f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_565 N_A_193_47#_M1024_g N_A_1028_413#_c_1302_n 0.011666f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_566 N_A_193_47#_c_614_n N_VPWR_c_1518_n 0.0127345f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_567 N_A_193_47#_M1011_g N_VPWR_c_1519_n 0.00113058f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_568 N_A_193_47#_c_614_n N_VPWR_c_1519_n 0.0222599f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_569 N_A_193_47#_c_614_n N_VPWR_c_1527_n 0.0156296f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_570 N_A_193_47#_M1011_g N_VPWR_c_1528_n 0.00541732f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_571 N_A_193_47#_M1024_g N_VPWR_c_1529_n 0.00369426f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_572 N_A_193_47#_M1024_g N_VPWR_c_1537_n 0.00197636f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_573 N_A_193_47#_M1011_g N_VPWR_c_1517_n 0.00628966f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_574 N_A_193_47#_M1024_g N_VPWR_c_1517_n 0.00544628f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_575 N_A_193_47#_c_614_n N_VPWR_c_1517_n 0.00399922f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_576 N_A_193_47#_c_597_n N_A_381_47#_M1010_d 4.25819e-19 $X=2.845 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_577 N_A_193_47#_c_597_n N_A_381_47#_c_1688_n 0.0148575f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_578 N_A_193_47#_c_598_n N_A_381_47#_c_1688_n 0.0013578f $X=1.295 $Y=0.85
+ $X2=0 $Y2=0
cc_579 N_A_193_47#_c_602_n N_A_381_47#_c_1688_n 0.0663617f $X=1.15 $Y=0.85 $X2=0
+ $Y2=0
cc_580 N_A_193_47#_c_597_n N_A_381_47#_c_1693_n 0.0198802f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_581 N_A_193_47#_c_604_n N_A_381_47#_c_1693_n 0.00201969f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_582 N_A_193_47#_c_596_n N_A_381_47#_c_1689_n 0.00354307f $X=1.12 $Y=0.68
+ $X2=0 $Y2=0
cc_583 N_A_193_47#_c_597_n N_A_381_47#_c_1689_n 0.00436942f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_584 N_A_193_47#_c_598_n N_A_381_47#_c_1689_n 0.00140924f $X=1.295 $Y=0.85
+ $X2=0 $Y2=0
cc_585 N_A_193_47#_c_602_n N_A_381_47#_c_1689_n 0.00998611f $X=1.15 $Y=0.85
+ $X2=0 $Y2=0
cc_586 N_A_193_47#_c_602_n N_A_381_47#_c_1691_n 0.0111323f $X=1.15 $Y=0.85 $X2=0
+ $Y2=0
cc_587 N_A_193_47#_M1011_g N_A_381_47#_c_1698_n 0.0102511f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_588 N_A_193_47#_c_596_n N_VGND_c_1788_n 0.00812552f $X=1.12 $Y=0.68 $X2=0
+ $Y2=0
cc_589 N_A_193_47#_c_597_n N_VGND_c_1788_n 0.0012296f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_590 N_A_193_47#_c_596_n N_VGND_c_1796_n 0.00962729f $X=1.12 $Y=0.68 $X2=0
+ $Y2=0
cc_591 N_A_193_47#_M1018_g N_VGND_c_1797_n 0.00359964f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_592 N_A_193_47#_M1014_g N_VGND_c_1798_n 0.00437852f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_593 N_A_193_47#_M1019_d N_VGND_c_1807_n 0.00318434f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_594 N_A_193_47#_M1018_g N_VGND_c_1807_n 0.0056346f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_595 N_A_193_47#_M1014_g N_VGND_c_1807_n 0.00575719f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_596 N_A_193_47#_c_596_n N_VGND_c_1807_n 0.00381167f $X=1.12 $Y=0.68 $X2=0
+ $Y2=0
cc_597 N_A_193_47#_c_597_n N_VGND_c_1807_n 0.072327f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_598 N_A_193_47#_c_598_n N_VGND_c_1807_n 0.015082f $X=1.295 $Y=0.85 $X2=0
+ $Y2=0
cc_599 N_A_193_47#_c_603_n N_VGND_c_1807_n 0.0151785f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_600 N_A_193_47#_c_604_n A_586_47# 0.00109469f $X=2.99 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_601 N_A_652_21#_M1022_g N_SET_B_c_912_n 0.0189903f $X=3.335 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_602 N_A_652_21#_c_799_n N_SET_B_c_912_n 7.60504e-19 $X=4.625 $Y=1.835
+ $X2=-0.19 $Y2=-0.24
cc_603 N_A_652_21#_M1022_g N_SET_B_M1026_g 0.0137896f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_604 N_A_652_21#_M1009_g N_SET_B_M1026_g 0.0113783f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_605 N_A_652_21#_c_803_n N_SET_B_M1026_g 0.0139954f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_606 N_A_652_21#_c_806_n N_SET_B_M1026_g 0.00563707f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_607 N_A_652_21#_c_807_n N_SET_B_M1026_g 0.0201938f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_608 N_A_652_21#_M1022_g N_SET_B_M1004_g 0.0141659f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_609 N_A_652_21#_c_798_n N_SET_B_M1004_g 0.00124922f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_610 N_A_652_21#_c_800_n N_SET_B_M1004_g 3.79232e-19 $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_611 N_A_652_21#_M1022_g SET_B 0.00110794f $X=3.335 $Y=0.445 $X2=0 $Y2=0
cc_612 N_A_652_21#_c_800_n SET_B 0.0144281f $X=4.625 $Y=0.895 $X2=0 $Y2=0
cc_613 N_A_652_21#_c_798_n N_SET_B_c_920_n 9.52814e-19 $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_614 N_A_652_21#_c_800_n N_SET_B_c_920_n 0.0196649f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_615 N_A_652_21#_c_800_n N_SET_B_c_921_n 0.00250762f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_616 N_A_652_21#_c_798_n N_A_476_47#_c_1047_n 0.00809901f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_617 N_A_652_21#_c_800_n N_A_476_47#_c_1047_n 4.65467e-19 $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_618 N_A_652_21#_c_799_n N_A_476_47#_c_1048_n 0.00246574f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_619 N_A_652_21#_c_800_n N_A_476_47#_c_1048_n 0.0035345f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_620 N_A_652_21#_c_804_n N_A_476_47#_M1020_g 0.0138123f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_621 N_A_652_21#_c_799_n N_A_476_47#_M1020_g 0.00531645f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_622 N_A_652_21#_c_798_n N_A_476_47#_c_1049_n 0.00253676f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_623 N_A_652_21#_c_799_n N_A_476_47#_c_1049_n 2.06235e-19 $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_624 N_A_652_21#_c_800_n N_A_476_47#_c_1049_n 0.0148491f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_625 N_A_652_21#_c_804_n N_A_476_47#_M1016_g 0.00844681f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_626 N_A_652_21#_c_799_n N_A_476_47#_M1016_g 0.00507438f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_627 N_A_652_21#_c_798_n N_A_476_47#_c_1050_n 0.0042575f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_628 N_A_652_21#_c_800_n N_A_476_47#_c_1051_n 0.00182302f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_629 N_A_652_21#_M1009_g N_A_476_47#_c_1074_n 0.00202046f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_630 N_A_652_21#_M1022_g N_A_476_47#_c_1079_n 0.00854236f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_631 N_A_652_21#_M1022_g N_A_476_47#_c_1059_n 0.015293f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_632 N_A_652_21#_c_806_n N_A_476_47#_c_1059_n 0.0366983f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_633 N_A_652_21#_M1022_g N_A_476_47#_c_1052_n 0.0188229f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_634 N_A_652_21#_c_803_n N_A_476_47#_c_1053_n 0.00881126f $X=3.99 $Y=1.96
+ $X2=0 $Y2=0
cc_635 N_A_652_21#_c_808_n N_A_476_47#_c_1053_n 0.00337624f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_636 N_A_652_21#_M1022_g N_A_476_47#_c_1054_n 0.0109017f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_637 N_A_652_21#_c_806_n N_A_476_47#_c_1054_n 0.0171213f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_638 N_A_652_21#_c_807_n N_A_476_47#_c_1054_n 0.0011995f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_639 N_A_652_21#_c_804_n N_A_476_47#_c_1055_n 0.0079382f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_640 N_A_652_21#_c_799_n N_A_476_47#_c_1055_n 0.0229291f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_641 N_A_652_21#_c_808_n N_A_476_47#_c_1055_n 0.00169427f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_642 N_A_652_21#_c_800_n N_A_476_47#_c_1055_n 0.0037745f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_643 N_A_652_21#_c_804_n N_A_476_47#_c_1056_n 0.0029883f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_644 N_A_652_21#_c_799_n N_A_476_47#_c_1056_n 0.0130643f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_645 N_A_652_21#_c_800_n N_A_476_47#_c_1056_n 0.00437877f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_646 N_A_652_21#_c_803_n N_VPWR_M1009_d 0.00131929f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_647 N_A_652_21#_c_806_n N_VPWR_M1009_d 0.00154452f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_648 N_A_652_21#_c_804_n N_VPWR_M1020_d 0.00161389f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_649 N_A_652_21#_c_803_n N_VPWR_c_1520_n 0.00266175f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_650 N_A_652_21#_c_887_p N_VPWR_c_1520_n 0.0070924f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_651 N_A_652_21#_c_804_n N_VPWR_c_1520_n 0.00248431f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_652 N_A_652_21#_c_804_n N_VPWR_c_1521_n 0.0155298f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_653 N_A_652_21#_M1009_g N_VPWR_c_1528_n 0.00532975f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_654 N_A_652_21#_c_806_n N_VPWR_c_1528_n 0.00105935f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_655 N_A_652_21#_c_804_n N_VPWR_c_1529_n 8.80252e-19 $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_656 N_A_652_21#_M1009_g N_VPWR_c_1535_n 0.00326498f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_657 N_A_652_21#_c_803_n N_VPWR_c_1535_n 0.0101842f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_658 N_A_652_21#_c_806_n N_VPWR_c_1535_n 0.0109284f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_659 N_A_652_21#_c_807_n N_VPWR_c_1535_n 6.81742e-19 $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_660 N_A_652_21#_M1026_d N_VPWR_c_1517_n 0.00202389f $X=3.94 $Y=2.065 $X2=0
+ $Y2=0
cc_661 N_A_652_21#_M1009_g N_VPWR_c_1517_n 0.0066225f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_662 N_A_652_21#_c_803_n N_VPWR_c_1517_n 0.00255051f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_663 N_A_652_21#_c_887_p N_VPWR_c_1517_n 0.00288476f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_664 N_A_652_21#_c_804_n N_VPWR_c_1517_n 0.0034475f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_665 N_A_652_21#_c_806_n N_VPWR_c_1517_n 0.00138626f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_666 N_A_652_21#_M1022_g N_VGND_c_1789_n 0.0040279f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_667 N_A_652_21#_c_798_n N_VGND_c_1790_n 0.0118981f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_668 N_A_652_21#_c_800_n N_VGND_c_1790_n 0.00244068f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_669 N_A_652_21#_c_798_n N_VGND_c_1791_n 0.0177704f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_670 N_A_652_21#_M1022_g N_VGND_c_1797_n 0.0035977f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_671 N_A_652_21#_M1007_d N_VGND_c_1807_n 0.00186029f $X=4.34 $Y=0.235 $X2=0
+ $Y2=0
cc_672 N_A_652_21#_M1022_g N_VGND_c_1807_n 0.00580574f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_673 N_A_652_21#_c_798_n N_VGND_c_1807_n 0.00426169f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_674 N_A_652_21#_c_800_n N_VGND_c_1807_n 0.00183644f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_675 N_SET_B_M1004_g N_A_476_47#_c_1047_n 0.0270653f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_912_n N_A_476_47#_c_1048_n 0.0146844f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_920_n N_A_476_47#_c_1048_n 8.12862e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_921_n N_A_476_47#_c_1048_n 7.28461e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_679 N_SET_B_M1026_g N_A_476_47#_M1020_g 0.0336841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_680 N_SET_B_c_920_n N_A_476_47#_c_1049_n 0.00253697f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_912_n N_A_476_47#_c_1051_n 0.0270653f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_682 SET_B N_A_476_47#_c_1051_n 0.0021684f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_683 N_SET_B_c_920_n N_A_476_47#_c_1051_n 0.00277782f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_921_n N_A_476_47#_c_1051_n 7.28461e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_912_n N_A_476_47#_c_1052_n 0.00218199f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_686 N_SET_B_M1026_g N_A_476_47#_c_1052_n 6.04572e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_687 N_SET_B_M1004_g N_A_476_47#_c_1052_n 0.00184201f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_688 SET_B N_A_476_47#_c_1052_n 0.0243988f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_689 N_SET_B_c_921_n N_A_476_47#_c_1052_n 0.00116251f $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_912_n N_A_476_47#_c_1053_n 0.00307815f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_691 N_SET_B_M1026_g N_A_476_47#_c_1053_n 0.0103672f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_692 SET_B N_A_476_47#_c_1053_n 0.0263655f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_693 N_SET_B_c_920_n N_A_476_47#_c_1053_n 3.66303e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_921_n N_A_476_47#_c_1053_n 5.23607e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_695 N_SET_B_M1026_g N_A_476_47#_c_1054_n 5.20457e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_696 N_SET_B_M1026_g N_A_476_47#_c_1055_n 0.00354841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_920_n N_A_476_47#_c_1055_n 0.00236582f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_698 N_SET_B_M1026_g N_A_476_47#_c_1056_n 0.0205296f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_699 N_SET_B_M1002_g N_A_1178_261#_M1033_g 0.0639772f $X=6.785 $Y=0.445 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_916_n N_A_1178_261#_M1033_g 0.0127642f $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_918_n N_A_1178_261#_M1033_g 0.00163506f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_920_n N_A_1178_261#_M1033_g 9.67282e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_703 N_SET_B_M1001_g N_A_1178_261#_c_1210_n 0.00284189f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_704 N_SET_B_c_927_n N_A_1178_261#_c_1210_n 0.0023606f $X=6.895 $Y=1.685 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_916_n N_A_1178_261#_c_1211_n 0.0023606f $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_922_n N_A_1178_261#_c_1206_n 0.00140313f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_923_n N_A_1178_261#_c_1206_n 0.0108155f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_916_n N_A_1178_261#_c_1213_n 0.00344372f $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_709 N_SET_B_M1001_g N_A_1178_261#_c_1213_n 0.00935477f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_710 N_SET_B_c_927_n N_A_1178_261#_c_1213_n 0.00443217f $X=6.895 $Y=1.685
+ $X2=0 $Y2=0
cc_711 N_SET_B_c_916_n N_A_1028_413#_M1027_g 0.031627f $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_712 N_SET_B_M1002_g N_A_1028_413#_M1013_g 0.0159181f $X=6.785 $Y=0.445 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_917_n N_A_1028_413#_M1013_g 0.00955494f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_918_n N_A_1028_413#_M1013_g 0.00121343f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_923_n N_A_1028_413#_M1013_g 0.00822182f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_917_n N_A_1028_413#_c_1285_n 0.0221954f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_923_n N_A_1028_413#_c_1285_n 0.0035987f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_718 N_SET_B_M1002_g N_A_1028_413#_c_1313_n 2.03126e-19 $X=6.785 $Y=0.445
+ $X2=0 $Y2=0
cc_719 N_SET_B_c_920_n N_A_1028_413#_c_1313_n 0.00655731f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_920_n N_A_1028_413#_c_1288_n 0.0102663f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_721 N_SET_B_c_920_n N_A_1028_413#_c_1289_n 0.00391758f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_722 N_SET_B_M1001_g N_A_1028_413#_c_1300_n 0.00433068f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_723 N_SET_B_M1002_g N_A_1028_413#_c_1290_n 0.00166893f $X=6.785 $Y=0.445
+ $X2=0 $Y2=0
cc_724 N_SET_B_c_916_n N_A_1028_413#_c_1290_n 4.23658e-19 $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_917_n N_A_1028_413#_c_1290_n 5.59208e-19 $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_918_n N_A_1028_413#_c_1290_n 0.0244533f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_727 N_SET_B_c_920_n N_A_1028_413#_c_1290_n 0.0174654f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_922_n N_A_1028_413#_c_1290_n 3.0985e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_916_n N_A_1028_413#_c_1291_n 6.54137e-19 $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_730 N_SET_B_c_922_n N_A_1028_413#_c_1291_n 9.06304e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_923_n N_A_1028_413#_c_1291_n 0.0144638f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_916_n N_A_1028_413#_c_1292_n 0.0109426f $X=6.895 $Y=1.6 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_917_n N_A_1028_413#_c_1292_n 0.00289453f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_734 N_SET_B_c_918_n N_A_1028_413#_c_1292_n 0.0243347f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_920_n N_A_1028_413#_c_1292_n 0.00830763f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_SET_B_c_922_n N_A_1028_413#_c_1292_n 0.00100931f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_737 N_SET_B_c_923_n N_A_1028_413#_c_1292_n 0.00719073f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_738 N_SET_B_M1026_g N_VPWR_c_1520_n 0.00368415f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_739 N_SET_B_M1026_g N_VPWR_c_1521_n 7.26951e-19 $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_740 N_SET_B_M1001_g N_VPWR_c_1522_n 0.00325743f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_741 N_SET_B_M1001_g N_VPWR_c_1530_n 0.00585385f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_742 N_SET_B_M1026_g N_VPWR_c_1535_n 0.00699603f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_743 N_SET_B_M1001_g N_VPWR_c_1537_n 0.00306764f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_744 N_SET_B_M1026_g N_VPWR_c_1517_n 0.00406312f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_745 N_SET_B_M1001_g N_VPWR_c_1517_n 0.0121782f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_746 N_SET_B_c_922_n N_VGND_M1002_d 0.00131987f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_747 N_SET_B_c_923_n N_VGND_M1002_d 9.1061e-19 $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_748 N_SET_B_c_912_n N_VGND_c_1789_n 0.00103531f $X=3.865 $Y=1.145 $X2=0 $Y2=0
cc_749 N_SET_B_M1004_g N_VGND_c_1789_n 0.0134999f $X=3.905 $Y=0.445 $X2=0 $Y2=0
cc_750 SET_B N_VGND_c_1789_n 0.0213368f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_751 N_SET_B_c_921_n N_VGND_c_1789_n 0.00267196f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_752 N_SET_B_c_920_n N_VGND_c_1791_n 0.00496953f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_753 N_SET_B_c_918_n N_VGND_c_1798_n 4.72037e-19 $X=7.01 $Y=0.9 $X2=0 $Y2=0
cc_754 N_SET_B_M1002_g N_VGND_c_1805_n 0.0196039f $X=6.785 $Y=0.445 $X2=0 $Y2=0
cc_755 N_SET_B_c_917_n N_VGND_c_1805_n 6.13185e-19 $X=6.845 $Y=0.98 $X2=0 $Y2=0
cc_756 N_SET_B_c_918_n N_VGND_c_1805_n 0.0391684f $X=7.01 $Y=0.9 $X2=0 $Y2=0
cc_757 N_SET_B_c_920_n N_VGND_c_1805_n 0.00136328f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_758 N_SET_B_c_922_n N_VGND_c_1805_n 0.00338478f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_759 N_SET_B_c_918_n N_VGND_c_1807_n 0.00125475f $X=7.01 $Y=0.9 $X2=0 $Y2=0
cc_760 SET_B N_VGND_c_1807_n 9.94995e-19 $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_761 N_SET_B_c_920_n N_VGND_c_1807_n 0.134969f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_762 N_SET_B_c_921_n N_VGND_c_1807_n 0.0146581f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_763 N_SET_B_c_922_n N_VGND_c_1807_n 0.0145013f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_764 N_SET_B_c_923_n N_VGND_c_1807_n 4.46136e-19 $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_765 N_A_476_47#_M1016_g N_A_1028_413#_c_1305_n 8.84083e-19 $X=4.705 $Y=2.275
+ $X2=0 $Y2=0
cc_766 N_A_476_47#_M1020_g N_VPWR_c_1520_n 0.00339367f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_767 N_A_476_47#_M1020_g N_VPWR_c_1521_n 0.00730335f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_768 N_A_476_47#_M1016_g N_VPWR_c_1521_n 0.00909428f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_769 N_A_476_47#_c_1074_n N_VPWR_c_1528_n 0.0377433f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_770 N_A_476_47#_M1016_g N_VPWR_c_1529_n 0.00414121f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_771 N_A_476_47#_M1020_g N_VPWR_c_1535_n 7.14614e-19 $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_772 N_A_476_47#_M1011_d N_VPWR_c_1517_n 0.00172638f $X=2.39 $Y=2.065 $X2=0
+ $Y2=0
cc_773 N_A_476_47#_M1020_g N_VPWR_c_1517_n 0.00379591f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_774 N_A_476_47#_M1016_g N_VPWR_c_1517_n 0.00402125f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_775 N_A_476_47#_c_1074_n N_VPWR_c_1517_n 0.0132505f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_776 N_A_476_47#_c_1074_n N_A_381_47#_c_1698_n 0.0102747f $X=3.02 $Y=2.335
+ $X2=0 $Y2=0
cc_777 N_A_476_47#_c_1074_n A_562_413# 0.00859792f $X=3.02 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_778 N_A_476_47#_c_1059_n A_562_413# 0.00578953f $X=3.105 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_779 N_A_476_47#_c_1047_n N_VGND_c_1789_n 0.00301834f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_780 N_A_476_47#_c_1047_n N_VGND_c_1790_n 0.00541969f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_781 N_A_476_47#_c_1049_n N_VGND_c_1790_n 0.00143459f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_782 N_A_476_47#_c_1047_n N_VGND_c_1791_n 0.00362321f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_783 N_A_476_47#_c_1049_n N_VGND_c_1791_n 0.00600607f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_784 N_A_476_47#_c_1050_n N_VGND_c_1791_n 0.00456783f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_785 N_A_476_47#_c_1079_n N_VGND_c_1797_n 0.055608f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_786 N_A_476_47#_c_1050_n N_VGND_c_1798_n 0.00437852f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_787 N_A_476_47#_M1028_d N_VGND_c_1807_n 0.00275359f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_788 N_A_476_47#_c_1047_n N_VGND_c_1807_n 0.00742824f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_789 N_A_476_47#_c_1049_n N_VGND_c_1807_n 6.5555e-19 $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_790 N_A_476_47#_c_1050_n N_VGND_c_1807_n 0.00674913f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_791 N_A_476_47#_c_1079_n N_VGND_c_1807_n 0.0223868f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_792 N_A_476_47#_c_1079_n A_586_47# 0.00628999f $X=3.27 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_793 N_A_1178_261#_c_1213_n N_A_1028_413#_M1027_g 0.014379f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_794 N_A_1178_261#_c_1206_n N_A_1028_413#_M1013_g 0.0097853f $X=7.785 $Y=1.575
+ $X2=0 $Y2=0
cc_795 N_A_1178_261#_c_1206_n N_A_1028_413#_c_1284_n 0.024367f $X=7.785 $Y=1.575
+ $X2=0 $Y2=0
cc_796 N_A_1178_261#_c_1214_n N_A_1028_413#_c_1284_n 0.00658845f $X=7.785
+ $Y=1.67 $X2=0 $Y2=0
cc_797 N_A_1178_261#_c_1207_n N_A_1028_413#_c_1284_n 0.00425847f $X=7.785
+ $Y=0.515 $X2=0 $Y2=0
cc_798 N_A_1178_261#_c_1206_n N_A_1028_413#_c_1285_n 0.0053543f $X=7.785
+ $Y=1.575 $X2=0 $Y2=0
cc_799 N_A_1178_261#_c_1213_n N_A_1028_413#_c_1285_n 0.00263958f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_800 N_A_1178_261#_c_1206_n N_A_1028_413#_M1030_g 4.30058e-19 $X=7.785
+ $Y=1.575 $X2=0 $Y2=0
cc_801 N_A_1178_261#_c_1206_n N_A_1028_413#_c_1296_n 4.56062e-19 $X=7.785
+ $Y=1.575 $X2=0 $Y2=0
cc_802 N_A_1178_261#_c_1205_n N_A_1028_413#_c_1298_n 0.00400996f $X=6.425
+ $Y=1.38 $X2=0 $Y2=0
cc_803 N_A_1178_261#_c_1213_n N_A_1028_413#_c_1298_n 0.0133834f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_804 N_A_1178_261#_M1033_g N_A_1028_413#_c_1313_n 0.00613779f $X=6.425
+ $Y=0.445 $X2=0 $Y2=0
cc_805 N_A_1178_261#_c_1205_n N_A_1028_413#_c_1288_n 0.0138248f $X=6.425 $Y=1.38
+ $X2=0 $Y2=0
cc_806 N_A_1178_261#_c_1213_n N_A_1028_413#_c_1288_n 0.0281674f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_807 N_A_1178_261#_M1015_g N_A_1028_413#_c_1300_n 0.0119267f $X=5.965 $Y=2.275
+ $X2=0 $Y2=0
cc_808 N_A_1178_261#_c_1210_n N_A_1028_413#_c_1300_n 0.00460004f $X=6.05
+ $Y=1.825 $X2=0 $Y2=0
cc_809 N_A_1178_261#_c_1213_n N_A_1028_413#_c_1300_n 0.0654175f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_810 N_A_1178_261#_M1033_g N_A_1028_413#_c_1290_n 0.0184288f $X=6.425 $Y=0.445
+ $X2=0 $Y2=0
cc_811 N_A_1178_261#_M1015_g N_A_1028_413#_c_1301_n 0.00296198f $X=5.965
+ $Y=2.275 $X2=0 $Y2=0
cc_812 N_A_1178_261#_M1015_g N_A_1028_413#_c_1302_n 0.00444241f $X=5.965
+ $Y=2.275 $X2=0 $Y2=0
cc_813 N_A_1178_261#_c_1210_n N_A_1028_413#_c_1302_n 0.00400996f $X=6.05
+ $Y=1.825 $X2=0 $Y2=0
cc_814 N_A_1178_261#_M1033_g N_A_1028_413#_c_1384_n 0.0023431f $X=6.425 $Y=0.445
+ $X2=0 $Y2=0
cc_815 N_A_1178_261#_c_1205_n N_A_1028_413#_c_1384_n 0.00339988f $X=6.425
+ $Y=1.38 $X2=0 $Y2=0
cc_816 N_A_1178_261#_c_1213_n N_A_1028_413#_c_1384_n 0.0135849f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_817 N_A_1178_261#_c_1206_n N_A_1028_413#_c_1291_n 0.0151462f $X=7.785
+ $Y=1.575 $X2=0 $Y2=0
cc_818 N_A_1178_261#_M1033_g N_A_1028_413#_c_1292_n 0.00108423f $X=6.425
+ $Y=0.445 $X2=0 $Y2=0
cc_819 N_A_1178_261#_c_1205_n N_A_1028_413#_c_1292_n 0.00142532f $X=6.425
+ $Y=1.38 $X2=0 $Y2=0
cc_820 N_A_1178_261#_c_1213_n N_A_1028_413#_c_1292_n 0.0722425f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_821 N_A_1178_261#_c_1206_n N_A_1602_47#_c_1444_n 0.0236103f $X=7.785 $Y=1.575
+ $X2=0 $Y2=0
cc_822 N_A_1178_261#_c_1207_n N_A_1602_47#_c_1444_n 0.0258113f $X=7.785 $Y=0.515
+ $X2=0 $Y2=0
cc_823 N_A_1178_261#_c_1264_p N_A_1602_47#_c_1450_n 0.00631112f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_824 N_A_1178_261#_c_1206_n N_A_1602_47#_c_1450_n 0.0187258f $X=7.785 $Y=1.575
+ $X2=0 $Y2=0
cc_825 N_A_1178_261#_c_1214_n N_A_1602_47#_c_1450_n 0.0159581f $X=7.785 $Y=1.67
+ $X2=0 $Y2=0
cc_826 N_A_1178_261#_c_1264_p N_A_1602_47#_c_1452_n 0.0244707f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_827 N_A_1178_261#_c_1206_n N_A_1602_47#_c_1446_n 0.0261658f $X=7.785 $Y=1.575
+ $X2=0 $Y2=0
cc_828 N_A_1178_261#_c_1213_n N_VPWR_M1001_d 0.00219976f $X=7.51 $Y=1.67 $X2=0
+ $Y2=0
cc_829 N_A_1178_261#_c_1213_n N_VPWR_c_1522_n 0.0194966f $X=7.51 $Y=1.67 $X2=0
+ $Y2=0
cc_830 N_A_1178_261#_M1015_g N_VPWR_c_1529_n 8.50188e-19 $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_831 N_A_1178_261#_c_1264_p N_VPWR_c_1531_n 0.00737773f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_832 N_A_1178_261#_M1015_g N_VPWR_c_1537_n 0.0145664f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_833 N_A_1178_261#_M1027_d N_VPWR_c_1517_n 0.00556469f $X=7.455 $Y=1.645 $X2=0
+ $Y2=0
cc_834 N_A_1178_261#_M1015_g N_VPWR_c_1517_n 0.00145798f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_835 N_A_1178_261#_c_1264_p N_VPWR_c_1517_n 0.00613728f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_836 N_A_1178_261#_M1033_g N_VGND_c_1798_n 0.0038242f $X=6.425 $Y=0.445 $X2=0
+ $Y2=0
cc_837 N_A_1178_261#_c_1207_n N_VGND_c_1799_n 0.0144375f $X=7.785 $Y=0.515 $X2=0
+ $Y2=0
cc_838 N_A_1178_261#_M1033_g N_VGND_c_1805_n 0.00311464f $X=6.425 $Y=0.445 $X2=0
+ $Y2=0
cc_839 N_A_1178_261#_M1013_d N_VGND_c_1807_n 0.00391384f $X=7.48 $Y=0.235 $X2=0
+ $Y2=0
cc_840 N_A_1178_261#_M1033_g N_VGND_c_1807_n 0.00503783f $X=6.425 $Y=0.445 $X2=0
+ $Y2=0
cc_841 N_A_1178_261#_c_1207_n N_VGND_c_1807_n 0.0125017f $X=7.785 $Y=0.515 $X2=0
+ $Y2=0
cc_842 N_A_1028_413#_M1030_g N_A_1602_47#_c_1442_n 0.0110206f $X=8.345 $Y=0.56
+ $X2=0 $Y2=0
cc_843 N_A_1028_413#_c_1287_n N_A_1602_47#_M1025_g 0.0143036f $X=8.345 $Y=1.252
+ $X2=0 $Y2=0
cc_844 N_A_1028_413#_M1030_g N_A_1602_47#_c_1444_n 0.00772027f $X=8.345 $Y=0.56
+ $X2=0 $Y2=0
cc_845 N_A_1028_413#_M1027_g N_A_1602_47#_c_1450_n 5.88209e-19 $X=7.38 $Y=2.065
+ $X2=0 $Y2=0
cc_846 N_A_1028_413#_c_1284_n N_A_1602_47#_c_1450_n 0.00606446f $X=8.27 $Y=1.252
+ $X2=0 $Y2=0
cc_847 N_A_1028_413#_c_1296_n N_A_1602_47#_c_1450_n 0.00735044f $X=8.345 $Y=1.41
+ $X2=0 $Y2=0
cc_848 N_A_1028_413#_c_1287_n N_A_1602_47#_c_1450_n 0.00151929f $X=8.345
+ $Y=1.252 $X2=0 $Y2=0
cc_849 N_A_1028_413#_M1030_g N_A_1602_47#_c_1445_n 0.00668119f $X=8.345 $Y=0.56
+ $X2=0 $Y2=0
cc_850 N_A_1028_413#_c_1287_n N_A_1602_47#_c_1445_n 0.0103507f $X=8.345 $Y=1.252
+ $X2=0 $Y2=0
cc_851 N_A_1028_413#_M1027_g N_A_1602_47#_c_1452_n 0.00147349f $X=7.38 $Y=2.065
+ $X2=0 $Y2=0
cc_852 N_A_1028_413#_c_1284_n N_A_1602_47#_c_1452_n 0.00235755f $X=8.27 $Y=1.252
+ $X2=0 $Y2=0
cc_853 N_A_1028_413#_c_1296_n N_A_1602_47#_c_1452_n 0.00559869f $X=8.345 $Y=1.41
+ $X2=0 $Y2=0
cc_854 N_A_1028_413#_c_1284_n N_A_1602_47#_c_1446_n 0.0112725f $X=8.27 $Y=1.252
+ $X2=0 $Y2=0
cc_855 N_A_1028_413#_M1030_g N_A_1602_47#_c_1446_n 0.00369472f $X=8.345 $Y=0.56
+ $X2=0 $Y2=0
cc_856 N_A_1028_413#_c_1287_n N_A_1602_47#_c_1446_n 6.49734e-19 $X=8.345
+ $Y=1.252 $X2=0 $Y2=0
cc_857 N_A_1028_413#_M1030_g N_A_1602_47#_c_1447_n 0.0215122f $X=8.345 $Y=0.56
+ $X2=0 $Y2=0
cc_858 N_A_1028_413#_c_1300_n N_VPWR_M1015_d 0.00216018f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_859 N_A_1028_413#_c_1305_n N_VPWR_c_1521_n 0.00557448f $X=5.57 $Y=2.29 $X2=0
+ $Y2=0
cc_860 N_A_1028_413#_M1027_g N_VPWR_c_1522_n 0.0157666f $X=7.38 $Y=2.065 $X2=0
+ $Y2=0
cc_861 N_A_1028_413#_c_1300_n N_VPWR_c_1522_n 0.00850121f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_862 N_A_1028_413#_c_1296_n N_VPWR_c_1523_n 0.00268723f $X=8.345 $Y=1.41 $X2=0
+ $Y2=0
cc_863 N_A_1028_413#_c_1305_n N_VPWR_c_1529_n 0.0200526f $X=5.57 $Y=2.29 $X2=0
+ $Y2=0
cc_864 N_A_1028_413#_c_1300_n N_VPWR_c_1529_n 0.00267646f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_865 N_A_1028_413#_c_1302_n N_VPWR_c_1529_n 0.00720374f $X=5.655 $Y=2 $X2=0
+ $Y2=0
cc_866 N_A_1028_413#_c_1300_n N_VPWR_c_1530_n 0.0036467f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_867 N_A_1028_413#_c_1301_n N_VPWR_c_1530_n 0.0101929f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_868 N_A_1028_413#_M1027_g N_VPWR_c_1531_n 0.00447018f $X=7.38 $Y=2.065 $X2=0
+ $Y2=0
cc_869 N_A_1028_413#_c_1296_n N_VPWR_c_1531_n 0.00542953f $X=8.345 $Y=1.41 $X2=0
+ $Y2=0
cc_870 N_A_1028_413#_c_1300_n N_VPWR_c_1537_n 0.0270337f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_871 N_A_1028_413#_c_1301_n N_VPWR_c_1537_n 0.00887045f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_872 N_A_1028_413#_c_1302_n N_VPWR_c_1537_n 0.0115187f $X=5.655 $Y=2 $X2=0
+ $Y2=0
cc_873 N_A_1028_413#_M1005_d N_VPWR_c_1517_n 0.0026466f $X=5.14 $Y=2.065 $X2=0
+ $Y2=0
cc_874 N_A_1028_413#_M1001_s N_VPWR_c_1517_n 0.00394021f $X=6.57 $Y=2.065 $X2=0
+ $Y2=0
cc_875 N_A_1028_413#_M1027_g N_VPWR_c_1517_n 0.0090376f $X=7.38 $Y=2.065 $X2=0
+ $Y2=0
cc_876 N_A_1028_413#_c_1296_n N_VPWR_c_1517_n 0.0108575f $X=8.345 $Y=1.41 $X2=0
+ $Y2=0
cc_877 N_A_1028_413#_c_1305_n N_VPWR_c_1517_n 0.00987026f $X=5.57 $Y=2.29 $X2=0
+ $Y2=0
cc_878 N_A_1028_413#_c_1300_n N_VPWR_c_1517_n 0.0124969f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_879 N_A_1028_413#_c_1301_n N_VPWR_c_1517_n 0.0086238f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_880 N_A_1028_413#_c_1302_n N_VPWR_c_1517_n 0.00578252f $X=5.655 $Y=2 $X2=0
+ $Y2=0
cc_881 N_A_1028_413#_c_1300_n A_1136_413# 0.00166681f $X=6.54 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_882 N_A_1028_413#_c_1302_n A_1136_413# 0.00336335f $X=5.655 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_883 N_A_1028_413#_M1030_g N_VGND_c_1792_n 0.0152147f $X=8.345 $Y=0.56 $X2=0
+ $Y2=0
cc_884 N_A_1028_413#_c_1313_n N_VGND_c_1798_n 0.0363343f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_885 N_A_1028_413#_M1013_g N_VGND_c_1799_n 0.00575639f $X=7.405 $Y=0.505 $X2=0
+ $Y2=0
cc_886 N_A_1028_413#_M1030_g N_VGND_c_1799_n 0.0046653f $X=8.345 $Y=0.56 $X2=0
+ $Y2=0
cc_887 N_A_1028_413#_M1013_g N_VGND_c_1805_n 0.00610968f $X=7.405 $Y=0.505 $X2=0
+ $Y2=0
cc_888 N_A_1028_413#_M1014_d N_VGND_c_1807_n 0.00232124f $X=5.64 $Y=0.235 $X2=0
+ $Y2=0
cc_889 N_A_1028_413#_M1013_g N_VGND_c_1807_n 0.0120867f $X=7.405 $Y=0.505 $X2=0
+ $Y2=0
cc_890 N_A_1028_413#_M1030_g N_VGND_c_1807_n 0.00934473f $X=8.345 $Y=0.56 $X2=0
+ $Y2=0
cc_891 N_A_1028_413#_c_1313_n N_VGND_c_1807_n 0.0135337f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_892 N_A_1028_413#_c_1313_n A_1228_47# 0.00244121f $X=6.32 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_893 N_A_1602_47#_c_1452_n N_VPWR_c_1522_n 0.00146605f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_894 N_A_1602_47#_M1025_g N_VPWR_c_1523_n 0.00146448f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_895 N_A_1602_47#_c_1445_n N_VPWR_c_1523_n 0.0139885f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_896 N_A_1602_47#_M1032_g N_VPWR_c_1525_n 0.00322031f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_897 N_A_1602_47#_c_1452_n N_VPWR_c_1531_n 0.0166647f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_898 N_A_1602_47#_M1025_g N_VPWR_c_1532_n 0.00541562f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_899 N_A_1602_47#_M1032_g N_VPWR_c_1532_n 0.00541562f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_900 N_A_1602_47#_M1006_s N_VPWR_c_1517_n 0.00211564f $X=8.01 $Y=1.485 $X2=0
+ $Y2=0
cc_901 N_A_1602_47#_M1025_g N_VPWR_c_1517_n 0.00952891f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_902 N_A_1602_47#_M1032_g N_VPWR_c_1517_n 0.0104607f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_903 N_A_1602_47#_c_1452_n N_VPWR_c_1517_n 0.0121504f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_904 N_A_1602_47#_c_1443_n Q 0.0123161f $X=9.185 $Y=0.995 $X2=0 $Y2=0
cc_905 N_A_1602_47#_c_1442_n Q 0.00254238f $X=8.765 $Y=0.995 $X2=0 $Y2=0
cc_906 N_A_1602_47#_M1025_g Q 0.00305599f $X=8.765 $Y=1.985 $X2=0 $Y2=0
cc_907 N_A_1602_47#_c_1443_n Q 0.00392121f $X=9.185 $Y=0.995 $X2=0 $Y2=0
cc_908 N_A_1602_47#_M1032_g Q 0.00472146f $X=9.185 $Y=1.985 $X2=0 $Y2=0
cc_909 N_A_1602_47#_c_1445_n Q 0.0272055f $X=8.765 $Y=1.16 $X2=0 $Y2=0
cc_910 N_A_1602_47#_c_1447_n Q 0.0186982f $X=9.185 $Y=1.16 $X2=0 $Y2=0
cc_911 N_A_1602_47#_M1025_g N_Q_c_1758_n 0.00232678f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_912 N_A_1602_47#_M1032_g N_Q_c_1758_n 0.0123446f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_913 N_A_1602_47#_c_1450_n N_Q_c_1758_n 0.00140427f $X=8.135 $Y=1.66 $X2=0
+ $Y2=0
cc_914 N_A_1602_47#_c_1445_n N_Q_c_1758_n 0.00272962f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_915 N_A_1602_47#_c_1447_n N_Q_c_1758_n 0.00274767f $X=9.185 $Y=1.16 $X2=0
+ $Y2=0
cc_916 N_A_1602_47#_M1025_g N_Q_c_1771_n 0.00904859f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_917 N_A_1602_47#_M1032_g N_Q_c_1771_n 0.0150609f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_918 N_A_1602_47#_c_1442_n N_Q_c_1756_n 0.00190516f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_919 N_A_1602_47#_c_1443_n N_Q_c_1756_n 0.00812757f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_920 N_A_1602_47#_c_1447_n N_Q_c_1756_n 0.00272044f $X=9.185 $Y=1.16 $X2=0
+ $Y2=0
cc_921 N_A_1602_47#_c_1442_n N_VGND_c_1792_n 0.0106232f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_922 N_A_1602_47#_c_1443_n N_VGND_c_1792_n 7.90377e-19 $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_923 N_A_1602_47#_c_1445_n N_VGND_c_1792_n 0.0225891f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_924 N_A_1602_47#_c_1447_n N_VGND_c_1792_n 0.00122405f $X=9.185 $Y=1.16 $X2=0
+ $Y2=0
cc_925 N_A_1602_47#_c_1443_n N_VGND_c_1794_n 0.00353994f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_926 N_A_1602_47#_c_1444_n N_VGND_c_1799_n 0.00732874f $X=8.135 $Y=0.51 $X2=0
+ $Y2=0
cc_927 N_A_1602_47#_c_1442_n N_VGND_c_1800_n 0.0046653f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_928 N_A_1602_47#_c_1443_n N_VGND_c_1800_n 0.00549284f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_929 N_A_1602_47#_M1030_s N_VGND_c_1807_n 0.00535012f $X=8.01 $Y=0.235 $X2=0
+ $Y2=0
cc_930 N_A_1602_47#_c_1442_n N_VGND_c_1807_n 0.00796766f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_931 N_A_1602_47#_c_1443_n N_VGND_c_1807_n 0.00681022f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_932 N_A_1602_47#_c_1444_n N_VGND_c_1807_n 0.00616598f $X=8.135 $Y=0.51 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1517_n N_A_381_47#_M1023_d 0.00325229f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_934 N_VPWR_M1023_s N_A_381_47#_c_1688_n 0.00237137f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_935 N_VPWR_M1023_s N_A_381_47#_c_1695_n 0.00471078f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1519_n N_A_381_47#_c_1695_n 0.00880041f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1528_n N_A_381_47#_c_1695_n 0.0018545f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1517_n N_A_381_47#_c_1695_n 0.00198108f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_939 N_VPWR_M1023_s N_A_381_47#_c_1691_n 0.00187968f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1519_n N_A_381_47#_c_1691_n 0.0114817f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1527_n N_A_381_47#_c_1691_n 3.86777e-19 $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1517_n N_A_381_47#_c_1691_n 7.1462e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1528_n N_A_381_47#_c_1698_n 0.0115924f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1517_n N_A_381_47#_c_1698_n 0.00307944f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1517_n A_562_413# 0.00355877f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_946 N_VPWR_c_1517_n A_956_413# 0.00250248f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_947 N_VPWR_c_1517_n A_1136_413# 0.00223276f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_948 N_VPWR_c_1517_n N_Q_M1025_s 0.00215347f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_949 N_VPWR_M1032_d N_Q_c_1758_n 0.00282209f $X=9.26 $Y=1.485 $X2=0 $Y2=0
cc_950 N_VPWR_c_1525_n N_Q_c_1758_n 0.0233625f $X=9.395 $Y=1.955 $X2=0 $Y2=0
cc_951 N_VPWR_c_1532_n N_Q_c_1771_n 0.0183232f $X=9.31 $Y=2.72 $X2=0 $Y2=0
cc_952 N_VPWR_c_1517_n N_Q_c_1771_n 0.0121916f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_953 N_A_381_47#_c_1688_n N_VGND_M1010_s 0.00105184f $X=1.515 $Y=1.795 $X2=0
+ $Y2=0
cc_954 N_A_381_47#_c_1693_n N_VGND_M1010_s 0.00264874f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_955 N_A_381_47#_c_1689_n N_VGND_M1010_s 0.0019591f $X=1.6 $Y=0.73 $X2=0 $Y2=0
cc_956 N_A_381_47#_c_1693_n N_VGND_c_1788_n 0.00883988f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_957 N_A_381_47#_c_1689_n N_VGND_c_1788_n 0.0114461f $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_958 N_A_381_47#_c_1689_n N_VGND_c_1796_n 4.97798e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_959 N_A_381_47#_c_1693_n N_VGND_c_1797_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_960 N_A_381_47#_c_1697_n N_VGND_c_1797_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_961 N_A_381_47#_M1010_d N_VGND_c_1807_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_962 N_A_381_47#_c_1693_n N_VGND_c_1807_n 0.00232804f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_963 N_A_381_47#_c_1689_n N_VGND_c_1807_n 8.52239e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_964 N_A_381_47#_c_1697_n N_VGND_c_1807_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_965 N_Q_c_1756_n N_VGND_M1008_d 0.00273341f $X=9.297 $Y=0.895 $X2=0 $Y2=0
cc_966 N_Q_c_1756_n N_VGND_c_1794_n 0.022629f $X=9.297 $Y=0.895 $X2=0 $Y2=0
cc_967 Q N_VGND_c_1800_n 0.013861f $X=8.895 $Y=0.425 $X2=0 $Y2=0
cc_968 N_Q_M1003_s N_VGND_c_1807_n 0.0039413f $X=8.84 $Y=0.235 $X2=0 $Y2=0
cc_969 Q N_VGND_c_1807_n 0.00918227f $X=8.895 $Y=0.425 $X2=0 $Y2=0
cc_970 N_Q_c_1756_n N_VGND_c_1807_n 0.007194f $X=9.297 $Y=0.895 $X2=0 $Y2=0
cc_971 N_VGND_c_1807_n A_586_47# 0.00231384f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_972 N_VGND_c_1807_n A_796_47# 0.00240916f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_973 N_VGND_c_1807_n A_1056_47# 0.00198596f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_974 N_VGND_c_1807_n A_1228_47# 0.0014047f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_975 N_VGND_c_1807_n A_1300_47# 0.00257789f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o2bb2ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.625000 1.445000 ;
        RECT 0.090000 1.445000 1.945000 1.615000 ;
        RECT 1.615000 1.075000 1.945000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795000 1.075000 1.400000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.075000 3.740000 1.445000 ;
        RECT 3.410000 1.445000 5.435000 1.615000 ;
        RECT 4.730000 1.075000 5.435000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.960000 1.075000 4.500000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 0.645000 3.075000 1.075000 ;
        RECT 2.745000 1.075000 3.215000 1.785000 ;
        RECT 2.745000 1.785000 4.330000 1.955000 ;
        RECT 2.745000 1.955000 3.035000 2.465000 ;
        RECT 4.080000 1.955000 4.330000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.195000  0.085000 0.365000 0.895000 ;
        RECT 1.875000  0.085000 2.045000 0.555000 ;
        RECT 3.700000  0.085000 3.870000 0.555000 ;
        RECT 4.540000  0.085000 4.710000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.150000 1.795000 0.400000 2.635000 ;
        RECT 0.995000 2.135000 1.245000 2.635000 ;
        RECT 1.835000 2.135000 2.575000 2.635000 ;
        RECT 3.205000 2.125000 3.490000 2.635000 ;
        RECT 4.965000 1.795000 5.170000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.535000 0.305000 1.705000 0.475000 ;
      RECT 0.535000 0.475000 0.785000 0.895000 ;
      RECT 0.575000 1.785000 2.285000 1.965000 ;
      RECT 0.575000 1.965000 0.825000 2.465000 ;
      RECT 0.955000 0.645000 1.285000 0.725000 ;
      RECT 0.955000 0.725000 2.285000 0.905000 ;
      RECT 1.415000 1.965000 1.665000 2.125000 ;
      RECT 2.115000 0.905000 2.285000 0.995000 ;
      RECT 2.115000 0.995000 2.575000 1.325000 ;
      RECT 2.115000 1.325000 2.285000 1.785000 ;
      RECT 2.325000 0.255000 3.530000 0.475000 ;
      RECT 2.325000 0.475000 2.575000 0.555000 ;
      RECT 3.245000 0.475000 3.530000 0.735000 ;
      RECT 3.245000 0.735000 5.210000 0.905000 ;
      RECT 3.660000 2.125000 3.910000 2.295000 ;
      RECT 3.660000 2.295000 4.750000 2.465000 ;
      RECT 4.040000 0.255000 4.370000 0.725000 ;
      RECT 4.040000 0.725000 5.210000 0.735000 ;
      RECT 4.500000 1.785000 4.750000 2.295000 ;
      RECT 4.880000 0.255000 5.210000 0.725000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_2
END LIBRARY

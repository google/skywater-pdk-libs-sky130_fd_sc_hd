* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2.spice
* Created: Tue Sep  1 19:13:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2  VGND VPB VPWRIN A
+ VPWR X
* 
* X	X
* VPWR	VPWR
* A	A
* VPWRIN	VPWRIN
* VPB	VPB
* VGND	VGND
MM1012 N_A_505_297#_M1012_d N_A_M1012_g N_VGND_M1012_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_620_911#_M1002_d N_A_505_297#_M1002_g N_VGND_M1002_s N_VGND_M1012_b
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_620_911#_M1002_d N_A_505_297#_M1008_g N_VGND_M1008_s N_VGND_M1012_b
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75000.6 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1003 N_A_714_47#_M1003_d N_A_M1003_g N_VGND_M1003_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.65 AD=0.091 AS=0.18525 PD=0.93 PS=1.87 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1015 N_A_620_911#_M1015_d N_A_505_297#_M1015_g N_VGND_M1008_s N_VGND_M1012_b
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75001.1 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_A_714_47#_M1003_d N_A_M1004_g N_VGND_M1004_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1016 N_A_620_911#_M1015_d N_A_505_297#_M1016_g N_VGND_M1016_s N_VGND_M1012_b
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.2015 PD=0.93 PS=1.27 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75001.5 SB=75001 A=0.0975 P=1.6 MULT=1
MM1007 N_A_714_47#_M1007_d N_A_M1007_g N_VGND_M1004_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_714_47#_M1007_d N_A_M1010_g N_VGND_M1010_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.65 AD=0.091 AS=0.104 PD=0.93 PS=0.97 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1009 N_A_1032_911#_M1009_d N_A_620_911#_M1009_g N_VGND_M1016_s N_VGND_M1012_b
+ NSHORT L=0.15 W=0.65 AD=0.17225 AS=0.2015 PD=1.83 PS=1.27 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1005_d N_A_1032_911#_M1005_g N_VGND_M1010_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=0 NRS=7.38 M=1 R=4.33333
+ SA=75002 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_X_M1005_d N_A_1032_911#_M1014_g N_VGND_M1014_s N_VGND_M1012_b NSHORT
+ L=0.15 W=0.65 AD=0.12025 AS=0.18525 PD=1.02 PS=1.87 NRD=16.608 NRS=0 M=1
+ R=4.33333 SA=75002.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_505_297#_M1011_d N_A_M1011_g N_VPWRIN_M1011_s N_VPWRIN_M1011_b
+ PHIGHVT L=0.15 W=1 AD=0.275 AS=0.275 PD=2.55 PS=2.55 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A_714_47#_M1017_g N_A_620_911#_M1017_s N_VPB_M1017_b
+ PHIGHVT L=0.15 W=0.79 AD=0.136485 AS=0.21725 PD=1.16955 PS=2.13 NRD=2.4822
+ NRS=2.4822 M=1 R=5.26667 SA=75000.2 SB=75001.2 A=0.1185 P=1.88 MULT=1
MM1000 N_VPWR_M1000_d N_A_620_911#_M1000_g N_A_714_47#_M1000_s N_VPB_M1017_b
+ PHIGHVT L=0.15 W=0.79 AD=0.120475 AS=0.21725 PD=1.095 PS=2.13 NRD=2.4822
+ NRS=1.2411 M=1 R=5.26667 SA=75000.2 SB=75000.7 A=0.1185 P=1.88 MULT=1
MM1001 N_A_1032_911#_M1001_d N_A_620_911#_M1001_g N_VPWR_M1000_d N_VPB_M1017_b
+ PHIGHVT L=0.15 W=0.79 AD=0.2133 AS=0.120475 PD=2.12 PS=1.095 NRD=1.2411
+ NRS=3.7233 M=1 R=5.26667 SA=75000.7 SB=75000.2 A=0.1185 P=1.88 MULT=1
MM1006 N_VPWR_M1017_d N_A_1032_911#_M1006_g N_X_M1006_s N_VPB_M1017_b PHIGHVT
+ L=0.15 W=1 AD=0.172765 AS=0.185 PD=1.48045 PS=1.37 NRD=6.8753 NRS=0 M=1
+ R=6.66667 SA=75000.6 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_1032_911#_M1013_g N_X_M1006_s N_VPB_M1017_b PHIGHVT
+ L=0.15 W=1 AD=0.285 AS=0.185 PD=2.57 PS=1.37 NRD=0 NRS=17.73 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref N_VGND_M1012_b N_VPB_X18_noxref_D1 NWDIODE A=2.3772 P=7.34
DX19_noxref N_VGND_M1012_b N_VPWRIN_M1011_b NWDIODE A=2.9998 P=7.78
DX20_noxref N_VGND_M1012_b N_VPB_M1017_b NWDIODE A=6.7354 P=10.42
*
.include "sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__fah_1.pxi.spice
* Created: Tue Sep  1 19:08:56 2020
* 
x_PM_SKY130_FD_SC_HD__FAH_1%A_67_199# N_A_67_199#_M1031_d N_A_67_199#_M1007_d
+ N_A_67_199#_M1029_g N_A_67_199#_M1006_g N_A_67_199#_c_236_n
+ N_A_67_199#_c_237_n N_A_67_199#_c_238_n N_A_67_199#_c_239_n
+ N_A_67_199#_c_240_n PM_SKY130_FD_SC_HD__FAH_1%A_67_199#
x_PM_SKY130_FD_SC_HD__FAH_1%A N_A_M1007_g N_A_c_297_n N_A_M1031_g N_A_c_298_n
+ N_A_M1018_g N_A_M1015_g N_A_c_299_n N_A_c_300_n N_A_c_301_n A
+ PM_SKY130_FD_SC_HD__FAH_1%A
x_PM_SKY130_FD_SC_HD__FAH_1%B N_B_M1012_g N_B_c_357_n N_B_M1000_g N_B_c_358_n
+ N_B_c_359_n N_B_c_360_n N_B_M1027_g N_B_M1023_g N_B_M1020_g N_B_c_361_n
+ N_B_M1014_g N_B_c_362_n N_B_c_397_p B N_B_c_363_n N_B_c_364_n B N_B_c_415_p
+ N_B_c_365_n N_B_c_366_n N_B_c_367_n PM_SKY130_FD_SC_HD__FAH_1%B
x_PM_SKY130_FD_SC_HD__FAH_1%A_508_297# N_A_508_297#_M1000_d N_A_508_297#_M1021_d
+ N_A_508_297#_M1012_d N_A_508_297#_M1026_s N_A_508_297#_c_533_n
+ N_A_508_297#_M1013_g N_A_508_297#_M1010_g N_A_508_297#_c_534_n
+ N_A_508_297#_M1002_g N_A_508_297#_M1022_g N_A_508_297#_c_535_n
+ N_A_508_297#_c_536_n N_A_508_297#_c_537_n N_A_508_297#_c_538_n
+ N_A_508_297#_c_726_p N_A_508_297#_c_595_p N_A_508_297#_c_637_p
+ N_A_508_297#_c_547_n N_A_508_297#_c_539_n N_A_508_297#_c_548_n
+ N_A_508_297#_c_540_n N_A_508_297#_c_549_n N_A_508_297#_c_550_n
+ N_A_508_297#_c_551_n N_A_508_297#_c_552_n N_A_508_297#_c_553_n
+ N_A_508_297#_c_554_n N_A_508_297#_c_555_n PM_SKY130_FD_SC_HD__FAH_1%A_508_297#
x_PM_SKY130_FD_SC_HD__FAH_1%A_719_47# N_A_719_47#_M1027_d N_A_719_47#_M1023_d
+ N_A_719_47#_M1026_g N_A_719_47#_c_737_n N_A_719_47#_M1004_g
+ N_A_719_47#_c_738_n N_A_719_47#_M1003_g N_A_719_47#_c_739_n
+ N_A_719_47#_c_740_n N_A_719_47#_M1016_g N_A_719_47#_c_742_n
+ N_A_719_47#_c_743_n N_A_719_47#_c_744_n N_A_719_47#_c_762_n
+ N_A_719_47#_c_763_n N_A_719_47#_c_758_n N_A_719_47#_c_745_n
+ N_A_719_47#_c_746_n N_A_719_47#_c_747_n N_A_719_47#_c_748_n
+ N_A_719_47#_c_749_n N_A_719_47#_c_750_n N_A_719_47#_c_751_n
+ N_A_719_47#_c_752_n N_A_719_47#_c_753_n PM_SKY130_FD_SC_HD__FAH_1%A_719_47#
x_PM_SKY130_FD_SC_HD__FAH_1%A_1008_47# N_A_1008_47#_M1002_d N_A_1008_47#_M1022_d
+ N_A_1008_47#_M1008_g N_A_1008_47#_c_958_n N_A_1008_47#_M1021_g
+ N_A_1008_47#_c_959_n N_A_1008_47#_M1009_g N_A_1008_47#_c_967_n
+ N_A_1008_47#_c_968_n N_A_1008_47#_M1019_g N_A_1008_47#_c_960_n
+ N_A_1008_47#_c_961_n N_A_1008_47#_c_971_n N_A_1008_47#_c_972_n
+ N_A_1008_47#_c_973_n N_A_1008_47#_c_962_n N_A_1008_47#_c_963_n
+ N_A_1008_47#_c_974_n N_A_1008_47#_c_975_n N_A_1008_47#_c_964_n
+ N_A_1008_47#_c_965_n PM_SKY130_FD_SC_HD__FAH_1%A_1008_47#
x_PM_SKY130_FD_SC_HD__FAH_1%CI N_CI_M1024_g N_CI_M1025_g N_CI_c_1128_n
+ N_CI_c_1129_n N_CI_c_1130_n CI N_CI_c_1132_n PM_SKY130_FD_SC_HD__FAH_1%CI
x_PM_SKY130_FD_SC_HD__FAH_1%A_1262_49# N_A_1262_49#_M1004_s N_A_1262_49#_M1009_s
+ N_A_1262_49#_M1024_s N_A_1262_49#_M1008_d N_A_1262_49#_M1016_d
+ N_A_1262_49#_M1028_g N_A_1262_49#_M1005_g N_A_1262_49#_c_1195_n
+ N_A_1262_49#_c_1216_n N_A_1262_49#_c_1203_n N_A_1262_49#_c_1204_n
+ N_A_1262_49#_c_1196_n N_A_1262_49#_c_1205_n N_A_1262_49#_c_1206_n
+ N_A_1262_49#_c_1274_n N_A_1262_49#_c_1233_n N_A_1262_49#_c_1277_n
+ N_A_1262_49#_c_1197_n N_A_1262_49#_c_1198_n N_A_1262_49#_c_1199_n
+ N_A_1262_49#_c_1258_n N_A_1262_49#_c_1217_n N_A_1262_49#_c_1200_n
+ N_A_1262_49#_c_1201_n PM_SKY130_FD_SC_HD__FAH_1%A_1262_49#
x_PM_SKY130_FD_SC_HD__FAH_1%A_1332_297# N_A_1332_297#_M1004_d
+ N_A_1332_297#_M1026_d N_A_1332_297#_M1011_g N_A_1332_297#_M1001_g
+ N_A_1332_297#_c_1369_n N_A_1332_297#_c_1370_n N_A_1332_297#_c_1377_n
+ N_A_1332_297#_c_1371_n N_A_1332_297#_c_1388_n N_A_1332_297#_c_1372_n
+ N_A_1332_297#_c_1442_p N_A_1332_297#_c_1373_n N_A_1332_297#_c_1374_n
+ N_A_1332_297#_c_1375_n PM_SKY130_FD_SC_HD__FAH_1%A_1332_297#
x_PM_SKY130_FD_SC_HD__FAH_1%A_1617_49# N_A_1617_49#_M1009_d N_A_1617_49#_M1019_d
+ N_A_1617_49#_c_1482_n N_A_1617_49#_M1017_g N_A_1617_49#_M1030_g
+ N_A_1617_49#_c_1483_n N_A_1617_49#_c_1484_n N_A_1617_49#_c_1489_n
+ N_A_1617_49#_c_1490_n N_A_1617_49#_c_1491_n N_A_1617_49#_c_1492_n
+ N_A_1617_49#_c_1485_n N_A_1617_49#_c_1486_n N_A_1617_49#_c_1495_n
+ PM_SKY130_FD_SC_HD__FAH_1%A_1617_49#
x_PM_SKY130_FD_SC_HD__FAH_1%A_27_47# N_A_27_47#_M1029_s N_A_27_47#_M1013_d
+ N_A_27_47#_M1014_d N_A_27_47#_M1006_s N_A_27_47#_M1023_s N_A_27_47#_M1022_s
+ N_A_27_47#_c_1601_n N_A_27_47#_c_1607_n N_A_27_47#_c_1608_n
+ N_A_27_47#_c_1609_n N_A_27_47#_c_1610_n N_A_27_47#_c_1611_n
+ N_A_27_47#_c_1649_n N_A_27_47#_c_1612_n N_A_27_47#_c_1602_n
+ N_A_27_47#_c_1652_n N_A_27_47#_c_1653_n N_A_27_47#_c_1680_n
+ N_A_27_47#_c_1603_n N_A_27_47#_c_1614_n N_A_27_47#_c_1604_n
+ N_A_27_47#_c_1616_n N_A_27_47#_c_1605_n N_A_27_47#_c_1606_n
+ PM_SKY130_FD_SC_HD__FAH_1%A_27_47#
x_PM_SKY130_FD_SC_HD__FAH_1%VPWR N_VPWR_M1006_d N_VPWR_M1015_d N_VPWR_M1025_d
+ N_VPWR_M1001_d N_VPWR_c_1770_n N_VPWR_c_1771_n N_VPWR_c_1772_n N_VPWR_c_1773_n
+ VPWR N_VPWR_c_1774_n N_VPWR_c_1775_n N_VPWR_c_1776_n N_VPWR_c_1777_n
+ N_VPWR_c_1778_n N_VPWR_c_1769_n N_VPWR_c_1780_n N_VPWR_c_1781_n
+ N_VPWR_c_1782_n N_VPWR_c_1783_n PM_SKY130_FD_SC_HD__FAH_1%VPWR
x_PM_SKY130_FD_SC_HD__FAH_1%A_310_49# N_A_310_49#_M1018_s N_A_310_49#_M1027_s
+ N_A_310_49#_M1002_s N_A_310_49#_M1015_s N_A_310_49#_M1010_d
+ N_A_310_49#_M1020_d N_A_310_49#_c_1884_n N_A_310_49#_c_1885_n
+ N_A_310_49#_c_1886_n N_A_310_49#_c_1911_n N_A_310_49#_c_1887_n
+ N_A_310_49#_c_1929_n N_A_310_49#_c_1888_n N_A_310_49#_c_1889_n
+ N_A_310_49#_c_1938_n N_A_310_49#_c_1894_n N_A_310_49#_c_1890_n
+ N_A_310_49#_c_1891_n N_A_310_49#_c_1961_n N_A_310_49#_c_1895_n
+ N_A_310_49#_c_1943_n N_A_310_49#_c_1896_n N_A_310_49#_c_1975_n
+ N_A_310_49#_c_1897_n PM_SKY130_FD_SC_HD__FAH_1%A_310_49#
x_PM_SKY130_FD_SC_HD__FAH_1%A_1640_380# N_A_1640_380#_M1003_d
+ N_A_1640_380#_M1028_d N_A_1640_380#_M1019_s N_A_1640_380#_M1005_d
+ N_A_1640_380#_c_2063_n N_A_1640_380#_c_2057_n N_A_1640_380#_c_2058_n
+ N_A_1640_380#_c_2059_n N_A_1640_380#_c_2064_n N_A_1640_380#_c_2060_n
+ N_A_1640_380#_c_2094_n N_A_1640_380#_c_2083_n N_A_1640_380#_c_2061_n
+ N_A_1640_380#_c_2066_n N_A_1640_380#_c_2062_n
+ PM_SKY130_FD_SC_HD__FAH_1%A_1640_380#
x_PM_SKY130_FD_SC_HD__FAH_1%COUT N_COUT_M1011_s N_COUT_M1001_s N_COUT_c_2173_n
+ N_COUT_c_2175_n N_COUT_c_2174_n COUT COUT PM_SKY130_FD_SC_HD__FAH_1%COUT
x_PM_SKY130_FD_SC_HD__FAH_1%SUM N_SUM_M1017_d N_SUM_M1030_d SUM SUM SUM SUM SUM
+ SUM N_SUM_c_2213_n PM_SKY130_FD_SC_HD__FAH_1%SUM
x_PM_SKY130_FD_SC_HD__FAH_1%VGND N_VGND_M1029_d N_VGND_M1018_d N_VGND_M1024_d
+ N_VGND_M1011_d N_VGND_c_2228_n N_VGND_c_2229_n N_VGND_c_2230_n N_VGND_c_2231_n
+ N_VGND_c_2232_n N_VGND_c_2233_n N_VGND_c_2234_n N_VGND_c_2235_n
+ N_VGND_c_2236_n VGND N_VGND_c_2237_n N_VGND_c_2238_n N_VGND_c_2239_n
+ N_VGND_c_2240_n N_VGND_c_2241_n PM_SKY130_FD_SC_HD__FAH_1%VGND
cc_1 VNB N_A_67_199#_c_236_n 0.00473073f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.82
cc_2 VNB N_A_67_199#_c_237_n 0.00449106f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_3 VNB N_A_67_199#_c_238_n 0.00578488f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_4 VNB N_A_67_199#_c_239_n 0.025437f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_5 VNB N_A_67_199#_c_240_n 0.019934f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_6 VNB N_A_c_297_n 0.0220617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_c_298_n 0.0222126f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_8 VNB N_A_c_299_n 0.0104647f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.735
cc_9 VNB N_A_c_300_n 0.0456507f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_10 VNB N_A_c_301_n 0.00979158f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_11 VNB N_B_c_357_n 0.0214995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_358_n 0.0452407f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_B_c_359_n 0.0256266f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_14 VNB N_B_c_360_n 0.0203774f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_15 VNB N_B_c_361_n 0.0222625f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.16
cc_16 VNB N_B_c_362_n 0.0102087f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.63
cc_17 VNB N_B_c_363_n 0.00471789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_364_n 0.00161826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_c_365_n 0.0347984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_c_366_n 0.00351047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B_c_367_n 0.00189585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_508_297#_c_533_n 0.021089f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_508_297#_c_534_n 0.0224318f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_24 VNB N_A_508_297#_c_535_n 0.0101917f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_25 VNB N_A_508_297#_c_536_n 0.0450407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_508_297#_c_537_n 0.0127717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_508_297#_c_538_n 0.00175838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_508_297#_c_539_n 0.00115395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_508_297#_c_540_n 0.00223243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_719_47#_c_737_n 0.0193631f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_31 VNB N_A_719_47#_c_738_n 0.0181023f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.82
cc_32 VNB N_A_719_47#_c_739_n 0.0222884f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_33 VNB N_A_719_47#_c_740_n 0.00652134f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_34 VNB N_A_719_47#_M1016_g 0.0119097f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.16
cc_35 VNB N_A_719_47#_c_742_n 0.0267992f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_36 VNB N_A_719_47#_c_743_n 0.0119196f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.63
cc_37 VNB N_A_719_47#_c_744_n 0.0155494f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_38 VNB N_A_719_47#_c_745_n 0.00785073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_719_47#_c_746_n 0.00174703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_719_47#_c_747_n 0.0084749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_719_47#_c_748_n 0.00357305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_719_47#_c_749_n 5.8293e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_719_47#_c_750_n 0.00682565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_719_47#_c_751_n 9.48022e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_719_47#_c_752_n 0.00535186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_719_47#_c_753_n 0.0315789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1008_47#_c_958_n 0.0201133f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_48 VNB N_A_1008_47#_c_959_n 0.0202539f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.82
cc_49 VNB N_A_1008_47#_c_960_n 0.0136199f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_50 VNB N_A_1008_47#_c_961_n 0.0600698f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.63
cc_51 VNB N_A_1008_47#_c_962_n 5.47017e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1008_47#_c_963_n 0.00255102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1008_47#_c_964_n 0.00189971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1008_47#_c_965_n 0.00346724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_CI_c_1128_n 0.0291297f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_56 VNB N_CI_c_1129_n 0.0018411f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_57 VNB N_CI_c_1130_n 0.00122315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB CI 0.00253582f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_59 VNB N_CI_c_1132_n 0.01917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1262_49#_c_1195_n 0.00582653f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_61 VNB N_A_1262_49#_c_1196_n 0.0203425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1262_49#_c_1197_n 6.94034e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1262_49#_c_1198_n 0.0277155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1262_49#_c_1199_n 0.00325149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1262_49#_c_1200_n 0.00115013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1262_49#_c_1201_n 0.0203229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1332_297#_c_1369_n 7.89673e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.82
cc_68 VNB N_A_1332_297#_c_1370_n 0.00126719f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_69 VNB N_A_1332_297#_c_1371_n 0.0266084f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_70 VNB N_A_1332_297#_c_1372_n 4.97394e-19 $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.16
cc_71 VNB N_A_1332_297#_c_1373_n 0.0320391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1332_297#_c_1374_n 0.00278304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1332_297#_c_1375_n 0.0195123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1617_49#_c_1482_n 0.0192654f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_75 VNB N_A_1617_49#_c_1483_n 0.00331773f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_76 VNB N_A_1617_49#_c_1484_n 5.08649e-19 $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_77 VNB N_A_1617_49#_c_1485_n 0.0235286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1617_49#_c_1486_n 0.00334846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_27_47#_c_1601_n 0.0152202f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.16
cc_80 VNB N_A_27_47#_c_1602_n 0.00159198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_27_47#_c_1603_n 0.00666696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_27_47#_c_1604_n 0.0225868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_27_47#_c_1605_n 0.00941237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_27_47#_c_1606_n 0.00403606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VPWR_c_1769_n 0.516438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_310_49#_c_1884_n 0.00454299f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.16
cc_87 VNB N_A_310_49#_c_1885_n 5.7052e-19 $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.63
cc_88 VNB N_A_310_49#_c_1886_n 4.28853e-19 $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.63
cc_89 VNB N_A_310_49#_c_1887_n 0.00375033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_310_49#_c_1888_n 0.00657402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_310_49#_c_1889_n 0.00595273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_310_49#_c_1890_n 0.00246601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_310_49#_c_1891_n 0.00268537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1640_380#_c_2057_n 6.19416e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_1640_380#_c_2058_n 0.00283907f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.16
cc_96 VNB N_A_1640_380#_c_2059_n 0.00183067f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_97 VNB N_A_1640_380#_c_2060_n 0.00855279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1640_380#_c_2061_n 5.16421e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_1640_380#_c_2062_n 0.00835108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_COUT_c_2173_n 0.0115301f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_101 VNB N_COUT_c_2174_n 0.00951395f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_102 VNB SUM 0.0307748f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_103 VNB N_SUM_c_2213_n 0.0161344f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_104 VNB N_VGND_c_2228_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_105 VNB N_VGND_c_2229_n 0.0315531f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=0.38
cc_106 VNB N_VGND_c_2230_n 0.00481171f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.16
cc_107 VNB N_VGND_c_2231_n 0.00484319f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.63
cc_108 VNB N_VGND_c_2232_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2233_n 0.175669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2234_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2235_n 0.0356572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2236_n 0.00439458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2237_n 0.0177718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2238_n 0.017187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2239_n 0.614213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2240_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2241_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VPB N_A_67_199#_M1006_g 0.0234826f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_119 VPB N_A_67_199#_c_238_n 0.00938921f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_120 VPB N_A_67_199#_c_239_n 0.00589649f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_121 VPB N_A_M1007_g 0.023946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_M1015_g 0.0235498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_c_299_n 6.67008e-19 $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.735
cc_124 VPB N_A_c_300_n 0.0185897f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.38
cc_125 VPB N_A_c_301_n 6.96258e-19 $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.38
cc_126 VPB N_B_M1012_g 0.0236212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_B_c_358_n 0.0239136f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_128 VPB N_B_c_359_n 0.00754796f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_129 VPB N_B_M1023_g 0.0215662f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_130 VPB N_B_M1020_g 0.0365122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_B_c_362_n 7.14365e-19 $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.63
cc_132 VPB B 0.0010349f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_B_c_364_n 2.61637e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_B_c_365_n 0.0115596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_B_c_366_n 0.00271253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_B_c_367_n 0.00188957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_508_297#_M1010_g 0.0207219f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.38
cc_138 VPB N_A_508_297#_M1022_g 0.0218528f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.63
cc_139 VPB N_A_508_297#_c_535_n 7.12844e-19 $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.325
cc_140 VPB N_A_508_297#_c_536_n 0.023824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_508_297#_c_537_n 7.97857e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_508_297#_c_538_n 0.00185703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_508_297#_c_547_n 0.00146805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_508_297#_c_548_n 0.00504274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_508_297#_c_549_n 0.00912644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_508_297#_c_550_n 0.0014202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_508_297#_c_551_n 0.0156531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_508_297#_c_552_n 0.0034335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_508_297#_c_553_n 0.00756233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_508_297#_c_554_n 0.00663457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_508_297#_c_555_n 0.00590851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_719_47#_M1026_g 0.0232126f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_153 VPB N_A_719_47#_M1016_g 0.0286488f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.16
cc_154 VPB N_A_719_47#_c_742_n 0.0104235f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_155 VPB N_A_719_47#_c_743_n 0.00274674f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.63
cc_156 VPB N_A_719_47#_c_758_n 0.00285592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_719_47#_c_749_n 0.00136505f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_1008_47#_M1008_g 0.0216864f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_159 VPB N_A_1008_47#_c_967_n 0.0276163f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.38
cc_160 VPB N_A_1008_47#_c_968_n 0.017473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1008_47#_c_960_n 0.00264917f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_162 VPB N_A_1008_47#_c_961_n 0.0508096f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.63
cc_163 VPB N_A_1008_47#_c_971_n 0.00358662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_1008_47#_c_972_n 0.0329404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1008_47#_c_973_n 0.00224836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1008_47#_c_974_n 8.35121e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1008_47#_c_975_n 0.00360404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1008_47#_c_965_n 0.00167687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_CI_M1025_g 0.0226253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_CI_c_1128_n 0.00674174f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.325
cc_171 VPB N_CI_c_1129_n 3.68234e-19 $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_172 VPB N_A_1262_49#_M1005_g 0.0229075f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.16
cc_173 VPB N_A_1262_49#_c_1203_n 9.62191e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_1262_49#_c_1204_n 0.00790951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1262_49#_c_1205_n 0.0144673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1262_49#_c_1206_n 0.00401851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1262_49#_c_1197_n 0.00132556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1262_49#_c_1198_n 0.00624554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1262_49#_c_1200_n 0.00274162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1332_297#_M1001_g 0.0228117f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_181 VPB N_A_1332_297#_c_1377_n 0.00217356f $X=-0.19 $Y=1.305 $X2=1.155
+ $Y2=0.38
cc_182 VPB N_A_1332_297#_c_1373_n 0.00770164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1332_297#_c_1374_n 0.00110252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1617_49#_M1030_g 0.0220957f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_185 VPB N_A_1617_49#_c_1483_n 8.39611e-19 $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_186 VPB N_A_1617_49#_c_1489_n 8.32785e-19 $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_187 VPB N_A_1617_49#_c_1490_n 0.0178267f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.16
cc_188 VPB N_A_1617_49#_c_1491_n 5.76018e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_189 VPB N_A_1617_49#_c_1492_n 6.72297e-19 $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.325
cc_190 VPB N_A_1617_49#_c_1485_n 0.00581389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1617_49#_c_1486_n 0.00304809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1617_49#_c_1495_n 0.00129733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_27_47#_c_1607_n 0.00840926f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_194 VPB N_A_27_47#_c_1608_n 0.0158366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_27_47#_c_1609_n 0.00979517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_27_47#_c_1610_n 0.00296262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_27_47#_c_1611_n 0.02618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_27_47#_c_1612_n 7.80393e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_27_47#_c_1602_n 0.00205529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_27_47#_c_1614_n 0.00710642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_27_47#_c_1604_n 0.00908389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_27_47#_c_1616_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1770_n 0.00280515f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_204 VPB N_VPWR_c_1771_n 0.00295613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1772_n 4.89207e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_206 VPB N_VPWR_c_1773_n 0.00231609f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_207 VPB N_VPWR_c_1774_n 0.0164904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1775_n 0.03017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1776_n 0.170605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1777_n 0.0347372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1778_n 0.0170749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1769_n 0.105106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1780_n 0.00553667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1781_n 0.00522083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1782_n 0.00442675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1783_n 0.0036033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_310_49#_c_1885_n 0.006035f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.63
cc_218 VPB N_A_310_49#_c_1888_n 0.00670127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_310_49#_c_1894_n 0.00215183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_310_49#_c_1895_n 0.00362529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_310_49#_c_1896_n 0.00402196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_310_49#_c_1897_n 0.00510342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1640_380#_c_2063_n 0.00309006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1640_380#_c_2064_n 0.00766219f $X=-0.19 $Y=1.305 $X2=0.51
+ $Y2=1.16
cc_225 VPB N_A_1640_380#_c_2061_n 0.00520199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1640_380#_c_2066_n 0.00288509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1640_380#_c_2062_n 0.00715997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_COUT_c_2175_n 0.00430967f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.735
cc_229 VPB N_COUT_c_2174_n 0.00416321f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.38
cc_230 VPB COUT 0.0127784f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=0.38
cc_231 VPB SUM 0.0210468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_232 VPB SUM 0.00733941f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_233 VPB SUM 0.022004f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_234 N_A_67_199#_M1006_g N_A_M1007_g 0.0376908f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_67_199#_c_238_n N_A_M1007_g 0.013914f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_67_199#_c_236_n N_A_c_297_n 0.0107959f $X=0.99 $Y=0.82 $X2=0 $Y2=0
cc_237 N_A_67_199#_c_237_n N_A_c_297_n 0.00717571f $X=1.155 $Y=0.38 $X2=0 $Y2=0
cc_238 N_A_67_199#_c_238_n N_A_c_297_n 0.00214026f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_67_199#_c_240_n N_A_c_297_n 0.0190051f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_67_199#_c_236_n N_A_c_298_n 3.48092e-19 $X=0.99 $Y=0.82 $X2=0 $Y2=0
cc_241 N_A_67_199#_c_238_n N_A_c_299_n 0.00627521f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_67_199#_c_239_n N_A_c_299_n 0.0216279f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_67_199#_c_236_n N_A_c_300_n 0.00537066f $X=0.99 $Y=0.82 $X2=0 $Y2=0
cc_244 N_A_67_199#_c_238_n N_A_c_300_n 0.00507301f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_67_199#_c_236_n A 0.0294319f $X=0.99 $Y=0.82 $X2=0 $Y2=0
cc_246 N_A_67_199#_c_238_n A 0.0437161f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_67_199#_c_237_n N_A_27_47#_c_1601_n 0.00528965f $X=1.155 $Y=0.38
+ $X2=0 $Y2=0
cc_248 N_A_67_199#_c_240_n N_A_27_47#_c_1601_n 0.00494523f $X=0.495 $Y=0.995
+ $X2=0 $Y2=0
cc_249 N_A_67_199#_M1006_g N_A_27_47#_c_1607_n 0.00403188f $X=0.49 $Y=1.985
+ $X2=0 $Y2=0
cc_250 N_A_67_199#_M1007_d N_A_27_47#_c_1609_n 0.00640233f $X=1.015 $Y=1.485
+ $X2=0 $Y2=0
cc_251 N_A_67_199#_M1006_g N_A_27_47#_c_1609_n 0.00990848f $X=0.49 $Y=1.985
+ $X2=0 $Y2=0
cc_252 N_A_67_199#_c_238_n N_A_27_47#_c_1609_n 0.0393279f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_253 N_A_67_199#_c_239_n N_A_27_47#_c_1603_n 0.00125578f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_254 N_A_67_199#_c_240_n N_A_27_47#_c_1603_n 0.00395003f $X=0.495 $Y=0.995
+ $X2=0 $Y2=0
cc_255 N_A_67_199#_M1006_g N_A_27_47#_c_1614_n 0.00310888f $X=0.49 $Y=1.985
+ $X2=0 $Y2=0
cc_256 N_A_67_199#_c_238_n N_A_27_47#_c_1614_n 0.00438642f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_257 N_A_67_199#_c_239_n N_A_27_47#_c_1614_n 0.00224305f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_258 N_A_67_199#_M1006_g N_A_27_47#_c_1604_n 0.00265765f $X=0.49 $Y=1.985
+ $X2=0 $Y2=0
cc_259 N_A_67_199#_c_238_n N_A_27_47#_c_1604_n 0.0366692f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_260 N_A_67_199#_c_239_n N_A_27_47#_c_1604_n 0.00817554f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_261 N_A_67_199#_c_240_n N_A_27_47#_c_1604_n 0.002508f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_67_199#_M1006_g N_A_27_47#_c_1616_n 0.00112032f $X=0.49 $Y=1.985
+ $X2=0 $Y2=0
cc_263 N_A_67_199#_c_238_n N_VPWR_M1006_d 0.00295338f $X=0.51 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_264 N_A_67_199#_M1006_g N_VPWR_c_1770_n 0.00321262f $X=0.49 $Y=1.985 $X2=0
+ $Y2=0
cc_265 N_A_67_199#_M1006_g N_VPWR_c_1774_n 0.00427264f $X=0.49 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_A_67_199#_M1007_d N_VPWR_c_1769_n 0.00315303f $X=1.015 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_67_199#_M1006_g N_VPWR_c_1769_n 0.00665585f $X=0.49 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A_67_199#_c_237_n N_A_310_49#_c_1884_n 0.036834f $X=1.155 $Y=0.38 $X2=0
+ $Y2=0
cc_269 N_A_67_199#_c_238_n N_A_310_49#_c_1885_n 0.0231436f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_270 N_A_67_199#_c_236_n N_A_310_49#_c_1890_n 0.0151952f $X=0.99 $Y=0.82 $X2=0
+ $Y2=0
cc_271 N_A_67_199#_c_237_n N_A_310_49#_c_1890_n 0.00165876f $X=1.155 $Y=0.38
+ $X2=0 $Y2=0
cc_272 N_A_67_199#_c_236_n N_VGND_M1029_d 6.20362e-19 $X=0.99 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_273 N_A_67_199#_c_238_n N_VGND_M1029_d 0.0025199f $X=0.51 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_274 N_A_67_199#_c_237_n N_VGND_c_2228_n 0.0172577f $X=1.155 $Y=0.38 $X2=0
+ $Y2=0
cc_275 N_A_67_199#_c_238_n N_VGND_c_2228_n 0.0127321f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_67_199#_c_239_n N_VGND_c_2228_n 2.49941e-19 $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_277 N_A_67_199#_c_240_n N_VGND_c_2228_n 0.00276849f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_67_199#_c_236_n N_VGND_c_2229_n 0.00245983f $X=0.99 $Y=0.82 $X2=0
+ $Y2=0
cc_279 N_A_67_199#_c_237_n N_VGND_c_2229_n 0.0209752f $X=1.155 $Y=0.38 $X2=0
+ $Y2=0
cc_280 N_A_67_199#_c_238_n N_VGND_c_2229_n 2.28683e-19 $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_281 N_A_67_199#_c_240_n N_VGND_c_2237_n 0.00541359f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_67_199#_M1031_d N_VGND_c_2239_n 0.00209319f $X=1.02 $Y=0.235 $X2=0
+ $Y2=0
cc_283 N_A_67_199#_c_236_n N_VGND_c_2239_n 0.00486164f $X=0.99 $Y=0.82 $X2=0
+ $Y2=0
cc_284 N_A_67_199#_c_237_n N_VGND_c_2239_n 0.0124119f $X=1.155 $Y=0.38 $X2=0
+ $Y2=0
cc_285 N_A_67_199#_c_238_n N_VGND_c_2239_n 0.00121564f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_286 N_A_67_199#_c_240_n N_VGND_c_2239_n 0.0106124f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_M1015_g N_B_M1012_g 0.0290054f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A_c_298_n N_B_c_357_n 0.0136738f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_c_301_n N_B_c_359_n 0.0223327f $X=1.892 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_M1015_g B 0.00215184f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_c_301_n N_B_c_364_n 0.00445593f $X=1.892 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_c_301_n N_B_c_367_n 0.00250242f $X=1.892 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A_c_297_n N_A_27_47#_c_1601_n 5.86324e-19 $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_M1007_g N_A_27_47#_c_1609_n 0.0139841f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A_M1015_g N_A_27_47#_c_1609_n 0.0178369f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A_c_300_n N_A_27_47#_c_1609_n 0.00408214f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_297 A N_A_27_47#_c_1609_n 0.00337405f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_298 N_A_M1007_g N_A_27_47#_c_1614_n 0.00125857f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_M1007_g N_VPWR_c_1770_n 0.017204f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A_M1015_g N_VPWR_c_1771_n 0.00967141f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A_M1007_g N_VPWR_c_1775_n 0.00241817f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_302 N_A_M1015_g N_VPWR_c_1775_n 0.00428022f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A_M1007_g N_VPWR_c_1769_n 0.00442857f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A_M1015_g N_VPWR_c_1769_n 0.00763561f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A_c_298_n N_A_310_49#_c_1884_n 0.00647197f $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_A_M1007_g N_A_310_49#_c_1885_n 0.00205822f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A_c_297_n N_A_310_49#_c_1885_n 8.89572e-19 $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_c_298_n N_A_310_49#_c_1885_n 0.00378738f $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_M1015_g N_A_310_49#_c_1885_n 0.0066041f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_c_300_n N_A_310_49#_c_1885_n 0.0235234f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_c_301_n N_A_310_49#_c_1885_n 0.00351964f $X=1.892 $Y=1.16 $X2=0 $Y2=0
cc_312 A N_A_310_49#_c_1885_n 0.0139893f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_313 N_A_c_298_n N_A_310_49#_c_1886_n 0.0123227f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_c_298_n N_A_310_49#_c_1911_n 0.0013711f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A_c_297_n N_A_310_49#_c_1890_n 4.08403e-19 $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_c_298_n N_A_310_49#_c_1890_n 0.00178391f $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_c_300_n N_A_310_49#_c_1890_n 0.00363608f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_c_297_n N_VGND_c_2228_n 0.00374985f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_c_297_n N_VGND_c_2229_n 0.00424416f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_c_298_n N_VGND_c_2229_n 0.00414015f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_c_298_n N_VGND_c_2230_n 0.00300458f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_c_297_n N_VGND_c_2239_n 0.00734157f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_c_298_n N_VGND_c_2239_n 0.00746784f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B_c_360_n N_A_508_297#_c_533_n 0.0269232f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_325 N_B_M1023_g N_A_508_297#_M1010_g 0.0269232f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_326 N_B_c_361_n N_A_508_297#_c_534_n 0.010929f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B_M1020_g N_A_508_297#_M1022_g 0.0301633f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_328 N_B_c_362_n N_A_508_297#_c_535_n 0.0269232f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_329 N_B_c_363_n N_A_508_297#_c_535_n 0.00434948f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_330 N_B_c_363_n N_A_508_297#_c_536_n 0.00297979f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_331 N_B_c_363_n N_A_508_297#_c_537_n 0.00422577f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_332 N_B_c_365_n N_A_508_297#_c_537_n 0.0128937f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_333 N_B_M1012_g N_A_508_297#_c_538_n 0.00265384f $X=2.465 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_B_c_357_n N_A_508_297#_c_538_n 0.00425383f $X=2.565 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_B_c_358_n N_A_508_297#_c_538_n 0.0217688f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_336 N_B_c_397_p N_A_508_297#_c_538_n 0.0113805f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_337 N_B_c_363_n N_A_508_297#_c_538_n 0.0163206f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_338 N_B_c_364_n N_A_508_297#_c_538_n 8.1681e-19 $X=2.22 $Y=1.19 $X2=0 $Y2=0
cc_339 N_B_c_367_n N_A_508_297#_c_538_n 0.00492309f $X=2.09 $Y=1.175 $X2=0 $Y2=0
cc_340 N_B_M1012_g N_A_508_297#_c_548_n 0.0101487f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_341 N_B_c_359_n N_A_508_297#_c_548_n 0.0031993f $X=2.64 $Y=1.16 $X2=0 $Y2=0
cc_342 N_B_c_397_p N_A_508_297#_c_548_n 0.0083703f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_343 B N_A_508_297#_c_548_n 0.0102706f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_344 N_B_c_363_n N_A_508_297#_c_548_n 0.00207715f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_345 N_B_c_358_n N_A_508_297#_c_549_n 0.00511709f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_346 N_B_c_363_n N_A_508_297#_c_549_n 0.12617f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_347 N_B_M1012_g N_A_508_297#_c_550_n 0.00130903f $X=2.465 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_B_c_359_n N_A_508_297#_c_550_n 9.72169e-19 $X=2.64 $Y=1.16 $X2=0 $Y2=0
cc_349 N_B_c_397_p N_A_508_297#_c_550_n 5.50246e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_350 B N_A_508_297#_c_550_n 0.00224172f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_351 N_B_c_363_n N_A_508_297#_c_550_n 0.0269983f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_352 N_B_M1020_g N_A_508_297#_c_551_n 0.00641348f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_353 N_B_c_363_n N_A_508_297#_c_551_n 0.0803776f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_354 N_B_c_415_p N_A_508_297#_c_551_n 0.0265446f $X=5.765 $Y=1.19 $X2=0 $Y2=0
cc_355 N_B_c_365_n N_A_508_297#_c_551_n 0.00211522f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_356 N_B_c_366_n N_A_508_297#_c_551_n 0.00324777f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_357 N_B_c_363_n N_A_508_297#_c_552_n 0.0255102f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_358 N_B_M1020_g N_A_508_297#_c_553_n 0.0017367f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_359 N_B_c_362_n N_A_508_297#_c_554_n 7.91898e-19 $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_360 N_B_c_363_n N_A_508_297#_c_554_n 0.0208077f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_361 N_B_M1020_g N_A_508_297#_c_555_n 0.00259507f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_362 N_B_c_365_n N_A_719_47#_c_742_n 0.0182536f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_363 N_B_c_366_n N_A_719_47#_c_742_n 0.00194158f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_364 N_B_c_360_n N_A_719_47#_c_762_n 0.00554204f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_365 N_B_c_360_n N_A_719_47#_c_763_n 0.00260989f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_366 N_B_c_363_n N_A_719_47#_c_763_n 0.00174126f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_367 N_B_M1023_g N_A_719_47#_c_758_n 0.0137413f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_368 N_B_c_363_n N_A_719_47#_c_758_n 0.00365267f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_369 N_B_c_361_n N_A_719_47#_c_745_n 0.00608225f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_370 N_B_c_363_n N_A_719_47#_c_745_n 0.159786f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_371 N_B_c_415_p N_A_719_47#_c_745_n 0.0263847f $X=5.765 $Y=1.19 $X2=0 $Y2=0
cc_372 N_B_c_365_n N_A_719_47#_c_745_n 0.00195555f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_373 N_B_c_366_n N_A_719_47#_c_745_n 0.00294584f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_374 N_B_c_358_n N_A_719_47#_c_746_n 7.46445e-19 $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_375 N_B_c_360_n N_A_719_47#_c_746_n 6.74404e-19 $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_376 N_B_c_363_n N_A_719_47#_c_746_n 0.0260189f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_377 N_B_c_361_n N_A_719_47#_c_748_n 0.00197478f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_378 N_B_c_358_n N_A_719_47#_c_749_n 0.00592709f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_379 N_B_c_360_n N_A_719_47#_c_749_n 0.00696619f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_380 N_B_M1023_g N_A_719_47#_c_749_n 0.00515949f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_381 N_B_c_362_n N_A_719_47#_c_749_n 0.00673989f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_382 N_B_c_363_n N_A_719_47#_c_749_n 0.0110245f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_383 N_B_c_361_n N_A_719_47#_c_750_n 0.00407965f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_384 N_B_c_415_p N_A_719_47#_c_750_n 0.00148832f $X=5.765 $Y=1.19 $X2=0 $Y2=0
cc_385 N_B_c_365_n N_A_719_47#_c_750_n 8.94532e-19 $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_386 N_B_c_366_n N_A_719_47#_c_750_n 0.0203469f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_387 N_B_M1020_g N_A_1008_47#_c_971_n 0.0161157f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_388 N_B_c_363_n N_A_1008_47#_c_971_n 2.63373e-19 $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_389 N_B_c_366_n N_A_1008_47#_c_971_n 2.01658e-19 $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_390 N_B_M1020_g N_A_1008_47#_c_972_n 0.0122079f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_391 N_B_c_361_n N_A_1008_47#_c_962_n 0.00409168f $X=5.705 $Y=0.995 $X2=0
+ $Y2=0
cc_392 N_B_c_363_n N_A_1008_47#_c_962_n 4.24552e-19 $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_393 N_B_c_365_n N_A_1008_47#_c_962_n 7.43354e-19 $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_394 N_B_c_361_n N_A_1008_47#_c_963_n 9.71077e-19 $X=5.705 $Y=0.995 $X2=0
+ $Y2=0
cc_395 N_B_c_363_n N_A_1008_47#_c_963_n 0.00438276f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_396 N_B_c_415_p N_A_1008_47#_c_963_n 0.00117336f $X=5.765 $Y=1.19 $X2=0 $Y2=0
cc_397 N_B_c_365_n N_A_1008_47#_c_963_n 0.00662516f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_398 N_B_c_366_n N_A_1008_47#_c_963_n 0.0102629f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_399 N_B_c_363_n N_A_1008_47#_c_965_n 0.0131096f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_400 N_B_c_415_p N_A_1008_47#_c_965_n 0.00119585f $X=5.765 $Y=1.19 $X2=0 $Y2=0
cc_401 N_B_c_365_n N_A_1008_47#_c_965_n 0.00678943f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_402 N_B_c_366_n N_A_1008_47#_c_965_n 0.0110529f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_403 N_B_c_361_n N_A_1262_49#_c_1199_n 5.09174e-19 $X=5.705 $Y=0.995 $X2=0
+ $Y2=0
cc_404 N_B_M1012_g N_A_27_47#_c_1609_n 0.0137507f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_405 N_B_c_358_n N_A_27_47#_c_1609_n 4.94926e-19 $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_406 N_B_c_359_n N_A_27_47#_c_1609_n 0.00266837f $X=2.64 $Y=1.16 $X2=0 $Y2=0
cc_407 N_B_M1023_g N_A_27_47#_c_1609_n 5.01419e-19 $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_408 N_B_c_397_p N_A_27_47#_c_1609_n 0.00361677f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_409 B N_A_27_47#_c_1609_n 0.012441f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_410 N_B_c_364_n N_A_27_47#_c_1609_n 0.00295284f $X=2.22 $Y=1.19 $X2=0 $Y2=0
cc_411 N_B_M1012_g N_A_27_47#_c_1610_n 0.00760191f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_412 N_B_M1023_g N_A_27_47#_c_1610_n 0.00376126f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_413 N_B_M1023_g N_A_27_47#_c_1611_n 0.0120506f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_414 N_B_M1012_g N_A_27_47#_c_1649_n 0.00394612f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_415 N_B_c_363_n N_A_27_47#_c_1602_n 0.0113527f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_416 N_B_c_365_n N_A_27_47#_c_1602_n 3.12132e-19 $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_417 N_B_c_361_n N_A_27_47#_c_1652_n 0.00153536f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_418 N_B_c_361_n N_A_27_47#_c_1653_n 0.00938736f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_419 N_B_c_365_n N_A_27_47#_c_1653_n 0.00252609f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_420 N_B_c_366_n N_A_27_47#_c_1653_n 8.20847e-19 $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_421 N_B_c_363_n N_A_27_47#_c_1605_n 0.0121232f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_422 N_B_c_361_n N_A_27_47#_c_1606_n 0.00533994f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_423 N_B_c_365_n N_A_27_47#_c_1606_n 5.06281e-19 $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_424 N_B_c_366_n N_A_27_47#_c_1606_n 0.0025959f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_425 B N_VPWR_M1015_d 0.00571503f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_426 N_B_M1012_g N_VPWR_c_1771_n 0.00761866f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_427 N_B_M1012_g N_VPWR_c_1776_n 0.00413026f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_428 N_B_M1023_g N_VPWR_c_1776_n 9.44495e-19 $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_429 N_B_M1020_g N_VPWR_c_1776_n 0.00335164f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_430 N_B_M1012_g N_VPWR_c_1769_n 0.0061246f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_431 N_B_M1020_g N_VPWR_c_1769_n 0.00686384f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_432 N_B_c_357_n N_A_310_49#_c_1885_n 3.70633e-19 $X=2.565 $Y=0.995 $X2=0
+ $Y2=0
cc_433 N_B_c_359_n N_A_310_49#_c_1885_n 4.45154e-19 $X=2.64 $Y=1.16 $X2=0 $Y2=0
cc_434 B N_A_310_49#_c_1885_n 0.00521252f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_435 N_B_c_364_n N_A_310_49#_c_1885_n 0.00671803f $X=2.22 $Y=1.19 $X2=0 $Y2=0
cc_436 N_B_c_367_n N_A_310_49#_c_1885_n 0.0226508f $X=2.09 $Y=1.175 $X2=0 $Y2=0
cc_437 N_B_c_357_n N_A_310_49#_c_1886_n 0.00569f $X=2.565 $Y=0.995 $X2=0 $Y2=0
cc_438 N_B_c_359_n N_A_310_49#_c_1886_n 0.00752215f $X=2.64 $Y=1.16 $X2=0 $Y2=0
cc_439 N_B_c_397_p N_A_310_49#_c_1886_n 0.0167607f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_440 N_B_c_363_n N_A_310_49#_c_1886_n 0.00262634f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_441 N_B_c_364_n N_A_310_49#_c_1886_n 0.00482262f $X=2.22 $Y=1.19 $X2=0 $Y2=0
cc_442 N_B_c_367_n N_A_310_49#_c_1886_n 0.0110728f $X=2.09 $Y=1.175 $X2=0 $Y2=0
cc_443 N_B_c_357_n N_A_310_49#_c_1911_n 0.00798792f $X=2.565 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_B_c_357_n N_A_310_49#_c_1887_n 0.0122179f $X=2.565 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_358_n N_A_310_49#_c_1887_n 0.0046212f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_446 N_B_c_357_n N_A_310_49#_c_1929_n 0.0027342f $X=2.565 $Y=0.995 $X2=0 $Y2=0
cc_447 N_B_M1012_g N_A_310_49#_c_1888_n 0.0038286f $X=2.465 $Y=1.985 $X2=0 $Y2=0
cc_448 N_B_c_357_n N_A_310_49#_c_1888_n 0.00241694f $X=2.565 $Y=0.995 $X2=0
+ $Y2=0
cc_449 N_B_c_358_n N_A_310_49#_c_1888_n 0.0207424f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_450 N_B_c_360_n N_A_310_49#_c_1888_n 0.00575478f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_451 N_B_M1023_g N_A_310_49#_c_1888_n 0.00799567f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_452 N_B_c_363_n N_A_310_49#_c_1888_n 0.0168314f $X=5.62 $Y=1.19 $X2=0 $Y2=0
cc_453 N_B_c_358_n N_A_310_49#_c_1889_n 0.00407611f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_454 N_B_c_360_n N_A_310_49#_c_1889_n 0.00859636f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_455 N_B_c_358_n N_A_310_49#_c_1938_n 0.00360667f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_456 N_B_M1023_g N_A_310_49#_c_1938_n 0.0119888f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_457 N_B_M1012_g N_A_310_49#_c_1894_n 6.41871e-19 $X=2.465 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_B_c_357_n N_A_310_49#_c_1891_n 7.51894e-19 $X=2.565 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_B_M1020_g N_A_310_49#_c_1895_n 0.00221459f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_460 N_B_M1023_g N_A_310_49#_c_1943_n 8.19423e-19 $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_461 N_B_M1023_g N_A_310_49#_c_1896_n 0.00148651f $X=3.52 $Y=1.905 $X2=0 $Y2=0
cc_462 N_B_M1020_g N_A_310_49#_c_1897_n 0.0071488f $X=5.485 $Y=2.03 $X2=0 $Y2=0
cc_463 N_B_c_365_n N_A_310_49#_c_1897_n 0.00426611f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_464 N_B_c_366_n N_A_310_49#_c_1897_n 0.00437575f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_465 N_B_c_357_n N_VGND_c_2230_n 0.00302765f $X=2.565 $Y=0.995 $X2=0 $Y2=0
cc_466 N_B_c_357_n N_VGND_c_2233_n 0.00357835f $X=2.565 $Y=0.995 $X2=0 $Y2=0
cc_467 N_B_c_360_n N_VGND_c_2233_n 0.00357877f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_468 N_B_c_361_n N_VGND_c_2233_n 0.00352679f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_469 N_B_c_357_n N_VGND_c_2239_n 0.00726199f $X=2.565 $Y=0.995 $X2=0 $Y2=0
cc_470 N_B_c_360_n N_VGND_c_2239_n 0.00649167f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_471 N_B_c_361_n N_VGND_c_2239_n 0.00697496f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_472 N_A_508_297#_c_549_n N_A_719_47#_M1023_d 5.23922e-19 $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_473 N_A_508_297#_c_595_p N_A_719_47#_M1026_g 0.0160825f $X=7.05 $Y=2.04 $X2=0
+ $Y2=0
cc_474 N_A_508_297#_c_547_n N_A_719_47#_M1026_g 5.91045e-19 $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_475 N_A_508_297#_c_553_n N_A_719_47#_M1026_g 7.5634e-19 $X=6.235 $Y=1.53
+ $X2=0 $Y2=0
cc_476 N_A_508_297#_c_555_n N_A_719_47#_M1026_g 9.30889e-19 $X=6.375 $Y=1.53
+ $X2=0 $Y2=0
cc_477 N_A_508_297#_c_553_n N_A_719_47#_c_742_n 0.00450943f $X=6.235 $Y=1.53
+ $X2=0 $Y2=0
cc_478 N_A_508_297#_c_555_n N_A_719_47#_c_742_n 0.00802782f $X=6.375 $Y=1.53
+ $X2=0 $Y2=0
cc_479 N_A_508_297#_c_533_n N_A_719_47#_c_763_n 0.00316543f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_480 N_A_508_297#_M1010_g N_A_719_47#_c_758_n 4.39035e-19 $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_481 N_A_508_297#_c_549_n N_A_719_47#_c_758_n 0.0192201f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_482 N_A_508_297#_c_552_n N_A_719_47#_c_758_n 0.00126168f $X=4.595 $Y=1.53
+ $X2=0 $Y2=0
cc_483 N_A_508_297#_c_554_n N_A_719_47#_c_758_n 0.00430772f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_484 N_A_508_297#_c_533_n N_A_719_47#_c_745_n 0.00535763f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_485 N_A_508_297#_c_536_n N_A_719_47#_c_745_n 0.00601333f $X=4.89 $Y=1.16
+ $X2=0 $Y2=0
cc_486 N_A_508_297#_c_551_n N_A_719_47#_c_745_n 0.00881115f $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_487 N_A_508_297#_c_554_n N_A_719_47#_c_745_n 0.00271844f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_488 N_A_508_297#_c_533_n N_A_719_47#_c_746_n 6.37996e-19 $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_489 N_A_508_297#_M1021_d N_A_719_47#_c_747_n 9.13112e-19 $X=7.145 $Y=0.245
+ $X2=0 $Y2=0
cc_490 N_A_508_297#_c_539_n N_A_719_47#_c_747_n 0.0124714f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_491 N_A_508_297#_c_540_n N_A_719_47#_c_747_n 0.00666967f $X=7.28 $Y=0.68
+ $X2=0 $Y2=0
cc_492 N_A_508_297#_c_555_n N_A_719_47#_c_747_n 0.00104218f $X=6.375 $Y=1.53
+ $X2=0 $Y2=0
cc_493 N_A_508_297#_c_553_n N_A_719_47#_c_748_n 0.0151797f $X=6.235 $Y=1.53
+ $X2=0 $Y2=0
cc_494 N_A_508_297#_c_555_n N_A_719_47#_c_748_n 2.10012e-19 $X=6.375 $Y=1.53
+ $X2=0 $Y2=0
cc_495 N_A_508_297#_c_533_n N_A_719_47#_c_749_n 0.00300604f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_496 N_A_508_297#_c_549_n N_A_719_47#_c_749_n 0.00119423f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_497 N_A_508_297#_c_554_n N_A_719_47#_c_749_n 0.00939663f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_498 N_A_508_297#_c_553_n N_A_719_47#_c_750_n 0.00305584f $X=6.235 $Y=1.53
+ $X2=0 $Y2=0
cc_499 N_A_508_297#_c_555_n N_A_719_47#_c_750_n 0.0228485f $X=6.375 $Y=1.53
+ $X2=0 $Y2=0
cc_500 N_A_508_297#_c_551_n N_A_1008_47#_M1022_d 8.14763e-19 $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_501 N_A_508_297#_c_595_p N_A_1008_47#_M1008_g 0.01446f $X=7.05 $Y=2.04 $X2=0
+ $Y2=0
cc_502 N_A_508_297#_c_547_n N_A_1008_47#_M1008_g 0.0187496f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_503 N_A_508_297#_c_539_n N_A_1008_47#_c_958_n 0.00434065f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_504 N_A_508_297#_c_540_n N_A_1008_47#_c_958_n 0.00237431f $X=7.28 $Y=0.68
+ $X2=0 $Y2=0
cc_505 N_A_508_297#_c_539_n N_A_1008_47#_c_959_n 6.56313e-19 $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_506 N_A_508_297#_c_547_n N_A_1008_47#_c_960_n 0.00382338f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_507 N_A_508_297#_c_539_n N_A_1008_47#_c_960_n 0.0042083f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_508 N_A_508_297#_c_547_n N_A_1008_47#_c_961_n 0.00463605f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_509 N_A_508_297#_c_539_n N_A_1008_47#_c_961_n 0.00631949f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_510 N_A_508_297#_c_540_n N_A_1008_47#_c_961_n 0.00541353f $X=7.28 $Y=0.68
+ $X2=0 $Y2=0
cc_511 N_A_508_297#_c_537_n N_A_1008_47#_c_971_n 0.00401729f $X=4.982 $Y=1.16
+ $X2=0 $Y2=0
cc_512 N_A_508_297#_c_551_n N_A_1008_47#_c_971_n 0.0131883f $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_513 N_A_508_297#_M1026_s N_A_1008_47#_c_972_n 0.00517659f $X=6.205 $Y=1.485
+ $X2=0 $Y2=0
cc_514 N_A_508_297#_c_595_p N_A_1008_47#_c_972_n 0.0362681f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_515 N_A_508_297#_c_637_p N_A_1008_47#_c_972_n 0.0121511f $X=6.46 $Y=2.04
+ $X2=0 $Y2=0
cc_516 N_A_508_297#_M1022_g N_A_1008_47#_c_973_n 0.00116158f $X=5 $Y=1.905 $X2=0
+ $Y2=0
cc_517 N_A_508_297#_c_534_n N_A_1008_47#_c_962_n 9.00239e-19 $X=4.965 $Y=0.995
+ $X2=0 $Y2=0
cc_518 N_A_508_297#_c_534_n N_A_1008_47#_c_963_n 6.49711e-19 $X=4.965 $Y=0.995
+ $X2=0 $Y2=0
cc_519 N_A_508_297#_c_537_n N_A_1008_47#_c_963_n 0.00135233f $X=4.982 $Y=1.16
+ $X2=0 $Y2=0
cc_520 N_A_508_297#_c_595_p N_A_1008_47#_c_974_n 0.0138309f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_521 N_A_508_297#_c_547_n N_A_1008_47#_c_974_n 0.0385813f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_522 N_A_508_297#_c_547_n N_A_1008_47#_c_975_n 0.0111211f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_523 N_A_508_297#_c_540_n N_A_1008_47#_c_975_n 7.42397e-19 $X=7.28 $Y=0.68
+ $X2=0 $Y2=0
cc_524 N_A_508_297#_c_547_n N_A_1008_47#_c_964_n 0.00464869f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_525 N_A_508_297#_c_539_n N_A_1008_47#_c_964_n 0.0115864f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_526 N_A_508_297#_c_537_n N_A_1008_47#_c_965_n 0.00165366f $X=4.982 $Y=1.16
+ $X2=0 $Y2=0
cc_527 N_A_508_297#_c_551_n N_A_1008_47#_c_965_n 0.00500126f $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_528 N_A_508_297#_c_595_p N_A_1262_49#_M1008_d 0.0027538f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_529 N_A_508_297#_c_547_n N_A_1262_49#_M1008_d 0.00499771f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_530 N_A_508_297#_M1021_d N_A_1262_49#_c_1195_n 0.00455419f $X=7.145 $Y=0.245
+ $X2=0 $Y2=0
cc_531 N_A_508_297#_c_539_n N_A_1262_49#_c_1195_n 6.31887e-19 $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_532 N_A_508_297#_c_540_n N_A_1262_49#_c_1195_n 0.0177614f $X=7.28 $Y=0.68
+ $X2=0 $Y2=0
cc_533 N_A_508_297#_c_540_n N_A_1262_49#_c_1216_n 0.00996058f $X=7.28 $Y=0.68
+ $X2=0 $Y2=0
cc_534 N_A_508_297#_c_539_n N_A_1262_49#_c_1217_n 0.0016936f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_535 N_A_508_297#_c_539_n N_A_1262_49#_c_1200_n 0.00453329f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_536 N_A_508_297#_c_595_p N_A_1332_297#_M1026_d 0.00321262f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_537 N_A_508_297#_c_539_n N_A_1332_297#_c_1369_n 0.00861527f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_538 N_A_508_297#_c_539_n N_A_1332_297#_c_1370_n 0.0163078f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_539 N_A_508_297#_c_595_p N_A_1332_297#_c_1377_n 0.0126919f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_540 N_A_508_297#_c_553_n N_A_1332_297#_c_1377_n 0.00246917f $X=6.235 $Y=1.53
+ $X2=0 $Y2=0
cc_541 N_A_508_297#_c_555_n N_A_1332_297#_c_1377_n 0.00205581f $X=6.375 $Y=1.53
+ $X2=0 $Y2=0
cc_542 N_A_508_297#_c_547_n N_A_1332_297#_c_1371_n 0.0123499f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_543 N_A_508_297#_c_539_n N_A_1332_297#_c_1371_n 0.00622931f $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_544 N_A_508_297#_c_547_n N_A_1332_297#_c_1388_n 2.80315e-19 $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_545 N_A_508_297#_c_539_n N_A_1332_297#_c_1388_n 2.91774e-19 $X=7.195 $Y=1.01
+ $X2=0 $Y2=0
cc_546 N_A_508_297#_c_547_n N_A_1332_297#_c_1372_n 0.0316923f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_547 N_A_508_297#_c_549_n N_A_27_47#_M1023_s 0.00168051f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_548 N_A_508_297#_c_551_n N_A_27_47#_M1022_s 0.00139415f $X=6.09 $Y=1.53 $X2=0
+ $Y2=0
cc_549 N_A_508_297#_M1012_d N_A_27_47#_c_1609_n 0.00331642f $X=2.54 $Y=1.485
+ $X2=0 $Y2=0
cc_550 N_A_508_297#_c_548_n N_A_27_47#_c_1609_n 0.0246875f $X=2.69 $Y=1.58 $X2=0
+ $Y2=0
cc_551 N_A_508_297#_c_549_n N_A_27_47#_c_1609_n 8.01532e-19 $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_552 N_A_508_297#_c_550_n N_A_27_47#_c_1609_n 0.00179344f $X=2.68 $Y=1.53
+ $X2=0 $Y2=0
cc_553 N_A_508_297#_M1012_d N_A_27_47#_c_1610_n 0.0036772f $X=2.54 $Y=1.485
+ $X2=0 $Y2=0
cc_554 N_A_508_297#_M1010_g N_A_27_47#_c_1611_n 0.0120107f $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_555 N_A_508_297#_c_548_n N_A_27_47#_c_1611_n 0.00195927f $X=2.69 $Y=1.58
+ $X2=0 $Y2=0
cc_556 N_A_508_297#_M1012_d N_A_27_47#_c_1649_n 0.00482075f $X=2.54 $Y=1.485
+ $X2=0 $Y2=0
cc_557 N_A_508_297#_M1022_g N_A_27_47#_c_1612_n 0.00634093f $X=5 $Y=1.905 $X2=0
+ $Y2=0
cc_558 N_A_508_297#_c_533_n N_A_27_47#_c_1602_n 0.00139071f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_559 N_A_508_297#_M1010_g N_A_27_47#_c_1602_n 0.00642871f $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_560 N_A_508_297#_c_534_n N_A_27_47#_c_1602_n 0.0018622f $X=4.965 $Y=0.995
+ $X2=0 $Y2=0
cc_561 N_A_508_297#_M1022_g N_A_27_47#_c_1602_n 0.012964f $X=5 $Y=1.905 $X2=0
+ $Y2=0
cc_562 N_A_508_297#_c_536_n N_A_27_47#_c_1602_n 0.0207132f $X=4.89 $Y=1.16 $X2=0
+ $Y2=0
cc_563 N_A_508_297#_c_551_n N_A_27_47#_c_1602_n 0.0111644f $X=6.09 $Y=1.53 $X2=0
+ $Y2=0
cc_564 N_A_508_297#_c_552_n N_A_27_47#_c_1602_n 0.00339125f $X=4.595 $Y=1.53
+ $X2=0 $Y2=0
cc_565 N_A_508_297#_c_554_n N_A_27_47#_c_1602_n 0.0360565f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_566 N_A_508_297#_c_534_n N_A_27_47#_c_1652_n 0.00725862f $X=4.965 $Y=0.995
+ $X2=0 $Y2=0
cc_567 N_A_508_297#_c_534_n N_A_27_47#_c_1680_n 0.00539843f $X=4.965 $Y=0.995
+ $X2=0 $Y2=0
cc_568 N_A_508_297#_c_533_n N_A_27_47#_c_1605_n 0.00563716f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_569 N_A_508_297#_c_534_n N_A_27_47#_c_1605_n 0.0193615f $X=4.965 $Y=0.995
+ $X2=0 $Y2=0
cc_570 N_A_508_297#_c_536_n N_A_27_47#_c_1605_n 0.017666f $X=4.89 $Y=1.16 $X2=0
+ $Y2=0
cc_571 N_A_508_297#_c_537_n N_A_27_47#_c_1605_n 0.00187305f $X=4.982 $Y=1.16
+ $X2=0 $Y2=0
cc_572 N_A_508_297#_c_554_n N_A_27_47#_c_1605_n 0.0289067f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_573 N_A_508_297#_M1010_g N_VPWR_c_1776_n 9.44495e-19 $X=3.945 $Y=1.905 $X2=0
+ $Y2=0
cc_574 N_A_508_297#_M1022_g N_VPWR_c_1776_n 0.00482137f $X=5 $Y=1.905 $X2=0
+ $Y2=0
cc_575 N_A_508_297#_M1012_d N_VPWR_c_1769_n 0.00247534f $X=2.54 $Y=1.485 $X2=0
+ $Y2=0
cc_576 N_A_508_297#_M1022_g N_VPWR_c_1769_n 0.00318289f $X=5 $Y=1.905 $X2=0
+ $Y2=0
cc_577 N_A_508_297#_c_549_n N_A_310_49#_M1010_d 2.223e-19 $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_578 N_A_508_297#_c_554_n N_A_310_49#_M1010_d 0.00318459f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_579 N_A_508_297#_c_548_n N_A_310_49#_c_1886_n 3.21698e-19 $X=2.69 $Y=1.58
+ $X2=0 $Y2=0
cc_580 N_A_508_297#_M1000_d N_A_310_49#_c_1887_n 0.00456566f $X=2.64 $Y=0.235
+ $X2=0 $Y2=0
cc_581 N_A_508_297#_c_538_n N_A_310_49#_c_1887_n 0.0123437f $X=2.775 $Y=0.76
+ $X2=0 $Y2=0
cc_582 N_A_508_297#_M1010_g N_A_310_49#_c_1888_n 2.02818e-19 $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_583 N_A_508_297#_c_538_n N_A_310_49#_c_1888_n 0.0598458f $X=2.775 $Y=0.76
+ $X2=0 $Y2=0
cc_584 N_A_508_297#_c_548_n N_A_310_49#_c_1888_n 0.0205524f $X=2.69 $Y=1.58
+ $X2=0 $Y2=0
cc_585 N_A_508_297#_c_549_n N_A_310_49#_c_1888_n 0.0162999f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_586 N_A_508_297#_c_550_n N_A_310_49#_c_1888_n 3.77776e-19 $X=2.68 $Y=1.53
+ $X2=0 $Y2=0
cc_587 N_A_508_297#_c_533_n N_A_310_49#_c_1889_n 0.0141448f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_588 N_A_508_297#_M1010_g N_A_310_49#_c_1938_n 0.00822917f $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_589 N_A_508_297#_c_549_n N_A_310_49#_c_1938_n 0.0129773f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_590 N_A_508_297#_c_533_n N_A_310_49#_c_1961_n 0.00299875f $X=3.945 $Y=0.995
+ $X2=0 $Y2=0
cc_591 N_A_508_297#_c_536_n N_A_310_49#_c_1961_n 5.09382e-19 $X=4.89 $Y=1.16
+ $X2=0 $Y2=0
cc_592 N_A_508_297#_M1022_g N_A_310_49#_c_1895_n 0.00681165f $X=5 $Y=1.905 $X2=0
+ $Y2=0
cc_593 N_A_508_297#_c_549_n N_A_310_49#_c_1895_n 0.00657534f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_594 N_A_508_297#_c_551_n N_A_310_49#_c_1895_n 0.0716911f $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_595 N_A_508_297#_c_552_n N_A_310_49#_c_1895_n 0.0278905f $X=4.595 $Y=1.53
+ $X2=0 $Y2=0
cc_596 N_A_508_297#_c_554_n N_A_310_49#_c_1895_n 0.00185487f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_597 N_A_508_297#_M1010_g N_A_310_49#_c_1943_n 0.00445969f $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_598 N_A_508_297#_c_549_n N_A_310_49#_c_1943_n 0.0268239f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_599 N_A_508_297#_c_554_n N_A_310_49#_c_1943_n 9.93033e-19 $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_600 N_A_508_297#_M1010_g N_A_310_49#_c_1896_n 0.00722633f $X=3.945 $Y=1.905
+ $X2=0 $Y2=0
cc_601 N_A_508_297#_c_536_n N_A_310_49#_c_1896_n 7.60146e-19 $X=4.89 $Y=1.16
+ $X2=0 $Y2=0
cc_602 N_A_508_297#_c_549_n N_A_310_49#_c_1896_n 0.00136998f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_603 N_A_508_297#_c_554_n N_A_310_49#_c_1896_n 0.0171065f $X=4.235 $Y=1.16
+ $X2=0 $Y2=0
cc_604 N_A_508_297#_c_726_p N_A_310_49#_c_1975_n 0.00116733f $X=6.375 $Y=1.62
+ $X2=0 $Y2=0
cc_605 N_A_508_297#_c_637_p N_A_310_49#_c_1975_n 2.13547e-19 $X=6.46 $Y=2.04
+ $X2=0 $Y2=0
cc_606 N_A_508_297#_c_551_n N_A_310_49#_c_1975_n 0.0262329f $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_607 N_A_508_297#_c_726_p N_A_310_49#_c_1897_n 0.009387f $X=6.375 $Y=1.62
+ $X2=0 $Y2=0
cc_608 N_A_508_297#_c_637_p N_A_310_49#_c_1897_n 0.00320248f $X=6.46 $Y=2.04
+ $X2=0 $Y2=0
cc_609 N_A_508_297#_c_551_n N_A_310_49#_c_1897_n 0.00903048f $X=6.09 $Y=1.53
+ $X2=0 $Y2=0
cc_610 N_A_508_297#_c_533_n N_VGND_c_2233_n 0.00357877f $X=3.945 $Y=0.995 $X2=0
+ $Y2=0
cc_611 N_A_508_297#_c_534_n N_VGND_c_2233_n 0.00421297f $X=4.965 $Y=0.995 $X2=0
+ $Y2=0
cc_612 N_A_508_297#_M1000_d N_VGND_c_2239_n 0.00201948f $X=2.64 $Y=0.235 $X2=0
+ $Y2=0
cc_613 N_A_508_297#_c_533_n N_VGND_c_2239_n 0.00662925f $X=3.945 $Y=0.995 $X2=0
+ $Y2=0
cc_614 N_A_508_297#_c_534_n N_VGND_c_2239_n 0.00760426f $X=4.965 $Y=0.995 $X2=0
+ $Y2=0
cc_615 N_A_719_47#_c_745_n N_A_1008_47#_M1002_d 0.00239794f $X=6.09 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_616 N_A_719_47#_M1026_g N_A_1008_47#_M1008_g 0.036343f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_617 N_A_719_47#_c_737_n N_A_1008_47#_c_958_n 0.0262742f $X=6.645 $Y=0.995
+ $X2=0 $Y2=0
cc_618 N_A_719_47#_c_747_n N_A_1008_47#_c_958_n 0.00235448f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_619 N_A_719_47#_c_738_n N_A_1008_47#_c_959_n 0.0247411f $X=8.45 $Y=0.96 $X2=0
+ $Y2=0
cc_620 N_A_719_47#_c_747_n N_A_1008_47#_c_959_n 0.00282219f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_621 N_A_719_47#_c_740_n N_A_1008_47#_c_967_n 0.0141772f $X=8.525 $Y=1.035
+ $X2=0 $Y2=0
cc_622 N_A_719_47#_M1016_g N_A_1008_47#_c_967_n 0.0428165f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_623 N_A_719_47#_c_743_n N_A_1008_47#_c_960_n 0.0221166f $X=6.615 $Y=1.16
+ $X2=0 $Y2=0
cc_624 N_A_719_47#_c_747_n N_A_1008_47#_c_960_n 0.00110819f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_625 N_A_719_47#_c_740_n N_A_1008_47#_c_961_n 0.00755358f $X=8.525 $Y=1.035
+ $X2=0 $Y2=0
cc_626 N_A_719_47#_M1016_g N_A_1008_47#_c_961_n 0.00266609f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_627 N_A_719_47#_c_747_n N_A_1008_47#_c_961_n 0.0068725f $X=8.86 $Y=0.85 $X2=0
+ $Y2=0
cc_628 N_A_719_47#_M1026_g N_A_1008_47#_c_972_n 0.012022f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_629 N_A_719_47#_c_745_n N_A_1008_47#_c_962_n 0.0137231f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_630 N_A_719_47#_c_748_n N_A_1008_47#_c_962_n 0.00116274f $X=6.38 $Y=0.85
+ $X2=0 $Y2=0
cc_631 N_A_719_47#_c_750_n N_A_1008_47#_c_962_n 0.00318188f $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_632 N_A_719_47#_c_748_n N_A_1008_47#_c_963_n 8.72058e-19 $X=6.38 $Y=0.85
+ $X2=0 $Y2=0
cc_633 N_A_719_47#_c_750_n N_A_1008_47#_c_963_n 0.00168529f $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_634 N_A_719_47#_c_747_n N_A_1008_47#_c_964_n 0.00251559f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_635 N_A_719_47#_c_745_n N_A_1008_47#_c_965_n 0.00122832f $X=6.09 $Y=0.85
+ $X2=0 $Y2=0
cc_636 N_A_719_47#_M1016_g N_CI_M1025_g 0.0117779f $X=8.955 $Y=1.995 $X2=0 $Y2=0
cc_637 N_A_719_47#_c_744_n N_CI_c_1128_n 0.0111111f $X=8.88 $Y=0.96 $X2=0 $Y2=0
cc_638 N_A_719_47#_c_744_n N_CI_c_1129_n 0.00102903f $X=8.88 $Y=0.96 $X2=0 $Y2=0
cc_639 N_A_719_47#_c_744_n N_CI_c_1130_n 4.19788e-19 $X=8.88 $Y=0.96 $X2=0 $Y2=0
cc_640 N_A_719_47#_c_751_n N_CI_c_1130_n 9.09351e-19 $X=9.005 $Y=0.85 $X2=0
+ $Y2=0
cc_641 N_A_719_47#_c_753_n N_CI_c_1130_n 0.00103451f $X=9.12 $Y=0.77 $X2=0 $Y2=0
cc_642 N_A_719_47#_c_751_n CI 0.00112253f $X=9.005 $Y=0.85 $X2=0 $Y2=0
cc_643 N_A_719_47#_c_752_n CI 0.00555861f $X=9.005 $Y=0.85 $X2=0 $Y2=0
cc_644 N_A_719_47#_c_753_n CI 2.8322e-19 $X=9.12 $Y=0.77 $X2=0 $Y2=0
cc_645 N_A_719_47#_c_752_n N_CI_c_1132_n 0.00183115f $X=9.005 $Y=0.85 $X2=0
+ $Y2=0
cc_646 N_A_719_47#_c_753_n N_CI_c_1132_n 0.00958846f $X=9.12 $Y=0.77 $X2=0 $Y2=0
cc_647 N_A_719_47#_c_747_n N_A_1262_49#_M1004_s 9.92452e-19 $X=8.86 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_648 N_A_719_47#_c_748_n N_A_1262_49#_M1004_s 5.32036e-19 $X=6.38 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_649 N_A_719_47#_c_750_n N_A_1262_49#_M1004_s 0.00226752f $X=6.235 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_650 N_A_719_47#_c_747_n N_A_1262_49#_M1009_s 2.50805e-19 $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_651 N_A_719_47#_c_737_n N_A_1262_49#_c_1195_n 0.0076515f $X=6.645 $Y=0.995
+ $X2=0 $Y2=0
cc_652 N_A_719_47#_c_747_n N_A_1262_49#_c_1195_n 0.00903042f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_653 N_A_719_47#_c_738_n N_A_1262_49#_c_1216_n 9.20553e-19 $X=8.45 $Y=0.96
+ $X2=0 $Y2=0
cc_654 N_A_719_47#_c_738_n N_A_1262_49#_c_1196_n 0.0124254f $X=8.45 $Y=0.96
+ $X2=0 $Y2=0
cc_655 N_A_719_47#_c_739_n N_A_1262_49#_c_1196_n 0.00381612f $X=8.88 $Y=1.035
+ $X2=0 $Y2=0
cc_656 N_A_719_47#_c_747_n N_A_1262_49#_c_1196_n 0.0120747f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_657 N_A_719_47#_c_751_n N_A_1262_49#_c_1196_n 0.00255767f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_658 N_A_719_47#_c_752_n N_A_1262_49#_c_1196_n 0.0170689f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_659 N_A_719_47#_c_753_n N_A_1262_49#_c_1196_n 0.00688049f $X=9.12 $Y=0.77
+ $X2=0 $Y2=0
cc_660 N_A_719_47#_M1016_g N_A_1262_49#_c_1205_n 0.0107372f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_661 N_A_719_47#_M1016_g N_A_1262_49#_c_1233_n 0.0040769f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_662 N_A_719_47#_c_737_n N_A_1262_49#_c_1199_n 0.00510065f $X=6.645 $Y=0.995
+ $X2=0 $Y2=0
cc_663 N_A_719_47#_c_742_n N_A_1262_49#_c_1199_n 0.00415785f $X=6.51 $Y=1.16
+ $X2=0 $Y2=0
cc_664 N_A_719_47#_c_747_n N_A_1262_49#_c_1199_n 0.00537753f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_665 N_A_719_47#_c_748_n N_A_1262_49#_c_1199_n 0.00123323f $X=6.38 $Y=0.85
+ $X2=0 $Y2=0
cc_666 N_A_719_47#_c_750_n N_A_1262_49#_c_1199_n 0.0115331f $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_667 N_A_719_47#_c_747_n N_A_1262_49#_c_1217_n 0.0116665f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_668 N_A_719_47#_c_747_n N_A_1262_49#_c_1200_n 0.00744446f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_669 N_A_719_47#_c_747_n N_A_1332_297#_M1004_d 4.43088e-19 $X=8.86 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_670 N_A_719_47#_c_737_n N_A_1332_297#_c_1369_n 0.00473778f $X=6.645 $Y=0.995
+ $X2=0 $Y2=0
cc_671 N_A_719_47#_c_747_n N_A_1332_297#_c_1369_n 0.0175732f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_672 N_A_719_47#_c_748_n N_A_1332_297#_c_1369_n 4.83658e-19 $X=6.38 $Y=0.85
+ $X2=0 $Y2=0
cc_673 N_A_719_47#_c_750_n N_A_1332_297#_c_1369_n 0.0113597f $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_674 N_A_719_47#_c_737_n N_A_1332_297#_c_1370_n 0.00162425f $X=6.645 $Y=0.995
+ $X2=0 $Y2=0
cc_675 N_A_719_47#_c_743_n N_A_1332_297#_c_1370_n 0.00395545f $X=6.615 $Y=1.16
+ $X2=0 $Y2=0
cc_676 N_A_719_47#_c_748_n N_A_1332_297#_c_1370_n 2.48897e-19 $X=6.38 $Y=0.85
+ $X2=0 $Y2=0
cc_677 N_A_719_47#_c_750_n N_A_1332_297#_c_1370_n 0.0228214f $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_678 N_A_719_47#_M1026_g N_A_1332_297#_c_1377_n 0.00319689f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_679 N_A_719_47#_c_743_n N_A_1332_297#_c_1377_n 0.00204841f $X=6.615 $Y=1.16
+ $X2=0 $Y2=0
cc_680 N_A_719_47#_c_740_n N_A_1332_297#_c_1371_n 9.99078e-19 $X=8.525 $Y=1.035
+ $X2=0 $Y2=0
cc_681 N_A_719_47#_c_747_n N_A_1332_297#_c_1371_n 0.15806f $X=8.86 $Y=0.85 $X2=0
+ $Y2=0
cc_682 N_A_719_47#_c_751_n N_A_1332_297#_c_1371_n 0.0260293f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_683 N_A_719_47#_c_752_n N_A_1332_297#_c_1371_n 0.00344529f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_684 N_A_719_47#_c_743_n N_A_1332_297#_c_1388_n 0.00985134f $X=6.615 $Y=1.16
+ $X2=0 $Y2=0
cc_685 N_A_719_47#_c_747_n N_A_1332_297#_c_1388_n 0.0254504f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_686 N_A_719_47#_c_750_n N_A_1332_297#_c_1388_n 0.00597131f $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_687 N_A_719_47#_c_743_n N_A_1332_297#_c_1372_n 0.00528701f $X=6.615 $Y=1.16
+ $X2=0 $Y2=0
cc_688 N_A_719_47#_c_747_n N_A_1617_49#_M1009_d 5.85211e-19 $X=8.86 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_689 N_A_719_47#_c_738_n N_A_1617_49#_c_1483_n 6.05958e-19 $X=8.45 $Y=0.96
+ $X2=0 $Y2=0
cc_690 N_A_719_47#_c_740_n N_A_1617_49#_c_1483_n 0.00364278f $X=8.525 $Y=1.035
+ $X2=0 $Y2=0
cc_691 N_A_719_47#_M1016_g N_A_1617_49#_c_1483_n 0.00121035f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_692 N_A_719_47#_c_738_n N_A_1617_49#_c_1484_n 0.00380168f $X=8.45 $Y=0.96
+ $X2=0 $Y2=0
cc_693 N_A_719_47#_c_747_n N_A_1617_49#_c_1484_n 0.0144575f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_694 N_A_719_47#_M1016_g N_A_1617_49#_c_1490_n 0.00366662f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_695 N_A_719_47#_M1016_g N_A_1617_49#_c_1491_n 4.6374e-19 $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_696 N_A_719_47#_c_739_n N_A_1617_49#_c_1495_n 0.00136732f $X=8.88 $Y=1.035
+ $X2=0 $Y2=0
cc_697 N_A_719_47#_c_740_n N_A_1617_49#_c_1495_n 0.00172225f $X=8.525 $Y=1.035
+ $X2=0 $Y2=0
cc_698 N_A_719_47#_M1016_g N_A_1617_49#_c_1495_n 0.00546399f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_699 N_A_719_47#_c_745_n N_A_27_47#_M1013_d 3.94762e-19 $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_700 N_A_719_47#_c_745_n N_A_27_47#_M1014_d 0.00206828f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_701 N_A_719_47#_c_758_n N_A_27_47#_M1023_s 0.00275401f $X=3.73 $Y=1.62 $X2=0
+ $Y2=0
cc_702 N_A_719_47#_M1023_d N_A_27_47#_c_1611_n 0.00171563f $X=3.595 $Y=1.485
+ $X2=0 $Y2=0
cc_703 N_A_719_47#_c_745_n N_A_27_47#_c_1653_n 0.00864742f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_704 N_A_719_47#_c_763_n N_A_27_47#_c_1605_n 0.00674531f $X=3.735 $Y=0.72
+ $X2=0 $Y2=0
cc_705 N_A_719_47#_c_745_n N_A_27_47#_c_1605_n 0.0469999f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_706 N_A_719_47#_c_746_n N_A_27_47#_c_1605_n 2.00081e-19 $X=3.6 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_A_719_47#_c_749_n N_A_27_47#_c_1605_n 0.00138412f $X=3.455 $Y=0.85
+ $X2=0 $Y2=0
cc_708 N_A_719_47#_c_737_n N_A_27_47#_c_1606_n 5.45612e-19 $X=6.645 $Y=0.995
+ $X2=0 $Y2=0
cc_709 N_A_719_47#_c_745_n N_A_27_47#_c_1606_n 0.00766236f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_710 N_A_719_47#_c_748_n N_A_27_47#_c_1606_n 3.05956e-19 $X=6.38 $Y=0.85 $X2=0
+ $Y2=0
cc_711 N_A_719_47#_M1026_g N_VPWR_c_1776_n 9.44495e-19 $X=6.585 $Y=1.905 $X2=0
+ $Y2=0
cc_712 N_A_719_47#_M1016_g N_VPWR_c_1776_n 0.00313972f $X=8.955 $Y=1.995 $X2=0
+ $Y2=0
cc_713 N_A_719_47#_M1016_g N_VPWR_c_1769_n 0.00490077f $X=8.955 $Y=1.995 $X2=0
+ $Y2=0
cc_714 N_A_719_47#_c_762_n N_A_310_49#_M1027_s 0.00160811f $X=3.54 $Y=0.72 $X2=0
+ $Y2=0
cc_715 N_A_719_47#_c_746_n N_A_310_49#_M1027_s 0.0016187f $X=3.6 $Y=0.85 $X2=0
+ $Y2=0
cc_716 N_A_719_47#_c_749_n N_A_310_49#_M1027_s 3.27123e-19 $X=3.455 $Y=0.85
+ $X2=0 $Y2=0
cc_717 N_A_719_47#_c_762_n N_A_310_49#_c_1888_n 0.0124754f $X=3.54 $Y=0.72 $X2=0
+ $Y2=0
cc_718 N_A_719_47#_c_758_n N_A_310_49#_c_1888_n 0.0246367f $X=3.73 $Y=1.62 $X2=0
+ $Y2=0
cc_719 N_A_719_47#_c_746_n N_A_310_49#_c_1888_n 0.00772633f $X=3.6 $Y=0.85 $X2=0
+ $Y2=0
cc_720 N_A_719_47#_c_749_n N_A_310_49#_c_1888_n 0.0442505f $X=3.455 $Y=0.85
+ $X2=0 $Y2=0
cc_721 N_A_719_47#_M1027_d N_A_310_49#_c_1889_n 0.00315453f $X=3.595 $Y=0.235
+ $X2=0 $Y2=0
cc_722 N_A_719_47#_c_762_n N_A_310_49#_c_1889_n 0.00771986f $X=3.54 $Y=0.72
+ $X2=0 $Y2=0
cc_723 N_A_719_47#_c_763_n N_A_310_49#_c_1889_n 0.0155392f $X=3.735 $Y=0.72
+ $X2=0 $Y2=0
cc_724 N_A_719_47#_c_745_n N_A_310_49#_c_1889_n 0.00727415f $X=6.09 $Y=0.85
+ $X2=0 $Y2=0
cc_725 N_A_719_47#_c_746_n N_A_310_49#_c_1889_n 0.00245497f $X=3.6 $Y=0.85 $X2=0
+ $Y2=0
cc_726 N_A_719_47#_M1023_d N_A_310_49#_c_1938_n 0.00327408f $X=3.595 $Y=1.485
+ $X2=0 $Y2=0
cc_727 N_A_719_47#_c_758_n N_A_310_49#_c_1938_n 0.0230086f $X=3.73 $Y=1.62 $X2=0
+ $Y2=0
cc_728 N_A_719_47#_c_745_n N_A_310_49#_c_1961_n 8.80211e-19 $X=6.09 $Y=0.85
+ $X2=0 $Y2=0
cc_729 N_A_719_47#_c_758_n N_A_310_49#_c_1943_n 0.00154141f $X=3.73 $Y=1.62
+ $X2=0 $Y2=0
cc_730 N_A_719_47#_M1026_g N_A_310_49#_c_1897_n 0.00101069f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_731 N_A_719_47#_c_747_n N_A_1640_380#_M1003_d 9.11257e-19 $X=8.86 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_732 N_A_719_47#_M1016_g N_A_1640_380#_c_2063_n 0.0116278f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_733 N_A_719_47#_c_738_n N_A_1640_380#_c_2057_n 7.6892e-19 $X=8.45 $Y=0.96
+ $X2=0 $Y2=0
cc_734 N_A_719_47#_c_739_n N_A_1640_380#_c_2057_n 0.0127342f $X=8.88 $Y=1.035
+ $X2=0 $Y2=0
cc_735 N_A_719_47#_c_747_n N_A_1640_380#_c_2057_n 0.0110725f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_736 N_A_719_47#_c_751_n N_A_1640_380#_c_2057_n 0.003361f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_737 N_A_719_47#_c_752_n N_A_1640_380#_c_2057_n 0.0172383f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_738 N_A_719_47#_c_753_n N_A_1640_380#_c_2057_n 0.00292818f $X=9.12 $Y=0.77
+ $X2=0 $Y2=0
cc_739 N_A_719_47#_c_739_n N_A_1640_380#_c_2058_n 0.00421511f $X=8.88 $Y=1.035
+ $X2=0 $Y2=0
cc_740 N_A_719_47#_M1016_g N_A_1640_380#_c_2058_n 0.00946354f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_741 N_A_719_47#_c_744_n N_A_1640_380#_c_2058_n 0.0088663f $X=8.88 $Y=0.96
+ $X2=0 $Y2=0
cc_742 N_A_719_47#_c_747_n N_A_1640_380#_c_2058_n 0.00252963f $X=8.86 $Y=0.85
+ $X2=0 $Y2=0
cc_743 N_A_719_47#_c_751_n N_A_1640_380#_c_2058_n 0.00260267f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_744 N_A_719_47#_c_752_n N_A_1640_380#_c_2058_n 0.0216967f $X=9.005 $Y=0.85
+ $X2=0 $Y2=0
cc_745 N_A_719_47#_c_739_n N_A_1640_380#_c_2059_n 0.00277276f $X=8.88 $Y=1.035
+ $X2=0 $Y2=0
cc_746 N_A_719_47#_M1016_g N_A_1640_380#_c_2083_n 0.00550078f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_747 N_A_719_47#_M1016_g N_A_1640_380#_c_2061_n 0.00883479f $X=8.955 $Y=1.995
+ $X2=0 $Y2=0
cc_748 N_A_719_47#_c_737_n N_VGND_c_2233_n 0.00352679f $X=6.645 $Y=0.995 $X2=0
+ $Y2=0
cc_749 N_A_719_47#_c_738_n N_VGND_c_2233_n 0.00357877f $X=8.45 $Y=0.96 $X2=0
+ $Y2=0
cc_750 N_A_719_47#_c_750_n N_VGND_c_2233_n 0.0025152f $X=6.235 $Y=0.85 $X2=0
+ $Y2=0
cc_751 N_A_719_47#_M1027_d N_VGND_c_2239_n 0.00181549f $X=3.595 $Y=0.235 $X2=0
+ $Y2=0
cc_752 N_A_719_47#_c_737_n N_VGND_c_2239_n 0.00640984f $X=6.645 $Y=0.995 $X2=0
+ $Y2=0
cc_753 N_A_719_47#_c_738_n N_VGND_c_2239_n 0.00676309f $X=8.45 $Y=0.96 $X2=0
+ $Y2=0
cc_754 N_A_719_47#_c_745_n N_VGND_c_2239_n 0.117796f $X=6.09 $Y=0.85 $X2=0 $Y2=0
cc_755 N_A_719_47#_c_746_n N_VGND_c_2239_n 0.0146392f $X=3.6 $Y=0.85 $X2=0 $Y2=0
cc_756 N_A_719_47#_c_747_n N_VGND_c_2239_n 0.119073f $X=8.86 $Y=0.85 $X2=0 $Y2=0
cc_757 N_A_719_47#_c_748_n N_VGND_c_2239_n 0.0165515f $X=6.38 $Y=0.85 $X2=0
+ $Y2=0
cc_758 N_A_719_47#_c_750_n N_VGND_c_2239_n 0.00100315f $X=6.235 $Y=0.85 $X2=0
+ $Y2=0
cc_759 N_A_719_47#_c_751_n N_VGND_c_2239_n 0.0150329f $X=9.005 $Y=0.85 $X2=0
+ $Y2=0
cc_760 N_A_1008_47#_c_972_n N_A_1262_49#_M1008_d 0.0081413f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_761 N_A_1008_47#_c_974_n N_A_1262_49#_M1008_d 0.0238122f $X=7.475 $Y=2.295
+ $X2=0 $Y2=0
cc_762 N_A_1008_47#_c_958_n N_A_1262_49#_c_1195_n 0.0126688f $X=7.07 $Y=0.995
+ $X2=0 $Y2=0
cc_763 N_A_1008_47#_c_960_n N_A_1262_49#_c_1195_n 8.84822e-19 $X=7.037 $Y=1.16
+ $X2=0 $Y2=0
cc_764 N_A_1008_47#_c_961_n N_A_1262_49#_c_1195_n 0.0033133f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_765 N_A_1008_47#_c_964_n N_A_1262_49#_c_1195_n 0.00223644f $X=7.535 $Y=1.16
+ $X2=0 $Y2=0
cc_766 N_A_1008_47#_c_958_n N_A_1262_49#_c_1216_n 0.00283052f $X=7.07 $Y=0.995
+ $X2=0 $Y2=0
cc_767 N_A_1008_47#_c_959_n N_A_1262_49#_c_1216_n 0.0048637f $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_768 N_A_1008_47#_c_961_n N_A_1262_49#_c_1203_n 0.00257993f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_769 N_A_1008_47#_c_974_n N_A_1262_49#_c_1203_n 0.0582258f $X=7.475 $Y=2.295
+ $X2=0 $Y2=0
cc_770 N_A_1008_47#_c_968_n N_A_1262_49#_c_1204_n 0.00593355f $X=8.535 $Y=1.5
+ $X2=0 $Y2=0
cc_771 N_A_1008_47#_c_959_n N_A_1262_49#_c_1196_n 0.00738169f $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_772 N_A_1008_47#_c_961_n N_A_1262_49#_c_1196_n 0.00121295f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_773 N_A_1008_47#_c_968_n N_A_1262_49#_c_1205_n 0.011405f $X=8.535 $Y=1.5
+ $X2=0 $Y2=0
cc_774 N_A_1008_47#_M1008_g N_A_1262_49#_c_1206_n 4.93356e-19 $X=7.005 $Y=1.905
+ $X2=0 $Y2=0
cc_775 N_A_1008_47#_c_972_n N_A_1262_49#_c_1206_n 0.0158225f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_776 N_A_1008_47#_c_958_n N_A_1262_49#_c_1199_n 7.8676e-19 $X=7.07 $Y=0.995
+ $X2=0 $Y2=0
cc_777 N_A_1008_47#_c_959_n N_A_1262_49#_c_1258_n 0.00470392f $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_778 N_A_1008_47#_c_959_n N_A_1262_49#_c_1217_n 0.00120482f $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_779 N_A_1008_47#_c_961_n N_A_1262_49#_c_1217_n 0.00303507f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_780 N_A_1008_47#_c_958_n N_A_1262_49#_c_1200_n 5.42905e-19 $X=7.07 $Y=0.995
+ $X2=0 $Y2=0
cc_781 N_A_1008_47#_c_959_n N_A_1262_49#_c_1200_n 0.00399477f $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_782 N_A_1008_47#_c_968_n N_A_1262_49#_c_1200_n 0.00119931f $X=8.535 $Y=1.5
+ $X2=0 $Y2=0
cc_783 N_A_1008_47#_c_961_n N_A_1262_49#_c_1200_n 0.0231073f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_784 N_A_1008_47#_c_974_n N_A_1262_49#_c_1200_n 0.00505102f $X=7.475 $Y=2.295
+ $X2=0 $Y2=0
cc_785 N_A_1008_47#_c_975_n N_A_1262_49#_c_1200_n 0.0107161f $X=7.535 $Y=1.275
+ $X2=0 $Y2=0
cc_786 N_A_1008_47#_c_964_n N_A_1262_49#_c_1200_n 0.0185404f $X=7.535 $Y=1.16
+ $X2=0 $Y2=0
cc_787 N_A_1008_47#_c_972_n N_A_1332_297#_M1026_d 0.00166235f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_788 N_A_1008_47#_c_958_n N_A_1332_297#_c_1369_n 3.84657e-19 $X=7.07 $Y=0.995
+ $X2=0 $Y2=0
cc_789 N_A_1008_47#_c_960_n N_A_1332_297#_c_1369_n 4.95569e-19 $X=7.037 $Y=1.16
+ $X2=0 $Y2=0
cc_790 N_A_1008_47#_c_958_n N_A_1332_297#_c_1370_n 5.0065e-19 $X=7.07 $Y=0.995
+ $X2=0 $Y2=0
cc_791 N_A_1008_47#_c_960_n N_A_1332_297#_c_1370_n 0.0017213f $X=7.037 $Y=1.16
+ $X2=0 $Y2=0
cc_792 N_A_1008_47#_c_967_n N_A_1332_297#_c_1371_n 0.00207942f $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_793 N_A_1008_47#_c_960_n N_A_1332_297#_c_1371_n 0.00656446f $X=7.037 $Y=1.16
+ $X2=0 $Y2=0
cc_794 N_A_1008_47#_c_961_n N_A_1332_297#_c_1371_n 0.0237072f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_795 N_A_1008_47#_c_975_n N_A_1332_297#_c_1371_n 0.00215928f $X=7.535 $Y=1.275
+ $X2=0 $Y2=0
cc_796 N_A_1008_47#_c_964_n N_A_1332_297#_c_1371_n 0.0157136f $X=7.535 $Y=1.16
+ $X2=0 $Y2=0
cc_797 N_A_1008_47#_M1008_g N_A_1332_297#_c_1372_n 0.0017213f $X=7.005 $Y=1.905
+ $X2=0 $Y2=0
cc_798 N_A_1008_47#_c_959_n N_A_1617_49#_c_1483_n 4.95831e-19 $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_799 N_A_1008_47#_c_967_n N_A_1617_49#_c_1483_n 0.00837279f $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_800 N_A_1008_47#_c_961_n N_A_1617_49#_c_1483_n 0.00438911f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_801 N_A_1008_47#_c_959_n N_A_1617_49#_c_1484_n 0.00115711f $X=8.01 $Y=0.995
+ $X2=0 $Y2=0
cc_802 N_A_1008_47#_c_967_n N_A_1617_49#_c_1484_n 0.00169035f $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_803 N_A_1008_47#_c_961_n N_A_1617_49#_c_1484_n 4.27141e-19 $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_804 N_A_1008_47#_c_967_n N_A_1617_49#_c_1489_n 0.00521858f $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_805 N_A_1008_47#_c_967_n N_A_1617_49#_c_1491_n 7.8975e-19 $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_806 N_A_1008_47#_c_967_n N_A_1617_49#_c_1495_n 0.00598359f $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_807 N_A_1008_47#_c_968_n N_A_1617_49#_c_1495_n 0.012293f $X=8.535 $Y=1.5
+ $X2=0 $Y2=0
cc_808 N_A_1008_47#_c_973_n N_A_27_47#_c_1612_n 0.0134475f $X=5.295 $Y=2.38
+ $X2=0 $Y2=0
cc_809 N_A_1008_47#_c_971_n N_A_27_47#_c_1602_n 0.0151785f $X=5.21 $Y=2.145
+ $X2=0 $Y2=0
cc_810 N_A_1008_47#_c_963_n N_A_27_47#_c_1602_n 0.00773686f $X=5.412 $Y=1.15
+ $X2=0 $Y2=0
cc_811 N_A_1008_47#_c_965_n N_A_27_47#_c_1602_n 0.00841489f $X=5.412 $Y=1.235
+ $X2=0 $Y2=0
cc_812 N_A_1008_47#_M1002_d N_A_27_47#_c_1652_n 0.00304555f $X=5.04 $Y=0.235
+ $X2=0 $Y2=0
cc_813 N_A_1008_47#_c_962_n N_A_27_47#_c_1652_n 0.00434454f $X=5.412 $Y=0.925
+ $X2=0 $Y2=0
cc_814 N_A_1008_47#_M1002_d N_A_27_47#_c_1653_n 0.010455f $X=5.04 $Y=0.235 $X2=0
+ $Y2=0
cc_815 N_A_1008_47#_c_962_n N_A_27_47#_c_1653_n 0.0126956f $X=5.412 $Y=0.925
+ $X2=0 $Y2=0
cc_816 N_A_1008_47#_M1002_d N_A_27_47#_c_1680_n 8.08698e-19 $X=5.04 $Y=0.235
+ $X2=0 $Y2=0
cc_817 N_A_1008_47#_M1002_d N_A_27_47#_c_1605_n 0.00206521f $X=5.04 $Y=0.235
+ $X2=0 $Y2=0
cc_818 N_A_1008_47#_c_962_n N_A_27_47#_c_1605_n 0.0187876f $X=5.412 $Y=0.925
+ $X2=0 $Y2=0
cc_819 N_A_1008_47#_c_965_n N_A_27_47#_c_1605_n 0.00215467f $X=5.412 $Y=1.235
+ $X2=0 $Y2=0
cc_820 N_A_1008_47#_M1008_g N_VPWR_c_1776_n 9.44495e-19 $X=7.005 $Y=1.905 $X2=0
+ $Y2=0
cc_821 N_A_1008_47#_c_968_n N_VPWR_c_1776_n 0.00313972f $X=8.535 $Y=1.5 $X2=0
+ $Y2=0
cc_822 N_A_1008_47#_c_972_n N_VPWR_c_1776_n 0.146665f $X=7.39 $Y=2.38 $X2=0
+ $Y2=0
cc_823 N_A_1008_47#_c_973_n N_VPWR_c_1776_n 0.0121882f $X=5.295 $Y=2.38 $X2=0
+ $Y2=0
cc_824 N_A_1008_47#_c_968_n N_VPWR_c_1769_n 0.00519382f $X=8.535 $Y=1.5 $X2=0
+ $Y2=0
cc_825 N_A_1008_47#_c_972_n N_VPWR_c_1769_n 0.0738253f $X=7.39 $Y=2.38 $X2=0
+ $Y2=0
cc_826 N_A_1008_47#_c_973_n N_VPWR_c_1769_n 0.00311866f $X=5.295 $Y=2.38 $X2=0
+ $Y2=0
cc_827 N_A_1008_47#_c_972_n N_A_310_49#_M1020_d 0.00316065f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_828 N_A_1008_47#_M1022_d N_A_310_49#_c_1895_n 0.00282986f $X=5.075 $Y=1.485
+ $X2=0 $Y2=0
cc_829 N_A_1008_47#_c_971_n N_A_310_49#_c_1895_n 0.0132514f $X=5.21 $Y=2.145
+ $X2=0 $Y2=0
cc_830 N_A_1008_47#_c_972_n N_A_310_49#_c_1895_n 0.00427928f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_831 N_A_1008_47#_c_971_n N_A_310_49#_c_1975_n 6.13307e-19 $X=5.21 $Y=2.145
+ $X2=0 $Y2=0
cc_832 N_A_1008_47#_c_972_n N_A_310_49#_c_1975_n 0.00121888f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_833 N_A_1008_47#_c_971_n N_A_310_49#_c_1897_n 0.021846f $X=5.21 $Y=2.145
+ $X2=0 $Y2=0
cc_834 N_A_1008_47#_c_972_n N_A_310_49#_c_1897_n 0.0147926f $X=7.39 $Y=2.38
+ $X2=0 $Y2=0
cc_835 N_A_1008_47#_c_965_n N_A_310_49#_c_1897_n 5.61716e-19 $X=5.412 $Y=1.235
+ $X2=0 $Y2=0
cc_836 N_A_1008_47#_c_967_n N_A_1640_380#_c_2063_n 8.27809e-19 $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_837 N_A_1008_47#_c_968_n N_A_1640_380#_c_2063_n 0.00826657f $X=8.535 $Y=1.5
+ $X2=0 $Y2=0
cc_838 N_A_1008_47#_c_961_n N_A_1640_380#_c_2063_n 0.0020961f $X=7.935 $Y=1.16
+ $X2=0 $Y2=0
cc_839 N_A_1008_47#_c_967_n N_A_1640_380#_c_2059_n 3.04458e-19 $X=8.46 $Y=1.425
+ $X2=0 $Y2=0
cc_840 N_A_1008_47#_c_968_n N_A_1640_380#_c_2083_n 6.28063e-19 $X=8.535 $Y=1.5
+ $X2=0 $Y2=0
cc_841 N_A_1008_47#_c_958_n N_VGND_c_2233_n 0.00351226f $X=7.07 $Y=0.995 $X2=0
+ $Y2=0
cc_842 N_A_1008_47#_c_959_n N_VGND_c_2233_n 0.00351191f $X=8.01 $Y=0.995 $X2=0
+ $Y2=0
cc_843 N_A_1008_47#_M1002_d N_VGND_c_2239_n 0.00240833f $X=5.04 $Y=0.235 $X2=0
+ $Y2=0
cc_844 N_A_1008_47#_c_958_n N_VGND_c_2239_n 0.00640986f $X=7.07 $Y=0.995 $X2=0
+ $Y2=0
cc_845 N_A_1008_47#_c_959_n N_VGND_c_2239_n 0.00645344f $X=8.01 $Y=0.995 $X2=0
+ $Y2=0
cc_846 N_CI_M1025_g N_A_1262_49#_M1005_g 0.0455799f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_847 N_CI_c_1128_n N_A_1262_49#_c_1196_n 0.00328825f $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_848 N_CI_c_1129_n N_A_1262_49#_c_1196_n 0.00469766f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_849 CI N_A_1262_49#_c_1196_n 0.00146691f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_850 N_CI_c_1132_n N_A_1262_49#_c_1196_n 0.00339629f $X=9.687 $Y=0.995 $X2=0
+ $Y2=0
cc_851 N_CI_M1025_g N_A_1262_49#_c_1205_n 0.00215859f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_852 N_CI_c_1128_n N_A_1262_49#_c_1274_n 0.0033461f $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_853 N_CI_c_1129_n N_A_1262_49#_c_1274_n 0.011697f $X=9.777 $Y=1.2 $X2=0 $Y2=0
cc_854 N_CI_M1025_g N_A_1262_49#_c_1233_n 0.0154098f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_855 N_CI_M1025_g N_A_1262_49#_c_1277_n 0.00893192f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_856 N_CI_c_1128_n N_A_1262_49#_c_1277_n 0.00143764f $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_857 N_CI_c_1129_n N_A_1262_49#_c_1277_n 0.0119884f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_858 CI N_A_1262_49#_c_1277_n 0.00197546f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_859 N_CI_c_1128_n N_A_1262_49#_c_1197_n 0.00222296f $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_860 N_CI_c_1129_n N_A_1262_49#_c_1197_n 0.00925524f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_861 N_CI_c_1130_n N_A_1262_49#_c_1197_n 0.00331727f $X=9.777 $Y=1.075 $X2=0
+ $Y2=0
cc_862 N_CI_c_1128_n N_A_1262_49#_c_1198_n 0.0172886f $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_863 N_CI_c_1129_n N_A_1262_49#_c_1198_n 9.45569e-19 $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_864 N_CI_c_1130_n N_A_1262_49#_c_1198_n 3.05215e-19 $X=9.777 $Y=1.075 $X2=0
+ $Y2=0
cc_865 N_CI_c_1130_n N_A_1262_49#_c_1201_n 5.20069e-19 $X=9.777 $Y=1.075 $X2=0
+ $Y2=0
cc_866 CI N_A_1262_49#_c_1201_n 0.00255732f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_867 N_CI_c_1132_n N_A_1262_49#_c_1201_n 0.0248932f $X=9.687 $Y=0.995 $X2=0
+ $Y2=0
cc_868 N_CI_c_1128_n N_A_1332_297#_c_1371_n 8.96363e-19 $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_869 N_CI_c_1129_n N_A_1332_297#_c_1371_n 0.0184708f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_870 N_CI_c_1130_n N_A_1332_297#_c_1371_n 0.00196071f $X=9.777 $Y=1.075 $X2=0
+ $Y2=0
cc_871 CI N_A_1332_297#_c_1371_n 0.00438763f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_872 N_CI_M1025_g N_A_1617_49#_c_1490_n 0.00139082f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_873 N_CI_c_1128_n N_A_1617_49#_c_1490_n 0.00340059f $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_874 N_CI_c_1129_n N_A_1617_49#_c_1490_n 0.00240273f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_875 N_CI_M1025_g N_VPWR_c_1772_n 0.00849915f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_876 N_CI_M1025_g N_VPWR_c_1776_n 0.0046653f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_877 N_CI_M1025_g N_VPWR_c_1769_n 0.00553016f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_878 N_CI_c_1128_n N_A_1640_380#_c_2058_n 5.81381e-19 $X=9.64 $Y=1.16 $X2=0
+ $Y2=0
cc_879 N_CI_c_1129_n N_A_1640_380#_c_2058_n 0.0100465f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_880 CI N_A_1640_380#_c_2060_n 0.00551664f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_881 N_CI_c_1132_n N_A_1640_380#_c_2060_n 9.34967e-19 $X=9.687 $Y=0.995 $X2=0
+ $Y2=0
cc_882 N_CI_M1025_g N_A_1640_380#_c_2094_n 0.00621384f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_883 N_CI_M1025_g N_A_1640_380#_c_2061_n 0.00262376f $X=9.795 $Y=1.985 $X2=0
+ $Y2=0
cc_884 N_CI_c_1129_n N_A_1640_380#_c_2061_n 0.00321606f $X=9.777 $Y=1.2 $X2=0
+ $Y2=0
cc_885 N_CI_c_1130_n N_A_1640_380#_c_2062_n 0.00174672f $X=9.777 $Y=1.075 $X2=0
+ $Y2=0
cc_886 CI N_A_1640_380#_c_2062_n 0.0021384f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_887 CI N_VGND_M1024_d 0.00260925f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_888 CI N_VGND_c_2231_n 0.00752265f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_889 N_CI_c_1132_n N_VGND_c_2231_n 0.00285523f $X=9.687 $Y=0.995 $X2=0 $Y2=0
cc_890 CI N_VGND_c_2233_n 0.00197327f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_891 N_CI_c_1132_n N_VGND_c_2233_n 0.00423442f $X=9.687 $Y=0.995 $X2=0 $Y2=0
cc_892 CI N_VGND_c_2239_n 0.00442485f $X=9.84 $Y=0.765 $X2=0 $Y2=0
cc_893 N_CI_c_1132_n N_VGND_c_2239_n 0.00723947f $X=9.687 $Y=0.995 $X2=0 $Y2=0
cc_894 N_A_1262_49#_c_1195_n N_A_1332_297#_M1004_d 0.00313786f $X=7.705 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_895 N_A_1262_49#_c_1195_n N_A_1332_297#_c_1369_n 0.0147958f $X=7.705 $Y=0.34
+ $X2=0 $Y2=0
cc_896 N_A_1262_49#_c_1203_n N_A_1332_297#_c_1371_n 0.00265658f $X=7.845
+ $Y=1.625 $X2=0 $Y2=0
cc_897 N_A_1262_49#_c_1196_n N_A_1332_297#_c_1371_n 0.00378056f $X=9.4 $Y=0.34
+ $X2=0 $Y2=0
cc_898 N_A_1262_49#_c_1274_n N_A_1332_297#_c_1371_n 5.28357e-19 $X=9.537
+ $Y=1.705 $X2=0 $Y2=0
cc_899 N_A_1262_49#_c_1277_n N_A_1332_297#_c_1371_n 0.00236034f $X=10.18 $Y=1.6
+ $X2=0 $Y2=0
cc_900 N_A_1262_49#_c_1197_n N_A_1332_297#_c_1371_n 0.0128995f $X=10.265 $Y=1.16
+ $X2=0 $Y2=0
cc_901 N_A_1262_49#_c_1198_n N_A_1332_297#_c_1371_n 0.00616793f $X=10.265
+ $Y=1.16 $X2=0 $Y2=0
cc_902 N_A_1262_49#_c_1217_n N_A_1332_297#_c_1371_n 4.35348e-19 $X=7.832
+ $Y=0.825 $X2=0 $Y2=0
cc_903 N_A_1262_49#_c_1200_n N_A_1332_297#_c_1371_n 0.0174424f $X=7.845 $Y=1.51
+ $X2=0 $Y2=0
cc_904 N_A_1262_49#_c_1198_n N_A_1332_297#_c_1373_n 0.00379954f $X=10.265
+ $Y=1.16 $X2=0 $Y2=0
cc_905 N_A_1262_49#_c_1196_n N_A_1617_49#_M1009_d 0.00338309f $X=9.4 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_906 N_A_1262_49#_c_1205_n N_A_1617_49#_M1019_d 0.00166235f $X=9.42 $Y=2.38
+ $X2=0 $Y2=0
cc_907 N_A_1262_49#_c_1200_n N_A_1617_49#_c_1483_n 0.0254092f $X=7.845 $Y=1.51
+ $X2=0 $Y2=0
cc_908 N_A_1262_49#_c_1216_n N_A_1617_49#_c_1484_n 0.0208352f $X=7.8 $Y=0.66
+ $X2=0 $Y2=0
cc_909 N_A_1262_49#_c_1196_n N_A_1617_49#_c_1484_n 0.0133054f $X=9.4 $Y=0.34
+ $X2=0 $Y2=0
cc_910 N_A_1262_49#_c_1200_n N_A_1617_49#_c_1489_n 0.0195371f $X=7.845 $Y=1.51
+ $X2=0 $Y2=0
cc_911 N_A_1262_49#_M1016_d N_A_1617_49#_c_1490_n 0.00175995f $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_912 N_A_1262_49#_M1005_g N_A_1617_49#_c_1490_n 6.19441e-19 $X=10.215 $Y=1.985
+ $X2=0 $Y2=0
cc_913 N_A_1262_49#_c_1274_n N_A_1617_49#_c_1490_n 0.00889489f $X=9.537 $Y=1.705
+ $X2=0 $Y2=0
cc_914 N_A_1262_49#_c_1277_n N_A_1617_49#_c_1490_n 0.0207848f $X=10.18 $Y=1.6
+ $X2=0 $Y2=0
cc_915 N_A_1262_49#_c_1197_n N_A_1617_49#_c_1490_n 0.00451552f $X=10.265 $Y=1.16
+ $X2=0 $Y2=0
cc_916 N_A_1262_49#_c_1198_n N_A_1617_49#_c_1490_n 0.00154994f $X=10.265 $Y=1.16
+ $X2=0 $Y2=0
cc_917 N_A_1262_49#_c_1200_n N_A_1617_49#_c_1491_n 0.00116903f $X=7.845 $Y=1.51
+ $X2=0 $Y2=0
cc_918 N_A_1262_49#_c_1199_n N_A_27_47#_c_1606_n 0.0259285f $X=6.435 $Y=0.34
+ $X2=0 $Y2=0
cc_919 N_A_1262_49#_c_1277_n N_VPWR_M1025_d 0.00471447f $X=10.18 $Y=1.6 $X2=0
+ $Y2=0
cc_920 N_A_1262_49#_M1005_g N_VPWR_c_1772_n 0.00877469f $X=10.215 $Y=1.985 $X2=0
+ $Y2=0
cc_921 N_A_1262_49#_c_1205_n N_VPWR_c_1772_n 0.0131625f $X=9.42 $Y=2.38 $X2=0
+ $Y2=0
cc_922 N_A_1262_49#_c_1233_n N_VPWR_c_1772_n 0.00138304f $X=9.537 $Y=2.295 $X2=0
+ $Y2=0
cc_923 N_A_1262_49#_c_1277_n N_VPWR_c_1772_n 0.00288797f $X=10.18 $Y=1.6 $X2=0
+ $Y2=0
cc_924 N_A_1262_49#_c_1205_n N_VPWR_c_1776_n 0.109331f $X=9.42 $Y=2.38 $X2=0
+ $Y2=0
cc_925 N_A_1262_49#_c_1206_n N_VPWR_c_1776_n 0.0164899f $X=7.96 $Y=2.38 $X2=0
+ $Y2=0
cc_926 N_A_1262_49#_M1005_g N_VPWR_c_1777_n 0.00447018f $X=10.215 $Y=1.985 $X2=0
+ $Y2=0
cc_927 N_A_1262_49#_M1016_d N_VPWR_c_1769_n 0.00501982f $X=9.03 $Y=1.575 $X2=0
+ $Y2=0
cc_928 N_A_1262_49#_M1005_g N_VPWR_c_1769_n 0.00565512f $X=10.215 $Y=1.985 $X2=0
+ $Y2=0
cc_929 N_A_1262_49#_c_1205_n N_VPWR_c_1769_n 0.0490306f $X=9.42 $Y=2.38 $X2=0
+ $Y2=0
cc_930 N_A_1262_49#_c_1206_n N_VPWR_c_1769_n 0.0088577f $X=7.96 $Y=2.38 $X2=0
+ $Y2=0
cc_931 N_A_1262_49#_c_1196_n N_A_1640_380#_M1003_d 0.00493723f $X=9.4 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_932 N_A_1262_49#_c_1205_n N_A_1640_380#_M1019_s 0.00269012f $X=9.42 $Y=2.38
+ $X2=0 $Y2=0
cc_933 N_A_1262_49#_c_1277_n N_A_1640_380#_M1005_d 0.00166138f $X=10.18 $Y=1.6
+ $X2=0 $Y2=0
cc_934 N_A_1262_49#_M1016_d N_A_1640_380#_c_2063_n 0.00359954f $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_935 N_A_1262_49#_c_1204_n N_A_1640_380#_c_2063_n 0.0136454f $X=7.815 $Y=1.675
+ $X2=0 $Y2=0
cc_936 N_A_1262_49#_c_1205_n N_A_1640_380#_c_2063_n 0.0591377f $X=9.42 $Y=2.38
+ $X2=0 $Y2=0
cc_937 N_A_1262_49#_c_1233_n N_A_1640_380#_c_2063_n 0.0136207f $X=9.537 $Y=2.295
+ $X2=0 $Y2=0
cc_938 N_A_1262_49#_c_1196_n N_A_1640_380#_c_2057_n 0.011666f $X=9.4 $Y=0.34
+ $X2=0 $Y2=0
cc_939 N_A_1262_49#_M1005_g N_A_1640_380#_c_2064_n 0.00442386f $X=10.215
+ $Y=1.985 $X2=0 $Y2=0
cc_940 N_A_1262_49#_c_1198_n N_A_1640_380#_c_2064_n 0.00176465f $X=10.265
+ $Y=1.16 $X2=0 $Y2=0
cc_941 N_A_1262_49#_c_1197_n N_A_1640_380#_c_2060_n 0.00601595f $X=10.265
+ $Y=1.16 $X2=0 $Y2=0
cc_942 N_A_1262_49#_c_1198_n N_A_1640_380#_c_2060_n 0.00388354f $X=10.265
+ $Y=1.16 $X2=0 $Y2=0
cc_943 N_A_1262_49#_c_1201_n N_A_1640_380#_c_2060_n 0.00790867f $X=10.277
+ $Y=0.995 $X2=0 $Y2=0
cc_944 N_A_1262_49#_M1016_d N_A_1640_380#_c_2094_n 0.00313878f $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_945 N_A_1262_49#_M1005_g N_A_1640_380#_c_2094_n 0.00567318f $X=10.215
+ $Y=1.985 $X2=0 $Y2=0
cc_946 N_A_1262_49#_c_1205_n N_A_1640_380#_c_2094_n 0.00271419f $X=9.42 $Y=2.38
+ $X2=0 $Y2=0
cc_947 N_A_1262_49#_c_1233_n N_A_1640_380#_c_2094_n 0.019506f $X=9.537 $Y=2.295
+ $X2=0 $Y2=0
cc_948 N_A_1262_49#_c_1277_n N_A_1640_380#_c_2094_n 0.015116f $X=10.18 $Y=1.6
+ $X2=0 $Y2=0
cc_949 N_A_1262_49#_M1016_d N_A_1640_380#_c_2083_n 0.00198034f $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_950 N_A_1262_49#_c_1205_n N_A_1640_380#_c_2083_n 0.00230246f $X=9.42 $Y=2.38
+ $X2=0 $Y2=0
cc_951 N_A_1262_49#_c_1233_n N_A_1640_380#_c_2083_n 0.00277295f $X=9.537
+ $Y=2.295 $X2=0 $Y2=0
cc_952 N_A_1262_49#_M1016_d N_A_1640_380#_c_2061_n 0.00465651f $X=9.03 $Y=1.575
+ $X2=0 $Y2=0
cc_953 N_A_1262_49#_c_1274_n N_A_1640_380#_c_2061_n 0.0159794f $X=9.537 $Y=1.705
+ $X2=0 $Y2=0
cc_954 N_A_1262_49#_c_1233_n N_A_1640_380#_c_2061_n 0.0171989f $X=9.537 $Y=2.295
+ $X2=0 $Y2=0
cc_955 N_A_1262_49#_M1005_g N_A_1640_380#_c_2066_n 0.00107225f $X=10.215
+ $Y=1.985 $X2=0 $Y2=0
cc_956 N_A_1262_49#_M1005_g N_A_1640_380#_c_2062_n 0.00572913f $X=10.215
+ $Y=1.985 $X2=0 $Y2=0
cc_957 N_A_1262_49#_c_1277_n N_A_1640_380#_c_2062_n 0.0159139f $X=10.18 $Y=1.6
+ $X2=0 $Y2=0
cc_958 N_A_1262_49#_c_1197_n N_A_1640_380#_c_2062_n 0.035651f $X=10.265 $Y=1.16
+ $X2=0 $Y2=0
cc_959 N_A_1262_49#_c_1198_n N_A_1640_380#_c_2062_n 0.00373686f $X=10.265
+ $Y=1.16 $X2=0 $Y2=0
cc_960 N_A_1262_49#_c_1201_n N_A_1640_380#_c_2062_n 0.00237687f $X=10.277
+ $Y=0.995 $X2=0 $Y2=0
cc_961 N_A_1262_49#_M1005_g N_COUT_c_2175_n 0.00140575f $X=10.215 $Y=1.985 $X2=0
+ $Y2=0
cc_962 N_A_1262_49#_c_1201_n N_VGND_c_2231_n 0.00285523f $X=10.277 $Y=0.995
+ $X2=0 $Y2=0
cc_963 N_A_1262_49#_c_1195_n N_VGND_c_2233_n 0.0649838f $X=7.705 $Y=0.34 $X2=0
+ $Y2=0
cc_964 N_A_1262_49#_c_1196_n N_VGND_c_2233_n 0.106655f $X=9.4 $Y=0.34 $X2=0
+ $Y2=0
cc_965 N_A_1262_49#_c_1199_n N_VGND_c_2233_n 0.0200489f $X=6.435 $Y=0.34 $X2=0
+ $Y2=0
cc_966 N_A_1262_49#_c_1258_n N_VGND_c_2233_n 0.0158168f $X=7.832 $Y=0.34 $X2=0
+ $Y2=0
cc_967 N_A_1262_49#_c_1201_n N_VGND_c_2235_n 0.0054256f $X=10.277 $Y=0.995 $X2=0
+ $Y2=0
cc_968 N_A_1262_49#_c_1195_n N_VGND_c_2239_n 0.018303f $X=7.705 $Y=0.34 $X2=0
+ $Y2=0
cc_969 N_A_1262_49#_c_1196_n N_VGND_c_2239_n 0.0411952f $X=9.4 $Y=0.34 $X2=0
+ $Y2=0
cc_970 N_A_1262_49#_c_1199_n N_VGND_c_2239_n 0.00562289f $X=6.435 $Y=0.34 $X2=0
+ $Y2=0
cc_971 N_A_1262_49#_c_1258_n N_VGND_c_2239_n 0.0046092f $X=7.832 $Y=0.34 $X2=0
+ $Y2=0
cc_972 N_A_1262_49#_c_1201_n N_VGND_c_2239_n 0.0110232f $X=10.277 $Y=0.995 $X2=0
+ $Y2=0
cc_973 N_A_1332_297#_c_1375_n N_A_1617_49#_c_1482_n 0.0114842f $X=11.325
+ $Y=0.995 $X2=0 $Y2=0
cc_974 N_A_1332_297#_M1001_g N_A_1617_49#_M1030_g 0.0261027f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_975 N_A_1332_297#_c_1371_n N_A_1617_49#_c_1483_n 0.0131697f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_976 N_A_1332_297#_c_1371_n N_A_1617_49#_c_1484_n 0.0019843f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_977 N_A_1332_297#_M1001_g N_A_1617_49#_c_1490_n 0.00902238f $X=11.435
+ $Y=1.985 $X2=0 $Y2=0
cc_978 N_A_1332_297#_c_1371_n N_A_1617_49#_c_1490_n 0.194152f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_979 N_A_1332_297#_c_1442_p N_A_1617_49#_c_1490_n 0.0264434f $X=11.305 $Y=1.19
+ $X2=0 $Y2=0
cc_980 N_A_1332_297#_c_1373_n N_A_1617_49#_c_1490_n 0.00108685f $X=11.295
+ $Y=1.16 $X2=0 $Y2=0
cc_981 N_A_1332_297#_c_1374_n N_A_1617_49#_c_1490_n 0.00296854f $X=11.295
+ $Y=1.16 $X2=0 $Y2=0
cc_982 N_A_1332_297#_c_1371_n N_A_1617_49#_c_1491_n 0.0269664f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_983 N_A_1332_297#_M1001_g N_A_1617_49#_c_1492_n 0.00142548f $X=11.435
+ $Y=1.985 $X2=0 $Y2=0
cc_984 N_A_1332_297#_c_1373_n N_A_1617_49#_c_1485_n 0.0206397f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_985 N_A_1332_297#_c_1374_n N_A_1617_49#_c_1485_n 3.20034e-19 $X=11.295
+ $Y=1.16 $X2=0 $Y2=0
cc_986 N_A_1332_297#_c_1442_p N_A_1617_49#_c_1486_n 0.00174077f $X=11.305
+ $Y=1.19 $X2=0 $Y2=0
cc_987 N_A_1332_297#_c_1373_n N_A_1617_49#_c_1486_n 0.00459494f $X=11.295
+ $Y=1.16 $X2=0 $Y2=0
cc_988 N_A_1332_297#_c_1374_n N_A_1617_49#_c_1486_n 0.0237104f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_989 N_A_1332_297#_c_1371_n N_A_1617_49#_c_1495_n 0.00366444f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_990 N_A_1332_297#_M1001_g N_VPWR_c_1773_n 0.00280208f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_991 N_A_1332_297#_M1001_g N_VPWR_c_1777_n 0.00541359f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_992 N_A_1332_297#_M1001_g N_VPWR_c_1769_n 0.0108548f $X=11.435 $Y=1.985 $X2=0
+ $Y2=0
cc_993 N_A_1332_297#_c_1371_n N_A_1640_380#_c_2058_n 0.0176627f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_994 N_A_1332_297#_c_1371_n N_A_1640_380#_c_2059_n 0.00757261f $X=11.16
+ $Y=1.19 $X2=0 $Y2=0
cc_995 N_A_1332_297#_c_1371_n N_A_1640_380#_c_2064_n 2.35227e-19 $X=11.16
+ $Y=1.19 $X2=0 $Y2=0
cc_996 N_A_1332_297#_c_1371_n N_A_1640_380#_c_2060_n 0.00809787f $X=11.16
+ $Y=1.19 $X2=0 $Y2=0
cc_997 N_A_1332_297#_c_1375_n N_A_1640_380#_c_2060_n 8.37019e-19 $X=11.325
+ $Y=0.995 $X2=0 $Y2=0
cc_998 N_A_1332_297#_c_1371_n N_A_1640_380#_c_2062_n 0.0171467f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_999 N_A_1332_297#_c_1371_n N_COUT_c_2173_n 0.00405329f $X=11.16 $Y=1.19 $X2=0
+ $Y2=0
cc_1000 N_A_1332_297#_c_1442_p N_COUT_c_2173_n 0.00217065f $X=11.305 $Y=1.19
+ $X2=0 $Y2=0
cc_1001 N_A_1332_297#_c_1373_n N_COUT_c_2173_n 0.00284389f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_1002 N_A_1332_297#_c_1374_n N_COUT_c_2173_n 0.00711623f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_1003 N_A_1332_297#_M1001_g N_COUT_c_2175_n 0.00365711f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_1004 N_A_1332_297#_c_1371_n N_COUT_c_2175_n 5.00076e-19 $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_1005 N_A_1332_297#_c_1442_p N_COUT_c_2175_n 4.17299e-19 $X=11.305 $Y=1.19
+ $X2=0 $Y2=0
cc_1006 N_A_1332_297#_c_1373_n N_COUT_c_2175_n 0.00288941f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_1007 N_A_1332_297#_c_1374_n N_COUT_c_2175_n 0.0107518f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_1008 N_A_1332_297#_M1001_g N_COUT_c_2174_n 0.00297235f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_1009 N_A_1332_297#_c_1371_n N_COUT_c_2174_n 0.0104408f $X=11.16 $Y=1.19 $X2=0
+ $Y2=0
cc_1010 N_A_1332_297#_c_1442_p N_COUT_c_2174_n 0.00237204f $X=11.305 $Y=1.19
+ $X2=0 $Y2=0
cc_1011 N_A_1332_297#_c_1373_n N_COUT_c_2174_n 0.00376522f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_1012 N_A_1332_297#_c_1374_n N_COUT_c_2174_n 0.0224713f $X=11.295 $Y=1.16
+ $X2=0 $Y2=0
cc_1013 N_A_1332_297#_c_1375_n N_COUT_c_2174_n 0.0049454f $X=11.325 $Y=0.995
+ $X2=0 $Y2=0
cc_1014 N_A_1332_297#_M1001_g COUT 0.00789344f $X=11.435 $Y=1.985 $X2=0 $Y2=0
cc_1015 N_A_1332_297#_c_1371_n N_VGND_c_2231_n 0.00253105f $X=11.16 $Y=1.19
+ $X2=0 $Y2=0
cc_1016 N_A_1332_297#_c_1375_n N_VGND_c_2232_n 0.0138246f $X=11.325 $Y=0.995
+ $X2=0 $Y2=0
cc_1017 N_A_1332_297#_c_1375_n N_VGND_c_2235_n 0.0046653f $X=11.325 $Y=0.995
+ $X2=0 $Y2=0
cc_1018 N_A_1332_297#_c_1375_n N_VGND_c_2239_n 0.00934473f $X=11.325 $Y=0.995
+ $X2=0 $Y2=0
cc_1019 N_A_1617_49#_c_1490_n N_VPWR_M1001_d 0.00240467f $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_1020 N_A_1617_49#_c_1492_n N_VPWR_M1001_d 0.00169173f $X=11.765 $Y=1.53 $X2=0
+ $Y2=0
cc_1021 N_A_1617_49#_c_1486_n N_VPWR_M1001_d 0.0013457f $X=11.855 $Y=1.16 $X2=0
+ $Y2=0
cc_1022 N_A_1617_49#_M1030_g N_VPWR_c_1773_n 0.0135622f $X=11.855 $Y=1.985 $X2=0
+ $Y2=0
cc_1023 N_A_1617_49#_c_1490_n N_VPWR_c_1773_n 0.00304002f $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_1024 N_A_1617_49#_c_1492_n N_VPWR_c_1773_n 0.00584345f $X=11.765 $Y=1.53
+ $X2=0 $Y2=0
cc_1025 N_A_1617_49#_c_1486_n N_VPWR_c_1773_n 0.00992907f $X=11.855 $Y=1.16
+ $X2=0 $Y2=0
cc_1026 N_A_1617_49#_M1030_g N_VPWR_c_1778_n 0.00447018f $X=11.855 $Y=1.985
+ $X2=0 $Y2=0
cc_1027 N_A_1617_49#_M1030_g N_VPWR_c_1769_n 0.00861832f $X=11.855 $Y=1.985
+ $X2=0 $Y2=0
cc_1028 N_A_1617_49#_c_1489_n N_A_1640_380#_M1019_s 0.00513254f $X=8.405
+ $Y=1.615 $X2=0 $Y2=0
cc_1029 N_A_1617_49#_c_1490_n N_A_1640_380#_M1005_d 8.77155e-19 $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_1030 N_A_1617_49#_M1019_d N_A_1640_380#_c_2063_n 0.00316995f $X=8.61 $Y=1.575
+ $X2=0 $Y2=0
cc_1031 N_A_1617_49#_c_1489_n N_A_1640_380#_c_2063_n 0.0144674f $X=8.405
+ $Y=1.615 $X2=0 $Y2=0
cc_1032 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2063_n 0.00481802f $X=11.62
+ $Y=1.53 $X2=0 $Y2=0
cc_1033 N_A_1617_49#_c_1491_n N_A_1640_380#_c_2063_n 0.0015003f $X=8.69 $Y=1.53
+ $X2=0 $Y2=0
cc_1034 N_A_1617_49#_c_1495_n N_A_1640_380#_c_2063_n 0.0232624f $X=8.745 $Y=1.7
+ $X2=0 $Y2=0
cc_1035 N_A_1617_49#_c_1484_n N_A_1640_380#_c_2057_n 0.0266716f $X=8.24 $Y=0.76
+ $X2=0 $Y2=0
cc_1036 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2058_n 0.00443484f $X=11.62
+ $Y=1.53 $X2=0 $Y2=0
cc_1037 N_A_1617_49#_c_1495_n N_A_1640_380#_c_2058_n 0.0104812f $X=8.745 $Y=1.7
+ $X2=0 $Y2=0
cc_1038 N_A_1617_49#_c_1483_n N_A_1640_380#_c_2059_n 0.0126646f $X=8.315
+ $Y=1.445 $X2=0 $Y2=0
cc_1039 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2059_n 2.40622e-19 $X=11.62
+ $Y=1.53 $X2=0 $Y2=0
cc_1040 N_A_1617_49#_c_1491_n N_A_1640_380#_c_2059_n 7.9457e-19 $X=8.69 $Y=1.53
+ $X2=0 $Y2=0
cc_1041 N_A_1617_49#_c_1495_n N_A_1640_380#_c_2059_n 0.012339f $X=8.745 $Y=1.7
+ $X2=0 $Y2=0
cc_1042 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2064_n 9.91473e-19 $X=11.62
+ $Y=1.53 $X2=0 $Y2=0
cc_1043 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2094_n 0.0893964f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_1044 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2083_n 0.0259007f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_1045 N_A_1617_49#_c_1495_n N_A_1640_380#_c_2083_n 7.88829e-19 $X=8.745 $Y=1.7
+ $X2=0 $Y2=0
cc_1046 N_A_1617_49#_c_1483_n N_A_1640_380#_c_2061_n 0.00403906f $X=8.315
+ $Y=1.445 $X2=0 $Y2=0
cc_1047 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2061_n 0.0111104f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_1048 N_A_1617_49#_c_1491_n N_A_1640_380#_c_2061_n 0.00112999f $X=8.69 $Y=1.53
+ $X2=0 $Y2=0
cc_1049 N_A_1617_49#_c_1495_n N_A_1640_380#_c_2061_n 0.0182172f $X=8.745 $Y=1.7
+ $X2=0 $Y2=0
cc_1050 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2066_n 0.0261739f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_1051 N_A_1617_49#_c_1490_n N_A_1640_380#_c_2062_n 0.0103815f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_1052 N_A_1617_49#_M1030_g N_COUT_c_2175_n 9.10273e-19 $X=11.855 $Y=1.985
+ $X2=0 $Y2=0
cc_1053 N_A_1617_49#_c_1490_n N_COUT_c_2175_n 0.0386363f $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_1054 N_A_1617_49#_c_1492_n N_COUT_c_2175_n 0.00183855f $X=11.765 $Y=1.53
+ $X2=0 $Y2=0
cc_1055 N_A_1617_49#_c_1486_n N_COUT_c_2175_n 0.00559661f $X=11.855 $Y=1.16
+ $X2=0 $Y2=0
cc_1056 N_A_1617_49#_c_1490_n N_COUT_c_2174_n 0.00445883f $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_1057 N_A_1617_49#_c_1492_n N_COUT_c_2174_n 9.84887e-19 $X=11.765 $Y=1.53
+ $X2=0 $Y2=0
cc_1058 N_A_1617_49#_c_1486_n N_COUT_c_2174_n 0.00437291f $X=11.855 $Y=1.16
+ $X2=0 $Y2=0
cc_1059 N_A_1617_49#_c_1482_n SUM 0.00418494f $X=11.855 $Y=0.995 $X2=0 $Y2=0
cc_1060 N_A_1617_49#_M1030_g SUM 0.00625436f $X=11.855 $Y=1.985 $X2=0 $Y2=0
cc_1061 N_A_1617_49#_c_1492_n SUM 0.00273148f $X=11.765 $Y=1.53 $X2=0 $Y2=0
cc_1062 N_A_1617_49#_c_1485_n SUM 0.00783697f $X=11.855 $Y=1.16 $X2=0 $Y2=0
cc_1063 N_A_1617_49#_c_1486_n SUM 0.0416233f $X=11.855 $Y=1.16 $X2=0 $Y2=0
cc_1064 N_A_1617_49#_c_1482_n N_VGND_c_2232_n 0.0122731f $X=11.855 $Y=0.995
+ $X2=0 $Y2=0
cc_1065 N_A_1617_49#_c_1492_n N_VGND_c_2232_n 0.00106357f $X=11.765 $Y=1.53
+ $X2=0 $Y2=0
cc_1066 N_A_1617_49#_c_1485_n N_VGND_c_2232_n 3.02148e-19 $X=11.855 $Y=1.16
+ $X2=0 $Y2=0
cc_1067 N_A_1617_49#_c_1486_n N_VGND_c_2232_n 0.012897f $X=11.855 $Y=1.16 $X2=0
+ $Y2=0
cc_1068 N_A_1617_49#_c_1482_n N_VGND_c_2238_n 0.0046653f $X=11.855 $Y=0.995
+ $X2=0 $Y2=0
cc_1069 N_A_1617_49#_c_1482_n N_VGND_c_2239_n 0.00904108f $X=11.855 $Y=0.995
+ $X2=0 $Y2=0
cc_1070 N_A_27_47#_c_1609_n N_VPWR_M1006_d 0.00445488f $X=2.635 $Y=1.98
+ $X2=-0.19 $Y2=-0.24
cc_1071 N_A_27_47#_c_1609_n N_VPWR_M1015_d 0.00794204f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1072 N_A_27_47#_c_1609_n N_VPWR_c_1770_n 0.0166389f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1073 N_A_27_47#_c_1609_n N_VPWR_c_1771_n 0.0207433f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1074 N_A_27_47#_c_1610_n N_VPWR_c_1771_n 0.00337017f $X=2.72 $Y=2.295 $X2=0
+ $Y2=0
cc_1075 N_A_27_47#_c_1649_n N_VPWR_c_1771_n 0.0107656f $X=2.805 $Y=2.38 $X2=0
+ $Y2=0
cc_1076 N_A_27_47#_c_1608_n N_VPWR_c_1774_n 0.0204719f $X=0.28 $Y=2.3 $X2=0
+ $Y2=0
cc_1077 N_A_27_47#_c_1609_n N_VPWR_c_1774_n 0.00185965f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1078 N_A_27_47#_c_1616_n N_VPWR_c_1774_n 6.87305e-19 $X=0.265 $Y=1.98 $X2=0
+ $Y2=0
cc_1079 N_A_27_47#_c_1609_n N_VPWR_c_1775_n 0.0176679f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1080 N_A_27_47#_c_1609_n N_VPWR_c_1776_n 0.00341521f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1081 N_A_27_47#_c_1611_n N_VPWR_c_1776_n 0.121949f $X=4.705 $Y=2.38 $X2=0
+ $Y2=0
cc_1082 N_A_27_47#_c_1649_n N_VPWR_c_1776_n 0.0118082f $X=2.805 $Y=2.38 $X2=0
+ $Y2=0
cc_1083 N_A_27_47#_c_1612_n N_VPWR_c_1776_n 0.0168202f $X=4.79 $Y=2.295 $X2=0
+ $Y2=0
cc_1084 N_A_27_47#_M1006_s N_VPWR_c_1769_n 0.00232367f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_1085 N_A_27_47#_M1023_s N_VPWR_c_1769_n 0.00271997f $X=3.085 $Y=1.485 $X2=0
+ $Y2=0
cc_1086 N_A_27_47#_M1022_s N_VPWR_c_1769_n 0.00202964f $X=4.6 $Y=1.485 $X2=0
+ $Y2=0
cc_1087 N_A_27_47#_c_1608_n N_VPWR_c_1769_n 0.0118616f $X=0.28 $Y=2.3 $X2=0
+ $Y2=0
cc_1088 N_A_27_47#_c_1609_n N_VPWR_c_1769_n 0.0423287f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_1089 N_A_27_47#_c_1611_n N_VPWR_c_1769_n 0.0547868f $X=4.705 $Y=2.38 $X2=0
+ $Y2=0
cc_1090 N_A_27_47#_c_1649_n N_VPWR_c_1769_n 0.00651702f $X=2.805 $Y=2.38 $X2=0
+ $Y2=0
cc_1091 N_A_27_47#_c_1612_n N_VPWR_c_1769_n 0.00439667f $X=4.79 $Y=2.295 $X2=0
+ $Y2=0
cc_1092 N_A_27_47#_c_1616_n N_VPWR_c_1769_n 0.00126261f $X=0.265 $Y=1.98 $X2=0
+ $Y2=0
cc_1093 N_A_27_47#_c_1605_n N_A_310_49#_M1002_s 0.00247727f $X=4.79 $Y=0.785
+ $X2=0 $Y2=0
cc_1094 N_A_27_47#_c_1609_n N_A_310_49#_M1015_s 0.00690806f $X=2.635 $Y=1.98
+ $X2=0 $Y2=0
cc_1095 N_A_27_47#_c_1611_n N_A_310_49#_M1010_d 0.0021731f $X=4.705 $Y=2.38
+ $X2=0 $Y2=0
cc_1096 N_A_27_47#_c_1609_n N_A_310_49#_c_1885_n 0.0231036f $X=2.635 $Y=1.98
+ $X2=0 $Y2=0
cc_1097 N_A_27_47#_M1023_s N_A_310_49#_c_1888_n 0.00704053f $X=3.085 $Y=1.485
+ $X2=0 $Y2=0
cc_1098 N_A_27_47#_c_1609_n N_A_310_49#_c_1888_n 0.00413027f $X=2.635 $Y=1.98
+ $X2=0 $Y2=0
cc_1099 N_A_27_47#_M1013_d N_A_310_49#_c_1889_n 0.0071763f $X=4.02 $Y=0.235
+ $X2=0 $Y2=0
cc_1100 N_A_27_47#_c_1605_n N_A_310_49#_c_1889_n 0.0311499f $X=4.79 $Y=0.785
+ $X2=0 $Y2=0
cc_1101 N_A_27_47#_M1023_s N_A_310_49#_c_1938_n 0.00400608f $X=3.085 $Y=1.485
+ $X2=0 $Y2=0
cc_1102 N_A_27_47#_c_1611_n N_A_310_49#_c_1938_n 0.0404929f $X=4.705 $Y=2.38
+ $X2=0 $Y2=0
cc_1103 N_A_27_47#_M1023_s N_A_310_49#_c_1894_n 0.0022887f $X=3.085 $Y=1.485
+ $X2=0 $Y2=0
cc_1104 N_A_27_47#_c_1609_n N_A_310_49#_c_1894_n 0.00845416f $X=2.635 $Y=1.98
+ $X2=0 $Y2=0
cc_1105 N_A_27_47#_c_1610_n N_A_310_49#_c_1894_n 0.00413025f $X=2.72 $Y=2.295
+ $X2=0 $Y2=0
cc_1106 N_A_27_47#_c_1611_n N_A_310_49#_c_1894_n 0.0130729f $X=4.705 $Y=2.38
+ $X2=0 $Y2=0
cc_1107 N_A_27_47#_c_1605_n N_A_310_49#_c_1961_n 0.0133167f $X=4.79 $Y=0.785
+ $X2=0 $Y2=0
cc_1108 N_A_27_47#_M1022_s N_A_310_49#_c_1895_n 0.00257902f $X=4.6 $Y=1.485
+ $X2=0 $Y2=0
cc_1109 N_A_27_47#_c_1611_n N_A_310_49#_c_1895_n 0.00990029f $X=4.705 $Y=2.38
+ $X2=0 $Y2=0
cc_1110 N_A_27_47#_c_1612_n N_A_310_49#_c_1895_n 0.00173116f $X=4.79 $Y=2.295
+ $X2=0 $Y2=0
cc_1111 N_A_27_47#_c_1602_n N_A_310_49#_c_1895_n 0.0144995f $X=4.79 $Y=1.62
+ $X2=0 $Y2=0
cc_1112 N_A_27_47#_c_1611_n N_A_310_49#_c_1943_n 8.75617e-19 $X=4.705 $Y=2.38
+ $X2=0 $Y2=0
cc_1113 N_A_27_47#_c_1602_n N_A_310_49#_c_1943_n 0.00142025f $X=4.79 $Y=1.62
+ $X2=0 $Y2=0
cc_1114 N_A_27_47#_c_1611_n N_A_310_49#_c_1896_n 0.0186135f $X=4.705 $Y=2.38
+ $X2=0 $Y2=0
cc_1115 N_A_27_47#_c_1602_n N_A_310_49#_c_1896_n 0.0125381f $X=4.79 $Y=1.62
+ $X2=0 $Y2=0
cc_1116 N_A_27_47#_c_1653_n N_VGND_c_2233_n 0.0342774f $X=5.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1117 N_A_27_47#_c_1680_n N_VGND_c_2233_n 0.00985107f $X=5.18 $Y=0.34 $X2=0
+ $Y2=0
cc_1118 N_A_27_47#_c_1605_n N_VGND_c_2233_n 0.00202761f $X=4.79 $Y=0.785 $X2=0
+ $Y2=0
cc_1119 N_A_27_47#_c_1606_n N_VGND_c_2233_n 0.0213821f $X=5.925 $Y=0.34 $X2=0
+ $Y2=0
cc_1120 N_A_27_47#_c_1601_n N_VGND_c_2237_n 0.0216364f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_1121 N_A_27_47#_M1029_s N_VGND_c_2239_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_1122 N_A_27_47#_M1013_d N_VGND_c_2239_n 0.00227294f $X=4.02 $Y=0.235 $X2=0
+ $Y2=0
cc_1123 N_A_27_47#_c_1601_n N_VGND_c_2239_n 0.0127767f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_1124 N_A_27_47#_c_1653_n N_VGND_c_2239_n 0.00948054f $X=5.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1125 N_A_27_47#_c_1680_n N_VGND_c_2239_n 0.00304257f $X=5.18 $Y=0.34 $X2=0
+ $Y2=0
cc_1126 N_A_27_47#_c_1605_n N_VGND_c_2239_n 0.00234177f $X=4.79 $Y=0.785 $X2=0
+ $Y2=0
cc_1127 N_A_27_47#_c_1606_n N_VGND_c_2239_n 0.0060564f $X=5.925 $Y=0.34 $X2=0
+ $Y2=0
cc_1128 N_VPWR_c_1769_n N_A_310_49#_M1015_s 0.00330716f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1129 N_VPWR_c_1769_n N_A_310_49#_c_1895_n 0.0636206f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1130 N_VPWR_c_1769_n N_A_310_49#_c_1943_n 0.0146746f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1131 N_VPWR_c_1769_n N_A_310_49#_c_1975_n 0.0146266f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1132 N_VPWR_c_1769_n N_A_1640_380#_M1005_d 0.00227642f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1133 N_VPWR_c_1777_n N_A_1640_380#_c_2064_n 0.0240549f $X=11.56 $Y=2.72 $X2=0
+ $Y2=0
cc_1134 N_VPWR_c_1769_n N_A_1640_380#_c_2064_n 0.0060554f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1135 N_VPWR_M1025_d N_A_1640_380#_c_2094_n 0.00345818f $X=9.87 $Y=1.485 $X2=0
+ $Y2=0
cc_1136 N_VPWR_c_1772_n N_A_1640_380#_c_2094_n 0.00438804f $X=10.005 $Y=2.36
+ $X2=0 $Y2=0
cc_1137 N_VPWR_c_1769_n N_A_1640_380#_c_2094_n 0.0545207f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1138 N_VPWR_c_1769_n N_A_1640_380#_c_2083_n 0.0148685f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1139 N_VPWR_c_1769_n N_A_1640_380#_c_2066_n 0.0151164f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1140 N_VPWR_c_1769_n N_COUT_M1001_s 0.00209319f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1141 N_VPWR_c_1777_n COUT 0.0346602f $X=11.56 $Y=2.72 $X2=0 $Y2=0
cc_1142 N_VPWR_c_1769_n COUT 0.019744f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1143 N_VPWR_c_1769_n N_SUM_M1030_d 0.0042075f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1144 N_VPWR_c_1778_n SUM 0.0246003f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1145 N_VPWR_c_1769_n SUM 0.0133969f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1146 N_A_310_49#_c_1886_n N_VGND_M1018_d 0.0101631f $X=2.35 $Y=0.8 $X2=0
+ $Y2=0
cc_1147 N_A_310_49#_c_1911_n N_VGND_M1018_d 0.00337392f $X=2.435 $Y=0.715 $X2=0
+ $Y2=0
cc_1148 N_A_310_49#_c_1929_n N_VGND_M1018_d 0.00242244f $X=2.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1149 N_A_310_49#_c_1884_n N_VGND_c_2229_n 0.0217208f $X=1.675 $Y=0.39 $X2=0
+ $Y2=0
cc_1150 N_A_310_49#_c_1886_n N_VGND_c_2229_n 0.0020257f $X=2.35 $Y=0.8 $X2=0
+ $Y2=0
cc_1151 N_A_310_49#_c_1886_n N_VGND_c_2230_n 0.0121971f $X=2.35 $Y=0.8 $X2=0
+ $Y2=0
cc_1152 N_A_310_49#_c_1911_n N_VGND_c_2230_n 0.00867962f $X=2.435 $Y=0.715 $X2=0
+ $Y2=0
cc_1153 N_A_310_49#_c_1929_n N_VGND_c_2230_n 0.0138309f $X=2.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1154 N_A_310_49#_c_1886_n N_VGND_c_2233_n 0.00249715f $X=2.35 $Y=0.8 $X2=0
+ $Y2=0
cc_1155 N_A_310_49#_c_1887_n N_VGND_c_2233_n 0.0305912f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_1156 N_A_310_49#_c_1929_n N_VGND_c_2233_n 0.00986054f $X=2.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1157 N_A_310_49#_c_1889_n N_VGND_c_2233_n 0.0862741f $X=4.65 $Y=0.36 $X2=0
+ $Y2=0
cc_1158 N_A_310_49#_c_1891_n N_VGND_c_2233_n 0.0121676f $X=3.115 $Y=0.36 $X2=0
+ $Y2=0
cc_1159 N_A_310_49#_c_1961_n N_VGND_c_2233_n 0.0123665f $X=4.745 $Y=0.36 $X2=0
+ $Y2=0
cc_1160 N_A_310_49#_M1027_s N_VGND_c_2239_n 0.00187139f $X=3.185 $Y=0.235 $X2=0
+ $Y2=0
cc_1161 N_A_310_49#_M1002_s N_VGND_c_2239_n 0.00187067f $X=4.63 $Y=0.235 $X2=0
+ $Y2=0
cc_1162 N_A_310_49#_c_1884_n N_VGND_c_2239_n 0.0128678f $X=1.675 $Y=0.39 $X2=0
+ $Y2=0
cc_1163 N_A_310_49#_c_1886_n N_VGND_c_2239_n 0.00917247f $X=2.35 $Y=0.8 $X2=0
+ $Y2=0
cc_1164 N_A_310_49#_c_1887_n N_VGND_c_2239_n 0.0184421f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_1165 N_A_310_49#_c_1929_n N_VGND_c_2239_n 0.00639673f $X=2.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1166 N_A_310_49#_c_1889_n N_VGND_c_2239_n 0.0263312f $X=4.65 $Y=0.36 $X2=0
+ $Y2=0
cc_1167 N_A_310_49#_c_1891_n N_VGND_c_2239_n 0.006547f $X=3.115 $Y=0.36 $X2=0
+ $Y2=0
cc_1168 N_A_310_49#_c_1961_n N_VGND_c_2239_n 0.00331998f $X=4.745 $Y=0.36 $X2=0
+ $Y2=0
cc_1169 N_A_1640_380#_c_2060_n N_COUT_c_2173_n 0.045257f $X=10.41 $Y=0.4 $X2=0
+ $Y2=0
cc_1170 N_A_1640_380#_c_2064_n N_COUT_c_2175_n 0.0610562f $X=10.517 $Y=2.047
+ $X2=0 $Y2=0
cc_1171 N_A_1640_380#_c_2062_n N_COUT_c_2174_n 0.0610562f $X=10.605 $Y=1.87
+ $X2=0 $Y2=0
cc_1172 N_A_1640_380#_c_2066_n COUT 0.00786871f $X=10.605 $Y=1.87 $X2=0 $Y2=0
cc_1173 N_A_1640_380#_c_2060_n N_VGND_c_2235_n 0.0243803f $X=10.41 $Y=0.4 $X2=0
+ $Y2=0
cc_1174 N_A_1640_380#_c_2060_n N_VGND_c_2239_n 0.0165976f $X=10.41 $Y=0.4 $X2=0
+ $Y2=0
cc_1175 N_COUT_c_2173_n N_VGND_c_2235_n 0.0277127f $X=11.225 $Y=0.55 $X2=0 $Y2=0
cc_1176 N_COUT_M1011_s N_VGND_c_2239_n 0.00392402f $X=11.09 $Y=0.235 $X2=0 $Y2=0
cc_1177 N_COUT_c_2173_n N_VGND_c_2239_n 0.0167206f $X=11.225 $Y=0.55 $X2=0 $Y2=0
cc_1178 N_SUM_c_2213_n N_VGND_c_2238_n 0.0245914f $X=12.145 $Y=0.39 $X2=0 $Y2=0
cc_1179 N_SUM_M1017_d N_VGND_c_2239_n 0.00452756f $X=11.93 $Y=0.235 $X2=0 $Y2=0
cc_1180 N_SUM_c_2213_n N_VGND_c_2239_n 0.0135719f $X=12.145 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o221ai_2.pxi.spice
* Created: Tue Sep  1 19:22:52 2020
* 
x_PM_SKY130_FD_SC_HD__O221AI_2%C1 N_C1_c_87_n N_C1_M1005_g N_C1_M1004_g
+ N_C1_c_88_n N_C1_M1008_g N_C1_M1010_g C1 N_C1_c_90_n
+ PM_SKY130_FD_SC_HD__O221AI_2%C1
x_PM_SKY130_FD_SC_HD__O221AI_2%B1 N_B1_c_128_n N_B1_M1006_g N_B1_M1007_g
+ N_B1_c_129_n N_B1_M1016_g N_B1_M1015_g N_B1_c_137_n N_B1_c_130_n N_B1_c_131_n
+ N_B1_c_132_n N_B1_c_133_n N_B1_c_134_n B1 PM_SKY130_FD_SC_HD__O221AI_2%B1
x_PM_SKY130_FD_SC_HD__O221AI_2%B2 N_B2_c_210_n N_B2_M1000_g N_B2_M1009_g
+ N_B2_c_211_n N_B2_M1001_g N_B2_M1013_g B2 N_B2_c_213_n
+ PM_SKY130_FD_SC_HD__O221AI_2%B2
x_PM_SKY130_FD_SC_HD__O221AI_2%A1 N_A1_c_251_n N_A1_M1002_g N_A1_M1011_g
+ N_A1_c_252_n N_A1_M1003_g N_A1_M1012_g N_A1_c_253_n N_A1_c_254_n N_A1_c_263_n
+ N_A1_c_264_n N_A1_c_255_n N_A1_c_256_n A1 N_A1_c_258_n A1
+ PM_SKY130_FD_SC_HD__O221AI_2%A1
x_PM_SKY130_FD_SC_HD__O221AI_2%A2 N_A2_c_337_n N_A2_M1017_g N_A2_M1014_g
+ N_A2_c_338_n N_A2_M1019_g N_A2_M1018_g A2 N_A2_c_339_n
+ PM_SKY130_FD_SC_HD__O221AI_2%A2
x_PM_SKY130_FD_SC_HD__O221AI_2%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1015_d
+ N_VPWR_M1012_s N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n
+ N_VPWR_c_390_n N_VPWR_c_391_n VPWR N_VPWR_c_392_n N_VPWR_c_393_n
+ N_VPWR_c_385_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n
+ PM_SKY130_FD_SC_HD__O221AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O221AI_2%Y N_Y_M1005_s N_Y_M1004_s N_Y_M1009_s N_Y_M1014_s
+ N_Y_c_459_n N_Y_c_463_n N_Y_c_496_n N_Y_c_475_n N_Y_c_464_n N_Y_c_458_n
+ N_Y_c_472_n N_Y_c_479_n N_Y_c_473_n N_Y_c_490_n Y
+ PM_SKY130_FD_SC_HD__O221AI_2%Y
x_PM_SKY130_FD_SC_HD__O221AI_2%A_382_297# N_A_382_297#_M1007_s
+ N_A_382_297#_M1013_d N_A_382_297#_c_526_n N_A_382_297#_c_532_n
+ N_A_382_297#_c_534_n PM_SKY130_FD_SC_HD__O221AI_2%A_382_297#
x_PM_SKY130_FD_SC_HD__O221AI_2%A_734_297# N_A_734_297#_M1011_d
+ N_A_734_297#_M1018_d N_A_734_297#_c_548_n N_A_734_297#_c_547_n
+ N_A_734_297#_c_554_n PM_SKY130_FD_SC_HD__O221AI_2%A_734_297#
x_PM_SKY130_FD_SC_HD__O221AI_2%A_28_47# N_A_28_47#_M1005_d N_A_28_47#_M1008_d
+ N_A_28_47#_M1006_s N_A_28_47#_M1001_d N_A_28_47#_c_561_n N_A_28_47#_c_562_n
+ N_A_28_47#_c_569_n N_A_28_47#_c_563_n N_A_28_47#_c_564_n N_A_28_47#_c_565_n
+ PM_SKY130_FD_SC_HD__O221AI_2%A_28_47#
x_PM_SKY130_FD_SC_HD__O221AI_2%A_300_47# N_A_300_47#_M1006_d N_A_300_47#_M1000_s
+ N_A_300_47#_M1016_d N_A_300_47#_M1017_s N_A_300_47#_M1003_s
+ N_A_300_47#_c_610_n N_A_300_47#_c_624_n N_A_300_47#_c_625_n
+ N_A_300_47#_c_611_n N_A_300_47#_c_612_n N_A_300_47#_c_633_n
+ N_A_300_47#_c_613_n N_A_300_47#_c_614_n N_A_300_47#_c_615_n
+ PM_SKY130_FD_SC_HD__O221AI_2%A_300_47#
x_PM_SKY130_FD_SC_HD__O221AI_2%VGND N_VGND_M1002_d N_VGND_M1019_d N_VGND_c_683_n
+ N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ VGND N_VGND_c_689_n N_VGND_c_690_n PM_SKY130_FD_SC_HD__O221AI_2%VGND
cc_1 VNB N_C1_c_87_n 0.021691f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_C1_c_88_n 0.0209917f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_3 VNB C1 0.00869944f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_C1_c_90_n 0.0603133f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.16
cc_5 VNB N_B1_c_128_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_6 VNB N_B1_c_129_n 0.0170683f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_7 VNB N_B1_c_130_n 0.00349127f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_8 VNB N_B1_c_131_n 0.0196886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_132_n 0.0118806f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.16
cc_10 VNB N_B1_c_133_n 0.0259565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B1_c_134_n 0.00215682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B2_c_210_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_13 VNB N_B2_c_211_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_14 VNB B2 0.00141292f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_B2_c_213_n 0.0299865f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.16
cc_16 VNB N_A1_c_251_n 0.0169197f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_17 VNB N_A1_c_252_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_18 VNB N_A1_c_253_n 0.00358781f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_19 VNB N_A1_c_254_n 0.0192897f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_20 VNB N_A1_c_255_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A1_c_256_n 0.00189758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB A1 0.0298833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_c_258_n 0.0265824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A2_c_337_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_25 VNB N_A2_c_338_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_26 VNB N_A2_c_339_n 0.0313072f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.16
cc_27 VNB N_VPWR_c_385_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_458_n 0.00100968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_28_47#_c_561_n 0.0095692f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.985
cc_30 VNB N_A_28_47#_c_562_n 0.0173145f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_31 VNB N_A_28_47#_c_563_n 0.00225907f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_32 VNB N_A_28_47#_c_564_n 0.00547341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_28_47#_c_565_n 0.0180191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_300_47#_c_610_n 0.00262034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_300_47#_c_611_n 0.00332606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_300_47#_c_612_n 0.00807318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_300_47#_c_613_n 0.0132865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_300_47#_c_614_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_300_47#_c_615_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_683_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.56
cc_41 VNB N_VGND_c_684_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.985
cc_42 VNB N_VGND_c_685_n 0.0875329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_686_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_44 VNB N_VGND_c_687_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_45 VNB N_VGND_c_688_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_689_n 0.0234308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_690_n 0.287693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VPB N_C1_M1004_g 0.025159f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_49 VPB N_C1_M1010_g 0.0211808f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_50 VPB N_C1_c_90_n 0.0142791f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.16
cc_51 VPB N_B1_M1007_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_52 VPB N_B1_M1015_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_53 VPB N_B1_c_137_n 0.00723927f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_54 VPB N_B1_c_130_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_55 VPB N_B1_c_131_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_B1_c_132_n 0.00432715f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.16
cc_57 VPB N_B1_c_133_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_B1_c_134_n 0.00156682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B2_M1009_g 0.0183345f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_60 VPB N_B2_M1013_g 0.0183375f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_61 VPB N_B2_c_213_n 0.00400361f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.16
cc_62 VPB N_A1_M1011_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_63 VPB N_A1_M1012_g 0.0245822f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_64 VPB N_A1_c_253_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_65 VPB N_A1_c_254_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_66 VPB N_A1_c_263_n 0.00689724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A1_c_264_n 2.50157e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.16
cc_68 VPB N_A1_c_255_n 0.00130531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A1_c_258_n 0.00655427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A2_M1014_g 0.0183373f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_71 VPB N_A2_M1018_g 0.0183337f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_72 VPB N_A2_c_339_n 0.00400351f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.16
cc_73 VPB N_VPWR_c_386_n 0.0114496f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_74 VPB N_VPWR_c_387_n 0.00760733f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_75 VPB N_VPWR_c_388_n 0.00561441f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.16
cc_76 VPB N_VPWR_c_389_n 0.00830908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_390_n 0.0363617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_391_n 0.00391723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_392_n 0.0349357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_393_n 0.0126445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_385_n 0.0538809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_395_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_396_n 0.0222705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_397_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_Y_c_459_n 8.73568e-19 $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_86 VPB N_Y_c_458_n 0.0011304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 N_C1_c_90_n N_B1_c_132_n 0.0140117f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_88 N_C1_M1004_g N_VPWR_c_387_n 0.00408087f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_89 C1 N_VPWR_c_387_n 0.0193718f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_90 N_C1_c_90_n N_VPWR_c_387_n 0.00610779f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_91 N_C1_M1004_g N_VPWR_c_385_n 0.0113957f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_92 N_C1_M1010_g N_VPWR_c_385_n 0.00720795f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_93 N_C1_M1004_g N_VPWR_c_395_n 0.00585385f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_94 N_C1_M1010_g N_VPWR_c_395_n 0.00585385f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_95 N_C1_M1010_g N_VPWR_c_396_n 0.00353572f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_96 N_C1_M1004_g N_Y_c_459_n 5.13163e-19 $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_97 N_C1_M1010_g N_Y_c_459_n 0.00196368f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_98 N_C1_M1010_g N_Y_c_463_n 0.00758424f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_99 N_C1_c_87_n N_Y_c_464_n 0.00407862f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_100 N_C1_c_88_n N_Y_c_464_n 0.00281475f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_101 N_C1_c_87_n N_Y_c_458_n 0.00262178f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_102 N_C1_M1004_g N_Y_c_458_n 0.00302963f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_103 N_C1_c_88_n N_Y_c_458_n 0.00513669f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_104 N_C1_M1010_g N_Y_c_458_n 0.00232215f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_105 C1 N_Y_c_458_n 0.0146705f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_106 N_C1_c_90_n N_Y_c_458_n 0.0254224f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_107 N_C1_M1010_g N_Y_c_472_n 0.00117879f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_108 N_C1_M1010_g N_Y_c_473_n 0.0138008f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_109 N_C1_c_87_n N_A_28_47#_c_562_n 2.32395e-19 $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_110 C1 N_A_28_47#_c_562_n 0.0192857f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_111 N_C1_c_90_n N_A_28_47#_c_562_n 0.00621075f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C1_c_87_n N_A_28_47#_c_569_n 0.012123f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_113 N_C1_c_88_n N_A_28_47#_c_569_n 0.0127333f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_114 C1 N_A_28_47#_c_569_n 0.00146328f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_115 N_C1_c_90_n N_A_28_47#_c_569_n 3.07604e-19 $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C1_c_88_n N_A_28_47#_c_564_n 4.59762e-19 $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C1_c_87_n N_VGND_c_685_n 0.00357877f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_118 N_C1_c_88_n N_VGND_c_685_n 0.00357877f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_119 N_C1_c_87_n N_VGND_c_690_n 0.00618415f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_120 N_C1_c_88_n N_VGND_c_690_n 0.00655123f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_128_n N_B2_c_210_n 0.0270078f $X=1.835 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_122 N_B1_M1007_g N_B2_M1009_g 0.0439701f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_c_137_n N_B2_M1009_g 0.0106267f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_124 N_B1_c_129_n N_B2_c_211_n 0.0267413f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B1_M1015_g N_B2_M1013_g 0.0440009f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_c_137_n N_B2_M1013_g 0.0103235f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_127 N_B1_c_137_n B2 0.0391837f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_128 N_B1_c_130_n B2 0.0172311f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B1_c_131_n B2 6.66616e-19 $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B1_c_133_n B2 2.07308e-19 $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B1_c_134_n B2 0.0173969f $X=2.035 $Y=1.345 $X2=0 $Y2=0
cc_132 N_B1_c_137_n N_B2_c_213_n 0.00214031f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_133 N_B1_c_130_n N_B2_c_213_n 0.00458063f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B1_c_131_n N_B2_c_213_n 0.0223771f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B1_c_133_n N_B2_c_213_n 0.0223199f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B1_c_134_n N_B2_c_213_n 0.00620106f $X=2.035 $Y=1.345 $X2=0 $Y2=0
cc_137 N_B1_c_129_n N_A1_c_251_n 0.00937759f $X=3.095 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_138 N_B1_M1015_g N_A1_M1011_g 0.0387452f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B1_c_137_n N_A1_M1011_g 5.77655e-19 $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_140 N_B1_c_130_n N_A1_M1011_g 3.59226e-19 $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B1_M1015_g N_A1_c_253_n 3.59226e-19 $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B1_c_130_n N_A1_c_253_n 0.0307171f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B1_c_131_n N_A1_c_253_n 7.80994e-19 $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B1_c_130_n N_A1_c_254_n 7.80994e-19 $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B1_c_131_n N_A1_c_254_n 0.0197715f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B1_M1015_g N_A1_c_264_n 5.77655e-19 $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_147 N_B1_c_137_n N_A1_c_264_n 0.0154679f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_148 N_B1_c_132_n N_VPWR_M1010_d 0.0112782f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_149 N_B1_c_137_n N_VPWR_M1015_d 0.00151212f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_150 N_B1_M1015_g N_VPWR_c_388_n 0.00323788f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B1_M1007_g N_VPWR_c_392_n 0.00585385f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B1_M1015_g N_VPWR_c_392_n 0.00585385f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B1_M1007_g N_VPWR_c_385_n 0.00723564f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B1_M1015_g N_VPWR_c_385_n 0.0061234f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B1_M1007_g N_VPWR_c_396_n 0.00518337f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B1_c_137_n N_Y_M1009_s 0.00165831f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B1_M1015_g N_Y_c_475_n 0.0119464f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_158 N_B1_c_137_n N_Y_c_475_n 0.0355123f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B1_c_131_n N_Y_c_475_n 3.01349e-19 $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B1_c_132_n N_Y_c_458_n 0.0384493f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_161 N_B1_c_137_n N_Y_c_479_n 0.0120079f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_162 N_B1_M1007_g N_Y_c_473_n 0.0136605f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_163 N_B1_c_132_n N_Y_c_473_n 0.0867304f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_164 N_B1_c_133_n N_Y_c_473_n 3.01392e-19 $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_137_n N_A_382_297#_M1007_s 9.27081e-19 $X=2.93 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_166 N_B1_c_134_n N_A_382_297#_M1007_s 7.50819e-19 $X=2.035 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_167 N_B1_c_137_n N_A_382_297#_M1013_d 0.00165255f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_168 N_B1_c_128_n N_A_28_47#_c_564_n 0.00300006f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B1_c_132_n N_A_28_47#_c_564_n 0.0228439f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_170 N_B1_c_128_n N_A_28_47#_c_565_n 0.0141874f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B1_c_129_n N_A_28_47#_c_565_n 0.00375446f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_137_n N_A_28_47#_c_565_n 0.0116483f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_173 N_B1_c_130_n N_A_28_47#_c_565_n 0.00964534f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_c_131_n N_A_28_47#_c_565_n 0.00149384f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B1_c_132_n N_A_28_47#_c_565_n 0.0631652f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_176 N_B1_c_133_n N_A_28_47#_c_565_n 0.00298952f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B1_c_128_n N_A_300_47#_c_610_n 0.00886996f $X=1.835 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_B1_c_129_n N_A_300_47#_c_610_n 0.0105068f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B1_c_130_n N_A_300_47#_c_610_n 0.00390962f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_c_129_n N_A_300_47#_c_612_n 2.00828e-19 $X=3.095 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_B1_c_130_n N_A_300_47#_c_612_n 0.00353546f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B1_c_131_n N_A_300_47#_c_612_n 2.55742e-19 $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B1_c_128_n N_VGND_c_685_n 0.00357877f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_c_129_n N_VGND_c_685_n 0.00357877f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B1_c_128_n N_VGND_c_690_n 0.00657948f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_129_n N_VGND_c_690_n 0.00546478f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B2_M1009_g N_VPWR_c_392_n 0.00357877f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B2_M1013_g N_VPWR_c_392_n 0.00357877f $X=2.675 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B2_M1009_g N_VPWR_c_385_n 0.00525237f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B2_M1013_g N_VPWR_c_385_n 0.00525237f $X=2.675 $Y=1.985 $X2=0 $Y2=0
cc_191 N_B2_M1013_g N_Y_c_475_n 0.00924026f $X=2.675 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B2_M1009_g N_Y_c_473_n 0.00924026f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B2_M1009_g N_A_382_297#_c_526_n 0.00851673f $X=2.255 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_B2_M1013_g N_A_382_297#_c_526_n 0.00851673f $X=2.675 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_B2_c_210_n N_A_28_47#_c_565_n 0.0112673f $X=2.255 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B2_c_211_n N_A_28_47#_c_565_n 0.0109578f $X=2.675 $Y=0.995 $X2=0 $Y2=0
cc_197 B2 N_A_28_47#_c_565_n 0.0405144f $X=2.465 $Y=1.105 $X2=0 $Y2=0
cc_198 N_B2_c_213_n N_A_28_47#_c_565_n 0.00224214f $X=2.675 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B2_c_210_n N_A_300_47#_c_610_n 0.00886996f $X=2.255 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_B2_c_211_n N_A_300_47#_c_610_n 0.00886996f $X=2.675 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_B2_c_210_n N_VGND_c_685_n 0.00357877f $X=2.255 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B2_c_211_n N_VGND_c_685_n 0.00357877f $X=2.675 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B2_c_210_n N_VGND_c_690_n 0.00525341f $X=2.255 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B2_c_211_n N_VGND_c_690_n 0.00525341f $X=2.675 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A1_c_251_n N_A2_c_337_n 0.0258191f $X=3.595 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A1_M1011_g N_A2_M1014_g 0.0440009f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A1_c_263_n N_A2_M1014_g 0.0108086f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_208 N_A1_c_252_n N_A2_c_338_n 0.0258694f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_M1012_g N_A2_M1018_g 0.0270786f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A1_c_263_n N_A2_M1018_g 0.0153291f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_211 N_A1_c_253_n A2 0.0133594f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A1_c_254_n A2 2.2122e-19 $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A1_c_263_n A2 0.0349894f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_214 N_A1_c_256_n A2 0.0172564f $X=4.815 $Y=1.175 $X2=0 $Y2=0
cc_215 N_A1_c_258_n A2 2.00336e-19 $X=4.855 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A1_c_253_n N_A2_c_339_n 0.00527477f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A1_c_254_n N_A2_c_339_n 0.022397f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A1_c_263_n N_A2_c_339_n 0.00214031f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_219 N_A1_c_255_n N_A2_c_339_n 0.00362491f $X=4.73 $Y=1.445 $X2=0 $Y2=0
cc_220 N_A1_c_256_n N_A2_c_339_n 0.00144374f $X=4.815 $Y=1.175 $X2=0 $Y2=0
cc_221 N_A1_c_258_n N_A2_c_339_n 0.0222902f $X=4.855 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A1_c_264_n N_VPWR_M1015_d 0.00151212f $X=3.76 $Y=1.53 $X2=0 $Y2=0
cc_223 N_A1_M1011_g N_VPWR_c_388_n 0.00525229f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A1_M1012_g N_VPWR_c_389_n 0.00505805f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A1_c_263_n N_VPWR_c_389_n 0.00786716f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_226 A1 N_VPWR_c_389_n 0.0166332f $X=5.225 $Y=1.105 $X2=0 $Y2=0
cc_227 N_A1_M1011_g N_VPWR_c_390_n 0.00585385f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A1_M1012_g N_VPWR_c_390_n 0.00585385f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A1_M1011_g N_VPWR_c_385_n 0.00617642f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_M1012_g N_VPWR_c_385_n 0.0116728f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_c_263_n N_Y_M1014_s 0.00165831f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_232 N_A1_M1011_g N_Y_c_475_n 0.0119464f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_c_254_n N_Y_c_475_n 3.01349e-19 $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A1_c_263_n N_Y_c_475_n 0.0190307f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_235 N_A1_c_264_n N_Y_c_475_n 0.0164816f $X=3.76 $Y=1.53 $X2=0 $Y2=0
cc_236 N_A1_c_263_n N_Y_c_490_n 0.0120079f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_237 N_A1_c_263_n N_A_734_297#_M1011_d 0.00130005f $X=4.645 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_238 N_A1_c_264_n N_A_734_297#_M1011_d 3.52503e-19 $X=3.76 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_239 N_A1_c_263_n N_A_734_297#_M1018_d 0.00167564f $X=4.645 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A1_c_263_n N_A_734_297#_c_547_n 0.0132239f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_241 N_A1_c_251_n N_A_300_47#_c_624_n 0.00255288f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A1_c_251_n N_A_300_47#_c_625_n 0.00393886f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A1_c_251_n N_A_300_47#_c_611_n 0.00845282f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A1_c_253_n N_A_300_47#_c_611_n 0.0160434f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A1_c_254_n N_A_300_47#_c_611_n 0.001478f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A1_c_263_n N_A_300_47#_c_611_n 0.0071189f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_247 N_A1_c_251_n N_A_300_47#_c_612_n 0.00111376f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A1_c_253_n N_A_300_47#_c_612_n 0.010391f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A1_c_254_n N_A_300_47#_c_612_n 0.00153445f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A1_c_251_n N_A_300_47#_c_633_n 5.22228e-19 $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A1_c_252_n N_A_300_47#_c_633_n 5.22228e-19 $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A1_c_252_n N_A_300_47#_c_613_n 0.00995081f $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A1_c_263_n N_A_300_47#_c_613_n 0.00549032f $X=4.645 $Y=1.53 $X2=0 $Y2=0
cc_254 N_A1_c_256_n N_A_300_47#_c_613_n 0.0135931f $X=4.815 $Y=1.175 $X2=0 $Y2=0
cc_255 A1 N_A_300_47#_c_613_n 0.0333889f $X=5.225 $Y=1.105 $X2=0 $Y2=0
cc_256 N_A1_c_258_n N_A_300_47#_c_613_n 0.00301563f $X=4.855 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A1_c_252_n N_A_300_47#_c_614_n 0.00630972f $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A1_c_251_n N_VGND_c_683_n 0.00268723f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_252_n N_VGND_c_684_n 0.00268723f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A1_c_251_n N_VGND_c_685_n 0.00422898f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A1_c_252_n N_VGND_c_689_n 0.00423334f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A1_c_251_n N_VGND_c_690_n 0.00598371f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_c_252_n N_VGND_c_690_n 0.00683939f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A2_M1014_g N_VPWR_c_390_n 0.00357877f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A2_M1018_g N_VPWR_c_390_n 0.00357877f $X=4.435 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A2_M1014_g N_VPWR_c_385_n 0.00525237f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A2_M1018_g N_VPWR_c_385_n 0.00525237f $X=4.435 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A2_M1014_g N_Y_c_475_n 0.00924026f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A2_M1014_g N_A_734_297#_c_548_n 0.00851673f $X=4.015 $Y=1.985 $X2=0
+ $Y2=0
cc_270 N_A2_M1018_g N_A_734_297#_c_548_n 0.0121306f $X=4.435 $Y=1.985 $X2=0
+ $Y2=0
cc_271 N_A2_c_337_n N_A_300_47#_c_625_n 4.86433e-19 $X=4.015 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A2_c_337_n N_A_300_47#_c_611_n 0.00894278f $X=4.015 $Y=0.995 $X2=0
+ $Y2=0
cc_273 A2 N_A_300_47#_c_611_n 0.00545718f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_274 N_A2_c_337_n N_A_300_47#_c_633_n 0.00630972f $X=4.015 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A2_c_338_n N_A_300_47#_c_633_n 0.00630972f $X=4.435 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A2_c_338_n N_A_300_47#_c_613_n 0.00908248f $X=4.435 $Y=0.995 $X2=0
+ $Y2=0
cc_277 A2 N_A_300_47#_c_613_n 0.00582553f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_278 N_A2_c_338_n N_A_300_47#_c_614_n 5.22228e-19 $X=4.435 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A2_c_337_n N_A_300_47#_c_615_n 0.00128009f $X=4.015 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A2_c_338_n N_A_300_47#_c_615_n 0.00113286f $X=4.435 $Y=0.995 $X2=0
+ $Y2=0
cc_281 A2 N_A_300_47#_c_615_n 0.0265405f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_282 N_A2_c_339_n N_A_300_47#_c_615_n 0.00230339f $X=4.435 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A2_c_337_n N_VGND_c_683_n 0.00146448f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A2_c_338_n N_VGND_c_684_n 0.00146448f $X=4.435 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A2_c_337_n N_VGND_c_687_n 0.00424416f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A2_c_338_n N_VGND_c_687_n 0.00423334f $X=4.435 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A2_c_337_n N_VGND_c_690_n 0.00576327f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A2_c_338_n N_VGND_c_690_n 0.0057435f $X=4.435 $Y=0.995 $X2=0 $Y2=0
cc_289 N_VPWR_c_385_n N_Y_M1004_s 0.00254112f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_c_385_n N_Y_M1009_s 0.00215227f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_c_385_n N_Y_M1014_s 0.0021603f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_387_n N_Y_c_459_n 0.00234f $X=0.265 $Y=1.65 $X2=0 $Y2=0
cc_293 N_VPWR_c_385_n N_Y_c_496_n 0.00955092f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_395_n N_Y_c_496_n 0.0142343f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_295 N_VPWR_M1015_d N_Y_c_475_n 0.0095835f $X=3.17 $Y=1.485 $X2=0 $Y2=0
cc_296 N_VPWR_c_388_n N_Y_c_475_n 0.0186532f $X=3.305 $Y=2.3 $X2=0 $Y2=0
cc_297 N_VPWR_c_385_n N_Y_c_475_n 0.0130817f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_c_385_n N_Y_c_472_n 0.00134725f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_M1010_d N_Y_c_473_n 0.0182311f $X=0.97 $Y=1.485 $X2=0 $Y2=0
cc_300 N_VPWR_c_385_n N_Y_c_473_n 0.0125007f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_396_n N_Y_c_473_n 0.0531577f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_302 N_VPWR_c_385_n N_A_382_297#_M1007_s 0.00219968f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_303 N_VPWR_c_385_n N_A_382_297#_M1013_d 0.00219968f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_392_n N_A_382_297#_c_526_n 0.0330174f $X=3.18 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_385_n N_A_382_297#_c_526_n 0.0204707f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_392_n N_A_382_297#_c_532_n 0.0137033f $X=3.18 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_385_n N_A_382_297#_c_532_n 0.00938745f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_392_n N_A_382_297#_c_534_n 0.0137033f $X=3.18 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_385_n N_A_382_297#_c_534_n 0.00938745f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_385_n N_A_734_297#_M1011_d 0.00219968f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_311 N_VPWR_c_385_n N_A_734_297#_M1018_d 0.00246446f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_390_n N_A_734_297#_c_548_n 0.0473226f $X=4.985 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_385_n N_A_734_297#_c_548_n 0.0300947f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_390_n N_A_734_297#_c_554_n 0.0137033f $X=4.985 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_385_n N_A_734_297#_c_554_n 0.00938745f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_Y_c_473_n N_A_382_297#_M1007_s 0.00325599f $X=2.34 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_317 N_Y_c_475_n N_A_382_297#_M1013_d 0.00325521f $X=4.1 $Y=1.87 $X2=0 $Y2=0
cc_318 N_Y_M1009_s N_A_382_297#_c_526_n 0.00312348f $X=2.33 $Y=1.485 $X2=0 $Y2=0
cc_319 N_Y_c_475_n N_A_382_297#_c_526_n 0.00506389f $X=4.1 $Y=1.87 $X2=0 $Y2=0
cc_320 N_Y_c_479_n N_A_382_297#_c_526_n 0.0112811f $X=2.465 $Y=1.87 $X2=0 $Y2=0
cc_321 N_Y_c_473_n N_A_382_297#_c_526_n 0.00506389f $X=2.34 $Y=1.87 $X2=0 $Y2=0
cc_322 N_Y_c_473_n N_A_382_297#_c_532_n 0.0116461f $X=2.34 $Y=1.87 $X2=0 $Y2=0
cc_323 N_Y_c_475_n N_A_382_297#_c_534_n 0.0116461f $X=4.1 $Y=1.87 $X2=0 $Y2=0
cc_324 N_Y_c_475_n N_A_734_297#_M1011_d 0.00325521f $X=4.1 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_325 N_Y_M1014_s N_A_734_297#_c_548_n 0.00312348f $X=4.09 $Y=1.485 $X2=0 $Y2=0
cc_326 N_Y_c_475_n N_A_734_297#_c_548_n 0.00506389f $X=4.1 $Y=1.87 $X2=0 $Y2=0
cc_327 N_Y_c_490_n N_A_734_297#_c_548_n 0.0112811f $X=4.225 $Y=1.87 $X2=0 $Y2=0
cc_328 N_Y_c_475_n N_A_734_297#_c_554_n 0.0116461f $X=4.1 $Y=1.87 $X2=0 $Y2=0
cc_329 N_Y_c_458_n N_A_28_47#_c_562_n 5.40026e-19 $X=0.705 $Y=1.445 $X2=0 $Y2=0
cc_330 N_Y_M1005_s N_A_28_47#_c_569_n 0.00304656f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_331 N_Y_c_464_n N_A_28_47#_c_569_n 0.0162479f $X=0.685 $Y=0.73 $X2=0 $Y2=0
cc_332 N_Y_c_464_n N_A_28_47#_c_564_n 0.0105846f $X=0.685 $Y=0.73 $X2=0 $Y2=0
cc_333 N_Y_M1005_s N_VGND_c_690_n 0.00216833f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_334 N_A_28_47#_c_565_n N_A_300_47#_M1006_d 0.0031705f $X=2.885 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_335 N_A_28_47#_c_565_n N_A_300_47#_M1000_s 0.00162317f $X=2.885 $Y=0.73 $X2=0
+ $Y2=0
cc_336 N_A_28_47#_M1006_s N_A_300_47#_c_610_n 0.00312026f $X=1.91 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_A_28_47#_M1001_d N_A_300_47#_c_610_n 0.00312026f $X=2.75 $Y=0.235 $X2=0
+ $Y2=0
cc_338 N_A_28_47#_c_563_n N_A_300_47#_c_610_n 0.0188707f $X=1.145 $Y=0.475 $X2=0
+ $Y2=0
cc_339 N_A_28_47#_c_565_n N_A_300_47#_c_610_n 0.0840906f $X=2.885 $Y=0.73 $X2=0
+ $Y2=0
cc_340 N_A_28_47#_c_565_n N_A_300_47#_c_612_n 0.00799569f $X=2.885 $Y=0.73 $X2=0
+ $Y2=0
cc_341 N_A_28_47#_c_561_n N_VGND_c_685_n 0.0173151f $X=0.225 $Y=0.475 $X2=0
+ $Y2=0
cc_342 N_A_28_47#_c_569_n N_VGND_c_685_n 0.0363282f $X=1.02 $Y=0.365 $X2=0 $Y2=0
cc_343 N_A_28_47#_c_563_n N_VGND_c_685_n 0.0173343f $X=1.145 $Y=0.475 $X2=0
+ $Y2=0
cc_344 N_A_28_47#_c_565_n N_VGND_c_685_n 0.00349681f $X=2.885 $Y=0.73 $X2=0
+ $Y2=0
cc_345 N_A_28_47#_M1005_d N_VGND_c_690_n 0.00209324f $X=0.14 $Y=0.235 $X2=0
+ $Y2=0
cc_346 N_A_28_47#_M1008_d N_VGND_c_690_n 0.00209324f $X=0.97 $Y=0.235 $X2=0
+ $Y2=0
cc_347 N_A_28_47#_M1006_s N_VGND_c_690_n 0.00216833f $X=1.91 $Y=0.235 $X2=0
+ $Y2=0
cc_348 N_A_28_47#_M1001_d N_VGND_c_690_n 0.00216833f $X=2.75 $Y=0.235 $X2=0
+ $Y2=0
cc_349 N_A_28_47#_c_561_n N_VGND_c_690_n 0.00961275f $X=0.225 $Y=0.475 $X2=0
+ $Y2=0
cc_350 N_A_28_47#_c_569_n N_VGND_c_690_n 0.023578f $X=1.02 $Y=0.365 $X2=0 $Y2=0
cc_351 N_A_28_47#_c_563_n N_VGND_c_690_n 0.00961652f $X=1.145 $Y=0.475 $X2=0
+ $Y2=0
cc_352 N_A_28_47#_c_565_n N_VGND_c_690_n 0.00853783f $X=2.885 $Y=0.73 $X2=0
+ $Y2=0
cc_353 N_A_300_47#_c_611_n N_VGND_M1002_d 0.00165819f $X=4.06 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_354 N_A_300_47#_c_613_n N_VGND_M1019_d 0.00162089f $X=4.9 $Y=0.815 $X2=0
+ $Y2=0
cc_355 N_A_300_47#_c_611_n N_VGND_c_683_n 0.0116528f $X=4.06 $Y=0.82 $X2=0 $Y2=0
cc_356 N_A_300_47#_c_613_n N_VGND_c_684_n 0.0122559f $X=4.9 $Y=0.815 $X2=0 $Y2=0
cc_357 N_A_300_47#_c_610_n N_VGND_c_685_n 0.0991765f $X=3.22 $Y=0.365 $X2=0
+ $Y2=0
cc_358 N_A_300_47#_c_624_n N_VGND_c_685_n 0.0208178f $X=3.385 $Y=0.475 $X2=0
+ $Y2=0
cc_359 N_A_300_47#_c_611_n N_VGND_c_685_n 0.00193763f $X=4.06 $Y=0.82 $X2=0
+ $Y2=0
cc_360 N_A_300_47#_c_611_n N_VGND_c_687_n 0.00193763f $X=4.06 $Y=0.82 $X2=0
+ $Y2=0
cc_361 N_A_300_47#_c_633_n N_VGND_c_687_n 0.0188551f $X=4.225 $Y=0.39 $X2=0
+ $Y2=0
cc_362 N_A_300_47#_c_613_n N_VGND_c_687_n 0.00198695f $X=4.9 $Y=0.815 $X2=0
+ $Y2=0
cc_363 N_A_300_47#_c_613_n N_VGND_c_689_n 0.00198695f $X=4.9 $Y=0.815 $X2=0
+ $Y2=0
cc_364 N_A_300_47#_c_614_n N_VGND_c_689_n 0.0209752f $X=5.065 $Y=0.39 $X2=0
+ $Y2=0
cc_365 N_A_300_47#_M1006_d N_VGND_c_690_n 0.00209344f $X=1.5 $Y=0.235 $X2=0
+ $Y2=0
cc_366 N_A_300_47#_M1000_s N_VGND_c_690_n 0.00215227f $X=2.33 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_300_47#_M1016_d N_VGND_c_690_n 0.00279445f $X=3.17 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_300_47#_M1017_s N_VGND_c_690_n 0.00215201f $X=4.09 $Y=0.235 $X2=0
+ $Y2=0
cc_369 N_A_300_47#_M1003_s N_VGND_c_690_n 0.00209319f $X=4.93 $Y=0.235 $X2=0
+ $Y2=0
cc_370 N_A_300_47#_c_610_n N_VGND_c_690_n 0.0628989f $X=3.22 $Y=0.365 $X2=0
+ $Y2=0
cc_371 N_A_300_47#_c_624_n N_VGND_c_690_n 0.0124843f $X=3.385 $Y=0.475 $X2=0
+ $Y2=0
cc_372 N_A_300_47#_c_611_n N_VGND_c_690_n 0.00827287f $X=4.06 $Y=0.82 $X2=0
+ $Y2=0
cc_373 N_A_300_47#_c_633_n N_VGND_c_690_n 0.0122069f $X=4.225 $Y=0.39 $X2=0
+ $Y2=0
cc_374 N_A_300_47#_c_613_n N_VGND_c_690_n 0.00835832f $X=4.9 $Y=0.815 $X2=0
+ $Y2=0
cc_375 N_A_300_47#_c_614_n N_VGND_c_690_n 0.0124119f $X=5.065 $Y=0.39 $X2=0
+ $Y2=0

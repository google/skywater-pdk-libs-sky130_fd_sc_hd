* File: sky130_fd_sc_hd__o221ai_4.spice.SKY130_FD_SC_HD__O221AI_4.pxi
* Created: Thu Aug 27 14:37:23 2020
* 
x_PM_SKY130_FD_SC_HD__O221AI_4%C1 N_C1_c_125_n N_C1_M1013_g N_C1_M1010_g
+ N_C1_c_126_n N_C1_M1018_g N_C1_M1029_g N_C1_c_127_n N_C1_M1026_g N_C1_M1032_g
+ N_C1_c_128_n N_C1_M1027_g N_C1_M1036_g C1 N_C1_c_129_n N_C1_c_130_n
+ PM_SKY130_FD_SC_HD__O221AI_4%C1
x_PM_SKY130_FD_SC_HD__O221AI_4%B1 N_B1_c_184_n N_B1_M1003_g N_B1_M1001_g
+ N_B1_c_185_n N_B1_M1011_g N_B1_M1007_g N_B1_c_186_n N_B1_M1019_g N_B1_M1023_g
+ N_B1_c_187_n N_B1_M1038_g N_B1_M1025_g N_B1_c_196_n N_B1_c_206_p N_B1_c_204_p
+ N_B1_c_188_n N_B1_c_189_n N_B1_c_190_n B1 N_B1_c_191_n
+ PM_SKY130_FD_SC_HD__O221AI_4%B1
x_PM_SKY130_FD_SC_HD__O221AI_4%B2 N_B2_c_295_n N_B2_M1004_g N_B2_M1008_g
+ N_B2_c_296_n N_B2_M1014_g N_B2_M1012_g N_B2_c_297_n N_B2_M1016_g N_B2_M1033_g
+ N_B2_c_298_n N_B2_M1020_g N_B2_M1037_g B2 N_B2_c_299_n N_B2_c_300_n
+ PM_SKY130_FD_SC_HD__O221AI_4%B2
x_PM_SKY130_FD_SC_HD__O221AI_4%A1 N_A1_c_370_n N_A1_M1005_g N_A1_M1015_g
+ N_A1_c_371_n N_A1_M1017_g N_A1_M1024_g N_A1_c_372_n N_A1_M1022_g N_A1_M1030_g
+ N_A1_c_373_n N_A1_M1028_g N_A1_M1035_g N_A1_c_374_n N_A1_c_375_n N_A1_c_385_n
+ N_A1_c_386_n N_A1_c_376_n N_A1_c_387_n A1 N_A1_c_377_n N_A1_c_378_n
+ PM_SKY130_FD_SC_HD__O221AI_4%A1
x_PM_SKY130_FD_SC_HD__O221AI_4%A2 N_A2_c_498_n N_A2_M1000_g N_A2_M1002_g
+ N_A2_c_499_n N_A2_M1006_g N_A2_M1031_g N_A2_c_500_n N_A2_M1009_g N_A2_M1034_g
+ N_A2_c_501_n N_A2_M1021_g N_A2_M1039_g A2 N_A2_c_516_n N_A2_c_502_n
+ PM_SKY130_FD_SC_HD__O221AI_4%A2
x_PM_SKY130_FD_SC_HD__O221AI_4%VPWR N_VPWR_M1010_s N_VPWR_M1029_s N_VPWR_M1036_s
+ N_VPWR_M1007_d N_VPWR_M1025_d N_VPWR_M1024_s N_VPWR_M1035_s N_VPWR_c_582_n
+ N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n
+ N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_592_n
+ N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n VPWR N_VPWR_c_596_n
+ N_VPWR_c_597_n N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_581_n
+ PM_SKY130_FD_SC_HD__O221AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O221AI_4%Y N_Y_M1013_d N_Y_M1026_d N_Y_M1010_d N_Y_M1032_d
+ N_Y_M1008_s N_Y_M1033_s N_Y_M1002_d N_Y_M1034_d N_Y_c_717_n N_Y_c_791_n
+ N_Y_c_719_n N_Y_c_793_n N_Y_c_718_n N_Y_c_721_n N_Y_c_753_n N_Y_c_755_n
+ N_Y_c_757_n N_Y_c_776_n N_Y_c_760_n N_Y_c_722_n N_Y_c_723_n N_Y_c_762_n
+ N_Y_c_763_n N_Y_c_781_n Y PM_SKY130_FD_SC_HD__O221AI_4%Y
x_PM_SKY130_FD_SC_HD__O221AI_4%A_553_297# N_A_553_297#_M1001_s
+ N_A_553_297#_M1023_s N_A_553_297#_M1012_d N_A_553_297#_M1037_d
+ N_A_553_297#_c_862_n N_A_553_297#_c_849_n N_A_553_297#_c_876_n
+ N_A_553_297#_c_867_n N_A_553_297#_c_852_n N_A_553_297#_c_880_n
+ N_A_553_297#_c_851_n N_A_553_297#_c_856_n
+ PM_SKY130_FD_SC_HD__O221AI_4%A_553_297#
x_PM_SKY130_FD_SC_HD__O221AI_4%A_1241_297# N_A_1241_297#_M1015_d
+ N_A_1241_297#_M1031_s N_A_1241_297#_M1039_s N_A_1241_297#_M1030_d
+ N_A_1241_297#_c_903_n N_A_1241_297#_c_905_n N_A_1241_297#_c_891_n
+ N_A_1241_297#_c_896_n N_A_1241_297#_c_886_n N_A_1241_297#_c_919_n
+ N_A_1241_297#_c_902_n N_A_1241_297#_c_923_n
+ PM_SKY130_FD_SC_HD__O221AI_4%A_1241_297#
x_PM_SKY130_FD_SC_HD__O221AI_4%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1018_s
+ N_A_27_47#_M1027_s N_A_27_47#_M1003_d N_A_27_47#_M1019_d N_A_27_47#_M1014_s
+ N_A_27_47#_M1020_s N_A_27_47#_c_935_n N_A_27_47#_c_936_n N_A_27_47#_c_937_n
+ PM_SKY130_FD_SC_HD__O221AI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O221AI_4%A_471_47# N_A_471_47#_M1003_s N_A_471_47#_M1011_s
+ N_A_471_47#_M1004_d N_A_471_47#_M1016_d N_A_471_47#_M1038_s
+ N_A_471_47#_M1000_d N_A_471_47#_M1009_d N_A_471_47#_M1017_s
+ N_A_471_47#_M1028_s N_A_471_47#_c_1008_n N_A_471_47#_c_981_n
+ N_A_471_47#_c_1012_n N_A_471_47#_c_982_n N_A_471_47#_c_1013_n
+ N_A_471_47#_c_983_n N_A_471_47#_c_1017_n N_A_471_47#_c_984_n
+ N_A_471_47#_c_985_n N_A_471_47#_c_986_n N_A_471_47#_c_987_n
+ N_A_471_47#_c_988_n N_A_471_47#_c_989_n N_A_471_47#_c_990_n
+ PM_SKY130_FD_SC_HD__O221AI_4%A_471_47#
x_PM_SKY130_FD_SC_HD__O221AI_4%VGND N_VGND_M1005_d N_VGND_M1006_s N_VGND_M1021_s
+ N_VGND_M1022_d N_VGND_c_1112_n N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n
+ N_VGND_c_1116_n N_VGND_c_1117_n N_VGND_c_1118_n N_VGND_c_1119_n
+ N_VGND_c_1120_n N_VGND_c_1121_n N_VGND_c_1122_n VGND N_VGND_c_1123_n
+ N_VGND_c_1124_n N_VGND_c_1125_n PM_SKY130_FD_SC_HD__O221AI_4%VGND
cc_1 VNB N_C1_c_125_n 0.021723f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_C1_c_126_n 0.0160049f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_C1_c_127_n 0.0160018f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_C1_c_128_n 0.0191948f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_C1_c_129_n 0.0153245f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_6 VNB N_C1_c_130_n 0.0778761f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_B1_c_184_n 0.0199049f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B1_c_185_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_9 VNB N_B1_c_186_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_10 VNB N_B1_c_187_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_11 VNB N_B1_c_188_n 0.00338706f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_12 VNB N_B1_c_189_n 0.0192845f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.16
cc_13 VNB N_B1_c_190_n 0.0114212f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_14 VNB N_B1_c_191_n 0.0534754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B2_c_295_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_16 VNB N_B2_c_296_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_17 VNB N_B2_c_297_n 0.016005f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_18 VNB N_B2_c_298_n 0.0162448f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_19 VNB N_B2_c_299_n 0.00237444f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_20 VNB N_B2_c_300_n 0.0608214f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_21 VNB N_A1_c_370_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_22 VNB N_A1_c_371_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_23 VNB N_A1_c_372_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_24 VNB N_A1_c_373_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_25 VNB N_A1_c_374_n 0.00351686f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_26 VNB N_A1_c_375_n 0.0193115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A1_c_376_n 0.00150905f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.16
cc_28 VNB N_A1_c_377_n 0.0244268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A1_c_378_n 0.0558695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A2_c_498_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_31 VNB N_A2_c_499_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_32 VNB N_A2_c_500_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_33 VNB N_A2_c_501_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_34 VNB N_A2_c_502_n 0.0639937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_581_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_717_n 0.00266041f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.325
cc_37 VNB N_Y_c_718_n 0.0103547f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.175
cc_38 VNB N_A_27_47#_c_935_n 0.00926099f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_39 VNB N_A_27_47#_c_936_n 0.0177907f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_40 VNB N_A_27_47#_c_937_n 0.0115835f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_41 VNB N_A_471_47#_c_981_n 0.00332606f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.175
cc_42 VNB N_A_471_47#_c_982_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_471_47#_c_983_n 0.00406612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_471_47#_c_984_n 0.0124737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_471_47#_c_985_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_471_47#_c_986_n 0.00253999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_471_47#_c_987_n 0.00830265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_471_47#_c_988_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_471_47#_c_989_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_471_47#_c_990_n 0.00222331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1112_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_52 VNB N_VGND_c_1113_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_53 VNB N_VGND_c_1114_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1115_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.325
cc_55 VNB N_VGND_c_1116_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_56 VNB N_VGND_c_1117_n 0.143733f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_57 VNB N_VGND_c_1118_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1119_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_59 VNB N_VGND_c_1120_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_60 VNB N_VGND_c_1121_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_61 VNB N_VGND_c_1122_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.16
cc_62 VNB N_VGND_c_1123_n 0.0210442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1124_n 0.455846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1125_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VPB N_C1_M1010_g 0.0259721f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_66 VPB N_C1_M1029_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_67 VPB N_C1_M1032_g 0.0181172f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_68 VPB N_C1_M1036_g 0.0219547f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_69 VPB N_C1_c_130_n 0.0136143f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_70 VPB N_B1_M1001_g 0.0227299f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_71 VPB N_B1_M1007_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_72 VPB N_B1_M1023_g 0.0184042f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_73 VPB N_B1_M1025_g 0.0181418f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_74 VPB N_B1_c_196_n 0.00158091f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B1_c_188_n 0.00292946f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_76 VPB N_B1_c_189_n 0.00442005f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_77 VPB N_B1_c_191_n 0.00852838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_B2_M1008_g 0.018386f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_79 VPB N_B2_M1012_g 0.0178055f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_80 VPB N_B2_M1033_g 0.0184733f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_81 VPB N_B2_M1037_g 0.0187972f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_82 VPB N_B2_c_300_n 0.010339f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.16
cc_83 VPB N_A1_M1015_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_84 VPB N_A1_M1024_g 0.0178828f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_85 VPB N_A1_M1030_g 0.0184569f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_86 VPB N_A1_M1035_g 0.0249322f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_87 VPB N_A1_c_374_n 0.00233133f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_88 VPB N_A1_c_375_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A1_c_385_n 0.0135863f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_90 VPB N_A1_c_386_n 2.57027e-19 $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_91 VPB N_A1_c_387_n 0.00119441f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.16
cc_92 VPB N_A1_c_378_n 0.00982609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A2_M1002_g 0.0183572f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_94 VPB N_A2_M1031_g 0.018119f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_95 VPB N_A2_M1034_g 0.01812f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_96 VPB N_A2_M1039_g 0.0183663f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_97 VPB N_A2_c_502_n 0.0100831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_582_n 0.011928f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.995
cc_99 VPB N_VPWR_c_583_n 0.00648869f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_100 VPB N_VPWR_c_584_n 0.0039289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_585_n 0.00454637f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_102 VPB N_VPWR_c_586_n 0.00506929f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.16
cc_103 VPB N_VPWR_c_587_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.175
cc_104 VPB N_VPWR_c_588_n 0.0151179f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_105 VPB N_VPWR_c_589_n 0.00873736f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.175
cc_106 VPB N_VPWR_c_590_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_591_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_592_n 0.0536884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_593_n 0.00477419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_594_n 0.0536819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_595_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_596_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_597_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_598_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_599_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_600_n 0.0216322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_581_n 0.050795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_719_n 0.00255113f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.16
cc_119 VPB N_Y_c_718_n 0.00432553f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_120 VPB N_Y_c_721_n 0.0180673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_Y_c_722_n 0.00234891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_Y_c_723_n 0.00420142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_1241_297#_c_886_n 0.00281045f $X=-0.19 $Y=1.305 $X2=1.75
+ $Y2=1.325
cc_124 N_C1_M1010_g N_VPWR_c_583_n 0.00338128f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_125 N_C1_c_129_n N_VPWR_c_583_n 0.015717f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C1_c_130_n N_VPWR_c_583_n 0.00174167f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_127 N_C1_M1029_g N_VPWR_c_584_n 0.00157837f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_128 N_C1_M1032_g N_VPWR_c_584_n 0.00157702f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_129 N_C1_M1010_g N_VPWR_c_596_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_130 N_C1_M1029_g N_VPWR_c_596_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_131 N_C1_M1032_g N_VPWR_c_599_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_132 N_C1_M1036_g N_VPWR_c_599_n 0.00585385f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C1_M1036_g N_VPWR_c_600_n 0.00353572f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C1_M1010_g N_VPWR_c_581_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C1_M1029_g N_VPWR_c_581_n 0.0104367f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_136 N_C1_M1032_g N_VPWR_c_581_n 0.0104367f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_137 N_C1_M1036_g N_VPWR_c_581_n 0.00720844f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_138 N_C1_c_125_n N_Y_c_717_n 0.00325185f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C1_c_126_n N_Y_c_717_n 0.00992642f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_140 N_C1_c_127_n N_Y_c_717_n 0.00992642f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_141 N_C1_c_128_n N_Y_c_717_n 0.012595f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C1_c_129_n N_Y_c_717_n 0.0627014f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_143 N_C1_c_130_n N_Y_c_717_n 0.00652975f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_144 N_C1_M1010_g N_Y_c_719_n 0.00130369f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_145 N_C1_c_129_n N_Y_c_719_n 0.0203891f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_146 N_C1_c_130_n N_Y_c_719_n 0.00222737f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_147 N_C1_c_128_n N_Y_c_718_n 0.0212082f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_148 N_C1_c_129_n N_Y_c_718_n 0.0160378f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_149 N_C1_M1029_g N_Y_c_722_n 0.0133089f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_150 N_C1_M1032_g N_Y_c_722_n 0.0133439f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_151 N_C1_c_129_n N_Y_c_722_n 0.0677173f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_152 N_C1_c_130_n N_Y_c_722_n 0.00214031f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_153 N_C1_M1036_g N_Y_c_723_n 0.0251909f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_154 N_C1_c_130_n N_Y_c_723_n 0.00220302f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_155 N_C1_c_125_n N_A_27_47#_c_936_n 3.87022e-19 $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C1_c_129_n N_A_27_47#_c_936_n 0.0200862f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_157 N_C1_c_130_n N_A_27_47#_c_936_n 9.92702e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_158 N_C1_c_125_n N_A_27_47#_c_937_n 0.0105669f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_159 N_C1_c_126_n N_A_27_47#_c_937_n 0.00892725f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_160 N_C1_c_127_n N_A_27_47#_c_937_n 0.00892725f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_161 N_C1_c_128_n N_A_27_47#_c_937_n 0.00892725f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_162 N_C1_c_129_n N_A_27_47#_c_937_n 0.00356026f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_163 N_C1_c_128_n N_A_471_47#_c_986_n 7.32022e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_164 N_C1_c_125_n N_VGND_c_1117_n 0.00357877f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_165 N_C1_c_126_n N_VGND_c_1117_n 0.00357877f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_166 N_C1_c_127_n N_VGND_c_1117_n 0.00357877f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_167 N_C1_c_128_n N_VGND_c_1117_n 0.00357877f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_168 N_C1_c_125_n N_VGND_c_1124_n 0.00619805f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_169 N_C1_c_126_n N_VGND_c_1124_n 0.00522516f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_170 N_C1_c_127_n N_VGND_c_1124_n 0.00522516f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_171 N_C1_c_128_n N_VGND_c_1124_n 0.00655123f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_186_n N_B2_c_295_n 0.0245982f $X=3.53 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_173 N_B1_M1023_g N_B2_M1008_g 0.0245982f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B1_c_196_n N_B2_M1008_g 7.43577e-19 $X=4.42 $Y=1.495 $X2=0 $Y2=0
cc_175 N_B1_c_196_n N_B2_M1012_g 0.00434944f $X=4.42 $Y=1.495 $X2=0 $Y2=0
cc_176 N_B1_c_204_p N_B2_M1012_g 0.00622646f $X=4.505 $Y=1.58 $X2=0 $Y2=0
cc_177 N_B1_c_196_n N_B2_M1033_g 0.0033124f $X=4.42 $Y=1.495 $X2=0 $Y2=0
cc_178 N_B1_c_206_p N_B2_M1033_g 0.0103677f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B1_c_187_n N_B2_c_298_n 0.0262556f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B1_M1025_g N_B2_M1037_g 0.0461811f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B1_c_206_p N_B2_M1037_g 0.0103235f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_182 N_B1_c_196_n N_B2_c_299_n 0.0036647f $X=4.42 $Y=1.495 $X2=0 $Y2=0
cc_183 N_B1_c_206_p N_B2_c_299_n 0.038721f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B1_c_188_n N_B2_c_299_n 0.0198443f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_185 N_B1_c_189_n N_B2_c_299_n 8.43231e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_186 N_B1_c_190_n N_B2_c_299_n 0.0167914f $X=4.335 $Y=1.175 $X2=0 $Y2=0
cc_187 N_B1_c_196_n N_B2_c_300_n 0.003462f $X=4.42 $Y=1.495 $X2=0 $Y2=0
cc_188 N_B1_c_206_p N_B2_c_300_n 0.0044825f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_189 N_B1_c_188_n N_B2_c_300_n 0.0047639f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B1_c_189_n N_B2_c_300_n 0.0212674f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B1_c_190_n N_B2_c_300_n 0.0348475f $X=4.335 $Y=1.175 $X2=0 $Y2=0
cc_192 N_B1_c_191_n N_B2_c_300_n 0.0245982f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B1_c_187_n N_A1_c_370_n 0.0187419f $X=5.63 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_194 N_B1_M1025_g N_A1_M1015_g 0.03475f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_c_206_p N_A1_M1015_g 0.00167791f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_196 N_B1_c_188_n N_A1_M1015_g 5.08505e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B1_M1025_g N_A1_c_374_n 3.56649e-19 $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B1_c_188_n N_A1_c_374_n 0.0307587f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_c_189_n N_A1_c_374_n 7.80994e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B1_c_188_n N_A1_c_375_n 7.80994e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B1_c_189_n N_A1_c_375_n 0.0197715f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_M1025_g N_A1_c_386_n 5.80938e-19 $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_c_206_p N_A1_c_386_n 0.0108192f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_204 N_B1_c_188_n N_A1_c_386_n 0.00434904f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B1_c_206_p N_VPWR_M1025_d 0.00215692f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B1_M1007_g N_VPWR_c_585_n 0.00157702f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1023_g N_VPWR_c_585_n 0.00302074f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_M1025_g N_VPWR_c_586_n 0.00291323f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1001_g N_VPWR_c_590_n 0.00585385f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1007_g N_VPWR_c_590_n 0.00585385f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1023_g N_VPWR_c_592_n 0.00585385f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1025_g N_VPWR_c_592_n 0.00420765f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1001_g N_VPWR_c_600_n 0.00353572f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1001_g N_VPWR_c_581_n 0.0117604f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1007_g N_VPWR_c_581_n 0.00588483f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_M1023_g N_VPWR_c_581_n 0.00591203f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B1_M1025_g N_VPWR_c_581_n 0.00594423f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_c_206_p N_Y_M1033_s 0.00311483f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B1_c_184_n N_Y_c_718_n 0.00298558f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B1_M1001_g N_Y_c_718_n 0.00298989f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B1_c_190_n N_Y_c_718_n 0.0134954f $X=4.335 $Y=1.175 $X2=0 $Y2=0
cc_222 N_B1_c_191_n N_Y_c_718_n 0.00502925f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B1_M1001_g N_Y_c_721_n 0.0170519f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B1_M1007_g N_Y_c_721_n 0.0103677f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B1_M1023_g N_Y_c_721_n 0.0103235f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B1_c_196_n N_Y_c_721_n 0.00398241f $X=4.42 $Y=1.495 $X2=0 $Y2=0
cc_227 N_B1_c_204_p N_Y_c_721_n 0.0104885f $X=4.505 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_c_190_n N_Y_c_721_n 0.131145f $X=4.335 $Y=1.175 $X2=0 $Y2=0
cc_229 N_B1_c_191_n N_Y_c_721_n 0.00535077f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B1_M1023_g N_Y_c_753_n 8.02934e-19 $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_231 N_B1_c_204_p N_Y_c_753_n 0.00389346f $X=4.505 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B1_c_206_p N_Y_c_755_n 0.0212097f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B1_c_204_p N_Y_c_755_n 0.0082755f $X=4.505 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B1_M1025_g N_Y_c_757_n 0.0120778f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_235 N_B1_c_206_p N_Y_c_757_n 0.035542f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B1_c_189_n N_Y_c_757_n 2.75745e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B1_M1025_g N_Y_c_760_n 0.00127015f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_238 N_B1_M1001_g N_Y_c_723_n 0.00796816f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B1_c_190_n N_Y_c_762_n 0.0039114f $X=4.335 $Y=1.175 $X2=0 $Y2=0
cc_240 N_B1_c_206_p N_Y_c_763_n 0.0118606f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B1_c_206_p N_A_553_297#_M1012_d 0.00426642f $X=5.465 $Y=1.58 $X2=0
+ $Y2=0
cc_242 N_B1_c_206_p N_A_553_297#_M1037_d 0.00423833f $X=5.465 $Y=1.58 $X2=0
+ $Y2=0
cc_243 N_B1_M1007_g N_A_553_297#_c_849_n 0.00956194f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_B1_M1023_g N_A_553_297#_c_849_n 0.00956194f $X=3.53 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_B1_M1025_g N_A_553_297#_c_851_n 0.00371016f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_B1_c_184_n N_A_27_47#_c_937_n 0.0116561f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B1_c_185_n N_A_27_47#_c_937_n 0.00892725f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_c_186_n N_A_27_47#_c_937_n 0.00892725f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B1_c_187_n N_A_27_47#_c_937_n 0.00296299f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_c_184_n N_A_471_47#_c_986_n 0.00898612f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B1_c_185_n N_A_471_47#_c_986_n 0.00898612f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_c_186_n N_A_471_47#_c_986_n 0.00894065f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B1_c_206_p N_A_471_47#_c_986_n 0.00704573f $X=5.465 $Y=1.58 $X2=0 $Y2=0
cc_254 N_B1_c_190_n N_A_471_47#_c_986_n 0.0972504f $X=4.335 $Y=1.175 $X2=0 $Y2=0
cc_255 N_B1_c_191_n N_A_471_47#_c_986_n 0.00419061f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_187_n N_A_471_47#_c_987_n 0.0149528f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B1_c_188_n N_A_471_47#_c_987_n 0.0264065f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_189_n N_A_471_47#_c_987_n 0.00298767f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B1_c_184_n N_VGND_c_1117_n 0.00357877f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B1_c_185_n N_VGND_c_1117_n 0.00357877f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B1_c_186_n N_VGND_c_1117_n 0.00357877f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B1_c_187_n N_VGND_c_1117_n 0.00412827f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_263 N_B1_c_184_n N_VGND_c_1124_n 0.00660224f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_264 N_B1_c_185_n N_VGND_c_1124_n 0.00522516f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B1_c_186_n N_VGND_c_1124_n 0.00525237f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_266 N_B1_c_187_n N_VGND_c_1124_n 0.00598156f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B2_M1008_g N_VPWR_c_592_n 0.00357877f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B2_M1012_g N_VPWR_c_592_n 0.00357877f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B2_M1033_g N_VPWR_c_592_n 0.00357877f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B2_M1037_g N_VPWR_c_592_n 0.00357877f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B2_M1008_g N_VPWR_c_581_n 0.00525237f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B2_M1012_g N_VPWR_c_581_n 0.00522516f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B2_M1033_g N_VPWR_c_581_n 0.00522516f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B2_M1037_g N_VPWR_c_581_n 0.00525237f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B2_M1008_g N_Y_c_721_n 0.0127446f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B2_M1012_g N_Y_c_721_n 0.0011553f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B2_c_300_n N_Y_c_721_n 0.00121587f $X=5.21 $Y=1.16 $X2=0 $Y2=0
cc_278 N_B2_M1008_g N_Y_c_753_n 0.00457096f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B2_M1012_g N_Y_c_753_n 0.00371906f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B2_M1012_g N_Y_c_755_n 0.00945997f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B2_M1033_g N_Y_c_755_n 0.0093114f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B2_M1037_g N_Y_c_757_n 0.0092042f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_283 N_B2_M1008_g N_Y_c_762_n 0.00349486f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B2_c_300_n N_Y_c_762_n 7.26014e-19 $X=5.21 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B2_M1008_g N_A_553_297#_c_852_n 0.0112448f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_286 N_B2_M1012_g N_A_553_297#_c_852_n 0.00824376f $X=4.37 $Y=1.985 $X2=0
+ $Y2=0
cc_287 N_B2_M1033_g N_A_553_297#_c_851_n 3.55797e-19 $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_B2_M1037_g N_A_553_297#_c_851_n 0.00327079f $X=5.21 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_B2_M1033_g N_A_553_297#_c_856_n 0.0075938f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_290 N_B2_M1037_g N_A_553_297#_c_856_n 0.00613019f $X=5.21 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_B2_c_295_n N_A_27_47#_c_937_n 0.00892725f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_296_n N_A_27_47#_c_937_n 0.00892725f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B2_c_297_n N_A_27_47#_c_937_n 0.00892725f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B2_c_298_n N_A_27_47#_c_937_n 0.00892725f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B2_c_295_n N_A_471_47#_c_986_n 0.00894065f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B2_c_296_n N_A_471_47#_c_986_n 0.00898205f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B2_c_297_n N_A_471_47#_c_986_n 0.00852218f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B2_c_298_n N_A_471_47#_c_986_n 0.00847671f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B2_c_299_n N_A_471_47#_c_986_n 0.0378422f $X=5.15 $Y=1.16 $X2=0 $Y2=0
cc_300 N_B2_c_300_n N_A_471_47#_c_986_n 0.00656134f $X=5.21 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B2_c_298_n N_A_471_47#_c_987_n 0.00227718f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B2_c_295_n N_VGND_c_1117_n 0.00357877f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B2_c_296_n N_VGND_c_1117_n 0.00357877f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B2_c_297_n N_VGND_c_1117_n 0.00357877f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B2_c_298_n N_VGND_c_1117_n 0.00357877f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B2_c_295_n N_VGND_c_1124_n 0.00525237f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B2_c_296_n N_VGND_c_1124_n 0.00522516f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_308 N_B2_c_297_n N_VGND_c_1124_n 0.00522516f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B2_c_298_n N_VGND_c_1124_n 0.00525237f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A1_c_370_n N_A2_c_498_n 0.0258234f $X=6.13 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_311 N_A1_M1015_g N_A2_M1002_g 0.0463944f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A1_c_385_n N_A2_M1002_g 0.0102975f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_313 N_A1_c_385_n N_A2_M1031_g 0.0103615f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_314 N_A1_c_385_n N_A2_M1034_g 0.0103615f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_315 N_A1_c_371_n N_A2_c_501_n 0.0240283f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A1_M1024_g N_A2_M1039_g 0.0240283f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A1_c_385_n N_A2_M1039_g 0.0148849f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_318 N_A1_c_374_n N_A2_c_516_n 0.0160038f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A1_c_375_n N_A2_c_516_n 2.34877e-19 $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A1_c_385_n N_A2_c_516_n 0.100214f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_321 N_A1_c_376_n N_A2_c_516_n 0.0116221f $X=8.287 $Y=1.275 $X2=0 $Y2=0
cc_322 N_A1_c_378_n N_A2_c_516_n 2.52028e-19 $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A1_c_374_n N_A2_c_502_n 0.00518416f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A1_c_375_n N_A2_c_502_n 0.0228076f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A1_c_385_n N_A2_c_502_n 0.00641737f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_326 N_A1_c_376_n N_A2_c_502_n 8.91817e-19 $X=8.287 $Y=1.275 $X2=0 $Y2=0
cc_327 N_A1_c_387_n N_A2_c_502_n 0.00112116f $X=8.287 $Y=1.445 $X2=0 $Y2=0
cc_328 N_A1_c_378_n N_A2_c_502_n 0.0240283f $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A1_c_386_n N_VPWR_M1025_d 0.00151145f $X=6.295 $Y=1.53 $X2=0 $Y2=0
cc_330 N_A1_c_385_n N_VPWR_M1024_s 0.00209238f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_331 N_A1_M1015_g N_VPWR_c_586_n 0.00291323f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A1_M1024_g N_VPWR_c_587_n 0.00302074f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A1_M1030_g N_VPWR_c_587_n 0.00157837f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A1_M1035_g N_VPWR_c_589_n 0.00431697f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A1_c_377_n N_VPWR_c_589_n 0.0210492f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A1_c_378_n N_VPWR_c_589_n 8.41451e-19 $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A1_M1015_g N_VPWR_c_594_n 0.00420655f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A1_M1024_g N_VPWR_c_594_n 0.00585385f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A1_M1030_g N_VPWR_c_597_n 0.00585385f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A1_M1035_g N_VPWR_c_597_n 0.00585385f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A1_M1015_g N_VPWR_c_581_n 0.00594226f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A1_M1024_g N_VPWR_c_581_n 0.00591203f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A1_M1030_g N_VPWR_c_581_n 0.00588483f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A1_M1035_g N_VPWR_c_581_n 0.0114878f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A1_c_385_n N_Y_M1002_d 0.00165831f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_346 N_A1_c_385_n N_Y_M1034_d 0.00165831f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_347 N_A1_c_385_n N_Y_c_776_n 0.0315971f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_348 N_A1_M1015_g N_Y_c_760_n 0.0138131f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A1_c_375_n N_Y_c_760_n 3.02339e-19 $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A1_c_385_n N_Y_c_760_n 0.0315216f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_351 N_A1_c_386_n N_Y_c_760_n 0.0168722f $X=6.295 $Y=1.53 $X2=0 $Y2=0
cc_352 N_A1_c_385_n N_Y_c_781_n 0.0120079f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_353 N_A1_c_385_n N_A_1241_297#_M1015_d 0.00129688f $X=8.155 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_354 N_A1_c_386_n N_A_1241_297#_M1015_d 3.51639e-19 $X=6.295 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_355 N_A1_c_385_n N_A_1241_297#_M1031_s 0.00166235f $X=8.155 $Y=1.53 $X2=0
+ $Y2=0
cc_356 N_A1_c_385_n N_A_1241_297#_M1039_s 0.00165831f $X=8.155 $Y=1.53 $X2=0
+ $Y2=0
cc_357 N_A1_M1024_g N_A_1241_297#_c_891_n 0.0095558f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A1_M1030_g N_A_1241_297#_c_891_n 0.0112521f $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A1_c_385_n N_A_1241_297#_c_891_n 0.0157651f $X=8.155 $Y=1.53 $X2=0
+ $Y2=0
cc_360 N_A1_c_377_n N_A_1241_297#_c_891_n 0.00808474f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_361 N_A1_c_378_n N_A_1241_297#_c_891_n 0.00129797f $X=9.07 $Y=1.16 $X2=0
+ $Y2=0
cc_362 N_A1_c_385_n N_A_1241_297#_c_896_n 0.0126919f $X=8.155 $Y=1.53 $X2=0
+ $Y2=0
cc_363 N_A1_M1030_g N_A_1241_297#_c_886_n 4.03862e-19 $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_364 N_A1_M1035_g N_A_1241_297#_c_886_n 3.09636e-19 $X=9.07 $Y=1.985 $X2=0
+ $Y2=0
cc_365 N_A1_c_385_n N_A_1241_297#_c_886_n 0.00592489f $X=8.155 $Y=1.53 $X2=0
+ $Y2=0
cc_366 N_A1_c_377_n N_A_1241_297#_c_886_n 0.020226f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_367 N_A1_c_378_n N_A_1241_297#_c_886_n 0.00222737f $X=9.07 $Y=1.16 $X2=0
+ $Y2=0
cc_368 N_A1_M1015_g N_A_1241_297#_c_902_n 0.00370893f $X=6.13 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_A1_c_370_n N_A_471_47#_c_1008_n 0.00502318f $X=6.13 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A1_c_370_n N_A_471_47#_c_981_n 0.00845282f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A1_c_375_n N_A_471_47#_c_981_n 0.001478f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_372 N_A1_c_385_n N_A_471_47#_c_981_n 0.00609408f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_373 N_A1_c_370_n N_A_471_47#_c_1012_n 5.24135e-19 $X=6.13 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A1_c_371_n N_A_471_47#_c_1013_n 5.22228e-19 $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A1_c_371_n N_A_471_47#_c_983_n 0.00845282f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A1_c_385_n N_A_471_47#_c_983_n 0.00913644f $X=8.155 $Y=1.53 $X2=0 $Y2=0
cc_377 N_A1_c_376_n N_A_471_47#_c_983_n 0.00893273f $X=8.287 $Y=1.275 $X2=0
+ $Y2=0
cc_378 N_A1_c_371_n N_A_471_47#_c_1017_n 0.00630972f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A1_c_372_n N_A_471_47#_c_1017_n 0.00630972f $X=8.65 $Y=0.995 $X2=0
+ $Y2=0
cc_380 N_A1_c_373_n N_A_471_47#_c_1017_n 5.22228e-19 $X=9.07 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A1_c_372_n N_A_471_47#_c_984_n 0.00870364f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A1_c_373_n N_A_471_47#_c_984_n 0.00999903f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_383 N_A1_c_377_n N_A_471_47#_c_984_n 0.0637671f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_384 N_A1_c_378_n N_A_471_47#_c_984_n 0.00337303f $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A1_c_372_n N_A_471_47#_c_985_n 5.22228e-19 $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A1_c_373_n N_A_471_47#_c_985_n 0.00630972f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A1_c_370_n N_A_471_47#_c_987_n 0.00284957f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A1_c_374_n N_A_471_47#_c_987_n 0.0256887f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A1_c_375_n N_A_471_47#_c_987_n 0.00149384f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A1_c_371_n N_A_471_47#_c_990_n 0.00127865f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_391 N_A1_c_372_n N_A_471_47#_c_990_n 0.00113286f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_392 N_A1_c_376_n N_A_471_47#_c_990_n 0.0125375f $X=8.287 $Y=1.275 $X2=0 $Y2=0
cc_393 N_A1_c_377_n N_A_471_47#_c_990_n 0.0148598f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_394 N_A1_c_378_n N_A_471_47#_c_990_n 0.00230291f $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_395 N_A1_c_370_n N_VGND_c_1112_n 0.00268723f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_396 N_A1_c_371_n N_VGND_c_1115_n 0.00146448f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A1_c_372_n N_VGND_c_1116_n 0.00146448f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A1_c_373_n N_VGND_c_1116_n 0.00268723f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A1_c_370_n N_VGND_c_1117_n 0.00423357f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A1_c_371_n N_VGND_c_1121_n 0.00424416f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A1_c_372_n N_VGND_c_1121_n 0.00423334f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A1_c_373_n N_VGND_c_1123_n 0.00423334f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A1_c_370_n N_VGND_c_1124_n 0.00597464f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A1_c_371_n N_VGND_c_1124_n 0.00576327f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A1_c_372_n N_VGND_c_1124_n 0.0057163f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A1_c_373_n N_VGND_c_1124_n 0.00676734f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A2_M1002_g N_VPWR_c_594_n 0.00357877f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A2_M1031_g N_VPWR_c_594_n 0.00357877f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_409 N_A2_M1034_g N_VPWR_c_594_n 0.00357877f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_410 N_A2_M1039_g N_VPWR_c_594_n 0.00357877f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_411 N_A2_M1002_g N_VPWR_c_581_n 0.00525237f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_412 N_A2_M1031_g N_VPWR_c_581_n 0.00522516f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_413 N_A2_M1034_g N_VPWR_c_581_n 0.00522516f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_414 N_A2_M1039_g N_VPWR_c_581_n 0.00525237f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_415 N_A2_M1031_g N_Y_c_776_n 0.00924026f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_416 N_A2_M1034_g N_Y_c_776_n 0.00928441f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_417 N_A2_M1002_g N_Y_c_760_n 0.0101984f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_418 N_A2_M1002_g N_A_1241_297#_c_903_n 0.00697687f $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_419 N_A2_M1031_g N_A_1241_297#_c_903_n 0.00856088f $X=6.97 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A2_M1034_g N_A_1241_297#_c_905_n 0.00851673f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_421 N_A2_M1039_g N_A_1241_297#_c_905_n 0.0121306f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_422 N_A2_M1002_g N_A_1241_297#_c_902_n 0.00327147f $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A2_M1031_g N_A_1241_297#_c_902_n 3.55948e-19 $X=6.97 $Y=1.985 $X2=0
+ $Y2=0
cc_424 N_A2_c_498_n N_A_471_47#_c_1008_n 2.88203e-19 $X=6.55 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_A2_c_498_n N_A_471_47#_c_981_n 0.00843917f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A2_c_516_n N_A_471_47#_c_981_n 0.00817906f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A2_c_498_n N_A_471_47#_c_1012_n 0.00629364f $X=6.55 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A2_c_499_n N_A_471_47#_c_1012_n 0.00630972f $X=6.97 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_A2_c_500_n N_A_471_47#_c_1012_n 5.22228e-19 $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A2_c_499_n N_A_471_47#_c_982_n 0.00869873f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A2_c_500_n N_A_471_47#_c_982_n 0.00869873f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_432 N_A2_c_516_n N_A_471_47#_c_982_n 0.0363039f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_433 N_A2_c_502_n N_A_471_47#_c_982_n 0.00222006f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A2_c_499_n N_A_471_47#_c_1013_n 5.22228e-19 $X=6.97 $Y=0.995 $X2=0
+ $Y2=0
cc_435 N_A2_c_500_n N_A_471_47#_c_1013_n 0.00630972f $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_436 N_A2_c_501_n N_A_471_47#_c_1013_n 0.00630972f $X=7.81 $Y=0.995 $X2=0
+ $Y2=0
cc_437 N_A2_c_501_n N_A_471_47#_c_983_n 0.00843917f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A2_c_516_n N_A_471_47#_c_983_n 0.00817906f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_439 N_A2_c_501_n N_A_471_47#_c_1017_n 5.22228e-19 $X=7.81 $Y=0.995 $X2=0
+ $Y2=0
cc_440 N_A2_c_498_n N_A_471_47#_c_987_n 2.60259e-19 $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_441 N_A2_c_498_n N_A_471_47#_c_988_n 0.00127865f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_442 N_A2_c_499_n N_A_471_47#_c_988_n 0.00113159f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_443 N_A2_c_516_n N_A_471_47#_c_988_n 0.0266779f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_444 N_A2_c_502_n N_A_471_47#_c_988_n 0.00230167f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_445 N_A2_c_500_n N_A_471_47#_c_989_n 0.00113159f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_446 N_A2_c_501_n N_A_471_47#_c_989_n 0.00127865f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_447 N_A2_c_516_n N_A_471_47#_c_989_n 0.0266779f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_448 N_A2_c_502_n N_A_471_47#_c_989_n 0.00230167f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_449 N_A2_c_498_n N_VGND_c_1112_n 0.00146448f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_450 N_A2_c_498_n N_VGND_c_1113_n 0.00424416f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_451 N_A2_c_499_n N_VGND_c_1113_n 0.00423334f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_452 N_A2_c_499_n N_VGND_c_1114_n 0.00146448f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_453 N_A2_c_500_n N_VGND_c_1114_n 0.00146448f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_454 N_A2_c_501_n N_VGND_c_1115_n 0.00146448f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_455 N_A2_c_500_n N_VGND_c_1119_n 0.00423334f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_456 N_A2_c_501_n N_VGND_c_1119_n 0.00424416f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_457 N_A2_c_498_n N_VGND_c_1124_n 0.00576327f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_458 N_A2_c_499_n N_VGND_c_1124_n 0.0057163f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_459 N_A2_c_500_n N_VGND_c_1124_n 0.0057163f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_460 N_A2_c_501_n N_VGND_c_1124_n 0.00576327f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_461 N_VPWR_c_581_n N_Y_M1010_d 0.00284632f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_462 N_VPWR_c_581_n N_Y_M1032_d 0.00251211f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_463 N_VPWR_c_581_n N_Y_M1008_s 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_464 N_VPWR_c_581_n N_Y_M1033_s 0.00215227f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_c_581_n N_Y_M1002_d 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_466 N_VPWR_c_581_n N_Y_M1034_d 0.0021603f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_467 N_VPWR_c_596_n N_Y_c_791_n 0.0142343f $X=0.995 $Y=2.72 $X2=0 $Y2=0
cc_468 N_VPWR_c_581_n N_Y_c_791_n 0.00955092f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_469 N_VPWR_c_599_n N_Y_c_793_n 0.0140073f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_470 N_VPWR_c_581_n N_Y_c_793_n 0.00948039f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_471 N_VPWR_M1036_s N_Y_c_721_n 0.0100922f $X=1.825 $Y=1.485 $X2=0 $Y2=0
cc_472 N_VPWR_M1007_d N_Y_c_721_n 0.00166235f $X=3.185 $Y=1.485 $X2=0 $Y2=0
cc_473 N_VPWR_c_600_n N_Y_c_721_n 0.0155161f $X=2.605 $Y=2.465 $X2=0 $Y2=0
cc_474 N_VPWR_M1025_d N_Y_c_757_n 0.00884898f $X=5.705 $Y=1.485 $X2=0 $Y2=0
cc_475 N_VPWR_c_586_n N_Y_c_757_n 0.0158147f $X=5.88 $Y=2.35 $X2=0 $Y2=0
cc_476 N_VPWR_c_592_n N_Y_c_757_n 0.00231767f $X=5.755 $Y=2.72 $X2=0 $Y2=0
cc_477 N_VPWR_c_581_n N_Y_c_757_n 0.00574489f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_478 N_VPWR_c_581_n N_Y_c_776_n 0.00127501f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_479 N_VPWR_M1025_d N_Y_c_760_n 0.00139829f $X=5.705 $Y=1.485 $X2=0 $Y2=0
cc_480 N_VPWR_c_586_n N_Y_c_760_n 0.00263443f $X=5.88 $Y=2.35 $X2=0 $Y2=0
cc_481 N_VPWR_c_594_n N_Y_c_760_n 0.0020648f $X=8.315 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_581_n N_Y_c_760_n 0.00508661f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_M1029_s N_Y_c_722_n 0.00181725f $X=0.985 $Y=1.485 $X2=0 $Y2=0
cc_484 N_VPWR_c_584_n N_Y_c_722_n 0.0108451f $X=1.12 $Y=1.99 $X2=0 $Y2=0
cc_485 N_VPWR_M1036_s N_Y_c_723_n 0.0118455f $X=1.825 $Y=1.485 $X2=0 $Y2=0
cc_486 N_VPWR_c_600_n N_Y_c_723_n 0.0205807f $X=2.605 $Y=2.465 $X2=0 $Y2=0
cc_487 N_VPWR_c_581_n N_Y_c_723_n 0.00685613f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_488 N_VPWR_c_581_n N_A_553_297#_M1001_s 0.00254126f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_489 N_VPWR_c_581_n N_A_553_297#_M1023_s 0.00220218f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_581_n N_A_553_297#_M1012_d 0.00215227f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_581_n N_A_553_297#_M1037_d 0.00215227f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_590_n N_A_553_297#_c_862_n 0.0142343f $X=3.195 $Y=2.72 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_581_n N_A_553_297#_c_862_n 0.00955092f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_494 N_VPWR_M1007_d N_A_553_297#_c_849_n 0.00317012f $X=3.185 $Y=1.485 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_585_n N_A_553_297#_c_849_n 0.0123301f $X=3.32 $Y=2.3 $X2=0 $Y2=0
cc_496 N_VPWR_c_581_n N_A_553_297#_c_849_n 0.0109281f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_592_n N_A_553_297#_c_867_n 0.012886f $X=5.755 $Y=2.72 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_581_n N_A_553_297#_c_867_n 0.00808747f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_592_n N_A_553_297#_c_852_n 0.0973478f $X=5.755 $Y=2.72 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_581_n N_A_553_297#_c_852_n 0.0626839f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_581_n N_A_1241_297#_M1015_d 0.00215227f $X=9.43 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_502 N_VPWR_c_581_n N_A_1241_297#_M1031_s 0.00213597f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_581_n N_A_1241_297#_M1039_s 0.00220214f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_581_n N_A_1241_297#_M1030_d 0.00254126f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_594_n N_A_1241_297#_c_905_n 0.0473226f $X=8.315 $Y=2.72 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_581_n N_A_1241_297#_c_905_n 0.0300947f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_507 N_VPWR_M1024_s N_A_1241_297#_c_891_n 0.00378557f $X=8.305 $Y=1.485 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_587_n N_A_1241_297#_c_891_n 0.0123301f $X=8.44 $Y=2.3 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_581_n N_A_1241_297#_c_891_n 0.0109281f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_589_n N_A_1241_297#_c_886_n 0.00311153f $X=9.28 $Y=1.62 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_597_n N_A_1241_297#_c_919_n 0.0142343f $X=9.155 $Y=2.72 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_581_n N_A_1241_297#_c_919_n 0.00955092f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_594_n N_A_1241_297#_c_902_n 0.048863f $X=8.315 $Y=2.72 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_581_n N_A_1241_297#_c_902_n 0.0312052f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_594_n N_A_1241_297#_c_923_n 0.0137033f $X=8.315 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_581_n N_A_1241_297#_c_923_n 0.00938745f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_Y_c_721_n N_A_553_297#_M1001_s 0.00165831f $X=3.995 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_518 N_Y_c_721_n N_A_553_297#_M1023_s 0.00165831f $X=3.995 $Y=1.53 $X2=0 $Y2=0
cc_519 N_Y_c_755_n N_A_553_297#_M1012_d 0.00312531f $X=4.875 $Y=1.92 $X2=0 $Y2=0
cc_520 N_Y_c_757_n N_A_553_297#_M1037_d 0.00323871f $X=5.965 $Y=1.92 $X2=0 $Y2=0
cc_521 N_Y_c_721_n N_A_553_297#_c_849_n 0.0442891f $X=3.995 $Y=1.53 $X2=0 $Y2=0
cc_522 N_Y_c_721_n N_A_553_297#_c_876_n 0.0126919f $X=3.995 $Y=1.53 $X2=0 $Y2=0
cc_523 N_Y_M1008_s N_A_553_297#_c_852_n 0.00311686f $X=4.025 $Y=1.485 $X2=0
+ $Y2=0
cc_524 N_Y_c_755_n N_A_553_297#_c_852_n 0.00585978f $X=4.875 $Y=1.92 $X2=0 $Y2=0
cc_525 N_Y_c_762_n N_A_553_297#_c_852_n 0.0130493f $X=4.285 $Y=1.98 $X2=0 $Y2=0
cc_526 N_Y_c_755_n N_A_553_297#_c_880_n 0.011218f $X=4.875 $Y=1.92 $X2=0 $Y2=0
cc_527 N_Y_c_757_n N_A_553_297#_c_851_n 0.0153733f $X=5.965 $Y=1.92 $X2=0 $Y2=0
cc_528 N_Y_M1033_s N_A_553_297#_c_856_n 0.00312348f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_529 N_Y_c_755_n N_A_553_297#_c_856_n 0.0043088f $X=4.875 $Y=1.92 $X2=0 $Y2=0
cc_530 N_Y_c_757_n N_A_553_297#_c_856_n 0.0027357f $X=5.965 $Y=1.92 $X2=0 $Y2=0
cc_531 N_Y_c_763_n N_A_553_297#_c_856_n 0.0111508f $X=5 $Y=1.96 $X2=0 $Y2=0
cc_532 N_Y_c_760_n N_A_1241_297#_M1015_d 0.00326812f $X=6.885 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_533 N_Y_c_776_n N_A_1241_297#_M1031_s 0.00317012f $X=7.475 $Y=1.87 $X2=0
+ $Y2=0
cc_534 N_Y_M1002_d N_A_1241_297#_c_903_n 0.00312348f $X=6.625 $Y=1.485 $X2=0
+ $Y2=0
cc_535 N_Y_c_776_n N_A_1241_297#_c_903_n 0.00506389f $X=7.475 $Y=1.87 $X2=0
+ $Y2=0
cc_536 N_Y_c_760_n N_A_1241_297#_c_903_n 0.016062f $X=6.885 $Y=1.87 $X2=0 $Y2=0
cc_537 N_Y_M1034_d N_A_1241_297#_c_905_n 0.00312348f $X=7.465 $Y=1.485 $X2=0
+ $Y2=0
cc_538 N_Y_c_776_n N_A_1241_297#_c_905_n 0.00506389f $X=7.475 $Y=1.87 $X2=0
+ $Y2=0
cc_539 N_Y_c_781_n N_A_1241_297#_c_905_n 0.0112811f $X=7.6 $Y=1.87 $X2=0 $Y2=0
cc_540 N_Y_c_760_n N_A_1241_297#_c_902_n 0.0157426f $X=6.885 $Y=1.87 $X2=0 $Y2=0
cc_541 N_Y_c_776_n N_A_1241_297#_c_923_n 0.0116461f $X=7.475 $Y=1.87 $X2=0 $Y2=0
cc_542 N_Y_c_717_n N_A_27_47#_M1018_s 0.00320532f $X=1.92 $Y=0.755 $X2=0 $Y2=0
cc_543 N_Y_c_717_n N_A_27_47#_M1027_s 0.00379863f $X=1.92 $Y=0.755 $X2=0 $Y2=0
cc_544 N_Y_c_718_n N_A_27_47#_M1027_s 3.00511e-19 $X=2.022 $Y=1.445 $X2=0 $Y2=0
cc_545 N_Y_M1013_d N_A_27_47#_c_937_n 0.00305026f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_546 N_Y_M1026_d N_A_27_47#_c_937_n 0.00305026f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_547 N_Y_c_717_n N_A_27_47#_c_937_n 0.0844245f $X=1.92 $Y=0.755 $X2=0 $Y2=0
cc_548 N_Y_c_717_n N_A_471_47#_c_986_n 0.0149754f $X=1.92 $Y=0.755 $X2=0 $Y2=0
cc_549 N_Y_c_721_n N_A_471_47#_c_986_n 0.00136402f $X=3.995 $Y=1.53 $X2=0 $Y2=0
cc_550 N_Y_M1013_d N_VGND_c_1124_n 0.00216833f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_551 N_Y_M1026_d N_VGND_c_1124_n 0.00216833f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_552 N_A_27_47#_c_937_n N_A_471_47#_M1003_s 0.00506759f $X=5.42 $Y=0.39
+ $X2=-0.19 $Y2=-0.24
cc_553 N_A_27_47#_c_937_n N_A_471_47#_M1011_s 0.00305026f $X=5.42 $Y=0.39 $X2=0
+ $Y2=0
cc_554 N_A_27_47#_c_937_n N_A_471_47#_M1004_d 0.00305026f $X=5.42 $Y=0.39 $X2=0
+ $Y2=0
cc_555 N_A_27_47#_c_937_n N_A_471_47#_M1016_d 0.00305026f $X=5.42 $Y=0.39 $X2=0
+ $Y2=0
cc_556 N_A_27_47#_M1003_d N_A_471_47#_c_986_n 0.00333526f $X=2.765 $Y=0.235
+ $X2=0 $Y2=0
cc_557 N_A_27_47#_M1019_d N_A_471_47#_c_986_n 0.0035985f $X=3.605 $Y=0.235 $X2=0
+ $Y2=0
cc_558 N_A_27_47#_M1014_s N_A_471_47#_c_986_n 0.00427696f $X=4.445 $Y=0.235
+ $X2=0 $Y2=0
cc_559 N_A_27_47#_M1020_s N_A_471_47#_c_986_n 0.00384155f $X=5.285 $Y=0.235
+ $X2=0 $Y2=0
cc_560 N_A_27_47#_c_937_n N_A_471_47#_c_986_n 0.165202f $X=5.42 $Y=0.39 $X2=0
+ $Y2=0
cc_561 N_A_27_47#_M1020_s N_A_471_47#_c_987_n 0.0012401f $X=5.285 $Y=0.235 $X2=0
+ $Y2=0
cc_562 N_A_27_47#_c_935_n N_VGND_c_1117_n 0.017288f $X=0.24 $Y=0.475 $X2=0 $Y2=0
cc_563 N_A_27_47#_c_937_n N_VGND_c_1117_n 0.295311f $X=5.42 $Y=0.39 $X2=0 $Y2=0
cc_564 N_A_27_47#_M1013_s N_VGND_c_1124_n 0.0022572f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_565 N_A_27_47#_M1018_s N_VGND_c_1124_n 0.00215227f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_566 N_A_27_47#_M1027_s N_VGND_c_1124_n 0.00209344f $X=1.825 $Y=0.235 $X2=0
+ $Y2=0
cc_567 N_A_27_47#_M1003_d N_VGND_c_1124_n 0.00215227f $X=2.765 $Y=0.235 $X2=0
+ $Y2=0
cc_568 N_A_27_47#_M1019_d N_VGND_c_1124_n 0.00215227f $X=3.605 $Y=0.235 $X2=0
+ $Y2=0
cc_569 N_A_27_47#_M1014_s N_VGND_c_1124_n 0.00215227f $X=4.445 $Y=0.235 $X2=0
+ $Y2=0
cc_570 N_A_27_47#_M1020_s N_VGND_c_1124_n 0.00215227f $X=5.285 $Y=0.235 $X2=0
+ $Y2=0
cc_571 N_A_27_47#_c_935_n N_VGND_c_1124_n 0.00961275f $X=0.24 $Y=0.475 $X2=0
+ $Y2=0
cc_572 N_A_27_47#_c_937_n N_VGND_c_1124_n 0.187004f $X=5.42 $Y=0.39 $X2=0 $Y2=0
cc_573 N_A_471_47#_c_981_n N_VGND_M1005_d 0.00165819f $X=6.595 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_574 N_A_471_47#_c_982_n N_VGND_M1006_s 0.00162089f $X=7.435 $Y=0.815 $X2=0
+ $Y2=0
cc_575 N_A_471_47#_c_983_n N_VGND_M1021_s 0.00165819f $X=8.275 $Y=0.82 $X2=0
+ $Y2=0
cc_576 N_A_471_47#_c_984_n N_VGND_M1022_d 0.00162089f $X=9.115 $Y=0.815 $X2=0
+ $Y2=0
cc_577 N_A_471_47#_c_981_n N_VGND_c_1112_n 0.0116528f $X=6.595 $Y=0.82 $X2=0
+ $Y2=0
cc_578 N_A_471_47#_c_981_n N_VGND_c_1113_n 0.00193763f $X=6.595 $Y=0.82 $X2=0
+ $Y2=0
cc_579 N_A_471_47#_c_1012_n N_VGND_c_1113_n 0.0188551f $X=6.76 $Y=0.39 $X2=0
+ $Y2=0
cc_580 N_A_471_47#_c_982_n N_VGND_c_1113_n 0.00198695f $X=7.435 $Y=0.815 $X2=0
+ $Y2=0
cc_581 N_A_471_47#_c_982_n N_VGND_c_1114_n 0.0122559f $X=7.435 $Y=0.815 $X2=0
+ $Y2=0
cc_582 N_A_471_47#_c_983_n N_VGND_c_1115_n 0.0116529f $X=8.275 $Y=0.82 $X2=0
+ $Y2=0
cc_583 N_A_471_47#_c_984_n N_VGND_c_1116_n 0.0122559f $X=9.115 $Y=0.815 $X2=0
+ $Y2=0
cc_584 N_A_471_47#_c_1008_n N_VGND_c_1117_n 0.0200505f $X=5.92 $Y=0.39 $X2=0
+ $Y2=0
cc_585 N_A_471_47#_c_981_n N_VGND_c_1117_n 0.00193763f $X=6.595 $Y=0.82 $X2=0
+ $Y2=0
cc_586 N_A_471_47#_c_987_n N_VGND_c_1117_n 0.00247354f $X=6.085 $Y=0.775 $X2=0
+ $Y2=0
cc_587 N_A_471_47#_c_982_n N_VGND_c_1119_n 0.00198695f $X=7.435 $Y=0.815 $X2=0
+ $Y2=0
cc_588 N_A_471_47#_c_1013_n N_VGND_c_1119_n 0.0188551f $X=7.6 $Y=0.39 $X2=0
+ $Y2=0
cc_589 N_A_471_47#_c_983_n N_VGND_c_1119_n 0.00193763f $X=8.275 $Y=0.82 $X2=0
+ $Y2=0
cc_590 N_A_471_47#_c_983_n N_VGND_c_1121_n 0.00193763f $X=8.275 $Y=0.82 $X2=0
+ $Y2=0
cc_591 N_A_471_47#_c_1017_n N_VGND_c_1121_n 0.0188551f $X=8.44 $Y=0.39 $X2=0
+ $Y2=0
cc_592 N_A_471_47#_c_984_n N_VGND_c_1121_n 0.00198695f $X=9.115 $Y=0.815 $X2=0
+ $Y2=0
cc_593 N_A_471_47#_c_984_n N_VGND_c_1123_n 0.00198695f $X=9.115 $Y=0.815 $X2=0
+ $Y2=0
cc_594 N_A_471_47#_c_985_n N_VGND_c_1123_n 0.0209752f $X=9.28 $Y=0.39 $X2=0
+ $Y2=0
cc_595 N_A_471_47#_M1003_s N_VGND_c_1124_n 0.00210147f $X=2.355 $Y=0.235 $X2=0
+ $Y2=0
cc_596 N_A_471_47#_M1011_s N_VGND_c_1124_n 0.00216833f $X=3.185 $Y=0.235 $X2=0
+ $Y2=0
cc_597 N_A_471_47#_M1004_d N_VGND_c_1124_n 0.00216833f $X=4.025 $Y=0.235 $X2=0
+ $Y2=0
cc_598 N_A_471_47#_M1016_d N_VGND_c_1124_n 0.00216833f $X=4.865 $Y=0.235 $X2=0
+ $Y2=0
cc_599 N_A_471_47#_M1038_s N_VGND_c_1124_n 0.00299586f $X=5.705 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_A_471_47#_M1000_d N_VGND_c_1124_n 0.00215201f $X=6.625 $Y=0.235 $X2=0
+ $Y2=0
cc_601 N_A_471_47#_M1009_d N_VGND_c_1124_n 0.00215201f $X=7.465 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_471_47#_M1017_s N_VGND_c_1124_n 0.00215201f $X=8.305 $Y=0.235 $X2=0
+ $Y2=0
cc_603 N_A_471_47#_M1028_s N_VGND_c_1124_n 0.00209319f $X=9.145 $Y=0.235 $X2=0
+ $Y2=0
cc_604 N_A_471_47#_c_1008_n N_VGND_c_1124_n 0.0122524f $X=5.92 $Y=0.39 $X2=0
+ $Y2=0
cc_605 N_A_471_47#_c_981_n N_VGND_c_1124_n 0.00827287f $X=6.595 $Y=0.82 $X2=0
+ $Y2=0
cc_606 N_A_471_47#_c_1012_n N_VGND_c_1124_n 0.0122069f $X=6.76 $Y=0.39 $X2=0
+ $Y2=0
cc_607 N_A_471_47#_c_982_n N_VGND_c_1124_n 0.00835832f $X=7.435 $Y=0.815 $X2=0
+ $Y2=0
cc_608 N_A_471_47#_c_1013_n N_VGND_c_1124_n 0.0122069f $X=7.6 $Y=0.39 $X2=0
+ $Y2=0
cc_609 N_A_471_47#_c_983_n N_VGND_c_1124_n 0.00827287f $X=8.275 $Y=0.82 $X2=0
+ $Y2=0
cc_610 N_A_471_47#_c_1017_n N_VGND_c_1124_n 0.0122069f $X=8.44 $Y=0.39 $X2=0
+ $Y2=0
cc_611 N_A_471_47#_c_984_n N_VGND_c_1124_n 0.00835832f $X=9.115 $Y=0.815 $X2=0
+ $Y2=0
cc_612 N_A_471_47#_c_985_n N_VGND_c_1124_n 0.0124119f $X=9.28 $Y=0.39 $X2=0
+ $Y2=0
cc_613 N_A_471_47#_c_986_n N_VGND_c_1124_n 0.0102047f $X=5.465 $Y=0.775 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__clkbuf_4.spice.pex
* Created: Thu Aug 27 14:11:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKBUF_4%A 3 7 9 10 14
c35 14 0 2.23144e-19 $X=0.51 $Y=1.16
r36 14 17 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=1.325
r37 14 16 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=0.995
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r39 10 15 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.16
r40 9 15 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.6 $Y=0.85 $X2=0.6
+ $Y2=1.16
r41 7 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r42 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 40 43
+ 45 48 49 54 60 62 71
c97 49 0 1.51549e-19 $X=1.115 $Y=1.16
c98 48 0 2.75502e-19 $X=1.03 $Y=1.495
r99 71 72 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=2.245 $Y=1.157
+ $X2=2.25 $Y2=1.157
r100 68 69 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=1.815 $Y=1.157
+ $X2=1.82 $Y2=1.157
r101 67 68 74.7628 $w=2.74e-07 $l=4.25e-07 $layer=POLY_cond $X=1.39 $Y=1.157
+ $X2=1.815 $Y2=1.157
r102 66 67 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=1.385 $Y=1.157
+ $X2=1.39 $Y2=1.157
r103 63 64 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=0.955 $Y=1.157
+ $X2=0.96 $Y2=1.157
r104 57 60 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r105 55 71 57.1715 $w=2.74e-07 $l=3.25e-07 $layer=POLY_cond $X=1.92 $Y=1.157
+ $X2=2.245 $Y2=1.157
r106 55 69 17.5912 $w=2.74e-07 $l=1e-07 $layer=POLY_cond $X=1.92 $Y=1.157
+ $X2=1.82 $Y2=1.157
r107 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r108 52 66 25.5073 $w=2.74e-07 $l=1.45e-07 $layer=POLY_cond $X=1.24 $Y=1.157
+ $X2=1.385 $Y2=1.157
r109 52 64 49.2555 $w=2.74e-07 $l=2.8e-07 $layer=POLY_cond $X=1.24 $Y=1.157
+ $X2=0.96 $Y2=1.157
r110 51 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.24 $Y=1.16
+ $X2=1.92 $Y2=1.16
r111 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.16 $X2=1.24 $Y2=1.16
r112 49 51 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.115 $Y=1.16
+ $X2=1.24 $Y2=1.16
r113 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=1.245
+ $X2=1.115 $Y2=1.16
r114 47 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.03 $Y=1.245
+ $X2=1.03 $Y2=1.495
r115 46 62 2.60907 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.58
+ $X2=0.24 $Y2=1.58
r116 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.945 $Y=1.58
+ $X2=1.03 $Y2=1.495
r117 45 46 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.945 $Y=1.58
+ $X2=0.395 $Y2=1.58
r118 41 62 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.58
r119 41 43 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.69
r120 40 62 3.84343 $w=2.4e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.17 $Y=1.495
+ $X2=0.24 $Y2=1.58
r121 39 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r122 39 40 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.495
r123 35 72 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=2.25 $Y=1.02
+ $X2=2.25 $Y2=1.157
r124 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.25 $Y=1.02
+ $X2=2.25 $Y2=0.445
r125 31 71 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=2.245 $Y=1.295
+ $X2=2.245 $Y2=1.157
r126 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.245 $Y=1.295
+ $X2=2.245 $Y2=1.985
r127 27 69 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=1.82 $Y=1.02
+ $X2=1.82 $Y2=1.157
r128 27 29 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.82 $Y=1.02
+ $X2=1.82 $Y2=0.445
r129 23 68 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=1.815 $Y=1.295
+ $X2=1.815 $Y2=1.157
r130 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.815 $Y=1.295
+ $X2=1.815 $Y2=1.985
r131 19 67 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=1.39 $Y=1.02
+ $X2=1.39 $Y2=1.157
r132 19 21 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.39 $Y=1.02
+ $X2=1.39 $Y2=0.445
r133 15 66 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=1.385 $Y=1.295
+ $X2=1.385 $Y2=1.157
r134 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.385 $Y=1.295
+ $X2=1.385 $Y2=1.985
r135 11 64 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=0.96 $Y=1.02
+ $X2=0.96 $Y2=1.157
r136 11 13 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.96 $Y=1.02
+ $X2=0.96 $Y2=0.445
r137 7 63 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=0.955 $Y=1.295
+ $X2=0.955 $Y2=1.157
r138 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.955 $Y=1.295
+ $X2=0.955 $Y2=1.985
r139 2 43 300 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.69
r140 1 60 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_4%VPWR 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r44 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r46 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 35 43 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.73 $Y=2.72
+ $X2=1.602 $Y2=2.72
r51 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.73 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 34 46 4.27389 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.547 $Y2=2.72
r53 34 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 30 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.72 $Y2=2.72
r58 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 29 43 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.602 $Y2=2.72
r60 29 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 24 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.72 $Y2=2.72
r62 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 22 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 18 46 3.12478 $w=2.85e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.477 $Y=2.635
+ $X2=2.547 $Y2=2.72
r66 18 20 28.5078 $w=2.83e-07 $l=7.05e-07 $layer=LI1_cond $X=2.477 $Y=2.635
+ $X2=2.477 $Y2=1.93
r67 14 43 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.602 $Y=2.635
+ $X2=1.602 $Y2=2.72
r68 14 16 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.602 $Y=2.635
+ $X2=1.602 $Y2=2.34
r69 10 40 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.72
r70 10 12 23.6065 $w=3.08e-07 $l=6.35e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2
r71 3 20 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.485 $X2=2.46 $Y2=1.93
r72 2 16 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.485 $X2=1.6 $Y2=2.34
r73 1 12 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_4%X 1 2 3 4 15 19 21 22 23 24 27 33 34 35 36
+ 46
c66 3 0 1.06215e-19 $X=1.03 $Y=1.485
r67 36 46 6.40246 $w=4.03e-07 $l=2.25e-07 $layer=LI1_cond $X=2.457 $Y=1.19
+ $X2=2.457 $Y2=1.415
r68 35 45 4.76257 $w=1.68e-07 $l=7.3e-08 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=2.457 $Y2=0.82
r69 35 36 7.68295 $w=4.03e-07 $l=2.7e-07 $layer=LI1_cond $X=2.457 $Y=0.92
+ $X2=2.457 $Y2=1.19
r70 35 45 0.426831 $w=4.03e-07 $l=1.5e-08 $layer=LI1_cond $X=2.457 $Y=0.92
+ $X2=2.457 $Y2=0.905
r71 34 46 25.2481 $w=1.68e-07 $l=3.87e-07 $layer=LI1_cond $X=2.07 $Y=1.5
+ $X2=2.457 $Y2=1.5
r72 34 42 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.07 $Y=1.5
+ $X2=2.035 $Y2=1.5
r73 34 42 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.035 $Y=1.6
+ $X2=2.035 $Y2=1.585
r74 31 34 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=2.035 $Y=1.835
+ $X2=2.035 $Y2=1.6
r75 31 33 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=1.835
+ $X2=2.035 $Y2=1.92
r76 25 45 27.5316 $w=1.68e-07 $l=4.22e-07 $layer=LI1_cond $X=2.035 $Y=0.82
+ $X2=2.457 $Y2=0.82
r77 25 27 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=2.035 $Y=0.735
+ $X2=2.035 $Y2=0.51
r78 23 33 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=1.92
+ $X2=2.035 $Y2=1.92
r79 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.905 $Y=1.92
+ $X2=1.305 $Y2=1.92
r80 21 25 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=0.82
+ $X2=2.035 $Y2=0.82
r81 21 22 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.905 $Y=0.82
+ $X2=1.305 $Y2=0.82
r82 17 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.175 $Y=2.005
+ $X2=1.305 $Y2=1.92
r83 17 19 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=1.175 $Y=2.005
+ $X2=1.175 $Y2=2.165
r84 13 22 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.157 $Y=0.735
+ $X2=1.305 $Y2=0.82
r85 13 15 8.78982 $w=2.93e-07 $l=2.25e-07 $layer=LI1_cond $X=1.157 $Y=0.735
+ $X2=1.157 $Y2=0.51
r86 4 34 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.03 $Y2=1.62
r87 4 33 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=1.485 $X2=2.03 $Y2=1.96
r88 3 19 600 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.17 $Y2=2.165
r89 2 27 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.035 $Y2=0.51
r90 1 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.175 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_4%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r45 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r47 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r49 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r50 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r51 35 43 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.602
+ $Y2=0
r52 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=2.07
+ $Y2=0
r53 34 46 4.22854 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.547
+ $Y2=0
r54 34 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.07
+ $Y2=0
r55 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r56 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r57 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 30 40 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r59 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.15
+ $Y2=0
r60 29 43 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.602
+ $Y2=0
r61 29 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.15
+ $Y2=0
r62 24 40 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r63 24 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.23
+ $Y2=0
r64 22 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 18 46 3.13151 $w=2.8e-07 $l=1.15521e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.547 $Y2=0
r67 18 20 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.4
r68 14 43 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0
r69 14 16 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0.4
r70 10 40 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r71 10 12 13.2007 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.4
r72 3 20 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.465 $Y2=0.4
r73 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.235 $X2=1.605 $Y2=0.4
r74 1 12 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.4
.ends


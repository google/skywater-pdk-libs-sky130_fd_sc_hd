* File: sky130_fd_sc_hd__a41o_1.pex.spice
* Created: Tue Sep  1 18:56:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A41O_1%A_79_21# 1 2 9 12 17 18 19 20 21 22 25 29 32
r66 27 29 9.7194 $w=4.13e-07 $l=3.5e-07 $layer=LI1_cond $X=1.322 $Y=0.735
+ $X2=1.322 $Y2=0.385
r67 23 25 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=1.995 $X2=1.2
+ $Y2=2
r68 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.035 $Y=1.91
+ $X2=1.2 $Y2=1.995
r69 21 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.035 $Y=1.91
+ $X2=0.685 $Y2=1.91
r70 19 27 28.1438 $w=8.8e-08 $l=2.45854e-07 $layer=LI1_cond $X=1.115 $Y=0.82
+ $X2=1.322 $Y2=0.735
r71 19 20 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.115 $Y=0.82
+ $X2=0.685 $Y2=0.82
r72 18 33 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.565 $Y2=1.325
r73 18 32 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.565 $Y2=0.995
r74 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r75 15 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=1.825
+ $X2=0.685 $Y2=1.91
r76 15 17 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=0.6 $Y=1.825 $X2=0.6
+ $Y2=1.16
r77 14 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.905
+ $X2=0.685 $Y2=0.82
r78 14 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.6 $Y=0.905
+ $X2=0.6 $Y2=1.16
r79 12 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r80 9 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
r81 2 25 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2
r82 1 29 91 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_NDIFF $count=2 $X=1.19
+ $Y=0.235 $X2=1.365 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%B1 1 3 6 8 9 17
c34 8 0 1.8994e-19 $X=1.175 $Y=1.19
r35 15 17 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.41 $Y2=1.16
r36 12 15 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=1.17 $Y2=1.16
r37 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.16 $X2=1.17
+ $Y2=1.53
r38 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r39 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r40 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325 $X2=1.41
+ $Y2=1.985
r41 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=0.995
+ $X2=1.115 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.115 $Y=0.995
+ $X2=1.115 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%A1 1 3 6 8 11
c34 11 0 2.19281e-19 $X=1.83 $Y=1.16
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.16 $X2=1.83 $Y2=1.16
r36 8 12 13.1988 $w=3.42e-07 $l=3.7e-07 $layer=LI1_cond $X=1.725 $Y=1.53
+ $X2=1.725 $Y2=1.16
r37 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.16
r38 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=1.985
r39 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.995 $X2=1.83
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%A2 3 6 10 11 13 14 18 20
r40 13 20 8.57297 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=2.095 $Y=0.507
+ $X2=2.225 $Y2=0.507
r41 11 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.16
+ $X2=2.31 $Y2=1.325
r42 11 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.16
+ $X2=2.31 $Y2=0.995
r43 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.16 $X2=2.31 $Y2=1.16
r44 8 14 13.1892 $w=1.83e-07 $l=2.2e-07 $layer=LI1_cond $X=2.335 $Y=0.507
+ $X2=2.555 $Y2=0.507
r45 8 20 6.59459 $w=1.83e-07 $l=1.1e-07 $layer=LI1_cond $X=2.335 $Y=0.507
+ $X2=2.225 $Y2=0.507
r46 8 10 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.335 $Y=0.6
+ $X2=2.335 $Y2=1.16
r47 6 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.985
+ $X2=2.25 $Y2=1.325
r48 3 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.25 $Y=0.56 $X2=2.25
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%A3 3 6 8 9 10 11 18 20 30
r38 28 30 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=2.895 $Y=1.185
+ $X2=2.895 $Y2=1.19
r39 19 28 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.895 $Y=1.16
+ $X2=2.895 $Y2=1.185
r40 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.16
+ $X2=2.79 $Y2=1.325
r41 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.16
+ $X2=2.79 $Y2=0.995
r42 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.16 $X2=2.79 $Y2=1.16
r43 10 19 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.895 $Y=1.145
+ $X2=2.895 $Y2=1.16
r44 10 36 6.97733 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.895 $Y=1.145
+ $X2=2.895 $Y2=0.995
r45 10 11 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=2.895 $Y=1.23
+ $X2=2.895 $Y2=1.53
r46 10 30 1.2131 $w=3.78e-07 $l=4e-08 $layer=LI1_cond $X=2.895 $Y=1.23 $X2=2.895
+ $Y2=1.19
r47 9 36 7.84479 $w=2.03e-07 $l=1.45e-07 $layer=LI1_cond $X=2.982 $Y=0.85
+ $X2=2.982 $Y2=0.995
r48 8 9 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=2.982 $Y=0.51
+ $X2=2.982 $Y2=0.85
r49 6 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.985
+ $X2=2.73 $Y2=1.325
r50 3 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.56 $X2=2.73
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%A4 1 3 6 8 9 15
r26 12 15 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.44 $Y2=1.16
r27 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.442 $Y=1.16
+ $X2=3.442 $Y2=1.53
r28 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r29 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.325 $X2=3.21
+ $Y2=1.985
r31 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995 $X2=3.21
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%X 1 2 7 8 9 10 11 12 38 42 45
r16 45 46 2.19202 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.255 $Y=2.21
+ $X2=0.255 $Y2=2.165
r17 42 43 2.36149 $w=3.38e-07 $l=5e-08 $layer=LI1_cond $X=0.255 $Y=0.51
+ $X2=0.255 $Y2=0.56
r18 12 49 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=0.255 $Y=2.23
+ $X2=0.255 $Y2=2.34
r19 12 45 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.255 $Y=2.23
+ $X2=0.255 $Y2=2.21
r20 12 46 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=0.215 $Y=2.145
+ $X2=0.215 $Y2=2.165
r21 11 12 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=2.145
r22 11 33 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=1.66
r23 10 33 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.53
+ $X2=0.215 $Y2=1.66
r24 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.215 $Y=1.19
+ $X2=0.215 $Y2=1.53
r25 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.215 $Y=0.85
+ $X2=0.215 $Y2=1.19
r26 8 25 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.85
+ $X2=0.215 $Y2=0.725
r27 7 42 0.610117 $w=3.38e-07 $l=1.8e-08 $layer=LI1_cond $X=0.255 $Y=0.492
+ $X2=0.255 $Y2=0.51
r28 7 38 3.62681 $w=3.38e-07 $l=1.07e-07 $layer=LI1_cond $X=0.255 $Y=0.492
+ $X2=0.255 $Y2=0.385
r29 7 25 6.56006 $w=2.58e-07 $l=1.48e-07 $layer=LI1_cond $X=0.215 $Y=0.577
+ $X2=0.215 $Y2=0.725
r30 7 43 0.75352 $w=2.58e-07 $l=1.7e-08 $layer=LI1_cond $X=0.215 $Y=0.577
+ $X2=0.215 $Y2=0.56
r31 2 49 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r32 2 33 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r33 1 38 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
r34 1 25 182 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%VPWR 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r66 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r71 39 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=2.72
+ $X2=2.97 $Y2=2.72
r72 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.095 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r76 35 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.04 $Y2=2.72
r77 35 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 34 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.97 $Y2=2.72
r79 34 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r81 33 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r83 30 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.72 $Y2=2.72
r84 30 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r85 29 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.04 $Y2=2.72
r86 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r87 24 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.72 $Y2=2.72
r88 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 18 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2.72
r92 18 20 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2.34
r93 14 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r94 14 16 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.34
r95 10 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.72
r96 10 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.34
r97 3 20 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.485 $X2=2.97 $Y2=2.34
r98 2 16 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2.34
r99 1 12 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%A_297_297# 1 2 3 12 16 21 23 25
c35 21 0 2.93415e-20 $X=1.62 $Y=1.96
r36 17 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.88
+ $X2=2.46 $Y2=1.88
r37 16 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.88
+ $X2=3.42 $Y2=1.88
r38 16 17 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.335 $Y=1.88
+ $X2=2.545 $Y2=1.88
r39 13 21 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.88
+ $X2=1.62 $Y2=1.88
r40 12 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=1.88
+ $X2=2.46 $Y2=1.88
r41 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.375 $Y=1.88
+ $X2=1.705 $Y2=1.88
r42 3 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.96
r43 2 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.96
r44 1 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_1%VGND 1 2 9 11 13 15 17 22 31 35
r48 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r50 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r51 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r53 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r54 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r55 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r56 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.76
+ $Y2=0
r57 23 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r58 22 34 4.90987 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r59 22 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r60 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.76
+ $Y2=0
r61 17 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r62 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r63 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r64 11 34 2.94129 $w=3.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.467 $Y2=0
r65 11 13 10.1686 $w=3.38e-07 $l=3e-07 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.425 $Y2=0.385
r66 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r67 7 9 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.48
r68 2 13 91 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.385
r69 1 9 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.76 $Y2=0.48
.ends


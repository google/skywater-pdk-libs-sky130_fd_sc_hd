* File: sky130_fd_sc_hd__or3_4.spice.pex
* Created: Thu Aug 27 14:43:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR3_4%C 1 3 6 8 14
c28 8 0 1.91457e-19 $X=0.235 $Y=1.19
r29 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r31 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r33 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_4%B 1 3 6 12 13 15 16
c39 13 0 1.91457e-19 $X=0.89 $Y=1.16
r40 15 16 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.712 $Y=1.53
+ $X2=0.712 $Y2=1.87
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r42 9 15 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.53
r43 8 12 8.20539 $w=2.48e-07 $l=1.78e-07 $layer=LI1_cond $X=0.712 $Y=1.2
+ $X2=0.89 $Y2=1.2
r44 8 9 1.11538 $w=2.35e-07 $l=1.25e-07 $layer=LI1_cond $X=0.712 $Y=1.2
+ $X2=0.712 $Y2=1.325
r45 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r46 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r47 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_4%A 3 6 8 11 13
c40 11 0 1.83425e-19 $X=1.39 $Y=1.16
r41 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.38 $Y2=1.325
r42 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.38 $Y2=0.995
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.16 $X2=1.39 $Y2=1.16
r44 8 12 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=1.615 $Y=1.2 $X2=1.39
+ $Y2=1.2
r45 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=1.325
r46 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.56 $X2=1.31
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_4%A_27_47# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 40 42 44 46 47 48 52 55 56 58 59 61 63 66 71 73 81
c159 63 0 1.83425e-19 $X=1.98 $Y=1.495
r160 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.68 $Y=1.16
+ $X2=3.1 $Y2=1.16
r161 77 78 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.68 $Y2=1.16
r162 74 77 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.065 $Y=1.16
+ $X2=2.26 $Y2=1.16
r163 73 74 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.065
+ $Y=1.16 $X2=2.065 $Y2=1.16
r164 67 81 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.425 $Y=1.16
+ $X2=3.52 $Y2=1.16
r165 67 79 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.425 $Y=1.16
+ $X2=3.1 $Y2=1.16
r166 66 67 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.425
+ $Y=1.16 $X2=3.425 $Y2=1.16
r167 64 73 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.09 $Y=1.16
+ $X2=1.98 $Y2=1.16
r168 64 66 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=2.09 $Y=1.16
+ $X2=3.425 $Y2=1.16
r169 62 73 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.245
+ $X2=1.98 $Y2=1.16
r170 62 63 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=1.98 $Y=1.245
+ $X2=1.98 $Y2=1.495
r171 61 73 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.075
+ $X2=1.98 $Y2=1.16
r172 60 61 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=1.98 $Y=0.905
+ $X2=1.98 $Y2=1.075
r173 58 63 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.87 $Y=1.58
+ $X2=1.98 $Y2=1.495
r174 58 59 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.87 $Y=1.58
+ $X2=1.265 $Y2=1.58
r175 57 71 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0.815
+ $X2=1.1 $Y2=0.815
r176 56 60 6.90553 $w=1.8e-07 $l=1.48324e-07 $layer=LI1_cond $X=1.87 $Y=0.815
+ $X2=1.98 $Y2=0.905
r177 56 57 37.2778 $w=1.78e-07 $l=6.05e-07 $layer=LI1_cond $X=1.87 $Y=0.815
+ $X2=1.265 $Y2=0.815
r178 54 59 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.132 $Y=1.665
+ $X2=1.265 $Y2=1.58
r179 54 55 27.3977 $w=2.63e-07 $l=6.3e-07 $layer=LI1_cond $X=1.132 $Y=1.665
+ $X2=1.132 $Y2=2.295
r180 50 71 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.1 $Y=0.725 $X2=1.1
+ $Y2=0.815
r181 50 52 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.1 $Y=0.725
+ $X2=1.1 $Y2=0.4
r182 49 70 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.255 $Y2=2.38
r183 48 55 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=1 $Y=2.38
+ $X2=1.132 $Y2=2.295
r184 48 49 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1 $Y=2.38
+ $X2=0.425 $Y2=2.38
r185 46 71 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.815
+ $X2=1.1 $Y2=0.815
r186 46 47 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.815
+ $X2=0.425 $Y2=0.815
r187 42 70 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.295
+ $X2=0.255 $Y2=2.38
r188 42 44 21.5236 $w=3.38e-07 $l=6.35e-07 $layer=LI1_cond $X=0.255 $Y=2.295
+ $X2=0.255 $Y2=1.66
r189 38 47 7.6914 $w=1.8e-07 $l=2.10238e-07 $layer=LI1_cond $X=0.255 $Y=0.725
+ $X2=0.425 $Y2=0.815
r190 38 40 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=0.255 $Y=0.725
+ $X2=0.255 $Y2=0.4
r191 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.16
r192 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.985
r193 31 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=0.995
+ $X2=3.52 $Y2=1.16
r194 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.52 $Y=0.995
+ $X2=3.52 $Y2=0.56
r195 27 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.325
+ $X2=3.1 $Y2=1.16
r196 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.1 $Y=1.325
+ $X2=3.1 $Y2=1.985
r197 24 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=0.995
+ $X2=3.1 $Y2=1.16
r198 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.1 $Y=0.995
+ $X2=3.1 $Y2=0.56
r199 20 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.325
+ $X2=2.68 $Y2=1.16
r200 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.68 $Y=1.325
+ $X2=2.68 $Y2=1.985
r201 17 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=0.995
+ $X2=2.68 $Y2=1.16
r202 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.68 $Y=0.995
+ $X2=2.68 $Y2=0.56
r203 13 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.325
+ $X2=2.26 $Y2=1.16
r204 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.26 $Y=1.325
+ $X2=2.26 $Y2=1.985
r205 10 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.995
+ $X2=2.26 $Y2=1.16
r206 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.26 $Y=0.995
+ $X2=2.26 $Y2=0.56
r207 3 70 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r208 3 44 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r209 2 52 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r210 1 40 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_4%VPWR 1 2 3 12 16 20 23 24 25 26 27 28 30 47 49
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r55 44 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 41 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 38 49 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=1.785 $Y2=2.72
r61 38 40 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 32 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 30 49 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.785 $Y2=2.72
r66 30 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 28 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 28 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 26 43 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.605 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.605 $Y=2.72
+ $X2=3.73 $Y2=2.72
r71 25 46 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.73 $Y2=2.72
r73 23 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.765 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=2.72
+ $X2=2.89 $Y2=2.72
r75 22 43 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.015 $Y=2.72
+ $X2=3.45 $Y2=2.72
r76 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=2.72
+ $X2=2.89 $Y2=2.72
r77 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=2.635
+ $X2=3.73 $Y2=2.72
r78 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.73 $Y=2.635
+ $X2=3.73 $Y2=1.96
r79 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=2.635
+ $X2=2.89 $Y2=2.72
r80 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.89 $Y=2.635
+ $X2=2.89 $Y2=1.96
r81 10 49 2.86223 $w=7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=2.635
+ $X2=1.785 $Y2=2.72
r82 10 12 10.8501 $w=6.98e-07 $l=6.35e-07 $layer=LI1_cond $X=1.785 $Y=2.635
+ $X2=1.785 $Y2=2
r83 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.595
+ $Y=1.485 $X2=3.73 $Y2=1.96
r84 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.755
+ $Y=1.485 $X2=2.89 $Y2=1.96
r85 1 12 150 $w=1.7e-07 $l=8.85833e-07 $layer=licon1_PDIFF $count=4 $X=1.385
+ $Y=1.485 $X2=2.05 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_4%X 1 2 3 4 15 17 19 21 23 24 27 31 33 35 39 41
+ 43 46
r77 43 46 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=0.82 $X2=3.91
+ $Y2=0.905
r78 43 46 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=3.91 $Y=0.92
+ $X2=3.91 $Y2=0.905
r79 42 43 21.2606 $w=2.88e-07 $l=5.35e-07 $layer=LI1_cond $X=3.91 $Y=1.455
+ $X2=3.91 $Y2=0.92
r80 36 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0.82
+ $X2=3.31 $Y2=0.82
r81 35 43 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.765 $Y=0.82
+ $X2=3.91 $Y2=0.82
r82 35 36 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.765 $Y=0.82
+ $X2=3.475 $Y2=0.82
r83 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.435 $Y=1.54
+ $X2=3.31 $Y2=1.54
r84 33 42 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.765 $Y=1.54
+ $X2=3.91 $Y2=1.455
r85 33 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.765 $Y=1.54
+ $X2=3.435 $Y2=1.54
r86 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=1.625
+ $X2=3.31 $Y2=1.54
r87 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.31 $Y=1.625
+ $X2=3.31 $Y2=2.3
r88 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=0.735
+ $X2=3.31 $Y2=0.82
r89 25 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.31 $Y=0.735
+ $X2=3.31 $Y2=0.39
r90 23 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0.82
+ $X2=3.31 $Y2=0.82
r91 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.145 $Y=0.82
+ $X2=2.635 $Y2=0.82
r92 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.595 $Y=1.54
+ $X2=2.47 $Y2=1.54
r93 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.185 $Y=1.54
+ $X2=3.31 $Y2=1.54
r94 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.185 $Y=1.54
+ $X2=2.595 $Y2=1.54
r95 17 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=1.625
+ $X2=2.47 $Y2=1.54
r96 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.47 $Y=1.625
+ $X2=2.47 $Y2=2.3
r97 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.47 $Y=0.735
+ $X2=2.635 $Y2=0.82
r98 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.47 $Y=0.735
+ $X2=2.47 $Y2=0.39
r99 4 41 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.485 $X2=3.31 $Y2=1.62
r100 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.485 $X2=3.31 $Y2=2.3
r101 3 38 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.47 $Y2=1.62
r102 3 19 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.47 $Y2=2.3
r103 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.175
+ $Y=0.235 $X2=3.31 $Y2=0.39
r104 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.335
+ $Y=0.235 $X2=2.47 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_4%VGND 1 2 3 4 15 19 23 26 27 29 30 32 33 34 52
+ 53 58 61
r70 60 61 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=0.235
+ $X2=2.135 $Y2=0.235
r71 56 60 8.22304 $w=6.38e-07 $l=4.4e-07 $layer=LI1_cond $X=1.61 $Y=0.235
+ $X2=2.05 $Y2=0.235
r72 56 58 10.6037 $w=6.38e-07 $l=1.75e-07 $layer=LI1_cond $X=1.61 $Y=0.235
+ $X2=1.435 $Y2=0.235
r73 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r75 50 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r76 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r77 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r78 47 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r79 46 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.135
+ $Y2=0
r80 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r81 43 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r82 42 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.435
+ $Y2=0
r83 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r84 34 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r85 34 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r86 32 49 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.45
+ $Y2=0
r87 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.73
+ $Y2=0
r88 31 52 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.91
+ $Y2=0
r89 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.73
+ $Y2=0
r90 29 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.53
+ $Y2=0
r91 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.89
+ $Y2=0
r92 28 49 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.45
+ $Y2=0
r93 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.89
+ $Y2=0
r94 26 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r95 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r96 25 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.15
+ $Y2=0
r97 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r98 21 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0
r99 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0.39
r100 17 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0
r101 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.89 $Y=0.085
+ $X2=2.89 $Y2=0.39
r102 13 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r103 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.39
r104 4 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.235 $X2=3.73 $Y2=0.39
r105 3 19 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.235 $X2=2.89 $Y2=0.39
r106 2 60 91 $w=1.7e-07 $l=7.38444e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=2.05 $Y2=0.39
r107 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends


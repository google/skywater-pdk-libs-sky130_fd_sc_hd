* File: sky130_fd_sc_hd__clkinvlp_2.pxi.spice
* Created: Thu Aug 27 14:12:58 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINVLP_2%A N_A_M1000_g N_A_c_29_n N_A_M1003_g N_A_c_30_n
+ N_A_c_31_n N_A_M1001_g N_A_M1002_g N_A_c_33_n N_A_c_34_n N_A_c_35_n A A
+ N_A_c_36_n PM_SKY130_FD_SC_HD__CLKINVLP_2%A
x_PM_SKY130_FD_SC_HD__CLKINVLP_2%VPWR N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_c_70_n N_VPWR_c_71_n N_VPWR_c_72_n N_VPWR_c_73_n VPWR N_VPWR_c_74_n
+ N_VPWR_c_69_n PM_SKY130_FD_SC_HD__CLKINVLP_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKINVLP_2%Y N_Y_M1001_d N_Y_M1000_d Y Y Y
+ PM_SKY130_FD_SC_HD__CLKINVLP_2%Y
x_PM_SKY130_FD_SC_HD__CLKINVLP_2%VGND N_VGND_M1003_s N_VGND_c_111_n
+ N_VGND_c_112_n N_VGND_c_113_n VGND N_VGND_c_114_n N_VGND_c_115_n
+ PM_SKY130_FD_SC_HD__CLKINVLP_2%VGND
cc_1 VNB N_A_c_29_n 0.0209738f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.995
cc_2 VNB N_A_c_30_n 0.00843475f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.082
cc_3 VNB N_A_c_31_n 0.0199958f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.99
cc_4 VNB N_A_M1002_g 0.0119835f $X=-0.19 $Y=-0.24 $X2=1.185 $Y2=1.985
cc_5 VNB N_A_c_33_n 0.0406229f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.155
cc_6 VNB N_A_c_34_n 0.0125088f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.155
cc_7 VNB N_A_c_35_n 0.0208311f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.08
cc_8 VNB N_A_c_36_n 0.00936522f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_9 VNB N_VPWR_c_69_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.372 $Y2=1.19
cc_10 VNB Y 0.0226948f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.61
cc_11 VNB Y 0.00600055f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.082
cc_12 VNB N_VGND_c_111_n 0.0239026f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.61
cc_13 VNB N_VGND_c_112_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.082
cc_14 VNB N_VGND_c_113_n 0.00589254f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.99
cc_15 VNB N_VGND_c_114_n 0.0351227f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_16 VNB N_VGND_c_115_n 0.149697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VPB N_A_M1000_g 0.0294005f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.985
cc_18 VPB N_A_M1002_g 0.0333682f $X=-0.19 $Y=1.305 $X2=1.185 $Y2=1.985
cc_19 VPB N_A_c_33_n 0.0119035f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.155
cc_20 VPB N_A_c_34_n 4.36774e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.155
cc_21 VPB N_A_c_36_n 0.0179329f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_22 VPB N_VPWR_c_70_n 0.0146623f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=0.61
cc_23 VPB N_VPWR_c_71_n 0.0278706f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.082
cc_24 VPB N_VPWR_c_72_n 0.0113758f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=0.61
cc_25 VPB N_VPWR_c_73_n 0.0570286f $X=-0.19 $Y=1.305 $X2=1.185 $Y2=1.17
cc_26 VPB N_VPWR_c_74_n 0.0231642f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.08
cc_27 VPB N_VPWR_c_69_n 0.0483895f $X=-0.19 $Y=1.305 $X2=0.372 $Y2=1.19
cc_28 VPB Y 0.00146391f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.082
cc_29 N_A_c_36_n N_VPWR_M1000_s 0.00310055f $X=0.515 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_30 N_A_M1000_g N_VPWR_c_71_n 0.0159201f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_31 N_A_M1002_g N_VPWR_c_71_n 0.00122857f $X=1.185 $Y=1.985 $X2=0 $Y2=0
cc_32 N_A_c_33_n N_VPWR_c_71_n 0.00106175f $X=0.53 $Y=1.155 $X2=0 $Y2=0
cc_33 N_A_c_36_n N_VPWR_c_71_n 0.0243702f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_34 N_A_M1002_g N_VPWR_c_73_n 0.028251f $X=1.185 $Y=1.985 $X2=0 $Y2=0
cc_35 N_A_M1000_g N_VPWR_c_74_n 0.00894766f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_36 N_A_M1002_g N_VPWR_c_74_n 0.00725938f $X=1.185 $Y=1.985 $X2=0 $Y2=0
cc_37 N_A_M1000_g N_VPWR_c_69_n 0.0143885f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_38 N_A_M1002_g N_VPWR_c_69_n 0.0115385f $X=1.185 $Y=1.985 $X2=0 $Y2=0
cc_39 N_A_c_29_n Y 0.0102147f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_40 N_A_c_31_n Y 0.0119755f $X=1.065 $Y=0.99 $X2=0 $Y2=0
cc_41 N_A_c_35_n Y 0.00318327f $X=1.15 $Y=1.08 $X2=0 $Y2=0
cc_42 N_A_c_30_n Y 0.00962668f $X=0.99 $Y=1.082 $X2=0 $Y2=0
cc_43 N_A_c_31_n Y 0.00850094f $X=1.065 $Y=0.99 $X2=0 $Y2=0
cc_44 N_A_M1002_g Y 0.0473616f $X=1.185 $Y=1.985 $X2=0 $Y2=0
cc_45 N_A_c_34_n Y 0.00415735f $X=0.655 $Y=1.155 $X2=0 $Y2=0
cc_46 N_A_c_35_n Y 0.0139081f $X=1.15 $Y=1.08 $X2=0 $Y2=0
cc_47 N_A_c_36_n Y 0.0397302f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_48 N_A_c_29_n N_VGND_c_111_n 0.0118628f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A_c_31_n N_VGND_c_111_n 9.92377e-19 $X=1.065 $Y=0.99 $X2=0 $Y2=0
cc_50 N_A_c_33_n N_VGND_c_111_n 0.00207251f $X=0.53 $Y=1.155 $X2=0 $Y2=0
cc_51 N_A_c_36_n N_VGND_c_111_n 0.0177327f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_c_29_n N_VGND_c_114_n 0.00407525f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_53 N_A_c_31_n N_VGND_c_114_n 0.00306164f $X=1.065 $Y=0.99 $X2=0 $Y2=0
cc_54 N_A_c_29_n N_VGND_c_115_n 0.00772944f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_55 N_A_c_31_n N_VGND_c_115_n 0.00436513f $X=1.065 $Y=0.99 $X2=0 $Y2=0
cc_56 N_VPWR_c_69_n N_Y_M1000_d 0.00332766f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_57 N_VPWR_c_73_n Y 0.0680398f $X=1.575 $Y=1.63 $X2=0 $Y2=0
cc_58 N_VPWR_c_74_n Y 0.0264844f $X=1.44 $Y=2.715 $X2=0 $Y2=0
cc_59 N_VPWR_c_69_n Y 0.0152919f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_60 Y N_VGND_c_111_n 0.0329647f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_61 Y N_VGND_c_114_n 0.0320436f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_62 Y N_VGND_c_115_n 0.0228211f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_63 Y A_150_67# 0.00365392f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_64 Y A_150_67# 0.00164634f $X=1.065 $Y=0.765 $X2=-0.19 $Y2=-0.24

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_1647_49# a_721_47# a_1636_315# VPB phighvt w=840000u l=150000u
+  ad=2.268e+11p pd=2.22e+06u as=4.834e+11p ps=4.73e+06u
M1001 VGND a_1636_315# a_1565_49# VNB nshort w=640000u l=150000u
+  ad=8.644e+11p pd=7.87e+06u as=3.392e+11p ps=3.62e+06u
M1002 VPWR a_1636_315# a_1565_49# VPB phighvt w=1e+06u l=150000u
+  ad=1.25e+12p pd=1.05e+07u as=8.984e+11p ps=3.96e+06u
M1003 a_67_199# a_489_21# a_434_49# VPB phighvt w=840000u l=150000u
+  ad=8.1155e+11p pd=7.43e+06u as=2.31e+11p ps=2.23e+06u
M1004 VPWR B a_489_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1005 a_434_49# B a_67_199# VNB nshort w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=8.10575e+11p ps=5.12e+06u
M1006 a_1142_49# a_489_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=7.652e+11p pd=3.58e+06u as=0p ps=0u
M1007 VGND a_67_199# a_27_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=5.3225e+11p ps=5.52e+06u
M1008 VGND CIN a_1251_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1009 a_1251_49# a_721_47# COUT VPB phighvt w=840000u l=150000u
+  ad=9.633e+11p pd=5.88e+06u as=2.268e+11p ps=2.22e+06u
M1010 a_67_199# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_67_199# B a_721_47# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=3.04525e+11p ps=2.6e+06u
M1012 a_27_47# B a_721_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.3135e+11p ps=2.33e+06u
M1013 VPWR a_67_199# a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=8.677e+11p ps=7.94e+06u
M1014 a_1142_49# a_721_47# COUT VNB nshort w=640000u l=150000u
+  ad=3.456e+11p pd=3.64e+06u as=1.76e+11p ps=1.83e+06u
M1015 VGND B a_489_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.65325e+11p ps=1.82e+06u
M1016 a_1636_315# CIN VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 SUM a_1647_49# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1018 a_67_199# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1636_315# a_434_49# a_1647_49# VNB nshort w=640000u l=150000u
+  ad=6.458e+11p pd=4.59e+06u as=1.856e+11p ps=1.86e+06u
M1020 a_721_47# a_489_21# a_27_47# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR CIN a_1251_49# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1636_315# CIN VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1565_49# a_434_49# a_1647_49# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1142_49# a_489_21# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 SUM a_1647_49# VGND VNB nshort w=650000u l=150000u
+  ad=1.8525e+11p pd=1.87e+06u as=0p ps=0u
M1026 a_27_47# a_489_21# a_434_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_434_49# B a_27_47# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_721_47# a_489_21# a_67_199# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1647_49# a_721_47# a_1565_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 COUT a_434_49# a_1142_49# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 COUT a_434_49# a_1251_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

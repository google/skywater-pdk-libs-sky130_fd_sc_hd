* File: sky130_fd_sc_hd__nand4bb_4.pxi.spice
* Created: Tue Sep  1 19:17:28 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4BB_4%A_N N_A_N_c_153_n N_A_N_M1031_g N_A_N_M1023_g
+ A_N A_N N_A_N_c_155_n PM_SKY130_FD_SC_HD__NAND4BB_4%A_N
x_PM_SKY130_FD_SC_HD__NAND4BB_4%B_N N_B_N_c_178_n N_B_N_M1015_g N_B_N_M1006_g
+ B_N B_N N_B_N_c_179_n N_B_N_c_180_n PM_SKY130_FD_SC_HD__NAND4BB_4%B_N
x_PM_SKY130_FD_SC_HD__NAND4BB_4%A_27_47# N_A_27_47#_M1031_s N_A_27_47#_M1023_s
+ N_A_27_47#_c_212_n N_A_27_47#_M1014_g N_A_27_47#_M1007_g N_A_27_47#_M1019_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1021_g N_A_27_47#_M1018_g N_A_27_47#_c_217_n
+ N_A_27_47#_M1027_g N_A_27_47#_M1024_g N_A_27_47#_c_220_n N_A_27_47#_c_229_n
+ N_A_27_47#_c_234_n N_A_27_47#_c_221_n N_A_27_47#_c_237_n N_A_27_47#_c_230_n
+ N_A_27_47#_c_222_n N_A_27_47#_c_273_p N_A_27_47#_c_223_n
+ PM_SKY130_FD_SC_HD__NAND4BB_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_4%A_193_47# N_A_193_47#_M1015_d
+ N_A_193_47#_M1006_d N_A_193_47#_M1017_g N_A_193_47#_M1000_g
+ N_A_193_47#_M1025_g N_A_193_47#_M1001_g N_A_193_47#_M1028_g
+ N_A_193_47#_M1011_g N_A_193_47#_M1034_g N_A_193_47#_M1030_g
+ N_A_193_47#_c_371_n N_A_193_47#_c_363_n N_A_193_47#_c_364_n
+ N_A_193_47#_c_372_n N_A_193_47#_c_395_n N_A_193_47#_c_365_n
+ N_A_193_47#_c_400_n N_A_193_47#_c_403_n N_A_193_47#_c_373_n
+ N_A_193_47#_c_405_n N_A_193_47#_c_366_n
+ PM_SKY130_FD_SC_HD__NAND4BB_4%A_193_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_4%C N_C_M1003_g N_C_M1012_g N_C_M1022_g
+ N_C_M1016_g N_C_M1032_g N_C_M1020_g N_C_M1033_g N_C_M1026_g C C C C
+ N_C_c_500_n N_C_c_501_n N_C_c_502_n PM_SKY130_FD_SC_HD__NAND4BB_4%C
x_PM_SKY130_FD_SC_HD__NAND4BB_4%D N_D_M1002_g N_D_M1004_g N_D_M1005_g
+ N_D_M1009_g N_D_M1008_g N_D_M1013_g N_D_M1029_g N_D_M1035_g D D D D
+ N_D_c_582_n N_D_c_583_n PM_SKY130_FD_SC_HD__NAND4BB_4%D
x_PM_SKY130_FD_SC_HD__NAND4BB_4%VPWR N_VPWR_M1023_d N_VPWR_M1007_d
+ N_VPWR_M1010_d N_VPWR_M1024_d N_VPWR_M1001_d N_VPWR_M1030_d N_VPWR_M1016_d
+ N_VPWR_M1026_d N_VPWR_M1009_s N_VPWR_M1035_s N_VPWR_c_652_n N_VPWR_c_653_n
+ N_VPWR_c_654_n N_VPWR_c_655_n N_VPWR_c_656_n N_VPWR_c_657_n N_VPWR_c_658_n
+ N_VPWR_c_659_n N_VPWR_c_660_n N_VPWR_c_661_n N_VPWR_c_662_n N_VPWR_c_663_n
+ N_VPWR_c_664_n N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n
+ N_VPWR_c_669_n N_VPWR_c_670_n N_VPWR_c_671_n N_VPWR_c_672_n VPWR
+ N_VPWR_c_673_n N_VPWR_c_674_n N_VPWR_c_675_n N_VPWR_c_676_n N_VPWR_c_677_n
+ N_VPWR_c_678_n N_VPWR_c_679_n N_VPWR_c_680_n N_VPWR_c_651_n
+ PM_SKY130_FD_SC_HD__NAND4BB_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND4BB_4%Y N_Y_M1014_d N_Y_M1021_d N_Y_M1007_s
+ N_Y_M1018_s N_Y_M1000_s N_Y_M1011_s N_Y_M1012_s N_Y_M1020_s N_Y_M1004_d
+ N_Y_M1013_d N_Y_c_801_n N_Y_c_825_n N_Y_c_803_n N_Y_c_804_n N_Y_c_833_n
+ N_Y_c_836_n N_Y_c_805_n N_Y_c_858_n N_Y_c_806_n N_Y_c_883_n N_Y_c_807_n
+ N_Y_c_890_n N_Y_c_808_n N_Y_c_894_n N_Y_c_809_n N_Y_c_810_n N_Y_c_916_n
+ N_Y_c_811_n N_Y_c_812_n N_Y_c_813_n N_Y_c_814_n N_Y_c_815_n N_Y_c_816_n Y Y
+ N_Y_c_846_n PM_SKY130_FD_SC_HD__NAND4BB_4%Y
x_PM_SKY130_FD_SC_HD__NAND4BB_4%VGND N_VGND_M1031_d N_VGND_M1002_s
+ N_VGND_M1008_s N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n VGND
+ N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n N_VGND_c_984_n
+ N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n
+ PM_SKY130_FD_SC_HD__NAND4BB_4%VGND
x_PM_SKY130_FD_SC_HD__NAND4BB_4%A_432_47# N_A_432_47#_M1014_s
+ N_A_432_47#_M1019_s N_A_432_47#_M1027_s N_A_432_47#_M1025_d
+ N_A_432_47#_M1034_d N_A_432_47#_c_1079_n N_A_432_47#_c_1091_n
+ N_A_432_47#_c_1080_n PM_SKY130_FD_SC_HD__NAND4BB_4%A_432_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_4%A_850_47# N_A_850_47#_M1017_s
+ N_A_850_47#_M1028_s N_A_850_47#_M1003_s N_A_850_47#_M1032_s
+ N_A_850_47#_c_1122_n N_A_850_47#_c_1123_n N_A_850_47#_c_1124_n
+ N_A_850_47#_c_1125_n N_A_850_47#_c_1126_n N_A_850_47#_c_1127_n
+ PM_SKY130_FD_SC_HD__NAND4BB_4%A_850_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_4%A_1266_47# N_A_1266_47#_M1003_d
+ N_A_1266_47#_M1022_d N_A_1266_47#_M1033_d N_A_1266_47#_M1005_d
+ N_A_1266_47#_M1029_d N_A_1266_47#_c_1175_n
+ PM_SKY130_FD_SC_HD__NAND4BB_4%A_1266_47#
cc_1 VNB N_A_N_c_153_n 0.0219513f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A_N 0.0132315f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_155_n 0.0365137f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B_N_c_178_n 0.0192654f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_B_N_c_179_n 0.0203603f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_B_N_c_180_n 0.00435695f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_7 VNB N_A_27_47#_c_212_n 0.0199068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1019_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_9 VNB N_A_27_47#_M1010_g 4.33051e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1021_g 0.0172724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1018_g 4.49026e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_217_n 0.0577432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_M1027_g 0.016843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_M1024_g 4.13233e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_220_n 0.0147604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_221_n 0.00802475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_222_n 0.00401002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_223_n 0.0847004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_193_47#_M1017_g 0.0176655f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_20 VNB N_A_193_47#_M1000_g 4.26703e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_21 VNB N_A_193_47#_M1025_g 0.0172847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_193_47#_M1001_g 4.49956e-19 $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_23 VNB N_A_193_47#_M1028_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_193_47#_M1011_g 4.50194e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_M1034_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_M1030_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_363_n 0.00944855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_364_n 0.0132578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_c_365_n 0.00471084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_366_n 0.0693236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_C_M1003_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_32 VNB N_C_M1012_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_C_M1022_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_C_M1016_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_C_M1032_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_C_M1020_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_C_M1033_g 0.0175697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_C_M1026_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_C_c_500_n 0.0345892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_C_c_501_n 0.00736492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_C_c_502_n 0.0582445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_D_M1002_g 0.0173425f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_43 VNB N_D_M1004_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_D_M1005_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_D_M1009_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_D_M1008_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_D_M1013_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_D_M1029_g 0.0228678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB D 0.00806404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_D_c_582_n 0.0589039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_D_c_583_n 0.0270804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VPWR_c_651_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_Y_c_801_n 0.0060158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB Y 0.00255022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_977_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_56 VNB N_VGND_c_978_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_57 VNB N_VGND_c_979_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_980_n 0.014294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_981_n 0.174493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_982_n 0.011903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_983_n 0.0160664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_984_n 0.490481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_985_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_986_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_987_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_432_47#_c_1079_n 0.00160946f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.16
cc_67 VNB N_A_432_47#_c_1080_n 0.00318621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_850_47#_c_1122_n 0.00532984f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_69 VNB N_A_850_47#_c_1123_n 0.0159739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_850_47#_c_1124_n 0.00711744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_850_47#_c_1125_n 0.0043247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_850_47#_c_1126_n 0.00542244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_850_47#_c_1127_n 8.6196e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1266_47#_c_1175_n 0.0349505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VPB N_A_N_M1023_g 0.0219202f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_76 VPB A_N 0.01258f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_77 VPB N_A_N_c_155_n 0.0102044f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_78 VPB N_B_N_M1006_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_79 VPB N_B_N_c_179_n 0.00459527f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_80 VPB N_B_N_c_180_n 0.00268628f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_81 VPB N_A_27_47#_M1007_g 0.0231885f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_82 VPB N_A_27_47#_M1010_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_M1018_g 0.019153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_217_n 6.59428e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_M1024_g 0.0186547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_229_n 0.0180063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_230_n 0.00912537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_222_n 0.0025799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_47#_c_223_n 0.0499399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_193_47#_M1000_g 0.0194271f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_91 VPB N_A_193_47#_M1001_g 0.0191804f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_92 VPB N_A_193_47#_M1011_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_193_47#_M1030_g 0.026721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_193_47#_c_371_n 0.0157519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_193_47#_c_372_n 0.0207544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_193_47#_c_373_n 0.0018142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_C_M1012_g 0.026721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_C_M1016_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_C_M1020_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_C_M1026_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_D_M1004_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_D_M1009_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_D_M1013_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_D_M1035_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_D_c_583_n 0.00847707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_652_n 0.00230843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_653_n 0.00407299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_654_n 0.0152056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_655_n 0.00171127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_656_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_657_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_658_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_659_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_660_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_661_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_662_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_663_n 0.0101727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_664_n 0.0467131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_665_n 0.0367988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_666_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_667_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_668_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_669_n 0.0189004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_670_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_671_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_672_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_673_n 0.0151232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_674_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_675_n 0.00320131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_676_n 0.00353672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_677_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_678_n 0.0195368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_679_n 0.0268977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_680_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_651_n 0.0621474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_Y_c_803_n 0.00227512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_Y_c_804_n 0.00151697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_Y_c_805_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_Y_c_806_n 0.0137645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_Y_c_807_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_Y_c_808_n 0.00408948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_Y_c_809_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_Y_c_810_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_Y_c_811_n 0.00125718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_Y_c_812_n 0.00181104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_Y_c_813_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_Y_c_814_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_Y_c_815_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_Y_c_816_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB Y 0.00183954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB Y 0.00272159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 N_A_N_c_153_n N_B_N_c_178_n 0.0263225f $X=0.47 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_N_M1023_g N_B_N_M1006_g 0.0449216f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_154 A_N N_B_N_c_179_n 2.39636e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_N_c_155_n N_B_N_c_179_n 0.0207686f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_156 A_N N_B_N_c_180_n 0.0321142f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A_N_c_155_n N_B_N_c_180_n 0.00505751f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_158 A_N N_A_27_47#_M1023_s 0.00453106f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A_N_c_153_n N_A_27_47#_c_234_n 0.0170415f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_160 A_N N_A_27_47#_c_221_n 0.0179334f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A_N_c_155_n N_A_27_47#_c_221_n 0.00222211f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_N_M1023_g N_A_27_47#_c_237_n 0.0192935f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_163 A_N N_A_27_47#_c_230_n 0.0204787f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A_N_c_155_n N_A_27_47#_c_230_n 0.00170498f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_N_M1023_g N_VPWR_c_652_n 0.00768947f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_N_M1023_g N_VPWR_c_673_n 0.00424408f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_N_M1023_g N_VPWR_c_651_n 0.00594309f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_N_c_153_n N_VGND_c_977_n 0.00831359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_N_c_153_n N_VGND_c_980_n 0.00339367f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_N_c_153_n N_VGND_c_984_n 0.00497794f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B_N_c_178_n N_A_27_47#_c_234_n 0.0133477f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B_N_c_179_n N_A_27_47#_c_234_n 0.00134087f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B_N_c_180_n N_A_27_47#_c_234_n 0.0251978f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_N_M1006_g N_A_27_47#_c_237_n 0.0147951f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B_N_c_179_n N_A_27_47#_c_237_n 9.50548e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B_N_c_180_n N_A_27_47#_c_237_n 0.024162f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B_N_c_178_n N_A_27_47#_c_222_n 0.00688199f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B_N_M1006_g N_A_27_47#_c_222_n 0.00827402f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_179 N_B_N_c_179_n N_A_27_47#_c_222_n 0.00199269f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B_N_c_180_n N_A_27_47#_c_222_n 0.0448178f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B_N_c_179_n N_A_27_47#_c_223_n 0.0202849f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B_N_c_180_n N_A_27_47#_c_223_n 3.14223e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B_N_M1006_g N_A_193_47#_c_371_n 0.00428252f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_B_N_c_178_n N_A_193_47#_c_364_n 0.00414979f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_B_N_M1006_g N_A_193_47#_c_372_n 0.00404608f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_B_N_c_180_n N_VPWR_M1023_d 0.00191019f $X=0.89 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_187 N_B_N_M1006_g N_VPWR_c_652_n 0.00276606f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B_N_M1006_g N_VPWR_c_665_n 0.00423478f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B_N_M1006_g N_VPWR_c_651_n 0.00710834f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B_N_c_178_n N_VGND_c_977_n 0.00833262f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B_N_c_178_n N_VGND_c_981_n 0.00339367f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B_N_c_178_n N_VGND_c_984_n 0.00536411f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_234_n N_A_193_47#_M1015_d 0.0139018f $X=1.145 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_194 N_A_27_47#_c_222_n N_A_193_47#_M1015_d 0.00200292f $X=1.37 $Y=1.16
+ $X2=-0.19 $Y2=-0.24
cc_195 N_A_27_47#_c_237_n N_A_193_47#_M1006_d 0.0147415f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_222_n N_A_193_47#_M1006_d 0.0112361f $X=1.37 $Y=1.16 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_M1027_g N_A_193_47#_M1017_g 0.0227611f $X=3.755 $Y=0.56 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_M1024_g N_A_193_47#_M1000_g 0.0227611f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_237_n N_A_193_47#_c_371_n 0.0364045f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_212_n N_A_193_47#_c_363_n 0.00102052f $X=2.495 $Y=0.995
+ $X2=0 $Y2=0
cc_201 N_A_27_47#_c_234_n N_A_193_47#_c_363_n 0.0327695f $X=1.145 $Y=0.72 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_223_n N_A_193_47#_c_363_n 0.00521991f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_212_n N_A_193_47#_c_364_n 0.00290407f $X=2.495 $Y=0.995
+ $X2=0 $Y2=0
cc_204 N_A_27_47#_c_234_n N_A_193_47#_c_364_n 0.0140572f $X=1.145 $Y=0.72 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_222_n N_A_193_47#_c_364_n 0.0204797f $X=1.37 $Y=1.16 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_223_n N_A_193_47#_c_364_n 0.00992468f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1007_g N_A_193_47#_c_372_n 0.00492478f $X=2.495 $Y=1.985
+ $X2=0 $Y2=0
cc_208 N_A_27_47#_c_237_n N_A_193_47#_c_372_n 0.0161245f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_222_n N_A_193_47#_c_372_n 0.0371854f $X=1.37 $Y=1.16 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_223_n N_A_193_47#_c_372_n 0.00552719f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_222_n N_A_193_47#_c_395_n 0.0173866f $X=1.37 $Y=1.16 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_223_n N_A_193_47#_c_395_n 0.00685844f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_217_n N_A_193_47#_c_365_n 0.0253382f $X=3.755 $Y=1.025 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_273_p N_A_193_47#_c_365_n 0.0247935f $X=3.12 $Y=1.16 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_223_n N_A_193_47#_c_365_n 0.00685773f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_222_n N_A_193_47#_c_400_n 8.60994e-19 $X=1.37 $Y=1.16 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_273_p N_A_193_47#_c_400_n 3.24364e-19 $X=3.12 $Y=1.16 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_223_n N_A_193_47#_c_400_n 0.0230996f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_273_p N_A_193_47#_c_403_n 0.00515123f $X=3.12 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_223_n N_A_193_47#_c_403_n 0.0321282f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_217_n N_A_193_47#_c_405_n 2.42253e-19 $X=3.755 $Y=1.025
+ $X2=0 $Y2=0
cc_222 N_A_27_47#_c_217_n N_A_193_47#_c_366_n 0.0227611f $X=3.755 $Y=1.025 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_237_n N_VPWR_M1023_d 0.00343054f $X=1.145 $Y=1.882 $X2=-0.19
+ $Y2=-0.24
cc_224 N_A_27_47#_c_237_n N_VPWR_c_652_n 0.0102755f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_M1007_g N_VPWR_c_653_n 0.0030732f $X=2.495 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_223_n N_VPWR_c_653_n 0.00480739f $X=2.42 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1007_g N_VPWR_c_654_n 0.00541359f $X=2.495 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1010_g N_VPWR_c_654_n 0.0046653f $X=2.915 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1007_g N_VPWR_c_655_n 7.17238e-19 $X=2.495 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_M1010_g N_VPWR_c_655_n 0.0108439f $X=2.915 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1018_g N_VPWR_c_655_n 0.00151363f $X=3.335 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1018_g N_VPWR_c_656_n 0.00541359f $X=3.335 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_M1024_g N_VPWR_c_656_n 0.00541359f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_M1024_g N_VPWR_c_657_n 0.00146448f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_237_n N_VPWR_c_665_n 0.00193599f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_229_n N_VPWR_c_673_n 0.0162479f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_237_n N_VPWR_c_673_n 0.00207649f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1023_s N_VPWR_c_651_n 0.00223307f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1007_g N_VPWR_c_651_n 0.0108276f $X=2.495 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1010_g N_VPWR_c_651_n 0.00789179f $X=2.915 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1018_g N_VPWR_c_651_n 0.00950154f $X=3.335 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1024_g N_VPWR_c_651_n 0.00952874f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_229_n N_VPWR_c_651_n 0.0107554f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_237_n N_VPWR_c_651_n 0.00886241f $X=1.145 $Y=1.882 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_212_n N_Y_c_801_n 0.00375135f $X=2.495 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_27_47#_M1019_g N_Y_c_801_n 0.0106345f $X=2.915 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1021_g N_Y_c_801_n 0.0118097f $X=3.335 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_217_n N_Y_c_801_n 0.0066355f $X=3.755 $Y=1.025 $X2=0 $Y2=0
cc_249 N_A_27_47#_M1027_g N_Y_c_801_n 0.00131391f $X=3.755 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_273_p N_Y_c_801_n 0.0492056f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_27_47#_M1007_g N_Y_c_825_n 0.0101262f $X=2.495 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1010_g N_Y_c_803_n 0.0152992f $X=2.915 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1018_g N_Y_c_803_n 0.0128842f $X=3.335 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_217_n N_Y_c_803_n 0.00203016f $X=3.755 $Y=1.025 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_273_p N_Y_c_803_n 0.0260603f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_27_47#_M1007_g N_Y_c_804_n 0.00639641f $X=2.495 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_217_n N_Y_c_804_n 0.00211055f $X=3.755 $Y=1.025 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_273_p N_Y_c_804_n 0.014659f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1010_g N_Y_c_833_n 4.51827e-19 $X=2.915 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_27_47#_M1018_g N_Y_c_833_n 0.0100737f $X=3.335 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A_27_47#_M1024_g N_Y_c_833_n 0.00985674f $X=3.755 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_27_47#_M1024_g N_Y_c_836_n 6.1949e-19 $X=3.755 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_27_47#_M1021_g Y 7.17425e-19 $X=3.335 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A_27_47#_M1018_g Y 9.02652e-19 $X=3.335 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_217_n Y 0.0126701f $X=3.755 $Y=1.025 $X2=0 $Y2=0
cc_266 N_A_27_47#_M1027_g Y 0.00393648f $X=3.755 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A_27_47#_M1024_g Y 0.00537732f $X=3.755 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_273_p Y 0.00436144f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1018_g Y 0.00180817f $X=3.335 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_217_n Y 0.0023737f $X=3.755 $Y=1.025 $X2=0 $Y2=0
cc_271 N_A_27_47#_M1024_g Y 0.0124238f $X=3.755 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_27_47#_M1027_g N_Y_c_846_n 0.00676775f $X=3.755 $Y=0.56 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_234_n N_VGND_M1031_d 0.00330044f $X=1.145 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_274 N_A_27_47#_c_234_n N_VGND_c_977_n 0.0159625f $X=1.145 $Y=0.72 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_220_n N_VGND_c_980_n 0.0177262f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_234_n N_VGND_c_980_n 0.00243651f $X=1.145 $Y=0.72 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_212_n N_VGND_c_981_n 0.00357877f $X=2.495 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1019_g N_VGND_c_981_n 0.00357877f $X=2.915 $Y=0.56 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1021_g N_VGND_c_981_n 0.00357877f $X=3.335 $Y=0.56 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1027_g N_VGND_c_981_n 0.00357877f $X=3.755 $Y=0.56 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_234_n N_VGND_c_981_n 0.00244309f $X=1.145 $Y=0.72 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1031_s N_VGND_c_984_n 0.0022756f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_212_n N_VGND_c_984_n 0.00664112f $X=2.495 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_M1019_g N_VGND_c_984_n 0.00522516f $X=2.915 $Y=0.56 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1021_g N_VGND_c_984_n 0.00522516f $X=3.335 $Y=0.56 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1027_g N_VGND_c_984_n 0.00525237f $X=3.755 $Y=0.56 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_220_n N_VGND_c_984_n 0.00988152f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_234_n N_VGND_c_984_n 0.0101727f $X=1.145 $Y=0.72 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_212_n N_A_432_47#_c_1079_n 0.0016109f $X=2.495 $Y=0.995
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_223_n N_A_432_47#_c_1079_n 0.00536536f $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_212_n N_A_432_47#_c_1080_n 0.0173415f $X=2.495 $Y=0.995
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_M1019_g N_A_432_47#_c_1080_n 0.00912735f $X=2.915 $Y=0.56
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_M1021_g N_A_432_47#_c_1080_n 0.00918728f $X=3.335 $Y=0.56
+ $X2=0 $Y2=0
cc_294 N_A_27_47#_M1027_g N_A_432_47#_c_1080_n 0.00918189f $X=3.755 $Y=0.56
+ $X2=0 $Y2=0
cc_295 N_A_27_47#_M1027_g N_A_850_47#_c_1122_n 2.08102e-19 $X=3.755 $Y=0.56
+ $X2=0 $Y2=0
cc_296 N_A_193_47#_c_366_n N_C_c_501_n 0.00606999f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_193_47#_c_371_n N_VPWR_c_653_n 0.014096f $X=1.625 $Y=2.307 $X2=0
+ $Y2=0
cc_298 N_A_193_47#_c_372_n N_VPWR_c_653_n 0.0260714f $X=1.71 $Y=2.15 $X2=0 $Y2=0
cc_299 N_A_193_47#_c_365_n N_VPWR_c_653_n 0.00433199f $X=4.22 $Y=1.19 $X2=0
+ $Y2=0
cc_300 N_A_193_47#_c_400_n N_VPWR_c_653_n 2.19293e-19 $X=2.21 $Y=1.19 $X2=0
+ $Y2=0
cc_301 N_A_193_47#_c_403_n N_VPWR_c_653_n 5.51824e-19 $X=2.065 $Y=1.19 $X2=0
+ $Y2=0
cc_302 N_A_193_47#_M1000_g N_VPWR_c_657_n 0.00146448f $X=4.175 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_193_47#_M1001_g N_VPWR_c_658_n 0.00146448f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A_193_47#_M1011_g N_VPWR_c_658_n 0.00268723f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_A_193_47#_c_371_n N_VPWR_c_665_n 0.0561203f $X=1.625 $Y=2.307 $X2=0
+ $Y2=0
cc_306 N_A_193_47#_M1000_g N_VPWR_c_667_n 0.00541359f $X=4.175 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_A_193_47#_M1001_g N_VPWR_c_667_n 0.00541359f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_308 N_A_193_47#_M1011_g N_VPWR_c_678_n 0.00541359f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_193_47#_M1030_g N_VPWR_c_678_n 0.00541359f $X=5.435 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_193_47#_M1030_g N_VPWR_c_679_n 0.00766777f $X=5.435 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_193_47#_M1006_d N_VPWR_c_651_n 0.00402019f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_312 N_A_193_47#_M1000_g N_VPWR_c_651_n 0.00948268f $X=4.175 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_193_47#_M1001_g N_VPWR_c_651_n 0.00950154f $X=4.595 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_193_47#_M1011_g N_VPWR_c_651_n 0.00950154f $X=5.015 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_193_47#_M1030_g N_VPWR_c_651_n 0.0109504f $X=5.435 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_193_47#_c_371_n N_VPWR_c_651_n 0.0323886f $X=1.625 $Y=2.307 $X2=0
+ $Y2=0
cc_317 N_A_193_47#_c_365_n N_Y_c_801_n 0.0156539f $X=4.22 $Y=1.19 $X2=0 $Y2=0
cc_318 N_A_193_47#_c_365_n N_Y_c_803_n 0.0215176f $X=4.22 $Y=1.19 $X2=0 $Y2=0
cc_319 N_A_193_47#_c_365_n N_Y_c_804_n 0.00564095f $X=4.22 $Y=1.19 $X2=0 $Y2=0
cc_320 N_A_193_47#_M1000_g N_Y_c_833_n 6.20279e-19 $X=4.175 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A_193_47#_M1000_g N_Y_c_836_n 0.00975139f $X=4.175 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_193_47#_M1001_g N_Y_c_836_n 0.00975139f $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_193_47#_M1011_g N_Y_c_836_n 6.1949e-19 $X=5.015 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A_193_47#_M1001_g N_Y_c_805_n 0.0120357f $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A_193_47#_M1011_g N_Y_c_805_n 0.0120357f $X=5.015 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_193_47#_c_405_n N_Y_c_805_n 0.0366837f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_193_47#_c_366_n N_Y_c_805_n 0.0019951f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_193_47#_M1001_g N_Y_c_858_n 6.1949e-19 $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_193_47#_M1011_g N_Y_c_858_n 0.00975139f $X=5.015 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A_193_47#_M1030_g N_Y_c_858_n 0.015395f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A_193_47#_M1030_g N_Y_c_806_n 0.0162259f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_193_47#_M1000_g N_Y_c_811_n 0.0120977f $X=4.175 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A_193_47#_c_365_n N_Y_c_811_n 0.0077781f $X=4.22 $Y=1.19 $X2=0 $Y2=0
cc_334 N_A_193_47#_c_405_n N_Y_c_811_n 0.00378334f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_193_47#_M1000_g N_Y_c_812_n 0.00147213f $X=4.175 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_193_47#_M1001_g N_Y_c_812_n 0.00149073f $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_193_47#_c_373_n N_Y_c_812_n 0.00839518f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_338 N_A_193_47#_c_405_n N_Y_c_812_n 0.0233462f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A_193_47#_c_366_n N_Y_c_812_n 0.00163629f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_193_47#_M1011_g N_Y_c_813_n 0.00149073f $X=5.015 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A_193_47#_M1030_g N_Y_c_813_n 0.00149073f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_193_47#_c_405_n N_Y_c_813_n 0.026643f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_193_47#_c_366_n N_Y_c_813_n 0.00206439f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A_193_47#_M1017_g Y 0.00976611f $X=4.175 $Y=0.56 $X2=0 $Y2=0
cc_345 N_A_193_47#_c_365_n Y 0.0260409f $X=4.22 $Y=1.19 $X2=0 $Y2=0
cc_346 N_A_193_47#_c_373_n Y 0.00174845f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_347 N_A_193_47#_c_405_n Y 0.0141073f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A_193_47#_c_365_n Y 0.00134533f $X=4.22 $Y=1.19 $X2=0 $Y2=0
cc_349 N_A_193_47#_M1017_g N_Y_c_846_n 0.00208455f $X=4.175 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A_193_47#_M1017_g N_VGND_c_981_n 0.00357877f $X=4.175 $Y=0.56 $X2=0
+ $Y2=0
cc_351 N_A_193_47#_M1025_g N_VGND_c_981_n 0.00357877f $X=4.595 $Y=0.56 $X2=0
+ $Y2=0
cc_352 N_A_193_47#_M1028_g N_VGND_c_981_n 0.00357877f $X=5.015 $Y=0.56 $X2=0
+ $Y2=0
cc_353 N_A_193_47#_M1034_g N_VGND_c_981_n 0.00357877f $X=5.435 $Y=0.56 $X2=0
+ $Y2=0
cc_354 N_A_193_47#_c_363_n N_VGND_c_981_n 0.0513547f $X=1.625 $Y=0.36 $X2=0
+ $Y2=0
cc_355 N_A_193_47#_M1015_d N_VGND_c_984_n 0.00421059f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_193_47#_M1017_g N_VGND_c_984_n 0.00525237f $X=4.175 $Y=0.56 $X2=0
+ $Y2=0
cc_357 N_A_193_47#_M1025_g N_VGND_c_984_n 0.00522516f $X=4.595 $Y=0.56 $X2=0
+ $Y2=0
cc_358 N_A_193_47#_M1028_g N_VGND_c_984_n 0.00522516f $X=5.015 $Y=0.56 $X2=0
+ $Y2=0
cc_359 N_A_193_47#_M1034_g N_VGND_c_984_n 0.00655123f $X=5.435 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_193_47#_c_363_n N_VGND_c_984_n 0.0293659f $X=1.625 $Y=0.36 $X2=0
+ $Y2=0
cc_361 N_A_193_47#_c_364_n N_A_432_47#_c_1079_n 0.0167417f $X=1.71 $Y=1.075
+ $X2=0 $Y2=0
cc_362 N_A_193_47#_c_365_n N_A_432_47#_c_1079_n 0.00443762f $X=4.22 $Y=1.19
+ $X2=0 $Y2=0
cc_363 N_A_193_47#_c_400_n N_A_432_47#_c_1079_n 2.20995e-19 $X=2.21 $Y=1.19
+ $X2=0 $Y2=0
cc_364 N_A_193_47#_c_403_n N_A_432_47#_c_1079_n 6.33188e-19 $X=2.065 $Y=1.19
+ $X2=0 $Y2=0
cc_365 N_A_193_47#_c_363_n N_A_432_47#_c_1091_n 0.010345f $X=1.625 $Y=0.36 $X2=0
+ $Y2=0
cc_366 N_A_193_47#_c_364_n N_A_432_47#_c_1091_n 8.65915e-19 $X=1.71 $Y=1.075
+ $X2=0 $Y2=0
cc_367 N_A_193_47#_M1017_g N_A_432_47#_c_1080_n 0.0118842f $X=4.175 $Y=0.56
+ $X2=0 $Y2=0
cc_368 N_A_193_47#_M1025_g N_A_432_47#_c_1080_n 0.00918728f $X=4.595 $Y=0.56
+ $X2=0 $Y2=0
cc_369 N_A_193_47#_M1028_g N_A_432_47#_c_1080_n 0.00918728f $X=5.015 $Y=0.56
+ $X2=0 $Y2=0
cc_370 N_A_193_47#_M1034_g N_A_432_47#_c_1080_n 0.00956495f $X=5.435 $Y=0.56
+ $X2=0 $Y2=0
cc_371 N_A_193_47#_c_405_n N_A_432_47#_c_1080_n 0.00150843f $X=5.225 $Y=1.16
+ $X2=0 $Y2=0
cc_372 N_A_193_47#_M1017_g N_A_850_47#_c_1122_n 0.00394364f $X=4.175 $Y=0.56
+ $X2=0 $Y2=0
cc_373 N_A_193_47#_M1025_g N_A_850_47#_c_1122_n 0.0107009f $X=4.595 $Y=0.56
+ $X2=0 $Y2=0
cc_374 N_A_193_47#_M1028_g N_A_850_47#_c_1122_n 0.0107009f $X=5.015 $Y=0.56
+ $X2=0 $Y2=0
cc_375 N_A_193_47#_c_373_n N_A_850_47#_c_1122_n 0.00691468f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_376 N_A_193_47#_c_405_n N_A_850_47#_c_1122_n 0.0830678f $X=5.225 $Y=1.16
+ $X2=0 $Y2=0
cc_377 N_A_193_47#_c_366_n N_A_850_47#_c_1122_n 0.00622116f $X=5.435 $Y=1.16
+ $X2=0 $Y2=0
cc_378 N_A_193_47#_M1034_g N_A_850_47#_c_1123_n 0.0108866f $X=5.435 $Y=0.56
+ $X2=0 $Y2=0
cc_379 N_A_193_47#_M1034_g N_A_850_47#_c_1124_n 0.00417358f $X=5.435 $Y=0.56
+ $X2=0 $Y2=0
cc_380 N_A_193_47#_M1034_g N_A_850_47#_c_1127_n 0.00315977f $X=5.435 $Y=0.56
+ $X2=0 $Y2=0
cc_381 N_C_M1033_g N_D_M1002_g 0.0246921f $X=7.955 $Y=0.56 $X2=0 $Y2=0
cc_382 N_C_M1026_g N_D_M1004_g 0.0246921f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_383 N_C_c_501_n D 0.00679138f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_384 N_C_c_502_n D 7.61915e-19 $X=7.955 $Y=1.16 $X2=0 $Y2=0
cc_385 N_C_c_501_n N_D_c_582_n 7.61915e-19 $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_386 N_C_c_502_n N_D_c_582_n 0.0246921f $X=7.955 $Y=1.16 $X2=0 $Y2=0
cc_387 N_C_M1016_g N_VPWR_c_659_n 0.00268723f $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_388 N_C_M1020_g N_VPWR_c_659_n 0.00146448f $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_389 N_C_M1026_g N_VPWR_c_660_n 0.00146448f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_390 N_C_M1012_g N_VPWR_c_669_n 0.00541359f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_391 N_C_M1016_g N_VPWR_c_669_n 0.00541359f $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_392 N_C_M1020_g N_VPWR_c_671_n 0.00541359f $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_393 N_C_M1026_g N_VPWR_c_671_n 0.00541359f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_394 N_C_M1012_g N_VPWR_c_679_n 0.00771316f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_395 N_C_M1012_g N_VPWR_c_651_n 0.0109004f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_396 N_C_M1016_g N_VPWR_c_651_n 0.00950154f $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_397 N_C_M1020_g N_VPWR_c_651_n 0.00950154f $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_398 N_C_M1026_g N_VPWR_c_651_n 0.00952874f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_399 N_C_M1012_g N_Y_c_806_n 0.0147646f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_400 N_C_c_500_n N_Y_c_806_n 0.00729564f $X=6.62 $Y=1.16 $X2=0 $Y2=0
cc_401 N_C_c_501_n N_Y_c_806_n 0.0459297f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_402 N_C_M1012_g N_Y_c_883_n 0.0150661f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_403 N_C_M1016_g N_Y_c_883_n 0.00975139f $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_404 N_C_M1020_g N_Y_c_883_n 6.1949e-19 $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_405 N_C_M1016_g N_Y_c_807_n 0.0120357f $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_406 N_C_M1020_g N_Y_c_807_n 0.0120357f $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_407 N_C_c_501_n N_Y_c_807_n 0.0366837f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_408 N_C_c_502_n N_Y_c_807_n 0.0019951f $X=7.955 $Y=1.16 $X2=0 $Y2=0
cc_409 N_C_M1016_g N_Y_c_890_n 6.1949e-19 $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_410 N_C_M1020_g N_Y_c_890_n 0.00975139f $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_411 N_C_M1026_g N_Y_c_890_n 0.00975139f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_412 N_C_M1026_g N_Y_c_808_n 0.0134397f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_413 N_C_M1026_g N_Y_c_894_n 6.1949e-19 $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_414 N_C_M1012_g N_Y_c_814_n 0.00149073f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_415 N_C_M1016_g N_Y_c_814_n 0.00149073f $X=7.115 $Y=1.985 $X2=0 $Y2=0
cc_416 N_C_c_501_n N_Y_c_814_n 0.026643f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_417 N_C_c_502_n N_Y_c_814_n 0.00206439f $X=7.955 $Y=1.16 $X2=0 $Y2=0
cc_418 N_C_M1020_g N_Y_c_815_n 0.00149073f $X=7.535 $Y=1.985 $X2=0 $Y2=0
cc_419 N_C_M1026_g N_Y_c_815_n 0.00149073f $X=7.955 $Y=1.985 $X2=0 $Y2=0
cc_420 N_C_c_501_n N_Y_c_815_n 0.026643f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_421 N_C_c_502_n N_Y_c_815_n 0.00206439f $X=7.955 $Y=1.16 $X2=0 $Y2=0
cc_422 N_C_M1033_g N_VGND_c_978_n 0.0018181f $X=7.955 $Y=0.56 $X2=0 $Y2=0
cc_423 N_C_M1003_g N_VGND_c_981_n 0.00357877f $X=6.695 $Y=0.56 $X2=0 $Y2=0
cc_424 N_C_M1022_g N_VGND_c_981_n 0.00357877f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_425 N_C_M1032_g N_VGND_c_981_n 0.00357877f $X=7.535 $Y=0.56 $X2=0 $Y2=0
cc_426 N_C_M1033_g N_VGND_c_981_n 0.00413993f $X=7.955 $Y=0.56 $X2=0 $Y2=0
cc_427 N_C_M1003_g N_VGND_c_984_n 0.00660224f $X=6.695 $Y=0.56 $X2=0 $Y2=0
cc_428 N_C_M1022_g N_VGND_c_984_n 0.00522516f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_429 N_C_M1032_g N_VGND_c_984_n 0.00522516f $X=7.535 $Y=0.56 $X2=0 $Y2=0
cc_430 N_C_M1033_g N_VGND_c_984_n 0.00578258f $X=7.955 $Y=0.56 $X2=0 $Y2=0
cc_431 N_C_M1003_g N_A_850_47#_c_1123_n 3.39797e-19 $X=6.695 $Y=0.56 $X2=0 $Y2=0
cc_432 N_C_c_501_n N_A_850_47#_c_1123_n 0.00255272f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_433 N_C_M1003_g N_A_850_47#_c_1124_n 0.00288969f $X=6.695 $Y=0.56 $X2=0 $Y2=0
cc_434 N_C_M1003_g N_A_850_47#_c_1126_n 0.0119076f $X=6.695 $Y=0.56 $X2=0 $Y2=0
cc_435 N_C_M1022_g N_A_850_47#_c_1126_n 0.00918728f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_436 N_C_M1032_g N_A_850_47#_c_1126_n 0.00918728f $X=7.535 $Y=0.56 $X2=0 $Y2=0
cc_437 N_C_M1033_g N_A_850_47#_c_1126_n 0.00463137f $X=7.955 $Y=0.56 $X2=0 $Y2=0
cc_438 N_C_c_500_n N_A_850_47#_c_1126_n 7.93922e-19 $X=6.62 $Y=1.16 $X2=0 $Y2=0
cc_439 N_C_c_501_n N_A_850_47#_c_1126_n 0.00545452f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_440 N_C_M1003_g N_A_1266_47#_c_1175_n 0.0108548f $X=6.695 $Y=0.56 $X2=0 $Y2=0
cc_441 N_C_M1022_g N_A_1266_47#_c_1175_n 0.0107009f $X=7.115 $Y=0.56 $X2=0 $Y2=0
cc_442 N_C_M1032_g N_A_1266_47#_c_1175_n 0.0107009f $X=7.535 $Y=0.56 $X2=0 $Y2=0
cc_443 N_C_M1033_g N_A_1266_47#_c_1175_n 0.0133309f $X=7.955 $Y=0.56 $X2=0 $Y2=0
cc_444 N_C_c_500_n N_A_1266_47#_c_1175_n 0.00689495f $X=6.62 $Y=1.16 $X2=0 $Y2=0
cc_445 N_C_c_501_n N_A_1266_47#_c_1175_n 0.116775f $X=7.745 $Y=1.16 $X2=0 $Y2=0
cc_446 N_C_c_502_n N_A_1266_47#_c_1175_n 0.00622382f $X=7.955 $Y=1.16 $X2=0
+ $Y2=0
cc_447 N_D_M1004_g N_VPWR_c_660_n 0.00146448f $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_448 N_D_M1004_g N_VPWR_c_661_n 0.00541359f $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_449 N_D_M1009_g N_VPWR_c_661_n 0.00541359f $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_450 N_D_M1009_g N_VPWR_c_662_n 0.00146448f $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_451 N_D_M1013_g N_VPWR_c_662_n 0.00146448f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_452 N_D_M1035_g N_VPWR_c_664_n 0.0041173f $X=9.635 $Y=1.985 $X2=0 $Y2=0
cc_453 D N_VPWR_c_664_n 0.0207117f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_454 N_D_c_583_n N_VPWR_c_664_n 0.00598079f $X=9.845 $Y=1.16 $X2=0 $Y2=0
cc_455 N_D_M1013_g N_VPWR_c_674_n 0.00541359f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_456 N_D_M1035_g N_VPWR_c_674_n 0.00541359f $X=9.635 $Y=1.985 $X2=0 $Y2=0
cc_457 N_D_M1004_g N_VPWR_c_651_n 0.00952874f $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_458 N_D_M1009_g N_VPWR_c_651_n 0.00950154f $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_459 N_D_M1013_g N_VPWR_c_651_n 0.00950154f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_460 N_D_M1035_g N_VPWR_c_651_n 0.0104699f $X=9.635 $Y=1.985 $X2=0 $Y2=0
cc_461 N_D_M1004_g N_Y_c_890_n 6.1949e-19 $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_462 N_D_M1004_g N_Y_c_808_n 0.0134397f $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_463 N_D_M1004_g N_Y_c_894_n 0.00975139f $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_464 N_D_M1009_g N_Y_c_894_n 0.00975139f $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_465 N_D_M1013_g N_Y_c_894_n 6.1949e-19 $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_466 N_D_M1009_g N_Y_c_809_n 0.0120357f $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_467 N_D_M1013_g N_Y_c_809_n 0.0120357f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_468 D N_Y_c_809_n 0.0366837f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_469 N_D_c_582_n N_Y_c_809_n 0.0019951f $X=9.71 $Y=1.16 $X2=0 $Y2=0
cc_470 N_D_M1013_g N_Y_c_810_n 0.00149073f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_471 N_D_M1035_g N_Y_c_810_n 0.00331821f $X=9.635 $Y=1.985 $X2=0 $Y2=0
cc_472 D N_Y_c_810_n 0.026643f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_473 N_D_c_582_n N_Y_c_810_n 0.00206439f $X=9.71 $Y=1.16 $X2=0 $Y2=0
cc_474 N_D_M1009_g N_Y_c_916_n 6.1949e-19 $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_475 N_D_M1013_g N_Y_c_916_n 0.00975139f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_476 N_D_M1035_g N_Y_c_916_n 0.00902485f $X=9.635 $Y=1.985 $X2=0 $Y2=0
cc_477 N_D_M1004_g N_Y_c_816_n 0.00149073f $X=8.375 $Y=1.985 $X2=0 $Y2=0
cc_478 N_D_M1009_g N_Y_c_816_n 0.00149073f $X=8.795 $Y=1.985 $X2=0 $Y2=0
cc_479 D N_Y_c_816_n 0.026643f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_480 N_D_c_582_n N_Y_c_816_n 0.00206439f $X=9.71 $Y=1.16 $X2=0 $Y2=0
cc_481 N_D_M1002_g N_VGND_c_978_n 0.00964559f $X=8.375 $Y=0.56 $X2=0 $Y2=0
cc_482 N_D_M1005_g N_VGND_c_978_n 0.00845732f $X=8.795 $Y=0.56 $X2=0 $Y2=0
cc_483 N_D_M1008_g N_VGND_c_978_n 0.00116151f $X=9.215 $Y=0.56 $X2=0 $Y2=0
cc_484 N_D_M1005_g N_VGND_c_979_n 0.00116151f $X=8.795 $Y=0.56 $X2=0 $Y2=0
cc_485 N_D_M1008_g N_VGND_c_979_n 0.00845732f $X=9.215 $Y=0.56 $X2=0 $Y2=0
cc_486 N_D_M1029_g N_VGND_c_979_n 0.0161007f $X=9.635 $Y=0.56 $X2=0 $Y2=0
cc_487 N_D_M1002_g N_VGND_c_981_n 0.00341689f $X=8.375 $Y=0.56 $X2=0 $Y2=0
cc_488 N_D_M1005_g N_VGND_c_982_n 0.00341689f $X=8.795 $Y=0.56 $X2=0 $Y2=0
cc_489 N_D_M1008_g N_VGND_c_982_n 0.00341689f $X=9.215 $Y=0.56 $X2=0 $Y2=0
cc_490 N_D_M1029_g N_VGND_c_983_n 0.00341689f $X=9.635 $Y=0.56 $X2=0 $Y2=0
cc_491 N_D_M1002_g N_VGND_c_984_n 0.00405445f $X=8.375 $Y=0.56 $X2=0 $Y2=0
cc_492 N_D_M1005_g N_VGND_c_984_n 0.0040262f $X=8.795 $Y=0.56 $X2=0 $Y2=0
cc_493 N_D_M1008_g N_VGND_c_984_n 0.0040262f $X=9.215 $Y=0.56 $X2=0 $Y2=0
cc_494 N_D_M1029_g N_VGND_c_984_n 0.00503176f $X=9.635 $Y=0.56 $X2=0 $Y2=0
cc_495 N_D_M1002_g N_A_850_47#_c_1126_n 6.66764e-19 $X=8.375 $Y=0.56 $X2=0 $Y2=0
cc_496 N_D_M1002_g N_A_1266_47#_c_1175_n 0.013302f $X=8.375 $Y=0.56 $X2=0 $Y2=0
cc_497 N_D_M1005_g N_A_1266_47#_c_1175_n 0.0118239f $X=8.795 $Y=0.56 $X2=0 $Y2=0
cc_498 N_D_M1008_g N_A_1266_47#_c_1175_n 0.0118239f $X=9.215 $Y=0.56 $X2=0 $Y2=0
cc_499 N_D_M1029_g N_A_1266_47#_c_1175_n 0.0119846f $X=9.635 $Y=0.56 $X2=0 $Y2=0
cc_500 D N_A_1266_47#_c_1175_n 0.117148f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_501 N_D_c_582_n N_A_1266_47#_c_1175_n 0.00622382f $X=9.71 $Y=1.16 $X2=0 $Y2=0
cc_502 N_D_c_583_n N_A_1266_47#_c_1175_n 0.00719798f $X=9.845 $Y=1.16 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_651_n N_Y_M1007_s 0.0038878f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_504 N_VPWR_c_651_n N_Y_M1018_s 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_505 N_VPWR_c_651_n N_Y_M1000_s 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_506 N_VPWR_c_651_n N_Y_M1011_s 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_507 N_VPWR_c_651_n N_Y_M1012_s 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_508 N_VPWR_c_651_n N_Y_M1020_s 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_509 N_VPWR_c_651_n N_Y_M1004_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_510 N_VPWR_c_651_n N_Y_M1013_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_511 N_VPWR_c_654_n N_Y_c_825_n 0.0151499f $X=2.96 $Y=2.72 $X2=0 $Y2=0
cc_512 N_VPWR_c_651_n N_Y_c_825_n 0.00934584f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_513 N_VPWR_M1010_d N_Y_c_803_n 0.00167154f $X=2.99 $Y=1.485 $X2=0 $Y2=0
cc_514 N_VPWR_c_655_n N_Y_c_803_n 0.01469f $X=3.125 $Y=2 $X2=0 $Y2=0
cc_515 N_VPWR_c_656_n N_Y_c_833_n 0.0189039f $X=3.88 $Y=2.72 $X2=0 $Y2=0
cc_516 N_VPWR_c_651_n N_Y_c_833_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_517 N_VPWR_c_667_n N_Y_c_836_n 0.0189039f $X=4.72 $Y=2.72 $X2=0 $Y2=0
cc_518 N_VPWR_c_651_n N_Y_c_836_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_519 N_VPWR_M1001_d N_Y_c_805_n 0.00167154f $X=4.67 $Y=1.485 $X2=0 $Y2=0
cc_520 N_VPWR_c_658_n N_Y_c_805_n 0.0129161f $X=4.805 $Y=2 $X2=0 $Y2=0
cc_521 N_VPWR_c_678_n N_Y_c_858_n 0.0189039f $X=5.61 $Y=2.32 $X2=0 $Y2=0
cc_522 N_VPWR_c_679_n N_Y_c_858_n 0.0425789f $X=6.54 $Y=2.32 $X2=0 $Y2=0
cc_523 N_VPWR_c_651_n N_Y_c_858_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_524 N_VPWR_M1030_d N_Y_c_806_n 0.0200182f $X=5.51 $Y=1.485 $X2=0 $Y2=0
cc_525 N_VPWR_c_679_n N_Y_c_806_n 0.0766622f $X=6.54 $Y=2.32 $X2=0 $Y2=0
cc_526 N_VPWR_c_669_n N_Y_c_883_n 0.0189039f $X=7.24 $Y=2.72 $X2=0 $Y2=0
cc_527 N_VPWR_c_679_n N_Y_c_883_n 0.0458126f $X=6.54 $Y=2.32 $X2=0 $Y2=0
cc_528 N_VPWR_c_651_n N_Y_c_883_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_529 N_VPWR_M1016_d N_Y_c_807_n 0.00167154f $X=7.19 $Y=1.485 $X2=0 $Y2=0
cc_530 N_VPWR_c_659_n N_Y_c_807_n 0.0129161f $X=7.325 $Y=2 $X2=0 $Y2=0
cc_531 N_VPWR_c_671_n N_Y_c_890_n 0.0189039f $X=8.08 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_c_651_n N_Y_c_890_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_533 N_VPWR_M1026_d N_Y_c_808_n 0.00167154f $X=8.03 $Y=1.485 $X2=0 $Y2=0
cc_534 N_VPWR_c_660_n N_Y_c_808_n 0.0129161f $X=8.165 $Y=2 $X2=0 $Y2=0
cc_535 N_VPWR_c_661_n N_Y_c_894_n 0.0189039f $X=8.92 $Y=2.72 $X2=0 $Y2=0
cc_536 N_VPWR_c_651_n N_Y_c_894_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_537 N_VPWR_M1009_s N_Y_c_809_n 0.00167154f $X=8.87 $Y=1.485 $X2=0 $Y2=0
cc_538 N_VPWR_c_662_n N_Y_c_809_n 0.0129161f $X=9.005 $Y=2 $X2=0 $Y2=0
cc_539 N_VPWR_c_664_n N_Y_c_810_n 0.0108524f $X=9.845 $Y=1.66 $X2=0 $Y2=0
cc_540 N_VPWR_c_674_n N_Y_c_916_n 0.0189039f $X=9.76 $Y=2.72 $X2=0 $Y2=0
cc_541 N_VPWR_c_651_n N_Y_c_916_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_542 N_VPWR_M1024_d N_Y_c_811_n 5.57182e-19 $X=3.83 $Y=1.485 $X2=0 $Y2=0
cc_543 N_VPWR_M1024_d Y 0.00110365f $X=3.83 $Y=1.485 $X2=0 $Y2=0
cc_544 N_VPWR_c_657_n Y 0.0125076f $X=3.965 $Y=2 $X2=0 $Y2=0
cc_545 N_VPWR_c_653_n N_A_432_47#_c_1079_n 0.00232699f $X=2.285 $Y=1.66 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_664_n N_A_1266_47#_c_1175_n 7.37744e-19 $X=9.845 $Y=1.66 $X2=0
+ $Y2=0
cc_547 N_Y_M1014_d N_VGND_c_984_n 0.00216833f $X=2.57 $Y=0.235 $X2=0 $Y2=0
cc_548 N_Y_M1021_d N_VGND_c_984_n 0.00216833f $X=3.41 $Y=0.235 $X2=0 $Y2=0
cc_549 N_Y_c_801_n N_A_432_47#_M1019_s 0.00162409f $X=3.7 $Y=0.78 $X2=0 $Y2=0
cc_550 N_Y_c_846_n N_A_432_47#_M1027_s 0.00330818f $X=3.845 $Y=0.905 $X2=0 $Y2=0
cc_551 N_Y_c_801_n N_A_432_47#_c_1079_n 0.0111269f $X=3.7 $Y=0.78 $X2=0 $Y2=0
cc_552 N_Y_M1014_d N_A_432_47#_c_1080_n 0.0030596f $X=2.57 $Y=0.235 $X2=0 $Y2=0
cc_553 N_Y_M1021_d N_A_432_47#_c_1080_n 0.0030596f $X=3.41 $Y=0.235 $X2=0 $Y2=0
cc_554 N_Y_c_801_n N_A_432_47#_c_1080_n 0.0576505f $X=3.7 $Y=0.78 $X2=0 $Y2=0
cc_555 N_Y_c_846_n N_A_432_47#_c_1080_n 0.0176783f $X=3.845 $Y=0.905 $X2=0 $Y2=0
cc_556 N_Y_c_846_n N_A_850_47#_c_1122_n 0.0171782f $X=3.845 $Y=0.905 $X2=0 $Y2=0
cc_557 N_Y_c_806_n N_A_850_47#_c_1123_n 0.0247465f $X=6.74 $Y=1.555 $X2=0 $Y2=0
cc_558 N_Y_c_808_n N_A_1266_47#_c_1175_n 0.0161838f $X=8.42 $Y=1.555 $X2=0 $Y2=0
cc_559 N_VGND_c_984_n N_A_432_47#_M1014_s 0.0034899f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_560 N_VGND_c_984_n N_A_432_47#_M1019_s 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_984_n N_A_432_47#_M1027_s 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_984_n N_A_432_47#_M1025_d 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_563 N_VGND_c_984_n N_A_432_47#_M1034_d 0.00209344f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_564 N_VGND_c_981_n N_A_432_47#_c_1091_n 0.011673f $X=8.42 $Y=0 $X2=0 $Y2=0
cc_565 N_VGND_c_984_n N_A_432_47#_c_1091_n 0.00653933f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_566 N_VGND_c_981_n N_A_432_47#_c_1080_n 0.193456f $X=8.42 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_984_n N_A_432_47#_c_1080_n 0.123001f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_984_n N_A_850_47#_M1017_s 0.00216833f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_569 N_VGND_c_984_n N_A_850_47#_M1028_s 0.00216833f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_c_984_n N_A_850_47#_M1003_s 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_984_n N_A_850_47#_M1032_s 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_981_n N_A_850_47#_c_1123_n 0.0025345f $X=8.42 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_984_n N_A_850_47#_c_1123_n 0.00538493f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_981_n N_A_850_47#_c_1125_n 0.0121466f $X=8.42 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_c_984_n N_A_850_47#_c_1125_n 0.00653924f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_c_978_n N_A_850_47#_c_1126_n 0.00739696f $X=8.585 $Y=0.4 $X2=0
+ $Y2=0
cc_577 N_VGND_c_981_n N_A_850_47#_c_1126_n 0.101254f $X=8.42 $Y=0 $X2=0 $Y2=0
cc_578 N_VGND_c_984_n N_A_850_47#_c_1126_n 0.0635093f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_579 N_VGND_c_984_n N_A_1266_47#_M1003_d 0.00234744f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_580 N_VGND_c_984_n N_A_1266_47#_M1022_d 0.00216833f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_c_984_n N_A_1266_47#_M1033_d 0.00323135f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_984_n N_A_1266_47#_M1005_d 0.00323135f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_984_n N_A_1266_47#_M1029_d 0.00330716f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_M1002_s N_A_1266_47#_c_1175_n 0.00162029f $X=8.45 $Y=0.235 $X2=0
+ $Y2=0
cc_585 N_VGND_M1008_s N_A_1266_47#_c_1175_n 0.00162029f $X=9.29 $Y=0.235 $X2=0
+ $Y2=0
cc_586 N_VGND_c_978_n N_A_1266_47#_c_1175_n 0.0164771f $X=8.585 $Y=0.4 $X2=0
+ $Y2=0
cc_587 N_VGND_c_979_n N_A_1266_47#_c_1175_n 0.0164771f $X=9.425 $Y=0.4 $X2=0
+ $Y2=0
cc_588 N_VGND_c_981_n N_A_1266_47#_c_1175_n 0.00756245f $X=8.42 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_982_n N_A_1266_47#_c_1175_n 0.00755316f $X=9.26 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_983_n N_A_1266_47#_c_1175_n 0.00708556f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_984_n N_A_1266_47#_c_1175_n 0.0444689f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_592 N_A_432_47#_c_1080_n N_A_850_47#_M1017_s 0.00303751f $X=5.645 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_593 N_A_432_47#_c_1080_n N_A_850_47#_M1028_s 0.0030596f $X=5.645 $Y=0.4 $X2=0
+ $Y2=0
cc_594 N_A_432_47#_M1025_d N_A_850_47#_c_1122_n 0.00162409f $X=4.67 $Y=0.235
+ $X2=0 $Y2=0
cc_595 N_A_432_47#_c_1080_n N_A_850_47#_c_1122_n 0.0579741f $X=5.645 $Y=0.4
+ $X2=0 $Y2=0
cc_596 N_A_432_47#_M1034_d N_A_850_47#_c_1123_n 0.0031542f $X=5.51 $Y=0.235
+ $X2=0 $Y2=0
cc_597 N_A_432_47#_c_1080_n N_A_850_47#_c_1123_n 0.0181731f $X=5.645 $Y=0.4
+ $X2=0 $Y2=0
cc_598 N_A_432_47#_c_1080_n N_A_850_47#_c_1125_n 0.0213628f $X=5.645 $Y=0.4
+ $X2=0 $Y2=0
cc_599 N_A_850_47#_c_1126_n N_A_1266_47#_M1003_d 0.00585151f $X=7.745 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_600 N_A_850_47#_c_1126_n N_A_1266_47#_M1022_d 0.0030596f $X=7.745 $Y=0.4
+ $X2=0 $Y2=0
cc_601 N_A_850_47#_M1003_s N_A_1266_47#_c_1175_n 0.00162409f $X=6.77 $Y=0.235
+ $X2=0 $Y2=0
cc_602 N_A_850_47#_M1032_s N_A_1266_47#_c_1175_n 0.00162409f $X=7.61 $Y=0.235
+ $X2=0 $Y2=0
cc_603 N_A_850_47#_c_1123_n N_A_1266_47#_c_1175_n 0.0158347f $X=5.98 $Y=0.82
+ $X2=0 $Y2=0
cc_604 N_A_850_47#_c_1124_n N_A_1266_47#_c_1175_n 0.0066345f $X=6.065 $Y=0.735
+ $X2=0 $Y2=0
cc_605 N_A_850_47#_c_1126_n N_A_1266_47#_c_1175_n 0.0842077f $X=7.745 $Y=0.4
+ $X2=0 $Y2=0

* File: sky130_fd_sc_hd__or4b_4.pxi.spice
* Created: Tue Sep  1 19:28:52 2020
* 
x_PM_SKY130_FD_SC_HD__OR4B_4%D_N N_D_N_M1017_g N_D_N_M1010_g D_N D_N D_N
+ N_D_N_c_96_n N_D_N_c_97_n N_D_N_c_98_n PM_SKY130_FD_SC_HD__OR4B_4%D_N
x_PM_SKY130_FD_SC_HD__OR4B_4%A_109_93# N_A_109_93#_M1017_d N_A_109_93#_M1010_d
+ N_A_109_93#_c_121_n N_A_109_93#_M1003_g N_A_109_93#_M1002_g
+ N_A_109_93#_c_122_n N_A_109_93#_c_123_n N_A_109_93#_c_124_n
+ N_A_109_93#_c_129_n N_A_109_93#_c_162_p N_A_109_93#_c_125_n
+ N_A_109_93#_c_131_n PM_SKY130_FD_SC_HD__OR4B_4%A_109_93#
x_PM_SKY130_FD_SC_HD__OR4B_4%C N_C_M1001_g N_C_M1014_g N_C_c_176_n N_C_c_177_n C
+ C N_C_c_178_n C PM_SKY130_FD_SC_HD__OR4B_4%C
x_PM_SKY130_FD_SC_HD__OR4B_4%B N_B_c_224_n N_B_M1006_g N_B_M1012_g N_B_c_225_n
+ N_B_c_226_n B B B PM_SKY130_FD_SC_HD__OR4B_4%B
x_PM_SKY130_FD_SC_HD__OR4B_4%A N_A_M1004_g N_A_M1005_g A N_A_c_264_n N_A_c_265_n
+ N_A_c_266_n PM_SKY130_FD_SC_HD__OR4B_4%A
x_PM_SKY130_FD_SC_HD__OR4B_4%A_215_297# N_A_215_297#_M1003_d
+ N_A_215_297#_M1006_d N_A_215_297#_M1002_s N_A_215_297#_c_305_n
+ N_A_215_297#_M1007_g N_A_215_297#_M1000_g N_A_215_297#_c_306_n
+ N_A_215_297#_M1008_g N_A_215_297#_M1013_g N_A_215_297#_c_307_n
+ N_A_215_297#_M1009_g N_A_215_297#_M1015_g N_A_215_297#_c_308_n
+ N_A_215_297#_M1011_g N_A_215_297#_M1016_g N_A_215_297#_c_317_n
+ N_A_215_297#_c_309_n N_A_215_297#_c_328_n N_A_215_297#_c_342_n
+ N_A_215_297#_c_329_n N_A_215_297#_c_434_p N_A_215_297#_c_356_n
+ N_A_215_297#_c_310_n N_A_215_297#_c_311_n N_A_215_297#_c_386_p
+ N_A_215_297#_c_319_n N_A_215_297#_c_351_n N_A_215_297#_c_312_n
+ PM_SKY130_FD_SC_HD__OR4B_4%A_215_297#
x_PM_SKY130_FD_SC_HD__OR4B_4%VPWR N_VPWR_M1010_s N_VPWR_M1005_d N_VPWR_M1013_d
+ N_VPWR_M1016_d N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n VPWR N_VPWR_c_456_n N_VPWR_c_457_n
+ N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_449_n
+ PM_SKY130_FD_SC_HD__OR4B_4%VPWR
x_PM_SKY130_FD_SC_HD__OR4B_4%X N_X_M1007_s N_X_M1009_s N_X_M1000_s N_X_M1015_s
+ N_X_c_531_n N_X_c_572_n N_X_c_540_n N_X_c_532_n N_X_c_525_n N_X_c_526_n
+ N_X_c_555_n N_X_c_576_n N_X_c_533_n N_X_c_527_n N_X_c_528_n N_X_c_534_n X
+ N_X_c_530_n PM_SKY130_FD_SC_HD__OR4B_4%X
x_PM_SKY130_FD_SC_HD__OR4B_4%VGND N_VGND_M1017_s N_VGND_M1003_s N_VGND_M1001_d
+ N_VGND_M1004_d N_VGND_M1008_d N_VGND_M1011_d N_VGND_c_599_n N_VGND_c_600_n
+ N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n N_VGND_c_605_n
+ N_VGND_c_606_n N_VGND_c_607_n VGND N_VGND_c_608_n N_VGND_c_609_n
+ N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n N_VGND_c_614_n
+ N_VGND_c_615_n N_VGND_c_616_n PM_SKY130_FD_SC_HD__OR4B_4%VGND
cc_1 VNB N_D_N_c_96_n 0.033414f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_2 VNB N_D_N_c_97_n 0.0159032f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_3 VNB N_D_N_c_98_n 0.0215995f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=0.995
cc_4 VNB N_A_109_93#_c_121_n 0.0205822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_109_93#_c_122_n 0.0276756f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_6 VNB N_A_109_93#_c_123_n 0.00880176f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_7 VNB N_A_109_93#_c_124_n 0.00251166f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_8 VNB N_A_109_93#_c_125_n 0.0195202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_c_176_n 6.47944e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.785
cc_10 VNB N_C_c_177_n 0.0229145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_C_c_178_n 0.0171358f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_12 VNB N_B_c_224_n 0.0162189f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_B_c_225_n 0.00583329f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.785
cc_14 VNB N_B_c_226_n 0.0186258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_c_264_n 0.0229306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_c_265_n 6.43385e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_c_266_n 0.0174079f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_18 VNB N_A_215_297#_c_305_n 0.0163299f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.785
cc_19 VNB N_A_215_297#_c_306_n 0.0157937f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=0.995
cc_20 VNB N_A_215_297#_c_307_n 0.0157971f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.87
cc_21 VNB N_A_215_297#_c_308_n 0.0191578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_215_297#_c_309_n 0.00293881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_215_297#_c_310_n 0.00157854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_215_297#_c_311_n 0.00376665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_215_297#_c_312_n 0.0647168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_449_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_525_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.53
cc_28 VNB N_X_c_526_n 0.00187124f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.87
cc_29 VNB N_X_c_527_n 0.00105843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_528_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB X 0.0201786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_530_n 0.00836446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_599_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_34 VNB N_VGND_c_600_n 0.035054f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.19
cc_35 VNB N_VGND_c_601_n 0.0122259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_602_n 4.04385e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_603_n 0.00239633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_604_n 0.0148447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_605_n 0.0035091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_606_n 0.011288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_607_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_608_n 0.0206507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_609_n 0.0181903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_610_n 0.0135943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_611_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_612_n 0.00478242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_613_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_614_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_615_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_616_n 0.274996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VPB N_D_N_M1010_g 0.0666737f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_52 VPB N_D_N_c_96_n 0.00765717f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_53 VPB N_D_N_c_97_n 0.029026f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_54 VPB N_A_109_93#_M1002_g 0.02369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_109_93#_c_122_n 0.0103765f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_56 VPB N_A_109_93#_c_123_n 5.67856e-19 $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_57 VPB N_A_109_93#_c_129_n 4.94811e-19 $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_58 VPB N_A_109_93#_c_125_n 0.0114982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_109_93#_c_131_n 0.0161695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_C_M1014_g 0.0193425f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_61 VPB N_C_c_176_n 0.00103465f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.785
cc_62 VPB N_C_c_177_n 0.00584707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B_M1012_g 0.0174093f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_64 VPB N_B_c_225_n 0.00536776f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.785
cc_65 VPB N_B_c_226_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB B 2.2598e-19 $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_67 VPB N_A_M1005_g 0.0193215f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_68 VPB A 0.00385897f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_69 VPB N_A_c_264_n 0.00445127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_c_265_n 0.00148828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_215_297#_M1000_g 0.0199018f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_72 VPB N_A_215_297#_M1013_g 0.0182214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_215_297#_M1015_g 0.0182002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_215_297#_M1016_g 0.0219116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_215_297#_c_317_n 0.00718014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_215_297#_c_309_n 0.00111305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_215_297#_c_319_n 0.00203375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_215_297#_c_312_n 0.0102664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_450_n 0.0102718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_451_n 0.0197393f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_81 VPB N_VPWR_c_452_n 0.00463796f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_82 VPB N_VPWR_c_453_n 0.00399514f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.53
cc_83 VPB N_VPWR_c_454_n 0.011928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_455_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_456_n 0.0713355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_457_n 0.0181285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_458_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_459_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_460_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_449_n 0.0554648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_X_c_531_n 0.00246856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_X_c_532_n 0.00252706f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.19
cc_93 VPB N_X_c_533_n 0.0109401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_X_c_534_n 0.00220075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB X 0.00752913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 N_D_N_c_96_n N_A_109_93#_c_122_n 0.00754566f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_97 N_D_N_c_97_n N_A_109_93#_c_122_n 2.13875e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_98 N_D_N_c_98_n N_A_109_93#_c_124_n 0.00223695f $X=0.395 $Y=0.995 $X2=0 $Y2=0
cc_99 N_D_N_c_96_n N_A_109_93#_c_125_n 0.0036779f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_100 N_D_N_c_97_n N_A_109_93#_c_125_n 0.027596f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_101 N_D_N_c_98_n N_A_109_93#_c_125_n 0.00419785f $X=0.395 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_D_N_M1010_g N_A_109_93#_c_131_n 0.0177249f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_103 N_D_N_c_97_n N_A_109_93#_c_131_n 0.0473758f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_104 N_D_N_M1010_g N_VPWR_c_451_n 0.00469082f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_105 N_D_N_c_97_n N_VPWR_c_451_n 0.0208024f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_106 N_D_N_M1010_g N_VPWR_c_456_n 0.00585385f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_107 N_D_N_M1010_g N_VPWR_c_449_n 0.011417f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_108 N_D_N_c_97_n N_VPWR_c_449_n 0.0039654f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_109 N_D_N_c_96_n N_VGND_c_600_n 9.23671e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_110 N_D_N_c_97_n N_VGND_c_600_n 0.0211216f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_111 N_D_N_c_98_n N_VGND_c_600_n 0.00481075f $X=0.395 $Y=0.995 $X2=0 $Y2=0
cc_112 N_D_N_c_98_n N_VGND_c_601_n 0.00284681f $X=0.395 $Y=0.995 $X2=0 $Y2=0
cc_113 N_D_N_c_98_n N_VGND_c_608_n 0.00510437f $X=0.395 $Y=0.995 $X2=0 $Y2=0
cc_114 N_D_N_c_98_n N_VGND_c_616_n 0.00512902f $X=0.395 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_109_93#_M1002_g N_C_M1014_g 0.038256f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_109_93#_M1002_g N_C_c_176_n 0.00106197f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_109_93#_c_123_n N_C_c_176_n 3.03197e-19 $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_109_93#_c_123_n N_C_c_177_n 0.0153576f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_109_93#_M1002_g C 0.00502403f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_109_93#_c_121_n N_C_c_178_n 0.0196894f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_109_93#_M1002_g N_A_215_297#_c_317_n 0.0121867f $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_122 N_A_109_93#_c_131_n N_A_215_297#_c_317_n 0.0422878f $X=0.69 $Y=2.065
+ $X2=0 $Y2=0
cc_123 N_A_109_93#_c_121_n N_A_215_297#_c_309_n 0.00550471f $X=1.41 $Y=0.995
+ $X2=0 $Y2=0
cc_124 N_A_109_93#_M1002_g N_A_215_297#_c_309_n 0.00807212f $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_125 N_A_109_93#_c_123_n N_A_215_297#_c_309_n 0.00851631f $X=1.41 $Y=1.16
+ $X2=0 $Y2=0
cc_126 N_A_109_93#_c_125_n N_A_215_297#_c_309_n 0.023066f $X=0.7 $Y=1.067 $X2=0
+ $Y2=0
cc_127 N_A_109_93#_c_131_n N_A_215_297#_c_309_n 0.00627081f $X=0.69 $Y=2.065
+ $X2=0 $Y2=0
cc_128 N_A_109_93#_c_121_n N_A_215_297#_c_328_n 0.00412485f $X=1.41 $Y=0.995
+ $X2=0 $Y2=0
cc_129 N_A_109_93#_c_121_n N_A_215_297#_c_329_n 0.0071144f $X=1.41 $Y=0.995
+ $X2=0 $Y2=0
cc_130 N_A_109_93#_c_124_n N_A_215_297#_c_329_n 0.00406625f $X=0.69 $Y=0.81
+ $X2=0 $Y2=0
cc_131 N_A_109_93#_c_125_n N_A_215_297#_c_329_n 3.7164e-19 $X=0.7 $Y=1.067 $X2=0
+ $Y2=0
cc_132 N_A_109_93#_M1002_g N_A_215_297#_c_319_n 0.0147557f $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_133 N_A_109_93#_c_122_n N_A_215_297#_c_319_n 0.00438149f $X=1.335 $Y=1.16
+ $X2=0 $Y2=0
cc_134 N_A_109_93#_c_125_n N_A_215_297#_c_319_n 0.00997443f $X=0.7 $Y=1.067
+ $X2=0 $Y2=0
cc_135 N_A_109_93#_c_131_n N_A_215_297#_c_319_n 0.0107041f $X=0.69 $Y=2.065
+ $X2=0 $Y2=0
cc_136 N_A_109_93#_M1002_g N_VPWR_c_456_n 0.00541964f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_109_93#_c_162_p N_VPWR_c_456_n 0.0121939f $X=0.68 $Y=2.275 $X2=0
+ $Y2=0
cc_138 N_A_109_93#_M1010_d N_VPWR_c_449_n 0.00460309f $X=0.545 $Y=2.065 $X2=0
+ $Y2=0
cc_139 N_A_109_93#_M1002_g N_VPWR_c_449_n 0.0113112f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_109_93#_c_162_p N_VPWR_c_449_n 0.00719548f $X=0.68 $Y=2.275 $X2=0
+ $Y2=0
cc_141 N_A_109_93#_c_124_n N_VGND_c_600_n 0.00173604f $X=0.69 $Y=0.81 $X2=0
+ $Y2=0
cc_142 N_A_109_93#_c_121_n N_VGND_c_601_n 0.00468801f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_109_93#_c_122_n N_VGND_c_601_n 0.00348948f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_109_93#_c_124_n N_VGND_c_601_n 0.00879004f $X=0.69 $Y=0.81 $X2=0
+ $Y2=0
cc_145 N_A_109_93#_c_125_n N_VGND_c_601_n 0.00759979f $X=0.7 $Y=1.067 $X2=0
+ $Y2=0
cc_146 N_A_109_93#_c_121_n N_VGND_c_602_n 0.0012701f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_109_93#_c_124_n N_VGND_c_608_n 0.00623684f $X=0.69 $Y=0.81 $X2=0
+ $Y2=0
cc_148 N_A_109_93#_c_121_n N_VGND_c_609_n 0.00553912f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_109_93#_c_121_n N_VGND_c_616_n 0.0112327f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A_109_93#_c_124_n N_VGND_c_616_n 0.0065085f $X=0.69 $Y=0.81 $X2=0 $Y2=0
cc_151 N_C_c_178_n N_B_c_224_n 0.0251622f $X=1.88 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_152 N_C_M1014_g N_B_M1012_g 0.0567371f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_153 N_C_c_176_n N_B_M1012_g 6.68774e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_154 C N_B_M1012_g 0.0048871f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_155 N_C_c_176_n N_B_c_225_n 0.0274089f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_156 N_C_c_177_n N_B_c_225_n 0.00284781f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_157 N_C_c_176_n N_B_c_226_n 3.68507e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_158 N_C_c_177_n N_B_c_226_n 0.0203414f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_159 N_C_M1014_g B 0.00125078f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_160 N_C_c_176_n B 0.00618476f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_161 C B 0.0277816f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_162 C B 0.0277816f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_163 N_C_M1014_g N_A_215_297#_c_317_n 9.75761e-19 $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_164 C N_A_215_297#_c_317_n 0.0240505f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_165 N_C_M1014_g N_A_215_297#_c_309_n 7.22404e-19 $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_166 N_C_c_176_n N_A_215_297#_c_309_n 0.0421841f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_167 N_C_c_177_n N_A_215_297#_c_309_n 0.0021031f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_168 N_C_c_178_n N_A_215_297#_c_309_n 0.00338056f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_169 N_C_c_176_n N_A_215_297#_c_342_n 0.0108856f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_170 N_C_c_177_n N_A_215_297#_c_342_n 3.62043e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_171 N_C_c_178_n N_A_215_297#_c_342_n 0.0131138f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_172 N_C_c_177_n N_A_215_297#_c_329_n 0.00189854f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_173 N_C_M1014_g N_A_215_297#_c_319_n 5.94654e-19 $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_174 N_C_c_176_n N_A_215_297#_c_319_n 0.0140115f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_175 N_C_M1014_g N_VPWR_c_456_n 0.00375793f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_176 C N_VPWR_c_456_n 0.0132182f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_177 N_C_M1014_g N_VPWR_c_449_n 0.0056317f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_178 C N_VPWR_c_449_n 0.0124185f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_179 N_C_c_176_n A_297_297# 0.00117377f $X=1.88 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_180 C A_297_297# 0.00185709f $X=1.985 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_181 C A_297_297# 0.00785243f $X=2.07 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_182 C A_403_297# 0.00525495f $X=1.985 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_183 C A_403_297# 0.0059265f $X=2.07 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_184 N_C_c_178_n N_VGND_c_602_n 0.00869343f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_185 N_C_c_178_n N_VGND_c_609_n 0.00341689f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_186 N_C_c_178_n N_VGND_c_616_n 0.00431054f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_M1012_g N_A_M1005_g 0.0564998f $X=2.36 $Y=1.985 $X2=0 $Y2=0
cc_188 B N_A_M1005_g 0.00907078f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_189 N_B_c_225_n A 0.0102002f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B_c_225_n N_A_c_264_n 0.00369534f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B_c_226_n N_A_c_264_n 0.0203414f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B_c_225_n N_A_c_265_n 0.0271074f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B_c_226_n N_A_c_265_n 3.68507e-19 $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B_c_224_n N_A_c_266_n 0.0243955f $X=2.36 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B_c_224_n N_A_215_297#_c_342_n 0.0110728f $X=2.36 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B_c_225_n N_A_215_297#_c_342_n 0.018226f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B_c_226_n N_A_215_297#_c_342_n 2.98597e-19 $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B_c_225_n N_A_215_297#_c_351_n 0.00316818f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_199 B N_VPWR_c_452_n 0.0308975f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_200 N_B_M1012_g N_VPWR_c_456_n 0.00447054f $X=2.36 $Y=1.985 $X2=0 $Y2=0
cc_201 B N_VPWR_c_456_n 0.0117985f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_202 N_B_M1012_g N_VPWR_c_449_n 0.00724306f $X=2.36 $Y=1.985 $X2=0 $Y2=0
cc_203 B N_VPWR_c_449_n 0.0104425f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_204 B A_487_297# 0.0163657f $X=2.445 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_205 N_B_c_224_n N_VGND_c_602_n 0.00732663f $X=2.36 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B_c_224_n N_VGND_c_610_n 0.00341689f $X=2.36 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B_c_224_n N_VGND_c_616_n 0.00405445f $X=2.36 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_c_266_n N_A_215_297#_c_305_n 0.0200495f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_M1005_g N_A_215_297#_M1000_g 0.0173803f $X=2.78 $Y=1.985 $X2=0 $Y2=0
cc_210 A N_A_215_297#_M1000_g 0.00128363f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_211 N_A_c_265_n N_A_215_297#_M1000_g 0.00219223f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_212 A N_A_215_297#_c_356_n 0.00495213f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_213 N_A_c_264_n N_A_215_297#_c_356_n 0.00173573f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_c_265_n N_A_215_297#_c_356_n 0.0104547f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_c_266_n N_A_215_297#_c_356_n 0.0134819f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_c_264_n N_A_215_297#_c_310_n 5.07416e-19 $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_c_265_n N_A_215_297#_c_310_n 0.00568393f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_c_266_n N_A_215_297#_c_310_n 0.00336447f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_219 A N_A_215_297#_c_311_n 0.00707041f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_220 N_A_c_264_n N_A_215_297#_c_311_n 0.00124527f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_c_265_n N_A_215_297#_c_311_n 0.0137152f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_c_264_n N_A_215_297#_c_312_n 0.0161964f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_c_265_n N_A_215_297#_c_312_n 7.74805e-19 $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_224 A N_VPWR_M1005_d 0.00433176f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_225 N_A_M1005_g N_VPWR_c_452_n 0.00789297f $X=2.78 $Y=1.985 $X2=0 $Y2=0
cc_226 A N_VPWR_c_452_n 0.0193325f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_227 N_A_M1005_g N_VPWR_c_456_n 0.00585385f $X=2.78 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_M1005_g N_VPWR_c_449_n 0.0109527f $X=2.78 $Y=1.985 $X2=0 $Y2=0
cc_229 A N_X_c_531_n 0.00229946f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_230 N_A_c_266_n N_VGND_c_602_n 6.8876e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_266_n N_VGND_c_603_n 0.00318791f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_266_n N_VGND_c_610_n 0.00428022f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_c_266_n N_VGND_c_616_n 0.00603983f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_215_297#_M1000_g N_VPWR_c_452_n 0.00430866f $X=3.31 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_215_297#_M1013_g N_VPWR_c_453_n 0.00165046f $X=3.73 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_215_297#_M1015_g N_VPWR_c_453_n 0.00157837f $X=4.15 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_215_297#_M1016_g N_VPWR_c_455_n 0.00338128f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_215_297#_c_317_n N_VPWR_c_456_n 0.0192488f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_239 N_A_215_297#_M1000_g N_VPWR_c_457_n 0.00585385f $X=3.31 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_215_297#_M1013_g N_VPWR_c_457_n 0.00585385f $X=3.73 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_215_297#_M1015_g N_VPWR_c_458_n 0.00585385f $X=4.15 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_215_297#_M1016_g N_VPWR_c_458_n 0.00585385f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_215_297#_M1002_s N_VPWR_c_449_n 0.00209863f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_244 N_A_215_297#_M1000_g N_VPWR_c_449_n 0.0108486f $X=3.31 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_A_215_297#_M1013_g N_VPWR_c_449_n 0.0104367f $X=3.73 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_A_215_297#_M1015_g N_VPWR_c_449_n 0.0104367f $X=4.15 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_215_297#_M1016_g N_VPWR_c_449_n 0.0114096f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_248 N_A_215_297#_c_317_n N_VPWR_c_449_n 0.0123483f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_249 N_A_215_297#_c_309_n A_297_297# 0.00101535f $X=1.54 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_250 N_A_215_297#_c_319_n A_297_297# 0.0048664f $X=1.54 $Y=1.66 $X2=-0.19
+ $Y2=-0.24
cc_251 N_A_215_297#_M1000_g N_X_c_531_n 2.80238e-19 $X=3.31 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_215_297#_c_386_p N_X_c_531_n 0.0172286f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_215_297#_c_312_n N_X_c_531_n 0.00226413f $X=4.57 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_215_297#_c_306_n N_X_c_540_n 0.00701434f $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_215_297#_c_307_n N_X_c_540_n 5.23786e-19 $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_215_297#_M1013_g N_X_c_532_n 0.0134538f $X=3.73 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A_215_297#_M1015_g N_X_c_532_n 0.013468f $X=4.15 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_215_297#_c_386_p N_X_c_532_n 0.03482f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_215_297#_c_312_n N_X_c_532_n 0.00216069f $X=4.57 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A_215_297#_c_306_n N_X_c_525_n 0.00870364f $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_215_297#_c_307_n N_X_c_525_n 0.00865686f $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_215_297#_c_386_p N_X_c_525_n 0.0356734f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_215_297#_c_312_n N_X_c_525_n 0.00222133f $X=4.57 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_215_297#_c_305_n N_X_c_526_n 8.16938e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_215_297#_c_306_n N_X_c_526_n 0.00250064f $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_215_297#_c_310_n N_X_c_526_n 0.00357582f $X=3.18 $Y=1.075 $X2=0 $Y2=0
cc_267 N_A_215_297#_c_386_p N_X_c_526_n 0.01996f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_215_297#_c_312_n N_X_c_526_n 0.00230339f $X=4.57 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_215_297#_c_306_n N_X_c_555_n 5.22228e-19 $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_215_297#_c_307_n N_X_c_555_n 0.00630972f $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_215_297#_c_308_n N_X_c_555_n 0.0109314f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_215_297#_M1016_g N_X_c_533_n 0.0159073f $X=4.57 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_215_297#_c_386_p N_X_c_533_n 0.00401279f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_215_297#_c_308_n N_X_c_527_n 0.0113288f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A_215_297#_c_386_p N_X_c_527_n 0.00200821f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_215_297#_c_307_n N_X_c_528_n 0.00113286f $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A_215_297#_c_308_n N_X_c_528_n 0.00113286f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_215_297#_c_386_p N_X_c_528_n 0.026256f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_215_297#_c_312_n N_X_c_528_n 0.00230339f $X=4.57 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_215_297#_c_386_p N_X_c_534_n 0.0172286f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_281 N_A_215_297#_c_312_n N_X_c_534_n 0.00226413f $X=4.57 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_215_297#_c_308_n X 0.0212036f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A_215_297#_c_386_p X 0.0137657f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_215_297#_c_342_n N_VGND_M1001_d 0.00664072f $X=2.485 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_215_297#_c_356_n N_VGND_M1004_d 0.00616911f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_215_297#_c_310_n N_VGND_M1004_d 7.20909e-19 $X=3.18 $Y=1.075 $X2=0
+ $Y2=0
cc_287 N_A_215_297#_c_328_n N_VGND_c_602_n 0.0117247f $X=1.7 $Y=0.49 $X2=0 $Y2=0
cc_288 N_A_215_297#_c_342_n N_VGND_c_602_n 0.0160613f $X=2.485 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_215_297#_c_305_n N_VGND_c_603_n 0.00675761f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_215_297#_c_306_n N_VGND_c_603_n 5.99174e-19 $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_215_297#_c_356_n N_VGND_c_603_n 0.0224385f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_215_297#_c_305_n N_VGND_c_604_n 0.00496106f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_215_297#_c_306_n N_VGND_c_604_n 0.00423334f $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_215_297#_c_306_n N_VGND_c_605_n 0.00138579f $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A_215_297#_c_307_n N_VGND_c_605_n 0.00146448f $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_215_297#_c_308_n N_VGND_c_607_n 0.00316354f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_215_297#_c_328_n N_VGND_c_609_n 0.00852533f $X=1.7 $Y=0.49 $X2=0
+ $Y2=0
cc_298 N_A_215_297#_c_329_n N_VGND_c_609_n 0.00502163f $X=1.785 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_215_297#_c_342_n N_VGND_c_610_n 0.00232396f $X=2.485 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_215_297#_c_434_p N_VGND_c_610_n 0.00846569f $X=2.57 $Y=0.49 $X2=0
+ $Y2=0
cc_301 N_A_215_297#_c_356_n N_VGND_c_610_n 0.0029785f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_302 N_A_215_297#_c_307_n N_VGND_c_611_n 0.00423334f $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_215_297#_c_308_n N_VGND_c_611_n 0.00423334f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_215_297#_M1003_d N_VGND_c_616_n 0.00390697f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_305 N_A_215_297#_M1006_d N_VGND_c_616_n 0.00256656f $X=2.435 $Y=0.235 $X2=0
+ $Y2=0
cc_306 N_A_215_297#_c_305_n N_VGND_c_616_n 0.00822344f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_215_297#_c_306_n N_VGND_c_616_n 0.00575518f $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_215_297#_c_307_n N_VGND_c_616_n 0.0057163f $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_215_297#_c_308_n N_VGND_c_616_n 0.00668918f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_A_215_297#_c_328_n N_VGND_c_616_n 0.00618681f $X=1.7 $Y=0.49 $X2=0
+ $Y2=0
cc_311 N_A_215_297#_c_342_n N_VGND_c_616_n 0.00554474f $X=2.485 $Y=0.74 $X2=0
+ $Y2=0
cc_312 N_A_215_297#_c_329_n N_VGND_c_616_n 0.00936859f $X=1.785 $Y=0.74 $X2=0
+ $Y2=0
cc_313 N_A_215_297#_c_434_p N_VGND_c_616_n 0.00625722f $X=2.57 $Y=0.49 $X2=0
+ $Y2=0
cc_314 N_A_215_297#_c_356_n N_VGND_c_616_n 0.00734097f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_449_n A_297_297# 0.0138706f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_316 N_VPWR_c_449_n A_403_297# 0.00676138f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_317 N_VPWR_c_449_n A_487_297# 0.0046981f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_318 N_VPWR_c_449_n N_X_M1000_s 0.00284632f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_c_449_n N_X_M1015_s 0.00284632f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_c_457_n N_X_c_572_n 0.0142343f $X=3.815 $Y=2.72 $X2=0 $Y2=0
cc_321 N_VPWR_c_449_n N_X_c_572_n 0.00955092f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_M1013_d N_X_c_532_n 0.00165831f $X=3.805 $Y=1.485 $X2=0 $Y2=0
cc_323 N_VPWR_c_453_n N_X_c_532_n 0.0126919f $X=3.94 $Y=1.96 $X2=0 $Y2=0
cc_324 N_VPWR_c_458_n N_X_c_576_n 0.0142343f $X=4.655 $Y=2.72 $X2=0 $Y2=0
cc_325 N_VPWR_c_449_n N_X_c_576_n 0.00955092f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_326 N_VPWR_M1016_d N_X_c_533_n 0.00283464f $X=4.645 $Y=1.485 $X2=0 $Y2=0
cc_327 N_VPWR_c_455_n N_X_c_533_n 0.0179737f $X=4.78 $Y=1.96 $X2=0 $Y2=0
cc_328 N_X_c_525_n N_VGND_M1008_d 0.00162089f $X=4.195 $Y=0.815 $X2=0 $Y2=0
cc_329 N_X_c_527_n N_VGND_M1011_d 2.28588e-19 $X=4.725 $Y=0.815 $X2=0 $Y2=0
cc_330 N_X_c_530_n N_VGND_M1011_d 0.00344973f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_331 N_X_c_540_n N_VGND_c_604_n 0.0151398f $X=3.52 $Y=0.485 $X2=0 $Y2=0
cc_332 N_X_c_525_n N_VGND_c_604_n 0.00198695f $X=4.195 $Y=0.815 $X2=0 $Y2=0
cc_333 N_X_c_525_n N_VGND_c_605_n 0.0122559f $X=4.195 $Y=0.815 $X2=0 $Y2=0
cc_334 N_X_c_530_n N_VGND_c_606_n 0.00165369f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_335 N_X_c_527_n N_VGND_c_607_n 0.00177288f $X=4.725 $Y=0.815 $X2=0 $Y2=0
cc_336 N_X_c_530_n N_VGND_c_607_n 0.0120207f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_337 N_X_c_525_n N_VGND_c_611_n 0.00198695f $X=4.195 $Y=0.815 $X2=0 $Y2=0
cc_338 N_X_c_555_n N_VGND_c_611_n 0.0188551f $X=4.36 $Y=0.39 $X2=0 $Y2=0
cc_339 N_X_c_527_n N_VGND_c_611_n 0.00198695f $X=4.725 $Y=0.815 $X2=0 $Y2=0
cc_340 N_X_M1007_s N_VGND_c_616_n 0.00393857f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_341 N_X_M1009_s N_VGND_c_616_n 0.00215201f $X=4.225 $Y=0.235 $X2=0 $Y2=0
cc_342 N_X_c_540_n N_VGND_c_616_n 0.00940698f $X=3.52 $Y=0.485 $X2=0 $Y2=0
cc_343 N_X_c_525_n N_VGND_c_616_n 0.00835832f $X=4.195 $Y=0.815 $X2=0 $Y2=0
cc_344 N_X_c_555_n N_VGND_c_616_n 0.0122069f $X=4.36 $Y=0.39 $X2=0 $Y2=0
cc_345 N_X_c_527_n N_VGND_c_616_n 0.00396723f $X=4.725 $Y=0.815 $X2=0 $Y2=0
cc_346 N_X_c_530_n N_VGND_c_616_n 0.00345847f $X=4.845 $Y=0.905 $X2=0 $Y2=0

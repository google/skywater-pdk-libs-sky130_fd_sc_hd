* NGSPICE file created from sky130_fd_sc_hd__o2111a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR C1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.88e+12p pd=1.776e+07u as=1.67e+12p ps=1.334e+07u
M1001 VGND A1 a_361_47# VNB nshort w=650000u l=150000u
+  ad=1.001e+12p pd=9.58e+06u as=6.2075e+11p ps=5.81e+06u
M1002 a_27_297# D1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_297# C1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_681_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1005 a_361_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_27_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1008 a_681_297# A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_47# D1 a_27_297# VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u
M1010 VPWR a_27_297# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_47# C1 a_445_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.365e+11p ps=1.72e+06u
M1012 a_361_47# B1 a_277_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1013 VGND a_27_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_277_47# C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR D1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_27_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A2 a_361_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_852_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.55e+11p pd=2.71e+06u as=0p ps=0u
M1020 a_445_47# B1 a_361_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_361_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_27_297# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_297# D1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_27_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_297# A2 a_852_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__einvn_1.spice
* Created: Thu Aug 27 14:20:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__einvn_1.spice.pex"
.subckt sky130_fd_sc_hd__einvn_1  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_TE_B_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.180757 AS=0.1092 PD=1.08729 PS=1.36 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1003 A_286_47# N_A_27_47#_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.279743 PD=0.975 PS=1.68271 NRD=19.836 NRS=11.076 M=1
+ R=4.33333 SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g A_286_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.105625 PD=1.82 PS=0.975 NRD=0 NRS=19.836 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=6.1464 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1000 A_204_297# N_TE_B_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.3675
+ AS=0.181707 PD=1.735 PS=1.61585 NRD=61.5428 NRS=4.9053 M=1 R=6.66667
+ SA=75000.5 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1004 N_Z_M1004_d N_A_M1004_g A_204_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.3675 PD=2.52 PS=1.735 NRD=0 NRS=61.5428 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_21 VNB 0 1.65488e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__einvn_1.spice.SKY130_FD_SC_HD__EINVN_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdfbbn_1.pex.spice
* Created: Thu Aug 27 14:45:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%CLK_N 4 5 7 8 10 13 17 19 20 24 26
c45 13 0 2.71124e-20 $X=0.47 $Y=0.805
r46 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r47 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r48 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r49 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r50 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r51 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r52 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r53 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r54 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r55 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r56 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r57 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r59 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_27_47# 1 2 9 13 17 19 20 23 26 27 29 32
+ 36 40 41 42 46 47 49 51 52 55 58 59 61 62 63 66 70 71 74 81 84
c286 84 0 9.50836e-20 $X=5.165 $Y=0.93
c287 70 0 1.98367e-19 $X=5.24 $Y=0.85
c288 63 0 8.87067e-20 $X=5.385 $Y=1.19
c289 61 0 9.24143e-20 $X=5.277 $Y=1.12
c290 49 0 1.22107e-19 $X=8.937 $Y=1.305
c291 47 0 1.7288e-19 $X=8.615 $Y=0.87
c292 17 0 4.75142e-20 $X=4.59 $Y=2.275
r293 84 87 39.0501 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=0.93
+ $X2=5.15 $Y2=1.095
r294 84 86 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=0.93
+ $X2=5.15 $Y2=0.765
r295 78 81 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=0.75 $Y=1.235
+ $X2=0.89 $Y2=1.235
r296 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.235 $X2=0.75 $Y2=1.235
r297 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.19
+ $X2=8.51 $Y2=1.19
r298 71 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.165
+ $Y=0.93 $X2=5.165 $Y2=0.93
r299 70 72 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=5.24 $Y=0.85
+ $X2=5.24 $Y2=0.965
r300 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.24 $Y=0.85
+ $X2=5.24 $Y2=0.85
r301 66 79 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.72 $Y=0.85
+ $X2=0.72 $Y2=1.235
r302 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0.85
+ $X2=0.69 $Y2=0.85
r303 62 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=8.51 $Y2=1.19
r304 62 63 3.68811 $w=1.4e-07 $l=2.98e-06 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=5.385 $Y2=1.19
r305 61 63 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=5.277 $Y=1.12
+ $X2=5.385 $Y2=1.19
r306 61 72 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=5.277 $Y=1.12
+ $X2=5.277 $Y2=0.965
r307 59 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=0.85
+ $X2=0.69 $Y2=0.85
r308 58 70 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=5.095 $Y=0.85
+ $X2=5.24 $Y2=0.85
r309 58 59 5.27227 $w=1.4e-07 $l=4.26e-06 $layer=MET1_cond $X=5.095 $Y=0.85
+ $X2=0.835 $Y2=0.85
r310 57 79 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.72 $Y=1.795
+ $X2=0.72 $Y2=1.235
r311 56 66 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.72 $Y=0.805
+ $X2=0.72 $Y2=0.85
r312 52 94 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.955 $Y=1.74
+ $X2=8.955 $Y2=1.875
r313 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.955
+ $Y=1.74 $X2=8.955 $Y2=1.74
r314 49 75 26.3101 $w=1.78e-07 $l=4.27e-07 $layer=LI1_cond $X=8.937 $Y=1.215
+ $X2=8.51 $Y2=1.215
r315 49 51 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=8.937 $Y=1.305
+ $X2=8.937 $Y2=1.74
r316 47 88 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=8.615 $Y=0.87
+ $X2=8.495 $Y2=0.87
r317 46 75 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=8.562 $Y=0.87
+ $X2=8.562 $Y2=1.125
r318 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.615
+ $Y=0.87 $X2=8.615 $Y2=0.87
r319 43 55 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.22 $Y2=1.88
r320 42 57 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.72 $Y2=1.795
r321 42 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.345 $Y2=1.88
r322 40 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.72 $Y2=0.805
r323 40 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.345 $Y2=0.72
r324 34 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=0.635
+ $X2=0.345 $Y2=0.72
r325 34 36 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.22 $Y=0.635
+ $X2=0.22 $Y2=0.51
r326 32 94 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.925 $Y=2.275
+ $X2=8.925 $Y2=1.875
r327 27 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.495 $Y=0.705
+ $X2=8.495 $Y2=0.87
r328 27 29 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.495 $Y=0.705
+ $X2=8.495 $Y2=0.415
r329 26 87 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=5.102 $Y=1.245
+ $X2=5.102 $Y2=1.095
r330 23 86 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.075 $Y=0.415
+ $X2=5.075 $Y2=0.765
r331 19 26 27.7801 $w=1.5e-07 $l=1.34365e-07 $layer=POLY_cond $X=5 $Y=1.32
+ $X2=5.102 $Y2=1.245
r332 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5 $Y=1.32
+ $X2=4.665 $Y2=1.32
r333 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.59 $Y=1.395
+ $X2=4.665 $Y2=1.32
r334 15 17 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.59 $Y=1.395
+ $X2=4.59 $Y2=2.275
r335 11 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r336 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r337 7 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r338 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r339 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r340 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%SCD 1 2 3 5 8 12 13 19
c52 12 0 1.76673e-19 $X=1.61 $Y=1.19
c53 8 0 1.50346e-19 $X=1.83 $Y=2.135
c54 1 0 1.68616e-20 $X=1.642 $Y=0.88
r55 17 19 5.86464 $w=2.63e-07 $l=3.2e-08 $layer=POLY_cond $X=1.61 $Y=1.49
+ $X2=1.642 $Y2=1.49
r56 13 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.49 $X2=1.61 $Y2=1.49
r57 12 13 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=1.555 $Y=1.19
+ $X2=1.555 $Y2=1.49
r58 6 19 34.4548 $w=2.63e-07 $l=2.57612e-07 $layer=POLY_cond $X=1.83 $Y=1.655
+ $X2=1.642 $Y2=1.49
r59 6 8 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.655 $X2=1.83
+ $Y2=2.135
r60 3 11 0.795936 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=0.73
+ $X2=1.83 $Y2=0.805
r61 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.73 $X2=1.83
+ $Y2=0.445
r62 2 19 12.4247 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.642 $Y=1.325
+ $X2=1.642 $Y2=1.49
r63 1 11 65.6638 $w=1.38e-07 $l=1.88e-07 $layer=POLY_cond $X=1.642 $Y=0.805
+ $X2=1.83 $Y2=0.805
r64 1 2 177.918 $w=1.75e-07 $l=4.45e-07 $layer=POLY_cond $X=1.642 $Y=0.88
+ $X2=1.642 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_423_315# 1 2 7 9 10 11 14 17 21 23 24 25
+ 27 28 34 38 39 42
c113 39 0 8.91744e-20 $X=2.845 $Y=1.65
c114 38 0 1.01009e-19 $X=3.615 $Y=0.93
c115 27 0 9.78226e-20 $X=3.517 $Y=1.095
c116 11 0 5.57791e-20 $X=2.265 $Y=1.65
r117 38 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.615 $Y=0.93
+ $X2=3.615 $Y2=0.765
r118 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=0.93 $X2=3.615 $Y2=0.93
r119 35 37 8.88742 $w=3.02e-07 $l=2.2e-07 $layer=LI1_cond $X=3.6 $Y=0.71 $X2=3.6
+ $Y2=0.93
r120 33 34 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=1.74
+ $X2=3.14 $Y2=1.74
r121 31 39 16.1264 $w=2.69e-07 $l=9e-08 $layer=POLY_cond $X=2.845 $Y=1.74
+ $X2=2.845 $Y2=1.65
r122 30 33 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.845 $Y=1.74
+ $X2=3.055 $Y2=1.74
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.74 $X2=2.845 $Y2=1.74
r124 27 37 8.80496 $w=3.02e-07 $l=2.02287e-07 $layer=LI1_cond $X=3.517 $Y=1.095
+ $X2=3.6 $Y2=0.93
r125 27 28 30.4208 $w=1.73e-07 $l=4.8e-07 $layer=LI1_cond $X=3.517 $Y=1.095
+ $X2=3.517 $Y2=1.575
r126 25 28 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.43 $Y=1.66
+ $X2=3.517 $Y2=1.575
r127 25 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.43 $Y=1.66
+ $X2=3.14 $Y2=1.66
r128 23 35 4.10007 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.43 $Y=0.71 $X2=3.6
+ $Y2=0.71
r129 23 24 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.43 $Y=0.71
+ $X2=3.04 $Y2=0.71
r130 19 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=1.905
+ $X2=3.055 $Y2=1.74
r131 19 21 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.055 $Y=1.905
+ $X2=3.055 $Y2=2.3
r132 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.955 $Y=0.625
+ $X2=3.04 $Y2=0.71
r133 15 17 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.955 $Y=0.625
+ $X2=2.955 $Y2=0.47
r134 14 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.6 $Y=0.445
+ $X2=3.6 $Y2=0.765
r135 10 39 16.4183 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.71 $Y=1.65
+ $X2=2.845 $Y2=1.65
r136 10 11 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.71 $Y=1.65
+ $X2=2.265 $Y2=1.65
r137 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.19 $Y=1.725
+ $X2=2.265 $Y2=1.65
r138 7 9 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.19 $Y=1.725
+ $X2=2.19 $Y2=2.135
r139 2 21 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=2.065 $X2=3.055 $Y2=2.3
r140 1 17 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.235 $X2=2.955 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%SCE 1 3 4 6 8 10 12 13 15 16 18 20 21 24 26
+ 27 28 29 34 37 44
c115 34 0 1.20894e-19 $X=2.242 $Y=0.81
r116 42 44 2.09535 $w=2.18e-07 $l=4e-08 $layer=LI1_cond $X=2.045 $Y=1.15
+ $X2=2.045 $Y2=1.19
r117 38 42 3.19822 $w=2.2e-07 $l=1.68e-07 $layer=LI1_cond $X=2.045 $Y=0.982
+ $X2=2.045 $Y2=1.15
r118 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=0.985 $X2=2.23 $Y2=0.985
r119 34 36 28.4007 $w=2.97e-07 $l=1.75e-07 $layer=POLY_cond $X=2.242 $Y=0.81
+ $X2=2.242 $Y2=0.985
r120 28 37 5.50421 $w=3.33e-07 $l=1.6e-07 $layer=LI1_cond $X=2.07 $Y=0.982
+ $X2=2.23 $Y2=0.982
r121 28 38 0.860032 $w=3.33e-07 $l=2.5e-08 $layer=LI1_cond $X=2.07 $Y=0.982
+ $X2=2.045 $Y2=0.982
r122 28 29 16.658 $w=2.18e-07 $l=3.18e-07 $layer=LI1_cond $X=2.045 $Y=1.212
+ $X2=2.045 $Y2=1.53
r123 28 44 1.15244 $w=2.18e-07 $l=2.2e-08 $layer=LI1_cond $X=2.045 $Y=1.212
+ $X2=2.045 $Y2=1.19
r124 27 38 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=2.045 $Y=0.51
+ $X2=2.045 $Y2=0.815
r125 22 24 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.165 $Y=1.33
+ $X2=3.265 $Y2=1.33
r126 18 20 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.685 $Y=1.985
+ $X2=3.685 $Y2=2.275
r127 17 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=1.91
+ $X2=3.265 $Y2=1.91
r128 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.61 $Y=1.91
+ $X2=3.685 $Y2=1.985
r129 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.61 $Y=1.91
+ $X2=3.34 $Y2=1.91
r130 13 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.985
+ $X2=3.265 $Y2=1.91
r131 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.265 $Y=1.985
+ $X2=3.265 $Y2=2.275
r132 12 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.835
+ $X2=3.265 $Y2=1.91
r133 11 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.405
+ $X2=3.265 $Y2=1.33
r134 11 12 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.265 $Y=1.405
+ $X2=3.265 $Y2=1.835
r135 10 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.255
+ $X2=3.165 $Y2=1.33
r136 9 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=0.885
+ $X2=3.165 $Y2=0.81
r137 9 10 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.165 $Y=0.885
+ $X2=3.165 $Y2=1.255
r138 6 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=0.735
+ $X2=3.165 $Y2=0.81
r139 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.165 $Y=0.735
+ $X2=3.165 $Y2=0.445
r140 5 34 18.7323 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=2.395 $Y=0.81
+ $X2=2.242 $Y2=0.81
r141 4 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.09 $Y=0.81
+ $X2=3.165 $Y2=0.81
r142 4 5 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.09 $Y=0.81
+ $X2=2.395 $Y2=0.81
r143 1 34 23.9601 $w=2.97e-07 $l=9.75961e-08 $layer=POLY_cond $X=2.19 $Y=0.735
+ $X2=2.242 $Y2=0.81
r144 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.19 $Y=0.735
+ $X2=2.19 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%D 3 7 9 10 18 20
r57 17 18 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=4.035 $Y=1.49
+ $X2=4.105 $Y2=1.49
r58 14 17 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.94 $Y=1.49
+ $X2=4.035 $Y2=1.49
r59 10 20 26.2365 $w=2.33e-07 $l=5.35e-07 $layer=LI1_cond $X=3.942 $Y=2.21
+ $X2=3.942 $Y2=1.675
r60 9 20 7.99605 $w=3.13e-07 $l=1.85997e-07 $layer=LI1_cond $X=3.94 $Y=1.49
+ $X2=3.942 $Y2=1.675
r61 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.49 $X2=3.94 $Y2=1.49
r62 5 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=1.49
r63 5 7 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=2.275
r64 1 17 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.035 $Y=1.355
+ $X2=4.035 $Y2=1.49
r65 1 3 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.035 $Y=1.355
+ $X2=4.035 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_193_47# 1 2 7 9 12 18 20 21 24 27 29 30
+ 33 34 35 36 45 53 54 58 59 60 63
c225 58 0 2.05666e-19 $X=8.445 $Y=1.74
c226 54 0 1.98367e-19 $X=5.04 $Y=1.74
c227 53 0 8.87067e-20 $X=5.04 $Y=1.74
c228 30 0 9.24143e-20 $X=4.655 $Y=0.87
c229 18 0 3.84972e-20 $X=8.505 $Y=2.275
r230 58 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.74
+ $X2=8.445 $Y2=1.905
r231 58 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.74
+ $X2=8.445 $Y2=1.575
r232 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.445
+ $Y=1.74 $X2=8.445 $Y2=1.74
r233 53 56 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.04 $Y=1.74
+ $X2=5.04 $Y2=1.875
r234 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.74 $X2=5.04 $Y2=1.74
r235 45 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.87
+ $X2=8.51 $Y2=1.87
r236 43 54 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=1.765
+ $X2=5.04 $Y2=1.765
r237 43 71 3.88191 $w=3.78e-07 $l=1.28e-07 $layer=LI1_cond $X=4.83 $Y=1.765
+ $X2=4.702 $Y2=1.765
r238 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.87
+ $X2=4.83 $Y2=1.87
r239 39 63 71.2419 $w=2.18e-07 $l=1.36e-06 $layer=LI1_cond $X=1.125 $Y=1.87
+ $X2=1.125 $Y2=0.51
r240 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r241 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=1.87
+ $X2=4.83 $Y2=1.87
r242 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.87
+ $X2=8.51 $Y2=1.87
r243 35 36 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=8.365 $Y=1.87
+ $X2=4.975 $Y2=1.87
r244 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r245 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=4.83 $Y2=1.87
r246 33 34 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=1.295 $Y2=1.87
r247 30 48 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.655 $Y=0.87
+ $X2=4.51 $Y2=0.87
r248 29 32 9.15829 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.68 $Y=0.87
+ $X2=4.68 $Y2=1.035
r249 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.655
+ $Y=0.87 $X2=4.655 $Y2=0.87
r250 27 71 5.30917 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=4.702 $Y=1.575
+ $X2=4.702 $Y2=1.765
r251 27 32 34.2234 $w=1.73e-07 $l=5.4e-07 $layer=LI1_cond $X=4.702 $Y=1.575
+ $X2=4.702 $Y2=1.035
r252 22 24 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.035 $Y=1.245
+ $X2=9.035 $Y2=0.415
r253 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.96 $Y=1.32
+ $X2=9.035 $Y2=1.245
r254 20 21 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=8.96 $Y=1.32
+ $X2=8.58 $Y2=1.32
r255 18 61 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.505 $Y=2.275
+ $X2=8.505 $Y2=1.905
r256 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.505 $Y=1.395
+ $X2=8.58 $Y2=1.32
r257 14 60 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.505 $Y=1.395
+ $X2=8.505 $Y2=1.575
r258 12 56 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.01 $Y=2.275
+ $X2=5.01 $Y2=1.875
r259 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.51 $Y=0.705
+ $X2=4.51 $Y2=0.87
r260 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.51 $Y=0.705
+ $X2=4.51 $Y2=0.415
r261 2 39 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r262 1 63 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_1102_21# 1 2 9 13 17 19 21 22 26 28 30 31
+ 32 35 36 41 45 49
c147 36 0 1.46668e-19 $X=5.72 $Y=1.74
r148 49 56 6.11232 $w=2.76e-07 $l=3.5e-08 $layer=POLY_cond $X=7.96 $Y=1.15
+ $X2=7.995 $Y2=1.15
r149 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.96
+ $Y=1.15 $X2=7.96 $Y2=1.15
r150 45 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.96 $Y=0.98
+ $X2=7.96 $Y2=1.15
r151 43 44 14.0202 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.845 $Y=0.695
+ $X2=6.845 $Y2=0.98
r152 36 53 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=5.682 $Y=1.74
+ $X2=5.682 $Y2=1.905
r153 36 52 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=5.682 $Y=1.74
+ $X2=5.682 $Y2=1.575
r154 35 38 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.76 $Y=1.74
+ $X2=5.76 $Y2=1.91
r155 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.72
+ $Y=1.74 $X2=5.72 $Y2=1.74
r156 33 44 2.94836 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.01 $Y=0.98
+ $X2=6.845 $Y2=0.98
r157 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=0.98
+ $X2=7.96 $Y2=0.98
r158 32 33 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.795 $Y=0.98
+ $X2=7.01 $Y2=0.98
r159 30 44 5.3975 $w=2.48e-07 $l=1.09087e-07 $layer=LI1_cond $X=6.9 $Y=1.065
+ $X2=6.845 $Y2=0.98
r160 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.9 $Y=1.065
+ $X2=6.9 $Y2=1.785
r161 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.91
+ $X2=6.47 $Y2=1.91
r162 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.815 $Y=1.91
+ $X2=6.9 $Y2=1.785
r163 28 29 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=6.815 $Y=1.91
+ $X2=6.555 $Y2=1.91
r164 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.47 $Y=2.035
+ $X2=6.47 $Y2=1.91
r165 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.47 $Y=2.035
+ $X2=6.47 $Y2=2.21
r166 23 38 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=1.91
+ $X2=5.76 $Y2=1.91
r167 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=6.47 $Y2=1.91
r168 22 23 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=5.885 $Y2=1.91
r169 19 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=0.985
+ $X2=7.995 $Y2=1.15
r170 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.995 $Y=0.985
+ $X2=7.995 $Y2=0.555
r171 15 49 30.5616 $w=2.76e-07 $l=2.43926e-07 $layer=POLY_cond $X=7.785 $Y=1.315
+ $X2=7.96 $Y2=1.15
r172 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=7.785 $Y=1.315
+ $X2=7.785 $Y2=2.065
r173 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.61 $Y=2.275
+ $X2=5.61 $Y2=1.905
r174 9 52 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=5.585 $Y=0.445
+ $X2=5.585 $Y2=1.575
r175 2 41 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.065 $X2=6.47 $Y2=1.87
r176 2 26 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.065 $X2=6.47 $Y2=2.21
r177 1 43 182 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_NDIFF $count=1 $X=6.71
+ $Y=0.235 $X2=6.845 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%SET_B 3 5 7 11 15 17 19 20 26 27 33
c130 33 0 1.34289e-19 $X=9.93 $Y=0.98
c131 15 0 1.0852e-19 $X=10.055 $Y=2.275
r132 33 36 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.962 $Y=0.98
+ $X2=9.962 $Y2=1.145
r133 33 35 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.962 $Y=0.98
+ $X2=9.962 $Y2=0.815
r134 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.035
+ $Y=0.98 $X2=6.035 $Y2=0.98
r135 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.93
+ $Y=0.98 $X2=9.93 $Y2=0.98
r136 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0.85
+ $X2=9.89 $Y2=0.85
r137 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.355 $Y=0.85
+ $X2=6.21 $Y2=0.85
r138 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.745 $Y=0.85
+ $X2=9.89 $Y2=0.85
r139 19 20 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=9.745 $Y=0.85
+ $X2=6.355 $Y2=0.85
r140 17 31 6.86495 $w=3.11e-07 $l=1.75e-07 $layer=LI1_cond $X=6.21 $Y=0.9
+ $X2=6.035 $Y2=0.9
r141 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0.85
+ $X2=6.21 $Y2=0.85
r142 15 36 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.055 $Y=2.275
+ $X2=10.055 $Y2=1.145
r143 11 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.945 $Y=0.445
+ $X2=9.945 $Y2=0.815
r144 5 30 38.6529 $w=3.37e-07 $l=2.08315e-07 $layer=POLY_cond $X=6.14 $Y=1.145
+ $X2=6.042 $Y2=0.98
r145 5 7 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.14 $Y=1.145
+ $X2=6.14 $Y2=2.275
r146 1 30 38.6529 $w=3.37e-07 $l=2.04316e-07 $layer=POLY_cond $X=6.13 $Y=0.815
+ $X2=6.042 $Y2=0.98
r147 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.13 $Y=0.815
+ $X2=6.13 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_917_47# 1 2 9 11 13 15 19 24 25 26 27 32
c113 32 0 1.42598e-19 $X=5.67 $Y=1.3
c114 27 0 1.57233e-19 $X=6.395 $Y=1.32
r115 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.56
+ $Y=1.32 $X2=6.56 $Y2=1.32
r116 31 32 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=1.3
+ $X2=5.67 $Y2=1.3
r117 29 31 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=5.38 $Y=1.3
+ $X2=5.585 $Y2=1.3
r118 27 35 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.32
+ $X2=6.56 $Y2=1.32
r119 27 32 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.395 $Y=1.32
+ $X2=5.67 $Y2=1.32
r120 26 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.585 $Y=1.195
+ $X2=5.585 $Y2=1.3
r121 25 26 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.585 $Y=0.655
+ $X2=5.585 $Y2=1.195
r122 23 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.38 $Y=1.405
+ $X2=5.38 $Y2=1.3
r123 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.38 $Y=1.405
+ $X2=5.38 $Y2=2.25
r124 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.295 $Y=2.335
+ $X2=5.38 $Y2=2.25
r125 19 21 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.295 $Y=2.335
+ $X2=4.8 $Y2=2.335
r126 15 25 20.5698 $w=1.72e-07 $l=2.93973e-07 $layer=LI1_cond $X=5.577 $Y=0.365
+ $X2=5.585 $Y2=0.655
r127 15 17 42.4227 $w=1.98e-07 $l=7.65e-07 $layer=LI1_cond $X=5.485 $Y=0.365
+ $X2=4.72 $Y2=0.365
r128 11 36 38.5481 $w=3.01e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.68 $Y=1.485
+ $X2=6.59 $Y2=1.32
r129 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.68 $Y=1.485
+ $X2=6.68 $Y2=2.065
r130 7 36 38.5481 $w=3.01e-07 $l=1.86145e-07 $layer=POLY_cond $X=6.635 $Y=1.155
+ $X2=6.59 $Y2=1.32
r131 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.635 $Y=1.155 $X2=6.635
+ $Y2=0.555
r132 2 21 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=2.065 $X2=4.8 $Y2=2.335
r133 1 17 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.235 $X2=4.72 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_1396_21# 1 2 9 13 17 21 23 24 25 27 31 34
+ 42 43 46 49 53 56 59
c161 56 0 6.74557e-20 $X=10.95 $Y=1.32
c162 53 0 1.57233e-19 $X=7.1 $Y=1.32
c163 42 0 2.58372e-20 $X=11.125 $Y=1.53
c164 27 0 1.52865e-19 $X=11.68 $Y=1.66
c165 9 0 1.18612e-19 $X=7.055 $Y=0.555
r166 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.165
+ $Y=1.32 $X2=11.165 $Y2=1.32
r167 56 58 33.5372 $w=3.09e-07 $l=2.15e-07 $layer=POLY_cond $X=10.95 $Y=1.32
+ $X2=11.165 $Y2=1.32
r168 55 56 8.57929 $w=3.09e-07 $l=5.5e-08 $layer=POLY_cond $X=10.895 $Y=1.32
+ $X2=10.95 $Y2=1.32
r169 52 53 6.97428 $w=3.11e-07 $l=4.5e-08 $layer=POLY_cond $X=7.055 $Y=1.32
+ $X2=7.1 $Y2=1.32
r170 50 59 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=11.217 $Y=1.53
+ $X2=11.217 $Y2=1.32
r171 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=1.53
+ $X2=11.27 $Y2=1.53
r172 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=1.53
+ $X2=8.05 $Y2=1.53
r173 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=1.53
+ $X2=8.05 $Y2=1.53
r174 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=1.53
+ $X2=11.27 $Y2=1.53
r175 42 43 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=1.53
+ $X2=8.195 $Y2=1.53
r176 41 50 1.88582 $w=2.73e-07 $l=4.5e-08 $layer=LI1_cond $X=11.217 $Y=1.575
+ $X2=11.217 $Y2=1.53
r177 40 59 16.5533 $w=2.73e-07 $l=3.95e-07 $layer=LI1_cond $X=11.217 $Y=0.925
+ $X2=11.217 $Y2=1.32
r178 38 46 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=7.485 $Y=1.535
+ $X2=8.05 $Y2=1.535
r179 37 38 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=1.535
+ $X2=7.485 $Y2=1.535
r180 35 53 34.0965 $w=3.11e-07 $l=2.2e-07 $layer=POLY_cond $X=7.32 $Y=1.32
+ $X2=7.1 $Y2=1.32
r181 34 37 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.32 $Y=1.32
+ $X2=7.32 $Y2=1.535
r182 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.32
+ $Y=1.32 $X2=7.32 $Y2=1.32
r183 29 31 17.1645 $w=2.08e-07 $l=3.25e-07 $layer=LI1_cond $X=11.67 $Y=0.755
+ $X2=11.67 $Y2=0.43
r184 25 41 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=11.355 $Y=1.66
+ $X2=11.217 $Y2=1.575
r185 25 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.355 $Y=1.66
+ $X2=11.68 $Y2=1.66
r186 24 40 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=11.355 $Y=0.84
+ $X2=11.217 $Y2=0.925
r187 23 29 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.67 $Y2=0.755
r188 23 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.355 $Y2=0.84
r189 19 56 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.95 $Y=1.155
+ $X2=10.95 $Y2=1.32
r190 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=10.95 $Y=1.155
+ $X2=10.95 $Y2=0.555
r191 15 55 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.895 $Y=1.485
+ $X2=10.895 $Y2=1.32
r192 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.895 $Y=1.485
+ $X2=10.895 $Y2=2.065
r193 11 53 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.1 $Y=1.485
+ $X2=7.1 $Y2=1.32
r194 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.1 $Y=1.485
+ $X2=7.1 $Y2=2.065
r195 7 52 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.055 $Y=1.155
+ $X2=7.055 $Y2=1.32
r196 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.055 $Y=1.155 $X2=7.055
+ $Y2=0.555
r197 2 27 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=11.555
+ $Y=1.505 $X2=11.68 $Y2=1.66
r198 1 31 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=11.555
+ $Y=0.235 $X2=11.68 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_1887_21# 1 2 9 13 15 17 20 22 25 27 28 30
+ 31 33 36 38 41 45 46 48 49 52 54 57 58 61 62 66 68 72 73
c181 46 0 1.29033e-19 $X=9.635 $Y=1.74
c182 20 0 1.52865e-19 $X=12.375 $Y=1.985
c183 9 0 8.93206e-20 $X=9.51 $Y=0.445
r184 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.34
+ $Y=1.16 $X2=12.34 $Y2=1.16
r185 69 72 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=12.245 $Y=1.16
+ $X2=12.34 $Y2=1.16
r186 64 66 4.61622 $w=1.83e-07 $l=7.7e-08 $layer=LI1_cond $X=10.74 $Y=0.687
+ $X2=10.817 $Y2=0.687
r187 60 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=1.325
+ $X2=12.245 $Y2=1.16
r188 60 61 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.245 $Y=1.325
+ $X2=12.245 $Y2=1.915
r189 59 68 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=10.905 $Y=2
+ $X2=10.817 $Y2=2
r190 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.16 $Y=2
+ $X2=12.245 $Y2=1.915
r191 58 59 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=12.16 $Y=2
+ $X2=10.905 $Y2=2
r192 57 68 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.817 $Y=1.915
+ $X2=10.817 $Y2=2
r193 56 66 1.08604 $w=1.75e-07 $l=9.3e-08 $layer=LI1_cond $X=10.817 $Y=0.78
+ $X2=10.817 $Y2=0.687
r194 56 57 71.9325 $w=1.73e-07 $l=1.135e-06 $layer=LI1_cond $X=10.817 $Y=0.78
+ $X2=10.817 $Y2=1.915
r195 55 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.41 $Y=2
+ $X2=10.325 $Y2=2
r196 54 68 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=10.73 $Y=2
+ $X2=10.817 $Y2=2
r197 54 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.73 $Y=2 $X2=10.41
+ $Y2=2
r198 50 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.325 $Y=2.085
+ $X2=10.325 $Y2=2
r199 50 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.325 $Y=2.085
+ $X2=10.325 $Y2=2.21
r200 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.24 $Y=2
+ $X2=10.325 $Y2=2
r201 48 49 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=10.24 $Y=2 $X2=9.8
+ $Y2=2
r202 46 77 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.602 $Y=1.74
+ $X2=9.602 $Y2=1.905
r203 46 76 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.602 $Y=1.74
+ $X2=9.602 $Y2=1.575
r204 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.635
+ $Y=1.74 $X2=9.635 $Y2=1.74
r205 43 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.675 $Y=1.915
+ $X2=9.8 $Y2=2
r206 43 45 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=9.675 $Y=1.915
+ $X2=9.675 $Y2=1.74
r207 39 41 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=13.19 $Y=1.61
+ $X2=13.315 $Y2=1.61
r208 34 36 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=13.19 $Y=0.805
+ $X2=13.315 $Y2=0.805
r209 31 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.315 $Y=1.685
+ $X2=13.315 $Y2=1.61
r210 31 33 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=13.315 $Y=1.685
+ $X2=13.315 $Y2=2.085
r211 28 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.315 $Y=0.73
+ $X2=13.315 $Y2=0.805
r212 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.315 $Y=0.73
+ $X2=13.315 $Y2=0.445
r213 27 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.19 $Y=1.535
+ $X2=13.19 $Y2=1.61
r214 26 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.19 $Y=1.295
+ $X2=13.19 $Y2=1.16
r215 26 27 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=13.19 $Y=1.295
+ $X2=13.19 $Y2=1.535
r216 25 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.19 $Y=1.025
+ $X2=13.19 $Y2=1.16
r217 24 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.19 $Y=0.88
+ $X2=13.19 $Y2=0.805
r218 24 25 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=13.19 $Y=0.88
+ $X2=13.19 $Y2=1.025
r219 23 73 2.60871 $w=2.7e-07 $l=1.23e-07 $layer=POLY_cond $X=12.45 $Y=1.16
+ $X2=12.327 $Y2=1.16
r220 22 38 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=13.115 $Y=1.16
+ $X2=13.19 $Y2=1.16
r221 22 23 147.746 $w=2.7e-07 $l=6.65e-07 $layer=POLY_cond $X=13.115 $Y=1.16
+ $X2=12.45 $Y2=1.16
r222 18 73 32.2453 $w=1.5e-07 $l=1.8747e-07 $layer=POLY_cond $X=12.375 $Y=1.325
+ $X2=12.327 $Y2=1.16
r223 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.375 $Y=1.325
+ $X2=12.375 $Y2=1.985
r224 15 73 32.2453 $w=1.5e-07 $l=1.8747e-07 $layer=POLY_cond $X=12.375 $Y=0.995
+ $X2=12.327 $Y2=1.16
r225 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.375 $Y=0.995
+ $X2=12.375 $Y2=0.56
r226 13 77 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.515 $Y=2.275
+ $X2=9.515 $Y2=1.905
r227 9 76 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=9.51 $Y=0.445
+ $X2=9.51 $Y2=1.575
r228 2 52 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.065 $X2=10.325 $Y2=2.21
r229 1 64 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=10.605
+ $Y=0.235 $X2=10.74 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_1714_47# 1 2 9 13 15 19 24 26 27 29 31 32
c99 32 0 2.58372e-20 $X=10.475 $Y=1.24
c100 31 0 1.75976e-19 $X=10.475 $Y=1.24
c101 26 0 3.84972e-20 $X=9.295 $Y=2.25
r102 32 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.475 $Y=1.24
+ $X2=10.475 $Y2=1.405
r103 32 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.475 $Y=1.24
+ $X2=10.475 $Y2=1.075
r104 31 34 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=10.45 $Y=1.24
+ $X2=10.45 $Y2=1.32
r105 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.475
+ $Y=1.24 $X2=10.475 $Y2=1.24
r106 28 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=1.32
+ $X2=9.295 $Y2=1.32
r107 27 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=10.34 $Y=1.32
+ $X2=10.45 $Y2=1.32
r108 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.34 $Y=1.32
+ $X2=9.38 $Y2=1.32
r109 25 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.405
+ $X2=9.295 $Y2=1.32
r110 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.295 $Y=1.405
+ $X2=9.295 $Y2=2.25
r111 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.235
+ $X2=9.295 $Y2=1.32
r112 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=9.295 $Y=0.465
+ $X2=9.295 $Y2=1.235
r113 19 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.21 $Y=0.365
+ $X2=9.295 $Y2=0.465
r114 19 21 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=9.21 $Y=0.365
+ $X2=8.78 $Y2=0.365
r115 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.21 $Y=2.335
+ $X2=9.295 $Y2=2.25
r116 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.21 $Y=2.335
+ $X2=8.715 $Y2=2.335
r117 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.535 $Y=2.065
+ $X2=10.535 $Y2=1.405
r118 9 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=10.53 $Y=0.555
+ $X2=10.53 $Y2=1.075
r119 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=8.58
+ $Y=2.065 $X2=8.715 $Y2=2.335
r120 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.57
+ $Y=0.235 $X2=8.78 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%RESET_B 3 7 9 15
r36 12 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=11.7 $Y=1.18
+ $X2=11.89 $Y2=1.18
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.7
+ $Y=1.18 $X2=11.7 $Y2=1.18
r38 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.89 $Y=1.345
+ $X2=11.89 $Y2=1.18
r39 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.89 $Y=1.345
+ $X2=11.89 $Y2=1.825
r40 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.89 $Y=1.015
+ $X2=11.89 $Y2=1.18
r41 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=11.89 $Y=1.015
+ $X2=11.89 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_2596_47# 1 2 9 12 16 20 24 25 27 29
c52 27 0 1.41074e-19 $X=13.117 $Y=1.16
r53 25 30 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=13.72 $Y=1.16
+ $X2=13.72 $Y2=1.325
r54 25 29 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=13.72 $Y=1.16
+ $X2=13.72 $Y2=0.995
r55 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.71
+ $Y=1.16 $X2=13.71 $Y2=1.16
r56 22 27 1.17559 $w=3.3e-07 $l=1.58e-07 $layer=LI1_cond $X=13.275 $Y=1.16
+ $X2=13.117 $Y2=1.16
r57 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=13.275 $Y=1.16
+ $X2=13.71 $Y2=1.16
r58 18 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=13.117 $Y=1.325
+ $X2=13.117 $Y2=1.16
r59 18 20 21.4025 $w=3.13e-07 $l=5.85e-07 $layer=LI1_cond $X=13.117 $Y=1.325
+ $X2=13.117 $Y2=1.91
r60 14 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=13.117 $Y=0.995
+ $X2=13.117 $Y2=1.16
r61 14 16 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=13.117 $Y=0.995
+ $X2=13.117 $Y2=0.51
r62 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.79 $Y=1.985
+ $X2=13.79 $Y2=1.325
r63 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.79 $Y=0.56
+ $X2=13.79 $Y2=0.995
r64 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.98
+ $Y=1.765 $X2=13.105 $Y2=1.91
r65 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=12.98
+ $Y=0.235 $X2=13.105 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 53
+ 54 55 59 60 62 64 70 75 83 95 106 110 117 118 121 124 127 130 133 144 146
c207 118 0 2.75701e-19 $X=14.03 $Y=2.72
r208 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r209 142 144 9.28831 $w=5.48e-07 $l=1.4e-07 $layer=LI1_cond $X=12.19 $Y=2.53
+ $X2=12.33 $Y2=2.53
r210 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r211 140 142 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=12.165 $Y=2.53
+ $X2=12.19 $Y2=2.53
r212 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r213 133 136 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=9.81 $Y=2.34
+ $X2=9.81 $Y2=2.72
r214 130 131 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r215 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r216 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r217 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r218 118 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=13.57 $Y2=2.72
r219 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r220 115 146 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=13.74 $Y=2.72
+ $X2=13.597 $Y2=2.72
r221 115 117 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.74 $Y=2.72
+ $X2=14.03 $Y2=2.72
r222 114 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r223 114 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=12.19 $Y2=2.72
r224 113 144 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.11 $Y=2.72
+ $X2=12.33 $Y2=2.72
r225 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r226 110 146 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=13.455 $Y=2.72
+ $X2=13.597 $Y2=2.72
r227 110 113 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.455 $Y=2.72
+ $X2=13.11 $Y2=2.72
r228 109 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r229 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r230 106 140 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=12.055 $Y=2.53
+ $X2=12.165 $Y2=2.53
r231 106 108 17.0713 $w=5.48e-07 $l=7.85e-07 $layer=LI1_cond $X=12.055 $Y=2.53
+ $X2=11.27 $Y2=2.53
r232 105 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r233 105 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=9.89 $Y2=2.72
r234 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r235 102 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10 $Y=2.72
+ $X2=9.81 $Y2=2.72
r236 102 104 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=10 $Y=2.72
+ $X2=10.81 $Y2=2.72
r237 101 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r238 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r239 98 101 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r240 97 100 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r241 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r242 95 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.81 $Y2=2.72
r243 95 100 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.43 $Y2=2.72
r244 94 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r245 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r246 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r247 91 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r248 90 93 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r249 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r250 88 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=5.895 $Y2=2.72
r251 88 90 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=6.21 $Y2=2.72
r252 87 131 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r253 87 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r254 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r255 84 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=2.72
+ $X2=3.475 $Y2=2.72
r256 84 86 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.64 $Y=2.72
+ $X2=3.91 $Y2=2.72
r257 83 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=5.895 $Y2=2.72
r258 83 86 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=3.91 $Y2=2.72
r259 82 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r260 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r261 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r262 79 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r263 78 81 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r264 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r265 76 124 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.607 $Y2=2.72
r266 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r267 75 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=3.475 $Y2=2.72
r268 75 81 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=2.99 $Y2=2.72
r269 74 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r270 74 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r271 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r272 71 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r273 71 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r274 70 124 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.607 $Y2=2.72
r275 70 73 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.15 $Y2=2.72
r276 64 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r277 62 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r278 60 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r279 60 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r280 59 104 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=10.94 $Y=2.72
+ $X2=10.81 $Y2=2.72
r281 58 59 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.105 $Y=2.53
+ $X2=10.94 $Y2=2.53
r282 55 108 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=11.215 $Y=2.53
+ $X2=11.27 $Y2=2.53
r283 55 58 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=11.215 $Y=2.53
+ $X2=11.105 $Y2=2.53
r284 53 93 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.13 $Y2=2.72
r285 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.34 $Y2=2.72
r286 52 97 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.59 $Y2=2.72
r287 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.34 $Y2=2.72
r288 48 146 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=13.597 $Y=2.635
+ $X2=13.597 $Y2=2.72
r289 48 50 28.1034 $w=2.83e-07 $l=6.95e-07 $layer=LI1_cond $X=13.597 $Y=2.635
+ $X2=13.597 $Y2=1.94
r290 44 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=2.635
+ $X2=7.34 $Y2=2.72
r291 44 46 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.34 $Y=2.635
+ $X2=7.34 $Y2=2
r292 40 130 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.895 $Y=2.635
+ $X2=5.895 $Y2=2.72
r293 40 42 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=5.895 $Y=2.635
+ $X2=5.895 $Y2=2.29
r294 36 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=2.635
+ $X2=3.475 $Y2=2.72
r295 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.475 $Y=2.635
+ $X2=3.475 $Y2=2.3
r296 32 124 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.72
r297 32 34 21.588 $w=3.53e-07 $l=6.65e-07 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=1.97
r298 28 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r299 28 30 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r300 9 50 300 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=2 $X=13.39
+ $Y=1.765 $X2=13.575 $Y2=1.94
r301 8 140 600 $w=1.7e-07 $l=9.29637e-07 $layer=licon1_PDIFF $count=1 $X=11.965
+ $Y=1.505 $X2=12.165 $Y2=2.34
r302 7 58 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=10.97
+ $Y=1.645 $X2=11.105 $Y2=2.34
r303 6 133 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=9.59
+ $Y=2.065 $X2=9.785 $Y2=2.34
r304 5 46 300 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_PDIFF $count=2 $X=7.175
+ $Y=1.645 $X2=7.34 $Y2=2
r305 4 42 600 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=2.065 $X2=5.87 $Y2=2.29
r306 3 38 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.065 $X2=3.475 $Y2=2.3
r307 2 34 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.815 $X2=1.62 $Y2=1.97
r308 1 30 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_453_47# 1 2 3 4 13 16 18 22 23 28 32 36
+ 37 39 40 43 46 47
c140 47 0 1.01009e-19 $X=4.315 $Y=1.19
c141 46 0 9.78226e-20 $X=4.315 $Y=1.19
c142 43 0 8.91744e-20 $X=2.99 $Y=1.19
c143 40 0 8.49446e-20 $X=3.135 $Y=1.19
c144 23 0 1.50346e-19 $X=2.395 $Y=1.875
c145 16 0 1.68616e-20 $X=2.57 $Y=1.075
r146 47 53 2.87435 $w=1.91e-07 $l=4.5e-08 $layer=LI1_cond $X=4.315 $Y=1.185
+ $X2=4.36 $Y2=1.185
r147 47 51 17.8848 $w=1.91e-07 $l=2.8e-07 $layer=LI1_cond $X=4.315 $Y=1.185
+ $X2=4.035 $Y2=1.185
r148 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.315 $Y=1.19
+ $X2=4.315 $Y2=1.19
r149 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.19
+ $X2=2.99 $Y2=1.19
r150 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.19
+ $X2=2.99 $Y2=1.19
r151 39 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.17 $Y=1.19
+ $X2=4.315 $Y2=1.19
r152 39 40 1.28094 $w=1.4e-07 $l=1.035e-06 $layer=MET1_cond $X=4.17 $Y=1.19
+ $X2=3.135 $Y2=1.19
r153 36 37 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.337 $Y=2.3
+ $X2=4.337 $Y2=2.135
r154 32 34 10.6307 $w=2.41e-07 $l=2.1e-07 $layer=LI1_cond $X=4.035 $Y=0.43
+ $X2=4.245 $Y2=0.43
r155 31 43 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.67 $Y=1.24
+ $X2=2.99 $Y2=1.24
r156 26 28 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.435 $Y=0.43
+ $X2=2.57 $Y2=0.43
r157 22 23 5.95004 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=1.96
+ $X2=2.395 $Y2=1.875
r158 19 53 1.41722 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.36 $Y=1.305
+ $X2=4.36 $Y2=1.185
r159 19 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.36 $Y=1.305
+ $X2=4.36 $Y2=2.135
r160 18 51 1.41722 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=1.185
r161 17 32 2.78154 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=0.595
+ $X2=4.035 $Y2=0.43
r162 17 18 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.035 $Y=0.595
+ $X2=4.035 $Y2=1.065
r163 16 31 9.88216 $w=2.17e-07 $l=1.80748e-07 $layer=LI1_cond $X=2.57 $Y=1.075
+ $X2=2.537 $Y2=1.24
r164 15 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0.595
+ $X2=2.57 $Y2=0.43
r165 15 16 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.57 $Y=0.595
+ $X2=2.57 $Y2=1.075
r166 13 31 15.5043 $w=2.17e-07 $l=2.87541e-07 $layer=LI1_cond $X=2.49 $Y=1.505
+ $X2=2.537 $Y2=1.24
r167 13 23 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.49 $Y=1.505
+ $X2=2.49 $Y2=1.875
r168 4 36 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=2.065 $X2=4.315 $Y2=2.3
r169 3 22 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.815 $X2=2.4 $Y2=1.96
r170 2 34 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=4.11
+ $Y=0.235 $X2=4.245 $Y2=0.43
r171 1 26 182 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.435 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%Q_N 1 2 9 10 11 12 13 18 21
r30 18 21 2.69684 $w=2.85e-07 $l=6.3e-08 $layer=LI1_cond $X=12.642 $Y=0.573
+ $X2=12.642 $Y2=0.51
r31 12 13 15.9725 $w=2.83e-07 $l=3.95e-07 $layer=LI1_cond $X=12.642 $Y=1.815
+ $X2=12.642 $Y2=2.21
r32 11 30 6.85431 $w=2.83e-07 $l=1.31e-07 $layer=LI1_cond $X=12.642 $Y=0.584
+ $X2=12.642 $Y2=0.715
r33 11 18 0.444803 $w=2.83e-07 $l=1.1e-08 $layer=LI1_cond $X=12.642 $Y=0.584
+ $X2=12.642 $Y2=0.573
r34 11 21 0.470877 $w=2.85e-07 $l=1.1e-08 $layer=LI1_cond $X=12.642 $Y=0.499
+ $X2=12.642 $Y2=0.51
r35 10 30 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=12.695 $Y=1.63
+ $X2=12.695 $Y2=0.715
r36 9 12 1.73877 $w=2.83e-07 $l=4.3e-08 $layer=LI1_cond $X=12.642 $Y=1.772
+ $X2=12.642 $Y2=1.815
r37 9 10 7.29911 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=12.642 $Y=1.772
+ $X2=12.642 $Y2=1.63
r38 2 12 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=12.45
+ $Y=1.485 $X2=12.585 $Y2=1.815
r39 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=12.45
+ $Y=0.235 $X2=12.585 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%Q 1 2 10 11 12 13 14 15
r16 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=14.045 $Y=1.82
+ $X2=14.045 $Y2=2.21
r17 11 14 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=14.045 $Y=1.6
+ $X2=14.045 $Y2=1.82
r18 11 12 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=14.045 $Y=1.6
+ $X2=14.045 $Y2=1.47
r19 10 12 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=14.07 $Y=0.785
+ $X2=14.07 $Y2=1.47
r20 9 13 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=14.045 $Y=0.655
+ $X2=14.045 $Y2=0.51
r21 9 10 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=14.045 $Y=0.655
+ $X2=14.045 $Y2=0.785
r22 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=13.865
+ $Y=1.485 $X2=14 $Y2=1.82
r23 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=13.865
+ $Y=0.235 $X2=14 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 66 68 70 76 81 108 115 122 123 126 129 132 135 138
c218 123 0 2.71124e-20 $X=14.03 $Y=0
c219 47 0 1.34289e-19 $X=9.735 $Y=0.36
r220 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r221 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r222 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r223 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r224 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r225 123 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=13.57 $Y2=0
r226 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r227 120 138 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.745 $Y=0
+ $X2=13.6 $Y2=0
r228 120 122 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.745 $Y=0
+ $X2=14.03 $Y2=0
r229 119 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r230 119 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=12.19 $Y2=0
r231 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r232 116 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.33 $Y=0
+ $X2=12.165 $Y2=0
r233 116 118 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=12.33 $Y=0
+ $X2=13.11 $Y2=0
r234 115 138 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.6 $Y2=0
r235 115 118 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.11 $Y2=0
r236 114 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r237 113 114 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r238 111 114 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r239 110 113 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r240 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r241 108 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12 $Y=0
+ $X2=12.165 $Y2=0
r242 108 113 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12 $Y=0 $X2=11.73
+ $Y2=0
r243 107 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r244 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r245 104 107 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.43 $Y2=0
r246 103 106 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=9.43 $Y2=0
r247 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r248 101 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r249 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r250 98 101 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r251 97 100 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r252 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r253 95 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r254 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r255 92 95 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r256 92 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=3.45 $Y2=0
r257 91 94 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.75
+ $Y2=0
r258 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r259 89 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.39 $Y2=0
r260 89 91 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.91 $Y2=0
r261 88 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.45 $Y2=0
r262 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r263 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r264 85 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r265 84 87 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r266 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r267 82 129 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=1.567 $Y2=0
r268 82 84 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r269 81 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=0
+ $X2=3.39 $Y2=0
r270 81 87 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.225 $Y=0
+ $X2=2.99 $Y2=0
r271 80 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r272 80 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r273 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r274 77 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r275 77 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r276 76 129 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.43 $Y=0
+ $X2=1.567 $Y2=0
r277 76 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.15
+ $Y2=0
r278 70 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r279 68 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r280 66 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r281 66 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r282 64 106 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=9.56 $Y=0 $X2=9.43
+ $Y2=0
r283 64 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.56 $Y=0 $X2=9.69
+ $Y2=0
r284 63 110 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=9.82 $Y=0 $X2=9.89
+ $Y2=0
r285 63 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.82 $Y=0 $X2=9.69
+ $Y2=0
r286 61 100 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.59
+ $Y2=0
r287 61 62 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.797
+ $Y2=0
r288 60 103 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.975 $Y=0
+ $X2=8.05 $Y2=0
r289 60 62 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=7.975 $Y=0
+ $X2=7.797 $Y2=0
r290 58 94 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.75
+ $Y2=0
r291 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.92
+ $Y2=0
r292 57 97 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.005 $Y=0
+ $X2=6.21 $Y2=0
r293 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0 $X2=5.92
+ $Y2=0
r294 53 138 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=13.6 $Y=0.085
+ $X2=13.6 $Y2=0
r295 53 55 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=13.6 $Y=0.085
+ $X2=13.6 $Y2=0.38
r296 49 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.165 $Y=0.085
+ $X2=12.165 $Y2=0
r297 49 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.165 $Y=0.085
+ $X2=12.165 $Y2=0.38
r298 45 65 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=0.085
+ $X2=9.69 $Y2=0
r299 45 47 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=9.69 $Y=0.085
+ $X2=9.69 $Y2=0.36
r300 41 62 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.797 $Y=0.085
+ $X2=7.797 $Y2=0
r301 41 43 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=7.797 $Y=0.085
+ $X2=7.797 $Y2=0.38
r302 37 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r303 37 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.36
r304 33 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0
r305 33 35 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0.36
r306 29 129 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.567 $Y=0.085
+ $X2=1.567 $Y2=0
r307 29 31 16.1342 $w=2.73e-07 $l=3.85e-07 $layer=LI1_cond $X=1.567 $Y=0.085
+ $X2=1.567 $Y2=0.47
r308 25 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r309 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r310 8 55 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=13.39
+ $Y=0.235 $X2=13.58 $Y2=0.38
r311 7 51 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=11.965
+ $Y=0.235 $X2=12.165 $Y2=0.38
r312 6 47 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=9.585
+ $Y=0.235 $X2=9.735 $Y2=0.36
r313 5 43 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.66
+ $Y=0.235 $X2=7.785 $Y2=0.38
r314 4 39 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=5.66
+ $Y=0.235 $X2=5.92 $Y2=0.36
r315 3 35 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.235 $X2=3.39 $Y2=0.36
r316 2 31 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.47
r317 1 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_1241_47# 1 2 7 11 16
c25 16 0 1.18612e-19 $X=6.59 $Y=0.36
r26 14 16 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=0.36
+ $X2=6.59 $Y2=0.36
r27 9 11 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=0.425
+ $X2=7.265 $Y2=0.55
r28 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.18 $Y=0.34
+ $X2=7.265 $Y2=0.425
r29 7 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.18 $Y=0.34 $X2=6.59
+ $Y2=0.34
r30 2 11 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.235 $X2=7.265 $Y2=0.55
r31 1 14 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=6.205
+ $Y=0.235 $X2=6.425 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_1%A_2004_47# 1 2 7 9
r20 9 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=10.245 $Y=0.34
+ $X2=10.245 $Y2=0.46
r21 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.41 $Y=0.34
+ $X2=10.245 $Y2=0.34
r22 7 8 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=11.075 $Y=0.34
+ $X2=10.41 $Y2=0.34
r23 2 7 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=11.025
+ $Y=0.235 $X2=11.16 $Y2=0.42
r24 1 12 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=10.02
+ $Y=0.235 $X2=10.245 $Y2=0.46
.ends


* File: sky130_fd_sc_hd__a32oi_2.pex.spice
* Created: Thu Aug 27 14:05:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A32OI_2%B2 1 3 6 8 10 13 15 16 17 26 28
c50 17 0 1.6358e-19 $X=0.695 $Y=1.19
r51 24 26 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.66 $Y=1.16
+ $X2=0.89 $Y2=1.16
r52 21 24 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.66 $Y2=1.16
r53 17 32 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=0.66 $Y=1.18
+ $X2=0.325 $Y2=1.18
r54 17 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.66
+ $Y=1.16 $X2=0.66 $Y2=1.16
r55 16 28 15.096 $w=1.78e-07 $l=2.45e-07 $layer=LI1_cond $X=0.235 $Y=1.53
+ $X2=0.235 $Y2=1.285
r56 15 28 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.235 $Y2=1.285
r57 15 32 3.17035 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=0.235 $Y=1.18 $X2=0.325
+ $Y2=1.18
r58 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r59 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r60 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r61 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r62 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r63 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r64 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r65 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%B1 1 3 6 8 10 13 15 16 24
c43 24 0 1.6358e-19 $X=1.73 $Y=1.135
c44 16 0 1.96155e-19 $X=1.615 $Y=1.19
r45 22 24 70.327 $w=3.2e-07 $l=3.9e-07 $layer=POLY_cond $X=1.34 $Y=1.135
+ $X2=1.73 $Y2=1.135
r46 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.16 $X2=1.34 $Y2=1.16
r47 19 22 5.40977 $w=3.2e-07 $l=3e-08 $layer=POLY_cond $X=1.31 $Y=1.135 $X2=1.34
+ $Y2=1.135
r48 16 23 16.2077 $w=2.07e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=1.34 $Y2=1.18
r49 15 23 10.9034 $w=2.07e-07 $l=1.85e-07 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=1.34 $Y2=1.18
r50 11 24 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.135
r51 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r52 8 24 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.73 $Y=0.975
+ $X2=1.73 $Y2=1.135
r53 8 10 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.73 $Y=0.975
+ $X2=1.73 $Y2=0.56
r54 4 19 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.135
r55 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295 $X2=1.31
+ $Y2=1.985
r56 1 19 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.31 $Y=0.975
+ $X2=1.31 $Y2=1.135
r57 1 3 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.31 $Y=0.975
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A1 3 5 6 9 13 17 19 21 30 31
c52 31 0 3.25977e-19 $X=3.145 $Y=1.16
c53 6 0 3.24478e-19 $X=2.225 $Y=1.16
r54 29 31 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=3.055 $Y=1.16
+ $X2=3.145 $Y2=1.16
r55 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.055
+ $Y=1.16 $X2=3.055 $Y2=1.16
r56 27 29 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.725 $Y=1.16
+ $X2=3.055 $Y2=1.16
r57 21 30 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=2.995 $Y=1.35
+ $X2=3.055 $Y2=1.35
r58 19 21 10.0036 $w=5.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.35
+ $X2=2.995 $Y2=1.35
r59 15 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.145 $Y=1.025
+ $X2=3.145 $Y2=1.16
r60 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.145 $Y=1.025
+ $X2=3.145 $Y2=0.56
r61 11 29 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.055 $Y=1.295
+ $X2=3.055 $Y2=1.16
r62 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.055 $Y=1.295
+ $X2=3.055 $Y2=1.985
r63 7 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.725 $Y=1.025
+ $X2=2.725 $Y2=1.16
r64 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.725 $Y=1.025
+ $X2=2.725 $Y2=0.56
r65 5 27 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=1.16 $X2=2.725
+ $Y2=1.16
r66 5 6 94.4238 $w=2.7e-07 $l=4.25e-07 $layer=POLY_cond $X=2.65 $Y=1.16
+ $X2=2.225 $Y2=1.16
r67 1 6 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.225 $Y2=1.16
r68 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295 $X2=2.15
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A2 3 7 11 15 17 19 29
c48 19 0 1.82667e-19 $X=4.375 $Y=1.53
r49 29 31 6.27138 $w=2.69e-07 $l=3.5e-08 $layer=POLY_cond $X=4.23 $Y=1.16
+ $X2=4.265 $Y2=1.16
r50 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.23
+ $Y=1.16 $X2=4.23 $Y2=1.16
r51 27 29 42.1078 $w=2.69e-07 $l=2.35e-07 $layer=POLY_cond $X=3.995 $Y=1.16
+ $X2=4.23 $Y2=1.16
r52 26 27 75.2565 $w=2.69e-07 $l=4.2e-07 $layer=POLY_cond $X=3.575 $Y=1.16
+ $X2=3.995 $Y2=1.16
r53 25 26 12.5428 $w=2.69e-07 $l=7e-08 $layer=POLY_cond $X=3.505 $Y=1.16
+ $X2=3.575 $Y2=1.16
r54 19 30 3.1533 $w=5.48e-07 $l=1.45e-07 $layer=LI1_cond $X=4.375 $Y=1.35
+ $X2=4.23 $Y2=1.35
r55 17 30 6.85027 $w=5.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=1.35
+ $X2=4.23 $Y2=1.35
r56 13 31 16.4183 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.265 $Y=1.295
+ $X2=4.265 $Y2=1.16
r57 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.265 $Y=1.295
+ $X2=4.265 $Y2=1.985
r58 9 27 16.4183 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.995 $Y=1.025
+ $X2=3.995 $Y2=1.16
r59 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.995 $Y=1.025
+ $X2=3.995 $Y2=0.56
r60 5 26 16.4183 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.575 $Y=1.025
+ $X2=3.575 $Y2=1.16
r61 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.575 $Y=1.025
+ $X2=3.575 $Y2=0.56
r62 1 25 16.4183 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.505 $Y=1.295
+ $X2=3.505 $Y2=1.16
r63 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.505 $Y=1.295
+ $X2=3.505 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A3 3 7 11 15 17 21 23 25 33 39
r46 37 39 38.2675 $w=2.9e-07 $l=1.85e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.695 $Y2=1.16
r47 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.355
+ $Y=1.16 $X2=5.355 $Y2=1.16
r48 33 37 15.8876 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=5.435 $Y=1.16
+ $X2=5.51 $Y2=1.16
r49 33 35 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=5.435 $Y=1.16
+ $X2=5.355 $Y2=1.16
r50 25 36 7.39394 $w=5.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.695 $Y=1.35
+ $X2=5.355 $Y2=1.35
r51 25 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.695
+ $Y=1.16 $X2=5.695 $Y2=1.16
r52 23 36 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=5.295 $Y=1.35
+ $X2=5.355 $Y2=1.35
r53 21 23 10.0036 $w=5.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.835 $Y=1.35
+ $X2=5.295 $Y2=1.35
r54 18 20 66.6521 $w=2.7e-07 $l=3e-07 $layer=POLY_cond $X=4.69 $Y=1.16 $X2=4.99
+ $Y2=1.16
r55 17 35 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=5.065 $Y=1.16
+ $X2=5.355 $Y2=1.16
r56 17 20 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.065 $Y=1.16
+ $X2=4.99 $Y2=1.16
r57 13 37 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.51 $Y=1.305
+ $X2=5.51 $Y2=1.16
r58 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.51 $Y=1.305
+ $X2=5.51 $Y2=1.985
r59 9 37 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.51 $Y=1.015
+ $X2=5.51 $Y2=1.16
r60 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.51 $Y=1.015
+ $X2=5.51 $Y2=0.56
r61 5 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.99 $Y=1.025
+ $X2=4.99 $Y2=1.16
r62 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.99 $Y=1.025
+ $X2=4.99 $Y2=0.56
r63 1 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.69 $Y=1.295
+ $X2=4.69 $Y2=1.16
r64 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.69 $Y=1.295 $X2=4.69
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A_27_297# 1 2 3 4 5 6 21 23 24 27 29 31 32
+ 33 37 39 43 45 47 49 51 57 59
c79 57 0 1.4331e-19 $X=3.265 $Y=1.96
r80 47 61 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.72 $Y=2.085
+ $X2=5.72 $Y2=1.94
r81 47 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.72 $Y=2.085
+ $X2=5.72 $Y2=2.3
r82 46 59 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.56 $Y=2
+ $X2=4.475 $Y2=1.94
r83 45 61 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.635 $Y=2
+ $X2=5.72 $Y2=1.94
r84 45 46 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=5.635 $Y=2
+ $X2=4.56 $Y2=2
r85 41 59 1.34256 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.475 $Y=2.085
+ $X2=4.475 $Y2=1.94
r86 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.475 $Y=2.085
+ $X2=4.475 $Y2=2.3
r87 40 57 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.35 $Y=2
+ $X2=3.265 $Y2=1.94
r88 39 59 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.39 $Y=2
+ $X2=4.475 $Y2=1.94
r89 39 40 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.39 $Y=2 $X2=3.35
+ $Y2=2
r90 35 57 1.34256 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=2.085
+ $X2=3.265 $Y2=1.94
r91 35 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.265 $Y=2.085
+ $X2=3.265 $Y2=2.3
r92 34 53 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.025 $Y=2
+ $X2=1.94 $Y2=1.94
r93 33 57 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.18 $Y=2
+ $X2=3.265 $Y2=1.94
r94 33 34 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=3.18 $Y=2
+ $X2=2.025 $Y2=2
r95 32 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=2.38
r96 31 53 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.94 $Y=2.085
+ $X2=1.94 $Y2=1.94
r97 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.94 $Y=2.085
+ $X2=1.94 $Y2=2.295
r98 30 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.38 $X2=1.1
+ $Y2=2.38
r99 29 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.38
+ $X2=1.94 $Y2=2.38
r100 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=2.38
+ $X2=1.185 $Y2=2.38
r101 25 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.295 $X2=1.1
+ $Y2=2.38
r102 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=2.295
+ $X2=1.1 $Y2=1.96
r103 23 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.38
+ $X2=1.1 $Y2=2.38
r104 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=2.38
+ $X2=0.345 $Y2=2.38
r105 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.345 $Y2=2.38
r106 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.96
r107 6 61 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=1.96
r108 6 49 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=2.3
r109 5 59 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.485 $X2=4.475 $Y2=1.96
r110 5 43 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.485 $X2=4.475 $Y2=2.3
r111 4 57 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.485 $X2=3.265 $Y2=1.96
r112 4 37 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.485 $X2=3.265 $Y2=2.3
r113 3 55 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.3
r114 3 53 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r115 2 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r116 1 21 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%Y 1 2 3 4 17 18 19 25 27 31 34 36 37 38 39
+ 46 48
r76 45 48 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.072 $Y=0.825
+ $X2=2.072 $Y2=0.85
r77 39 46 3.07165 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.072 $Y=1.54
+ $X2=2.072 $Y2=1.455
r78 39 46 0.26801 $w=2.13e-07 $l=5e-09 $layer=LI1_cond $X=2.072 $Y=1.45
+ $X2=2.072 $Y2=1.455
r79 38 39 13.9365 $w=2.13e-07 $l=2.6e-07 $layer=LI1_cond $X=2.072 $Y=1.19
+ $X2=2.072 $Y2=1.45
r80 37 45 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.072 $Y=0.74
+ $X2=2.072 $Y2=0.825
r81 37 38 16.6166 $w=2.13e-07 $l=3.1e-07 $layer=LI1_cond $X=2.072 $Y=0.88
+ $X2=2.072 $Y2=1.19
r82 37 48 1.60806 $w=2.13e-07 $l=3e-08 $layer=LI1_cond $X=2.072 $Y=0.88
+ $X2=2.072 $Y2=0.85
r83 29 37 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.18 $Y=0.74
+ $X2=2.072 $Y2=0.74
r84 29 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.18 $Y=0.74
+ $X2=2.935 $Y2=0.74
r85 28 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.54
+ $X2=1.52 $Y2=1.54
r86 27 39 3.86667 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.965 $Y=1.54
+ $X2=2.072 $Y2=1.54
r87 27 28 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.965 $Y=1.54
+ $X2=1.605 $Y2=1.54
r88 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.625
+ $X2=1.52 $Y2=1.54
r89 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=1.625
+ $X2=1.52 $Y2=1.96
r90 19 37 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.965 $Y=0.74
+ $X2=2.072 $Y2=0.74
r91 19 21 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.965 $Y=0.74
+ $X2=1.52 $Y2=0.74
r92 17 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=1.54
+ $X2=1.52 $Y2=1.54
r93 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=1.54
+ $X2=0.765 $Y2=1.54
r94 14 34 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.955
+ $X2=0.68 $Y2=2.04
r95 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.68 $Y=1.955
+ $X2=0.68 $Y2=1.7
r96 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=1.625
+ $X2=0.765 $Y2=1.54
r97 13 16 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.68 $Y=1.625
+ $X2=0.68 $Y2=1.7
r98 4 25 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r99 3 34 600 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.04
r100 3 16 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.7
r101 2 31 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.935 $Y2=0.74
r102 1 21 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%VPWR 1 2 3 12 29 30 35 38 42 45 49 55
r81 53 55 9.39704 $w=5.48e-07 $l=1.45e-07 $layer=LI1_cond $X=5.29 $Y=2.53
+ $X2=5.435 $Y2=2.53
r82 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r83 51 53 0.434938 $w=5.48e-07 $l=2e-08 $layer=LI1_cond $X=5.27 $Y=2.53 $X2=5.29
+ $Y2=2.53
r84 48 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r85 47 51 9.56863 $w=5.48e-07 $l=4.4e-07 $layer=LI1_cond $X=4.83 $Y=2.53
+ $X2=5.27 $Y2=2.53
r86 47 49 7.65729 $w=5.48e-07 $l=6.5e-08 $layer=LI1_cond $X=4.83 $Y=2.53
+ $X2=4.765 $Y2=2.53
r87 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r88 45 49 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.22 $Y=2.72
+ $X2=4.765 $Y2=2.72
r89 44 45 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=2.53
+ $X2=4.22 $Y2=2.53
r90 41 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r91 40 44 3.1533 $w=5.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=4.055 $Y2=2.53
r92 40 42 14.0726 $w=5.48e-07 $l=3.6e-07 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=3.55 $Y2=2.53
r93 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r94 37 38 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=2.53
+ $X2=2.94 $Y2=2.53
r95 33 37 5.32799 $w=5.48e-07 $l=2.45e-07 $layer=LI1_cond $X=2.53 $Y=2.53
+ $X2=2.775 $Y2=2.53
r96 33 35 11.8979 $w=5.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.53 $Y=2.53
+ $X2=2.27 $Y2=2.53
r97 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 30 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r99 29 55 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=5.435 $Y2=2.72
r100 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 26 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r102 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 25 42 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.45 $Y=2.72 $X2=3.55
+ $Y2=2.72
r104 25 38 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=2.94 $Y2=2.72
r105 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r106 21 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 20 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.07 $Y=2.72 $X2=2.27
+ $Y2=2.72
r108 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 16 20 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 12 21 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r111 12 16 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r112 3 51 300 $w=1.7e-07 $l=1.07833e-06 $layer=licon1_PDIFF $count=2 $X=4.765
+ $Y=1.485 $X2=5.27 $Y2=2.34
r113 2 44 300 $w=1.7e-07 $l=1.06637e-06 $layer=licon1_PDIFF $count=2 $X=3.58
+ $Y=1.485 $X2=4.055 $Y2=2.34
r114 1 37 300 $w=1.7e-07 $l=1.09603e-06 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.775 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A_27_47# 1 2 3 11 12 14 15 18 21
c43 18 0 1.28323e-19 $X=1.94 $Y=0.38
r44 16 26 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.185 $Y=0.38
+ $X2=1.06 $Y2=0.38
r45 16 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.185 $Y=0.38
+ $X2=1.94 $Y2=0.38
r46 15 28 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.715 $X2=1.1
+ $Y2=0.8
r47 14 26 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.1 $Y=0.465
+ $X2=1.06 $Y2=0.38
r48 14 15 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.1 $Y=0.465 $X2=1.1
+ $Y2=0.715
r49 13 24 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.8 $X2=0.26
+ $Y2=0.8
r50 12 28 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.8 $X2=1.1
+ $Y2=0.8
r51 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.8
+ $X2=0.345 $Y2=0.8
r52 11 24 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.26 $Y2=0.8
r53 10 21 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.465
+ $X2=0.26 $Y2=0.38
r54 10 11 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.26 $Y=0.465
+ $X2=0.26 $Y2=0.715
r55 3 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r56 2 28 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.72
r57 2 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r58 1 24 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
r59 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%VGND 1 2 3 12 16 18 20 23 24 25 27 36 41 45
r73 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r74 41 42 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r75 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r76 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r77 36 44 4.72899 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.56 $Y=0 $X2=5.77
+ $Y2=0
r78 36 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.56 $Y=0 $X2=5.29
+ $Y2=0
r79 35 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r80 35 42 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=0.69
+ $Y2=0
r81 34 35 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r82 32 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r83 32 34 235.193 $w=1.68e-07 $l=3.605e-06 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=4.37 $Y2=0
r84 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r85 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r86 25 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r87 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r88 23 34 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.37
+ $Y2=0
r89 23 24 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.722
+ $Y2=0
r90 22 38 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.89 $Y=0 $X2=5.29
+ $Y2=0
r91 22 24 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.89 $Y=0 $X2=4.722
+ $Y2=0
r92 18 44 2.99503 $w=3.25e-07 $l=1.06325e-07 $layer=LI1_cond $X=5.722 $Y=0.085
+ $X2=5.77 $Y2=0
r93 18 20 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=5.722 $Y=0.085
+ $X2=5.722 $Y2=0.38
r94 14 24 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.722 $Y=0.085
+ $X2=4.722 $Y2=0
r95 14 16 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=4.722 $Y=0.085
+ $X2=4.722 $Y2=0.38
r96 10 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r97 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r98 3 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.38
r99 2 16 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.235 $X2=4.725 $Y2=0.38
r100 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A_478_47# 1 2 3 16
r20 14 16 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.365 $Y=0.38
+ $X2=4.205 $Y2=0.38
r21 11 14 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.515 $Y=0.38
+ $X2=3.365 $Y2=0.38
r22 3 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.235 $X2=4.205 $Y2=0.38
r23 2 14 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.235 $X2=3.365 $Y2=0.38
r24 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.235 $X2=2.515 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_2%A_730_47# 1 2 7 13
r24 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.225 $Y=0.635
+ $X2=5.225 $Y2=0.36
r25 7 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.06 $Y=0.72
+ $X2=5.225 $Y2=0.635
r26 7 9 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=5.06 $Y=0.72
+ $X2=3.785 $Y2=0.72
r27 2 13 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=5.065
+ $Y=0.235 $X2=5.225 $Y2=0.36
r28 1 9 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.785 $Y2=0.72
.ends


* File: sky130_fd_sc_hd__mux2i_1.pex.spice
* Created: Thu Aug 27 14:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2I_1%A0 1 3 6 8 13
c26 6 0 6.40318e-20 $X=0.49 $Y=1.985
c27 1 0 1.08085e-19 $X=0.47 $Y=0.995
r28 13 14 2.93009 $w=3.29e-07 $l=2e-08 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.49
+ $Y2=1.16
r29 11 13 31.4985 $w=3.29e-07 $l=2.15e-07 $layer=POLY_cond $X=0.255 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r31 4 14 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r33 1 13 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%A1 3 6 8 9 14 16 18 26
c38 18 0 1.36568e-19 $X=1.135 $Y=1.545
c39 16 0 1.18867e-19 $X=0.995 $Y=0.995
r40 18 26 0.915 $w=2e-07 $l=4.69042e-08 $layer=LI1_cond $X=1.135 $Y=1.545
+ $X2=1.095 $Y2=1.53
r41 14 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=1.325
r42 14 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=0.995
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.16 $X2=1.04 $Y2=1.16
r44 8 26 2.135 $w=2e-07 $l=3.5e-08 $layer=LI1_cond $X=1.095 $Y=1.495 $X2=1.095
+ $Y2=1.53
r45 8 15 20.435 $w=2e-07 $l=3.35e-07 $layer=LI1_cond $X=1.095 $Y=1.495 $X2=1.095
+ $Y2=1.16
r46 8 9 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=1.135 $Y=1.58
+ $X2=1.135 $Y2=1.87
r47 8 18 1.94091 $w=1.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.135 $Y=1.58
+ $X2=1.135 $Y2=1.545
r48 6 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.945 $Y=1.985
+ $X2=0.945 $Y2=1.325
r49 3 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.56 $X2=0.89
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%A_283_205# 1 2 9 13 15 23 26 31 34 38
c65 38 0 7.6268e-20 $X=1.85 $Y=1.16
c66 13 0 1.36568e-19 $X=1.85 $Y=0.56
r67 31 33 3.26856 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.982 $Y=0.4
+ $X2=2.982 $Y2=0.485
r68 26 28 34.8294 $w=2.23e-07 $l=6.8e-07 $layer=LI1_cond $X=2.972 $Y=1.62
+ $X2=2.972 $Y2=2.3
r69 24 34 4.82399 $w=2.55e-07 $l=1.32151e-07 $layer=LI1_cond $X=2.972 $Y=1.31
+ $X2=2.942 $Y2=1.192
r70 24 26 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=2.972 $Y=1.31
+ $X2=2.972 $Y2=1.62
r71 23 33 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=2.942 $Y=0.74
+ $X2=2.942 $Y2=0.485
r72 21 34 4.82399 $w=2.55e-07 $l=1.17e-07 $layer=LI1_cond $X=2.942 $Y=1.075
+ $X2=2.942 $Y2=1.192
r73 21 23 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=2.942 $Y=1.075
+ $X2=2.942 $Y2=0.74
r74 18 38 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=1.58 $Y=1.16
+ $X2=1.85 $Y2=1.16
r75 18 35 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.58 $Y=1.16 $X2=1.49
+ $Y2=1.16
r76 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.16 $X2=1.58 $Y2=1.16
r77 15 34 1.63827 $w=2.35e-07 $l=1.42e-07 $layer=LI1_cond $X=2.8 $Y=1.192
+ $X2=2.942 $Y2=1.192
r78 15 17 59.829 $w=2.33e-07 $l=1.22e-06 $layer=LI1_cond $X=2.8 $Y=1.192
+ $X2=1.58 $Y2=1.192
r79 11 38 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.85 $Y=1.025
+ $X2=1.85 $Y2=1.16
r80 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.85 $Y=1.025
+ $X2=1.85 $Y2=0.56
r81 7 35 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.49 $Y=1.295
+ $X2=1.49 $Y2=1.16
r82 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.49 $Y=1.295 $X2=1.49
+ $Y2=1.985
r83 2 28 400 $w=1.7e-07 $l=8.89129e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.485 $X2=3 $Y2=2.3
r84 2 26 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.485 $X2=3 $Y2=1.62
r85 1 31 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.235 $X2=3 $Y2=0.4
r86 1 23 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.235 $X2=3 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%S 3 7 9 11 13 16 18 19 20 21 25
r57 25 27 31.6181 $w=3.43e-07 $l=2.25e-07 $layer=POLY_cond $X=3.21 $Y=1.17
+ $X2=3.435 $Y2=1.17
r58 20 21 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.427 $Y=1.16
+ $X2=3.427 $Y2=1.53
r59 20 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.435
+ $Y=1.16 $X2=3.435 $Y2=1.16
r60 19 20 10.6644 $w=3.33e-07 $l=3.1e-07 $layer=LI1_cond $X=3.427 $Y=0.85
+ $X2=3.427 $Y2=1.16
r61 14 25 22.1447 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.21 $Y=1.35
+ $X2=3.21 $Y2=1.17
r62 14 16 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.21 $Y=1.35
+ $X2=3.21 $Y2=1.985
r63 11 25 22.1447 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.21 $Y=0.99
+ $X2=3.21 $Y2=1.17
r64 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.21 $Y=0.99
+ $X2=3.21 $Y2=0.56
r65 10 18 2.36823 $w=1.85e-07 $l=9e-08 $layer=POLY_cond $X=2.345 $Y=1.257
+ $X2=2.255 $Y2=1.257
r66 9 25 20.7004 $w=3.43e-07 $l=1.18718e-07 $layer=POLY_cond $X=3.135 $Y=1.257
+ $X2=3.21 $Y2=1.17
r67 9 10 291.844 $w=1.85e-07 $l=7.9e-07 $layer=POLY_cond $X=3.135 $Y=1.257
+ $X2=2.345 $Y2=1.257
r68 5 18 24.2117 $w=1.5e-07 $l=9.92169e-08 $layer=POLY_cond $X=2.27 $Y=1.165
+ $X2=2.255 $Y2=1.257
r69 5 7 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.27 $Y=1.165
+ $X2=2.27 $Y2=0.56
r70 1 18 24.2117 $w=1.5e-07 $l=1.0022e-07 $layer=POLY_cond $X=2.24 $Y=1.35
+ $X2=2.255 $Y2=1.257
r71 1 3 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.24 $Y=1.35 $X2=2.24
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%A_27_297# 1 2 7 9 11 14 15 16 17 19
c41 16 0 2.31995e-19 $X=1.575 $Y=1.565
c42 7 0 6.40318e-20 $X=0.27 $Y=2.295
r43 17 24 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=1.65 $X2=2.45
+ $Y2=1.565
r44 17 19 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.45 $Y=1.65
+ $X2=2.45 $Y2=2.32
r45 15 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=1.565
+ $X2=2.45 $Y2=1.565
r46 15 16 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.285 $Y=1.565
+ $X2=1.575 $Y2=1.565
r47 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.49 $Y=1.65
+ $X2=1.575 $Y2=1.565
r48 13 14 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.49 $Y=1.65
+ $X2=1.49 $Y2=2.295
r49 12 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.42 $Y=2.38 $X2=0.27
+ $Y2=2.38
r50 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=2.38
+ $X2=1.49 $Y2=2.295
r51 11 12 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=1.405 $Y=2.38
+ $X2=0.42 $Y2=2.38
r52 7 22 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.295 $X2=0.27
+ $Y2=2.38
r53 7 9 25.93 $w=2.98e-07 $l=6.75e-07 $layer=LI1_cond $X=0.27 $Y=2.295 $X2=0.27
+ $Y2=1.62
r54 2 24 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.485 $X2=2.45 $Y2=1.64
r55 2 19 400 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.485 $X2=2.45 $Y2=2.32
r56 1 22 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r57 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%Y 1 2 7 8 15
r20 7 18 2.90416 $w=2.48e-07 $l=6.3e-08 $layer=LI1_cond $X=0.715 $Y=1.517
+ $X2=0.715 $Y2=1.58
r21 7 25 3.54971 $w=2.48e-07 $l=6.2e-08 $layer=LI1_cond $X=0.715 $Y=1.517
+ $X2=0.715 $Y2=1.455
r22 7 8 12.5847 $w=2.48e-07 $l=2.73e-07 $layer=LI1_cond $X=0.715 $Y=1.597
+ $X2=0.715 $Y2=1.87
r23 7 18 0.783661 $w=2.48e-07 $l=1.7e-08 $layer=LI1_cond $X=0.715 $Y=1.597
+ $X2=0.715 $Y2=1.58
r24 7 25 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=0.685 $Y=1.45
+ $X2=0.685 $Y2=1.455
r25 7 15 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=0.685 $Y=1.45
+ $X2=0.685 $Y2=0.76
r26 2 7 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.62
r27 1 15 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%VPWR 1 2 9 11 13 16 17 18 27 36
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r41 33 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r42 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 27 35 4.45865 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.487 $Y2=2.72
r47 27 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 26 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r49 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 21 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 18 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 18 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 16 25 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 16 17 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=1.86 $Y2=2.72
r55 15 29 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 15 17 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.86 $Y2=2.72
r57 11 35 3.01888 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.442 $Y=2.635
+ $X2=3.487 $Y2=2.72
r58 11 13 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=3.442 $Y=2.635
+ $X2=3.442 $Y2=2
r59 7 17 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=2.635
+ $X2=1.86 $Y2=2.72
r60 7 9 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.86 $Y=2.635
+ $X2=1.86 $Y2=2
r61 2 13 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=2
r62 1 9 300 $w=1.7e-07 $l=6.33798e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.485 $X2=1.83 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%A_27_47# 1 2 9 13 15 20 21
c26 20 0 1.18867e-19 $X=0.44 $Y=0.36
c27 13 0 1.08085e-19 $X=1.175 $Y=0.36
r28 20 21 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=0.44 $Y=0.34
+ $X2=0.965 $Y2=0.34
r29 13 21 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=1.175 $Y=0.36
+ $X2=0.965 $Y2=0.36
r30 13 15 24.5584 $w=2.08e-07 $l=4.65e-07 $layer=LI1_cond $X=1.175 $Y=0.36
+ $X2=1.64 $Y2=0.36
r31 7 20 12.318 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=0.215 $Y=0.36
+ $X2=0.44 $Y2=0.36
r32 7 9 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=0.465
+ $X2=0.215 $Y2=0.72
r33 2 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.235 $X2=1.64 $Y2=0.38
r34 1 7 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r35 1 9 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%A_193_47# 1 2 11 15 17 18
r33 17 18 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.295 $Y=0.77
+ $X2=1.52 $Y2=0.77
r34 13 15 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.502 $Y=0.715
+ $X2=2.502 $Y2=0.55
r35 11 13 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.385 $Y=0.8
+ $X2=2.502 $Y2=0.715
r36 11 18 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.385 $Y=0.8
+ $X2=1.52 $Y2=0.8
r37 9 17 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.12 $Y=0.74
+ $X2=1.295 $Y2=0.74
r38 2 15 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.48 $Y2=0.55
r39 1 9 182 $w=1.7e-07 $l=5.77321e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.12 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_1%VGND 1 2 9 11 13 15 17 25 31 35
r43 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r44 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r45 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r46 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r47 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r48 26 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.06
+ $Y2=0
r49 26 28 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.99
+ $Y2=0
r50 25 34 3.75447 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.507
+ $Y2=0
r51 25 28 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=2.99
+ $Y2=0
r52 24 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r53 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r54 19 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r55 17 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.06
+ $Y2=0
r56 17 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.61
+ $Y2=0
r57 15 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r58 15 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r59 11 34 3.20876 $w=2.2e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.445 $Y=0.085
+ $X2=3.507 $Y2=0
r60 11 13 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.445 $Y=0.085
+ $X2=3.445 $Y2=0.38
r61 7 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=0.085 $X2=2.06
+ $Y2=0
r62 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.06 $Y=0.085 $X2=2.06
+ $Y2=0.38
r63 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.38
r64 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.06 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.spice
* Created: Thu Aug 27 14:26:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.spice.pex"
.subckt sky130_fd_sc_hd__lpflow_isobufsrckapwr_16  VNB VPB A SLEEP VPWR KAPWR X
+ VGND
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1032 N_A_147_47#_M1032_d N_A_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.1755 PD=1.86 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_147_47#_M1002_g N_A_341_47#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_147_47#_M1009_g N_A_341_47#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1009_d N_A_147_47#_M1010_g N_A_341_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_147_47#_M1012_g N_A_341_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1012_d N_SLEEP_M1019_g N_A_341_47#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_SLEEP_M1025_g N_A_341_47#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1025_d N_SLEEP_M1026_g N_A_341_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1030 N_VGND_M1030_d N_SLEEP_M1030_g N_A_341_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_1122_47#_M1003_d N_A_341_47#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75008.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_1122_47#_M1003_d N_A_341_47#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75007.9 A=0.063 P=1.14 MULT=1
MM1028 N_A_1122_47#_M1028_d N_A_341_47#_M1028_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75007.5 A=0.063 P=1.14 MULT=1
MM1038 N_A_1122_47#_M1028_d N_A_341_47#_M1038_g N_VGND_M1038_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75007.1 A=0.063 P=1.14 MULT=1
MM1013 N_X_M1013_d N_A_1122_47#_M1013_g N_VGND_M1038_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75006.6
+ A=0.063 P=1.14 MULT=1
MM1014 N_X_M1013_d N_A_1122_47#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75006.2
+ A=0.063 P=1.14 MULT=1
MM1016 N_X_M1016_d N_A_1122_47#_M1016_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75005.8
+ A=0.063 P=1.14 MULT=1
MM1020 N_X_M1016_d N_A_1122_47#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75005.3
+ A=0.063 P=1.14 MULT=1
MM1023 N_X_M1023_d N_A_1122_47#_M1023_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.6 SB=75004.9
+ A=0.063 P=1.14 MULT=1
MM1024 N_X_M1023_d N_A_1122_47#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.1 SB=75004.5
+ A=0.063 P=1.14 MULT=1
MM1027 N_X_M1027_d N_A_1122_47#_M1027_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.5 SB=75004.1
+ A=0.063 P=1.14 MULT=1
MM1041 N_X_M1027_d N_A_1122_47#_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.05775 PD=0.7 PS=0.695 NRD=0 NRS=0 M=1 R=2.8 SA=75004.9
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1046 N_X_M1046_d N_A_1122_47#_M1046_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.05775 PD=0.7 PS=0.695 NRD=0 NRS=0 M=1 R=2.8 SA=75005.3
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1047 N_X_M1046_d N_A_1122_47#_M1047_g N_VGND_M1047_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.8 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1049 N_X_M1049_d N_A_1122_47#_M1049_g N_VGND_M1047_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1050 N_X_M1049_d N_A_1122_47#_M1050_g N_VGND_M1050_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1051 N_X_M1051_d N_A_1122_47#_M1051_g N_VGND_M1050_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.1 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1055 N_X_M1051_d N_A_1122_47#_M1055_g N_VGND_M1055_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.5 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1056 N_X_M1056_d N_A_1122_47#_M1056_g N_VGND_M1055_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.9 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1057 N_X_M1056_d N_A_1122_47#_M1057_g N_VGND_M1057_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75008.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_147_47#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.28 PD=2.54 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_A_255_297#_M1005_d N_A_147_47#_M1005_g N_A_341_47#_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1017 N_A_255_297#_M1017_d N_A_147_47#_M1017_g N_A_341_47#_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1029 N_A_255_297#_M1017_d N_A_147_47#_M1029_g N_A_341_47#_M1029_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1052 N_A_255_297#_M1052_d N_A_147_47#_M1052_g N_A_341_47#_M1029_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.5 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_A_255_297#_M1052_d N_SLEEP_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1034 N_A_255_297#_M1034_d N_SLEEP_M1034_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1039 N_A_255_297#_M1034_d N_SLEEP_M1039_g N_VPWR_M1039_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1053 N_A_255_297#_M1053_d N_SLEEP_M1053_g N_VPWR_M1039_s VPB PHIGHVT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1015 N_A_1122_47#_M1015_d N_A_341_47#_M1015_g N_KAPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75008.4 A=0.15 P=2.3 MULT=1
MM1037 N_A_1122_47#_M1015_d N_A_341_47#_M1037_g N_KAPWR_M1037_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75007.9 A=0.15 P=2.3 MULT=1
MM1042 N_A_1122_47#_M1042_d N_A_341_47#_M1042_g N_KAPWR_M1037_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75007.5 A=0.15 P=2.3 MULT=1
MM1054 N_A_1122_47#_M1042_d N_A_341_47#_M1054_g N_KAPWR_M1054_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.5 SB=75007.1 A=0.15 P=2.3 MULT=1
MM1001 N_KAPWR_M1054_s N_A_1122_47#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1004 N_KAPWR_M1004_d N_A_1122_47#_M1004_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75006.2 A=0.15 P=2.3 MULT=1
MM1008 N_KAPWR_M1004_d N_A_1122_47#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75005.8 A=0.15 P=2.3 MULT=1
MM1011 N_KAPWR_M1011_d N_A_1122_47#_M1011_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1018 N_KAPWR_M1011_d N_A_1122_47#_M1018_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1021 N_KAPWR_M1021_d N_A_1122_47#_M1021_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1022 N_KAPWR_M1021_d N_A_1122_47#_M1022_g N_X_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1031 N_KAPWR_M1031_d N_A_1122_47#_M1031_g N_X_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.14 PD=1.275 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.9
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1033 N_KAPWR_M1031_d N_A_1122_47#_M1033_g N_X_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.14 PD=1.275 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.3
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1035 N_KAPWR_M1035_d N_A_1122_47#_M1035_g N_X_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.8
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1036 N_KAPWR_M1035_d N_A_1122_47#_M1036_g N_X_M1036_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1040 N_KAPWR_M1040_d N_A_1122_47#_M1040_g N_X_M1036_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1043 N_KAPWR_M1040_d N_A_1122_47#_M1043_g N_X_M1043_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1044 N_KAPWR_M1044_d N_A_1122_47#_M1044_g N_X_M1043_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.5 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1045 N_KAPWR_M1044_d N_A_1122_47#_M1045_g N_X_M1045_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1048 N_KAPWR_M1048_d N_A_1122_47#_M1048_g N_X_M1045_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX58_noxref VNB VPB NWDIODE A=23.4972 P=32.49
c_129 VNB 0 1.68547e-19 $X=5.205 $Y=-0.085
*
.include "sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.spice.SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16.pxi"
*
.ends
*
*

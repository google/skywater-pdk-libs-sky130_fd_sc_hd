* File: sky130_fd_sc_hd__a2bb2o_1.spice.pex
* Created: Thu Aug 27 14:03:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%A_76_199# 1 2 9 12 15 16 17 19 20 21 23 26
+ 29 30 34 38 41
c97 38 0 7.28036e-20 $X=2.495 $Y=0.785
c98 34 0 1.61547e-19 $X=2.16 $Y=2.275
c99 29 0 1.32536e-19 $X=0.515 $Y=1.16
r100 36 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.315 $Y=0.785
+ $X2=2.495 $Y2=0.785
r101 34 35 0.405316 $w=3.01e-07 $l=1e-08 $layer=LI1_cond $X=2.195 $Y=2.275
+ $X2=2.195 $Y2=2.285
r102 30 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r103 30 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r104 29 32 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.557 $Y=1.16
+ $X2=0.557 $Y2=1.325
r105 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r106 24 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.7
+ $X2=2.495 $Y2=0.785
r107 24 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.495 $Y=0.7
+ $X2=2.495 $Y2=0.445
r108 23 34 17.6939 $w=3.01e-07 $l=4.3589e-07 $layer=LI1_cond $X=2.315 $Y=1.895
+ $X2=2.195 $Y2=2.275
r109 22 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=0.87
+ $X2=2.315 $Y2=0.785
r110 22 23 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.315 $Y=0.87
+ $X2=2.315 $Y2=1.895
r111 20 35 4.08057 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.99 $Y=2.285
+ $X2=2.195 $Y2=2.285
r112 20 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.99 $Y=2.285
+ $X2=1.275 $Y2=2.285
r113 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=2.2
+ $X2=1.275 $Y2=2.285
r114 18 19 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.19 $Y=1.975
+ $X2=1.19 $Y2=2.2
r115 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=1.89
+ $X2=1.19 $Y2=1.975
r116 16 17 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.105 $Y=1.89
+ $X2=0.685 $Y2=1.89
r117 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=1.805
+ $X2=0.685 $Y2=1.89
r118 15 32 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.6 $Y=1.805
+ $X2=0.6 $Y2=1.325
r119 12 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r120 9 41 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
r121 2 34 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=2.065 $X2=2.16 $Y2=2.275
r122 1 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.235 $X2=2.495 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%A1_N 3 7 9 10 14 15
r36 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=1.325
r37 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=0.995
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r39 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.075 $Y=1.19
+ $X2=1.075 $Y2=1.53
r40 9 15 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.075 $Y=1.19 $X2=1.075
+ $Y2=1.16
r41 7 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.055 $Y=1.695
+ $X2=1.055 $Y2=1.325
r42 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.055 $Y=0.445
+ $X2=1.055 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%A2_N 1 3 6 8
c31 6 0 7.28036e-20 $X=1.475 $Y=0.445
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r33 8 12 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=1.615 $Y=1.185
+ $X2=1.495 $Y2=1.185
r34 4 11 38.945 $w=2.68e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.485 $Y2=1.16
r35 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.445
r36 1 11 47.9375 $w=2.68e-07 $l=2.47538e-07 $layer=POLY_cond $X=1.415 $Y=1.375
+ $X2=1.485 $Y2=1.16
r37 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.415 $Y=1.375
+ $X2=1.415 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%A_226_47# 1 2 9 11 14 18 22 24 25 26 31 32
+ 35 38
c68 32 0 4.6512e-20 $X=1.975 $Y=1.07
c69 31 0 1.04517e-19 $X=1.975 $Y=1.07
r70 32 39 67.6946 $w=5.2e-07 $l=3.65e-07 $layer=POLY_cond $X=2.1 $Y=1.07 $X2=2.1
+ $Y2=1.435
r71 32 38 61.5212 $w=5.2e-07 $l=3.05e-07 $layer=POLY_cond $X=2.1 $Y=1.07 $X2=2.1
+ $Y2=0.765
r72 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=1.07 $X2=1.975 $Y2=1.07
r73 29 31 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.975 $Y=1.545
+ $X2=1.975 $Y2=1.07
r74 28 31 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.975 $Y=0.825
+ $X2=1.975 $Y2=1.07
r75 27 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.63
+ $X2=1.625 $Y2=1.63
r76 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.89 $Y=1.63
+ $X2=1.975 $Y2=1.545
r77 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.89 $Y=1.63
+ $X2=1.71 $Y2=1.63
r78 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.89 $Y=0.74
+ $X2=1.975 $Y2=0.825
r79 24 25 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.89 $Y=0.74
+ $X2=1.35 $Y2=0.74
r80 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.265 $Y=0.655
+ $X2=1.35 $Y2=0.74
r81 20 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.265 $Y=0.655
+ $X2=1.265 $Y2=0.445
r82 16 18 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=2.285 $Y=1.83
+ $X2=2.37 $Y2=1.83
r83 12 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.905
+ $X2=2.37 $Y2=1.83
r84 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.37 $Y=1.905
+ $X2=2.37 $Y2=2.275
r85 11 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=1.755
+ $X2=2.285 $Y2=1.83
r86 11 39 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.285 $Y=1.755
+ $X2=2.285 $Y2=1.435
r87 9 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.285 $Y=0.445
+ $X2=2.285 $Y2=0.765
r88 2 35 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.485 $X2=1.625 $Y2=1.71
r89 1 22 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.265 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%B2 3 7 11 14 20
c46 20 0 4.6512e-20 $X=2.95 $Y=1.505
c47 11 0 1.22353e-19 $X=2.995 $Y=1.53
c48 7 0 1.75342e-19 $X=2.79 $Y=2.275
c49 3 0 1.04517e-19 $X=2.705 $Y=0.445
r50 15 20 7.10673 $w=2.98e-07 $l=1.85e-07 $layer=LI1_cond $X=2.765 $Y=1.505
+ $X2=2.95 $Y2=1.505
r51 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.47
+ $X2=2.765 $Y2=1.635
r52 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.47
+ $X2=2.765 $Y2=1.305
r53 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.47 $X2=2.765 $Y2=1.47
r54 11 20 1.72866 $w=2.98e-07 $l=4.5e-08 $layer=LI1_cond $X=2.995 $Y=1.505
+ $X2=2.95 $Y2=1.505
r55 7 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.79 $Y=2.275 $X2=2.79
+ $Y2=1.635
r56 3 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.705 $Y=0.445
+ $X2=2.705 $Y2=1.305
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%B1 3 7 9 10 11 16
c30 16 0 1.22353e-19 $X=3.21 $Y=1.16
c31 9 0 1.37947e-20 $X=3.455 $Y=0.85
r32 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.365
+ $Y=1.16 $X2=3.365 $Y2=1.16
r33 16 18 25.2399 $w=2.96e-07 $l=1.55e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.365 $Y2=1.16
r34 10 11 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.41 $Y=1.19
+ $X2=3.41 $Y2=1.53
r35 10 19 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=3.41 $Y=1.19 $X2=3.41
+ $Y2=1.16
r36 9 19 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=3.41 $Y=0.85 $X2=3.41
+ $Y2=1.16
r37 5 16 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r38 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.21 $Y=1.325 $X2=3.21
+ $Y2=2.275
r39 1 16 13.8412 $w=2.96e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.125 $Y=0.995
+ $X2=3.21 $Y2=1.16
r40 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.125 $Y=0.995
+ $X2=3.125 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%X 1 2 10 11 12 13 14 15 24
r17 14 15 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=2.21
r18 14 24 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=1.76
r19 11 24 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=0.215 $Y=1.655
+ $X2=0.215 $Y2=1.76
r20 11 12 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.655
+ $X2=0.215 $Y2=1.525
r21 10 12 45.3143 $w=1.73e-07 $l=7.15e-07 $layer=LI1_cond $X=0.172 $Y=0.81
+ $X2=0.172 $Y2=1.525
r22 9 13 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.215 $Y=0.68
+ $X2=0.215 $Y2=0.51
r23 9 10 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=0.68
+ $X2=0.215 $Y2=0.81
r24 2 24 300 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.76
r25 1 13 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%VPWR 1 2 9 13 15 17 19 24 26 33 34 37 40
r52 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 34 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 31 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.04 $Y2=2.72
r57 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 30 41 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 30 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 27 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r62 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 26 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.04 $Y2=2.72
r64 26 29 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 19 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r66 17 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 17 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 15 19 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.515 $Y2=2.72
r69 15 24 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 11 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=2.635
+ $X2=3.04 $Y2=2.72
r71 11 13 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.04 $Y=2.635
+ $X2=3.04 $Y2=2.34
r72 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r73 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.32
r74 2 13 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=2.065 $X2=3 $Y2=2.34
r75 1 9 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%A_489_413# 1 2 8 9 10 13 16
r33 11 13 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.425 $Y=2.005
+ $X2=3.425 $Y2=2.275
r34 9 11 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.335 $Y=1.92
+ $X2=3.425 $Y2=2.005
r35 9 10 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.335 $Y=1.92
+ $X2=2.745 $Y2=1.92
r36 8 16 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.66 $Y=2.255
+ $X2=2.58 $Y2=2.34
r37 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.66 $Y=2.005
+ $X2=2.745 $Y2=1.92
r38 7 8 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.66 $Y=2.005 $X2=2.66
+ $Y2=2.255
r39 2 13 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=2.065 $X2=3.42 $Y2=2.275
r40 1 16 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=2.065 $X2=2.58 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_1%VGND 1 2 3 12 14 16 18 20 22 27 34 40 45 51
+ 54
r55 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 50 51 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=0.2
+ $X2=2.24 $Y2=0.2
r57 47 50 0.104919 $w=5.68e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=0.2 $X2=2.075
+ $Y2=0.2
r58 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r59 44 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r60 43 47 9.65256 $w=5.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=0.2 $X2=2.07
+ $Y2=0.2
r61 43 45 8.38723 $w=5.68e-07 $l=9e-08 $layer=LI1_cond $X=1.61 $Y=0.2 $X2=1.52
+ $Y2=0.2
r62 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r63 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r64 38 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r65 38 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r66 37 51 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.24
+ $Y2=0
r67 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r68 34 53 5.3623 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.417
+ $Y2=0
r69 34 37 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=2.99
+ $Y2=0
r70 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r71 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r72 32 45 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.52
+ $Y2=0
r73 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r74 30 40 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.73
+ $Y2=0
r75 30 32 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.15
+ $Y2=0
r76 22 40 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.73
+ $Y2=0
r77 20 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r78 20 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r79 18 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.515
+ $Y2=0
r80 18 27 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r81 14 53 3.00862 $w=4e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.417 $Y2=0
r82 14 16 9.93982 $w=3.98e-07 $l=3.45e-07 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0.43
r83 10 40 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r84 10 12 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.445
r85 3 16 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.235 $X2=3.335 $Y2=0.43
r86 2 50 91 $w=1.7e-07 $l=6.01872e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.235 $X2=2.075 $Y2=0.4
r87 1 12 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.445
.ends


* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR B1 a_730_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.94e+12p pd=1.388e+07u as=5.4e+11p ps=5.08e+06u
M1001 a_471_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=7.1825e+11p pd=7.41e+06u as=7.02e+11p ps=7.36e+06u
M1002 a_113_297# A1_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1003 a_730_297# B2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1004 a_113_47# A2_N a_113_297# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=1.755e+11p ps=1.84e+06u
M1005 a_113_297# A2_N a_113_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B1 a_471_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_471_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B2 a_730_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B2 a_471_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1_N a_113_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_113_47# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_113_297# a_471_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1013 VPWR A1_N a_113_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_113_297# A2_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_471_47# a_113_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_113_297# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A2_N a_113_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_730_297# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y a_113_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


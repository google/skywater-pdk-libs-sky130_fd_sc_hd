* File: sky130_fd_sc_hd__or4_4.pxi.spice
* Created: Tue Sep  1 19:28:33 2020
* 
x_PM_SKY130_FD_SC_HD__OR4_4%D N_D_c_80_n N_D_M1004_g N_D_M1002_g D D N_D_c_82_n
+ PM_SKY130_FD_SC_HD__OR4_4%D
x_PM_SKY130_FD_SC_HD__OR4_4%C N_C_M1012_g N_C_M1009_g N_C_c_113_n N_C_c_114_n C
+ C N_C_c_115_n C PM_SKY130_FD_SC_HD__OR4_4%C
x_PM_SKY130_FD_SC_HD__OR4_4%B N_B_c_161_n N_B_M1014_g N_B_M1008_g N_B_c_162_n
+ N_B_c_163_n B B B PM_SKY130_FD_SC_HD__OR4_4%B
x_PM_SKY130_FD_SC_HD__OR4_4%A N_A_M1000_g N_A_M1005_g A N_A_c_201_n N_A_c_202_n
+ N_A_c_203_n PM_SKY130_FD_SC_HD__OR4_4%A
x_PM_SKY130_FD_SC_HD__OR4_4%A_32_297# N_A_32_297#_M1004_d N_A_32_297#_M1014_d
+ N_A_32_297#_M1002_s N_A_32_297#_c_242_n N_A_32_297#_M1001_g
+ N_A_32_297#_M1007_g N_A_32_297#_c_243_n N_A_32_297#_M1003_g
+ N_A_32_297#_M1010_g N_A_32_297#_c_244_n N_A_32_297#_M1006_g
+ N_A_32_297#_M1011_g N_A_32_297#_c_245_n N_A_32_297#_M1015_g
+ N_A_32_297#_M1013_g N_A_32_297#_c_254_n N_A_32_297#_c_246_n
+ N_A_32_297#_c_263_n N_A_32_297#_c_274_n N_A_32_297#_c_264_n
+ N_A_32_297#_c_366_p N_A_32_297#_c_288_n N_A_32_297#_c_247_n
+ N_A_32_297#_c_248_n N_A_32_297#_c_318_p N_A_32_297#_c_256_n
+ N_A_32_297#_c_283_n N_A_32_297#_c_249_n PM_SKY130_FD_SC_HD__OR4_4%A_32_297#
x_PM_SKY130_FD_SC_HD__OR4_4%VPWR N_VPWR_M1005_d N_VPWR_M1010_d N_VPWR_M1013_d
+ N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n VPWR
+ N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n
+ N_VPWR_c_392_n VPWR PM_SKY130_FD_SC_HD__OR4_4%VPWR
x_PM_SKY130_FD_SC_HD__OR4_4%X N_X_M1001_d N_X_M1006_d N_X_M1007_s N_X_M1011_s
+ N_X_c_453_n N_X_c_494_n N_X_c_462_n N_X_c_454_n N_X_c_447_n N_X_c_448_n
+ N_X_c_477_n N_X_c_498_n N_X_c_455_n N_X_c_449_n N_X_c_450_n N_X_c_456_n X
+ N_X_c_452_n PM_SKY130_FD_SC_HD__OR4_4%X
x_PM_SKY130_FD_SC_HD__OR4_4%VGND N_VGND_M1004_s N_VGND_M1012_d N_VGND_M1000_d
+ N_VGND_M1003_s N_VGND_M1015_s N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n
+ N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n
+ N_VGND_c_529_n VGND N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n
+ N_VGND_c_533_n N_VGND_c_534_n N_VGND_c_535_n VGND
+ PM_SKY130_FD_SC_HD__OR4_4%VGND
cc_1 VNB N_D_c_80_n 0.0197158f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_2 VNB D 0.0217888f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=0.765
cc_3 VNB N_D_c_82_n 0.035408f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_4 VNB N_C_c_113_n 6.47944e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_C_c_114_n 0.0229145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_C_c_115_n 0.0171358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_161_n 0.0162189f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_8 VNB N_B_c_162_n 0.00583329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_163_n 0.0186258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_201_n 0.0229306f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_11 VNB N_A_c_202_n 6.43385e-19 $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_12 VNB N_A_c_203_n 0.0174079f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_13 VNB N_A_32_297#_c_242_n 0.0163299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_32_297#_c_243_n 0.0157937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_32_297#_c_244_n 0.0157971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_32_297#_c_245_n 0.0191578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_32_297#_c_246_n 0.00293881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_32_297#_c_247_n 0.00157854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_32_297#_c_248_n 0.00376665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_32_297#_c_249_n 0.0647168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_392_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_447_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_448_n 0.00187124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_449_n 0.00105843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_450_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0202945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_452_n 0.00847149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_521_n 0.0106918f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_29 VNB N_VGND_c_522_n 0.0185191f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=0.85
cc_30 VNB N_VGND_c_523_n 0.0181903f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_31 VNB N_VGND_c_524_n 4.04385e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_525_n 0.00239633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_526_n 0.0148447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_527_n 0.0035091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_528_n 0.0111098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_529_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_530_n 0.0135943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_531_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_532_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_533_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_534_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_535_n 0.218315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_D_M1002_g 0.0265308f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_44 VPB D 0.00425673f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=0.765
cc_45 VPB N_D_c_82_n 0.00920598f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_46 VPB N_C_M1009_g 0.019342f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_47 VPB N_C_c_113_n 0.00103465f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_C_c_114_n 0.00584707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_B_M1008_g 0.0174072f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_50 VPB N_B_c_162_n 0.00536776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_B_c_163_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB B 2.2639e-19 $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_53 VPB N_A_M1005_g 0.0193215f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_54 VPB A 0.00385897f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=0.765
cc_55 VPB N_A_c_201_n 0.00445127f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_56 VPB N_A_c_202_n 0.00148828f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_57 VPB N_A_32_297#_M1007_g 0.0199018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_32_297#_M1010_g 0.0182214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_32_297#_M1011_g 0.0182002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_32_297#_M1013_g 0.0219116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_32_297#_c_254_n 0.0310345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_32_297#_c_246_n 0.00111305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_32_297#_c_256_n 0.00750303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_32_297#_c_249_n 0.0102664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_393_n 0.00463796f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_66 VPB N_VPWR_c_394_n 0.00399514f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_67 VPB N_VPWR_c_395_n 0.0117686f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=0.85
cc_68 VPB N_VPWR_c_396_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.16
cc_69 VPB N_VPWR_c_397_n 0.0576502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_398_n 0.0181285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_399_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_400_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_401_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_392_n 0.046466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_X_c_453_n 0.00246856f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_76 VPB N_X_c_454_n 0.00252706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_X_c_455_n 0.0107161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_X_c_456_n 0.00220075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB X 0.00757383f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 N_D_M1002_g N_C_M1009_g 0.0380647f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_81 N_D_M1002_g N_C_c_113_n 8.39734e-19 $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_82 N_D_c_82_n N_C_c_113_n 3.03886e-19 $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_83 N_D_c_82_n N_C_c_114_n 0.0153445f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_84 N_D_M1002_g C 0.00563885f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_85 N_D_c_80_n N_C_c_115_n 0.0196848f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_86 N_D_M1002_g N_A_32_297#_c_254_n 0.0135008f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_87 N_D_c_80_n N_A_32_297#_c_246_n 0.00353f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_88 N_D_M1002_g N_A_32_297#_c_246_n 0.00854641f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_89 D N_A_32_297#_c_246_n 0.0334541f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_90 N_D_c_82_n N_A_32_297#_c_246_n 0.0076194f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_91 N_D_c_80_n N_A_32_297#_c_263_n 0.00412485f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_92 N_D_c_80_n N_A_32_297#_c_264_n 0.00875447f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_93 N_D_M1002_g N_A_32_297#_c_256_n 0.0147115f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_94 D N_A_32_297#_c_256_n 0.0196765f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_95 N_D_c_82_n N_A_32_297#_c_256_n 0.00153074f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_96 N_D_M1002_g N_VPWR_c_397_n 0.00541964f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_97 N_D_M1002_g N_VPWR_c_392_n 0.0109626f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_98 D N_VGND_M1004_s 0.00285205f $X=0.14 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_99 D N_VGND_c_521_n 5.41347e-19 $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_100 N_D_c_80_n N_VGND_c_522_n 0.0044954f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_101 D N_VGND_c_522_n 0.0209517f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_102 N_D_c_82_n N_VGND_c_522_n 9.93976e-19 $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_103 N_D_c_80_n N_VGND_c_523_n 0.00553912f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_104 N_D_c_80_n N_VGND_c_524_n 0.0012701f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_105 N_D_c_80_n N_VGND_c_535_n 0.010884f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_106 D N_VGND_c_535_n 0.00197281f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_107 N_C_c_115_n N_B_c_161_n 0.0251622f $X=0.965 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_108 N_C_M1009_g N_B_M1008_g 0.0567511f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_109 N_C_c_113_n N_B_M1008_g 6.62811e-19 $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_110 C N_B_M1008_g 0.00466387f $X=1.06 $Y=1.785 $X2=0 $Y2=0
cc_111 N_C_c_113_n N_B_c_162_n 0.0274089f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C_c_114_n N_B_c_162_n 0.00284781f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_113 N_C_c_113_n N_B_c_163_n 3.68507e-19 $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_114 N_C_c_114_n N_B_c_163_n 0.0203414f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C_M1009_g B 0.00129617f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_116 N_C_c_113_n B 0.00652405f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_117 C B 0.0291214f $X=1.06 $Y=1.785 $X2=0 $Y2=0
cc_118 C B 0.0291214f $X=1.145 $Y=1.87 $X2=0 $Y2=0
cc_119 N_C_M1009_g N_A_32_297#_c_254_n 0.00105448f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_120 C N_A_32_297#_c_254_n 0.0270752f $X=1.06 $Y=1.785 $X2=0 $Y2=0
cc_121 N_C_M1009_g N_A_32_297#_c_246_n 4.90921e-19 $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_122 N_C_c_113_n N_A_32_297#_c_246_n 0.0363735f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_123 N_C_c_114_n N_A_32_297#_c_246_n 0.0021031f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C_c_115_n N_A_32_297#_c_246_n 0.00338056f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_125 N_C_c_113_n N_A_32_297#_c_274_n 0.0108856f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C_c_114_n N_A_32_297#_c_274_n 3.62043e-19 $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_127 N_C_c_115_n N_A_32_297#_c_274_n 0.0131138f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C_c_114_n N_A_32_297#_c_264_n 0.00189854f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_129 N_C_M1009_g N_A_32_297#_c_256_n 5.95476e-19 $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_130 N_C_c_113_n N_A_32_297#_c_256_n 0.0136667f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_131 N_C_c_113_n A_114_297# 0.00117219f $X=0.965 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_132 C A_114_297# 0.00214124f $X=1.06 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_133 C A_114_297# 0.00791228f $X=1.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_134 C A_220_297# 0.00473131f $X=1.06 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_135 C A_220_297# 0.00575507f $X=1.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_136 N_C_M1009_g N_VPWR_c_397_n 0.00375793f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_137 C N_VPWR_c_397_n 0.0127745f $X=1.145 $Y=1.87 $X2=0 $Y2=0
cc_138 N_C_M1009_g N_VPWR_c_392_n 0.0056317f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_139 C N_VPWR_c_392_n 0.0120515f $X=1.145 $Y=1.87 $X2=0 $Y2=0
cc_140 N_C_c_115_n N_VGND_c_523_n 0.00341689f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_141 N_C_c_115_n N_VGND_c_524_n 0.00869343f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C_c_115_n N_VGND_c_535_n 0.00431054f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B_M1008_g N_A_M1005_g 0.0564998f $X=1.445 $Y=1.985 $X2=0 $Y2=0
cc_144 B N_A_M1005_g 0.00915664f $X=1.52 $Y=1.785 $X2=0 $Y2=0
cc_145 N_B_c_162_n A 0.0102741f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B_c_162_n N_A_c_201_n 0.00373575f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B_c_163_n N_A_c_201_n 0.0203414f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B_c_162_n N_A_c_202_n 0.0271074f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B_c_163_n N_A_c_202_n 3.68507e-19 $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_150 N_B_c_161_n N_A_c_203_n 0.0243955f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B_c_161_n N_A_32_297#_c_274_n 0.0110728f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B_c_162_n N_A_32_297#_c_274_n 0.018276f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_153 N_B_c_163_n N_A_32_297#_c_274_n 2.98597e-19 $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B_c_162_n N_A_32_297#_c_283_n 0.00316818f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_155 B A_304_297# 0.0164072f $X=1.52 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_156 B N_VPWR_c_393_n 0.031049f $X=1.52 $Y=1.785 $X2=0 $Y2=0
cc_157 N_B_M1008_g N_VPWR_c_397_n 0.00419108f $X=1.445 $Y=1.985 $X2=0 $Y2=0
cc_158 B N_VPWR_c_397_n 0.0126498f $X=1.52 $Y=1.785 $X2=0 $Y2=0
cc_159 N_B_M1008_g N_VPWR_c_392_n 0.00651073f $X=1.445 $Y=1.985 $X2=0 $Y2=0
cc_160 B N_VPWR_c_392_n 0.0110804f $X=1.52 $Y=1.785 $X2=0 $Y2=0
cc_161 N_B_c_161_n N_VGND_c_524_n 0.00732663f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B_c_161_n N_VGND_c_530_n 0.00341689f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B_c_161_n N_VGND_c_535_n 0.00405445f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_203_n N_A_32_297#_c_242_n 0.0200495f $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_M1005_g N_A_32_297#_M1007_g 0.0173803f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_166 A N_A_32_297#_M1007_g 0.00128363f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_167 N_A_c_202_n N_A_32_297#_M1007_g 0.00219223f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_168 A N_A_32_297#_c_288_n 0.00495213f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_169 N_A_c_201_n N_A_32_297#_c_288_n 0.00173573f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_202_n N_A_32_297#_c_288_n 0.0104547f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_203_n N_A_32_297#_c_288_n 0.0134819f $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_201_n N_A_32_297#_c_247_n 5.07416e-19 $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_202_n N_A_32_297#_c_247_n 0.00568393f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_203_n N_A_32_297#_c_247_n 0.00336447f $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_175 A N_A_32_297#_c_248_n 0.00707041f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_176 N_A_c_201_n N_A_32_297#_c_248_n 0.00124527f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_c_202_n N_A_32_297#_c_248_n 0.0137152f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_201_n N_A_32_297#_c_249_n 0.0161964f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_202_n N_A_32_297#_c_249_n 7.74805e-19 $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_180 A N_VPWR_M1005_d 0.00433176f $X=1.98 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_181 N_A_M1005_g N_VPWR_c_393_n 0.00789297f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_182 A N_VPWR_c_393_n 0.0193325f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_183 N_A_M1005_g N_VPWR_c_397_n 0.00585385f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_M1005_g N_VPWR_c_392_n 0.0109527f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_185 A N_X_c_453_n 0.00229946f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_186 N_A_c_203_n N_VGND_c_524_n 6.8876e-19 $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_203_n N_VGND_c_525_n 0.00318791f $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_203_n N_VGND_c_530_n 0.00428022f $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_203_n N_VGND_c_535_n 0.00603983f $X=1.925 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_32_297#_c_246_n A_114_297# 3.28342e-19 $X=0.625 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_32_297#_c_256_n A_114_297# 0.00486679f $X=0.625 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_192 N_A_32_297#_M1007_g N_VPWR_c_393_n 0.00430866f $X=2.395 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_32_297#_M1010_g N_VPWR_c_394_n 0.00165046f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_32_297#_M1011_g N_VPWR_c_394_n 0.00157837f $X=3.235 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_32_297#_M1013_g N_VPWR_c_396_n 0.00338128f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_32_297#_c_254_n N_VPWR_c_397_n 0.0195303f $X=0.285 $Y=2.34 $X2=0
+ $Y2=0
cc_197 N_A_32_297#_M1007_g N_VPWR_c_398_n 0.00585385f $X=2.395 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_32_297#_M1010_g N_VPWR_c_398_n 0.00585385f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_32_297#_M1011_g N_VPWR_c_399_n 0.00585385f $X=3.235 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_32_297#_M1013_g N_VPWR_c_399_n 0.00585385f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_32_297#_M1002_s N_VPWR_c_392_n 0.00209863f $X=0.16 $Y=1.485 $X2=0
+ $Y2=0
cc_202 N_A_32_297#_M1007_g N_VPWR_c_392_n 0.0108486f $X=2.395 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_32_297#_M1010_g N_VPWR_c_392_n 0.0104367f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_32_297#_M1011_g N_VPWR_c_392_n 0.0104367f $X=3.235 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_32_297#_M1013_g N_VPWR_c_392_n 0.0114051f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_32_297#_c_254_n N_VPWR_c_392_n 0.012527f $X=0.285 $Y=2.34 $X2=0 $Y2=0
cc_207 N_A_32_297#_M1007_g N_X_c_453_n 2.80238e-19 $X=2.395 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_32_297#_c_318_p N_X_c_453_n 0.0172286f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_32_297#_c_249_n N_X_c_453_n 0.00226413f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_32_297#_c_243_n N_X_c_462_n 0.00701434f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_32_297#_c_244_n N_X_c_462_n 5.23786e-19 $X=3.235 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_32_297#_M1010_g N_X_c_454_n 0.0134538f $X=2.815 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_32_297#_M1011_g N_X_c_454_n 0.013468f $X=3.235 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_32_297#_c_318_p N_X_c_454_n 0.03482f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_32_297#_c_249_n N_X_c_454_n 0.00216069f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_32_297#_c_243_n N_X_c_447_n 0.00870364f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_32_297#_c_244_n N_X_c_447_n 0.00865686f $X=3.235 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_32_297#_c_318_p N_X_c_447_n 0.0356734f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_32_297#_c_249_n N_X_c_447_n 0.00222133f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_32_297#_c_242_n N_X_c_448_n 8.16938e-19 $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_32_297#_c_243_n N_X_c_448_n 0.00250064f $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_32_297#_c_247_n N_X_c_448_n 0.00357582f $X=2.265 $Y=1.075 $X2=0 $Y2=0
cc_223 N_A_32_297#_c_318_p N_X_c_448_n 0.01996f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_32_297#_c_249_n N_X_c_448_n 0.00230339f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_32_297#_c_243_n N_X_c_477_n 5.22228e-19 $X=2.815 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_32_297#_c_244_n N_X_c_477_n 0.00630972f $X=3.235 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_32_297#_c_245_n N_X_c_477_n 0.0109314f $X=3.655 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_32_297#_M1013_g N_X_c_455_n 0.0159196f $X=3.655 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_32_297#_c_318_p N_X_c_455_n 0.00401279f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_32_297#_c_245_n N_X_c_449_n 0.0113418f $X=3.655 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_32_297#_c_318_p N_X_c_449_n 0.00200821f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_32_297#_c_244_n N_X_c_450_n 0.00113286f $X=3.235 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_32_297#_c_245_n N_X_c_450_n 0.00113286f $X=3.655 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_32_297#_c_318_p N_X_c_450_n 0.026256f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_32_297#_c_249_n N_X_c_450_n 0.00230339f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_32_297#_c_318_p N_X_c_456_n 0.0172286f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_32_297#_c_249_n N_X_c_456_n 0.00226413f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_32_297#_c_245_n X 0.0212433f $X=3.655 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_32_297#_c_318_p X 0.0137867f $X=3.475 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_32_297#_c_274_n N_VGND_M1012_d 0.00664072f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_32_297#_c_288_n N_VGND_M1000_d 0.00616911f $X=2.18 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_32_297#_c_247_n N_VGND_M1000_d 7.20909e-19 $X=2.265 $Y=1.075 $X2=0
+ $Y2=0
cc_243 N_A_32_297#_c_263_n N_VGND_c_523_n 0.00852533f $X=0.785 $Y=0.49 $X2=0
+ $Y2=0
cc_244 N_A_32_297#_c_264_n N_VGND_c_523_n 0.00502163f $X=0.87 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_32_297#_c_263_n N_VGND_c_524_n 0.0117247f $X=0.785 $Y=0.49 $X2=0
+ $Y2=0
cc_246 N_A_32_297#_c_274_n N_VGND_c_524_n 0.0160613f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_32_297#_c_242_n N_VGND_c_525_n 0.00675761f $X=2.395 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_32_297#_c_243_n N_VGND_c_525_n 5.99174e-19 $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_32_297#_c_288_n N_VGND_c_525_n 0.0224385f $X=2.18 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_32_297#_c_242_n N_VGND_c_526_n 0.00496106f $X=2.395 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_32_297#_c_243_n N_VGND_c_526_n 0.00423334f $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_32_297#_c_243_n N_VGND_c_527_n 0.00138579f $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A_32_297#_c_244_n N_VGND_c_527_n 0.00146448f $X=3.235 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A_32_297#_c_245_n N_VGND_c_529_n 0.00316354f $X=3.655 $Y=0.995 $X2=0
+ $Y2=0
cc_255 N_A_32_297#_c_274_n N_VGND_c_530_n 0.00232396f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_32_297#_c_366_p N_VGND_c_530_n 0.00846569f $X=1.655 $Y=0.49 $X2=0
+ $Y2=0
cc_257 N_A_32_297#_c_288_n N_VGND_c_530_n 0.0029785f $X=2.18 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_32_297#_c_244_n N_VGND_c_531_n 0.00423334f $X=3.235 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_32_297#_c_245_n N_VGND_c_531_n 0.00423334f $X=3.655 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_32_297#_M1004_d N_VGND_c_535_n 0.00390697f $X=0.57 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_32_297#_M1014_d N_VGND_c_535_n 0.00256656f $X=1.52 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_32_297#_c_242_n N_VGND_c_535_n 0.00822344f $X=2.395 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A_32_297#_c_243_n N_VGND_c_535_n 0.00575518f $X=2.815 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_32_297#_c_244_n N_VGND_c_535_n 0.0057163f $X=3.235 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_32_297#_c_245_n N_VGND_c_535_n 0.00668462f $X=3.655 $Y=0.995 $X2=0
+ $Y2=0
cc_266 N_A_32_297#_c_263_n N_VGND_c_535_n 0.00618681f $X=0.785 $Y=0.49 $X2=0
+ $Y2=0
cc_267 N_A_32_297#_c_274_n N_VGND_c_535_n 0.00554474f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_32_297#_c_264_n N_VGND_c_535_n 0.00936859f $X=0.87 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_32_297#_c_366_p N_VGND_c_535_n 0.00625722f $X=1.655 $Y=0.49 $X2=0
+ $Y2=0
cc_270 N_A_32_297#_c_288_n N_VGND_c_535_n 0.00734097f $X=2.18 $Y=0.74 $X2=0
+ $Y2=0
cc_271 A_114_297# N_VPWR_c_392_n 0.0138706f $X=0.57 $Y=1.485 $X2=0 $Y2=0
cc_272 A_220_297# N_VPWR_c_392_n 0.00710526f $X=1.1 $Y=1.485 $X2=0 $Y2=0
cc_273 A_304_297# N_VPWR_c_392_n 0.0046981f $X=1.52 $Y=1.485 $X2=0 $Y2=0
cc_274 N_VPWR_c_392_n N_X_M1007_s 0.00284632f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_c_392_n N_X_M1011_s 0.00284632f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_276 N_VPWR_c_398_n N_X_c_494_n 0.0142343f $X=2.9 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_392_n N_X_c_494_n 0.00955092f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_M1010_d N_X_c_454_n 0.00165831f $X=2.89 $Y=1.485 $X2=0 $Y2=0
cc_279 N_VPWR_c_394_n N_X_c_454_n 0.0126919f $X=3.025 $Y=1.96 $X2=0 $Y2=0
cc_280 N_VPWR_c_399_n N_X_c_498_n 0.0142343f $X=3.74 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_392_n N_X_c_498_n 0.00955092f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_M1013_d N_X_c_455_n 0.00340835f $X=3.73 $Y=1.485 $X2=0 $Y2=0
cc_283 N_VPWR_c_396_n N_X_c_455_n 0.0179737f $X=3.865 $Y=1.96 $X2=0 $Y2=0
cc_284 N_X_c_447_n N_VGND_M1003_s 0.00162089f $X=3.28 $Y=0.815 $X2=0 $Y2=0
cc_285 N_X_c_449_n N_VGND_M1015_s 2.28588e-19 $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_286 N_X_c_452_n N_VGND_M1015_s 0.00344973f $X=3.932 $Y=0.905 $X2=0 $Y2=0
cc_287 N_X_c_462_n N_VGND_c_526_n 0.0151398f $X=2.605 $Y=0.485 $X2=0 $Y2=0
cc_288 N_X_c_447_n N_VGND_c_526_n 0.00198695f $X=3.28 $Y=0.815 $X2=0 $Y2=0
cc_289 N_X_c_447_n N_VGND_c_527_n 0.0122559f $X=3.28 $Y=0.815 $X2=0 $Y2=0
cc_290 N_X_c_452_n N_VGND_c_528_n 0.00173903f $X=3.932 $Y=0.905 $X2=0 $Y2=0
cc_291 N_X_c_449_n N_VGND_c_529_n 0.00177288f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_292 N_X_c_452_n N_VGND_c_529_n 0.0120207f $X=3.932 $Y=0.905 $X2=0 $Y2=0
cc_293 N_X_c_447_n N_VGND_c_531_n 0.00198695f $X=3.28 $Y=0.815 $X2=0 $Y2=0
cc_294 N_X_c_477_n N_VGND_c_531_n 0.0188551f $X=3.445 $Y=0.39 $X2=0 $Y2=0
cc_295 N_X_c_449_n N_VGND_c_531_n 0.00198695f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_296 N_X_M1001_d N_VGND_c_535_n 0.00393857f $X=2.47 $Y=0.235 $X2=0 $Y2=0
cc_297 N_X_M1006_d N_VGND_c_535_n 0.00215201f $X=3.31 $Y=0.235 $X2=0 $Y2=0
cc_298 N_X_c_462_n N_VGND_c_535_n 0.00940698f $X=2.605 $Y=0.485 $X2=0 $Y2=0
cc_299 N_X_c_447_n N_VGND_c_535_n 0.00835832f $X=3.28 $Y=0.815 $X2=0 $Y2=0
cc_300 N_X_c_477_n N_VGND_c_535_n 0.0122069f $X=3.445 $Y=0.39 $X2=0 $Y2=0
cc_301 N_X_c_449_n N_VGND_c_535_n 0.00396723f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_302 N_X_c_452_n N_VGND_c_535_n 0.0035992f $X=3.932 $Y=0.905 $X2=0 $Y2=0

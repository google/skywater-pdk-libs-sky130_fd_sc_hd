* File: sky130_fd_sc_hd__or2b_1.spice.SKY130_FD_SC_HD__OR2B_1.pxi
* Created: Thu Aug 27 14:42:55 2020
* 
x_PM_SKY130_FD_SC_HD__OR2B_1%B_N N_B_N_M1003_g N_B_N_M1007_g B_N N_B_N_c_57_n
+ B_N PM_SKY130_FD_SC_HD__OR2B_1%B_N
x_PM_SKY130_FD_SC_HD__OR2B_1%A_27_53# N_A_27_53#_M1003_s N_A_27_53#_M1007_d
+ N_A_27_53#_M1002_g N_A_27_53#_M1005_g N_A_27_53#_c_82_n N_A_27_53#_c_83_n
+ N_A_27_53#_c_84_n N_A_27_53#_c_89_n N_A_27_53#_c_85_n N_A_27_53#_c_86_n
+ N_A_27_53#_c_87_n PM_SKY130_FD_SC_HD__OR2B_1%A_27_53#
x_PM_SKY130_FD_SC_HD__OR2B_1%A N_A_c_130_n N_A_M1001_g N_A_M1006_g A N_A_c_133_n
+ PM_SKY130_FD_SC_HD__OR2B_1%A
x_PM_SKY130_FD_SC_HD__OR2B_1%A_219_297# N_A_219_297#_M1002_d
+ N_A_219_297#_M1005_s N_A_219_297#_M1004_g N_A_219_297#_M1000_g
+ N_A_219_297#_c_177_n N_A_219_297#_c_216_p N_A_219_297#_c_165_n
+ N_A_219_297#_c_166_n N_A_219_297#_c_172_n N_A_219_297#_c_173_n
+ N_A_219_297#_c_167_n N_A_219_297#_c_168_n N_A_219_297#_c_169_n
+ N_A_219_297#_c_170_n PM_SKY130_FD_SC_HD__OR2B_1%A_219_297#
x_PM_SKY130_FD_SC_HD__OR2B_1%VPWR N_VPWR_M1007_s N_VPWR_M1006_d N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n VPWR N_VPWR_c_227_n N_VPWR_c_228_n
+ N_VPWR_c_223_n N_VPWR_c_230_n PM_SKY130_FD_SC_HD__OR2B_1%VPWR
x_PM_SKY130_FD_SC_HD__OR2B_1%X N_X_M1004_d N_X_M1000_d N_X_c_256_n N_X_c_258_n
+ N_X_c_257_n X PM_SKY130_FD_SC_HD__OR2B_1%X
x_PM_SKY130_FD_SC_HD__OR2B_1%VGND N_VGND_M1003_d N_VGND_M1001_d N_VGND_c_272_n
+ VGND N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n N_VGND_c_276_n
+ N_VGND_c_277_n N_VGND_c_278_n PM_SKY130_FD_SC_HD__OR2B_1%VGND
cc_1 VNB N_B_N_M1003_g 0.0404018f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB B_N 0.0092769f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_B_N_c_57_n 0.0401388f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_53#_M1002_g 0.0326337f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_53#_c_82_n 0.0195877f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_6 VNB N_A_27_53#_c_83_n 0.00282658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_53#_c_84_n 0.00888346f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_8 VNB N_A_27_53#_c_85_n 0.00460073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_86_n 0.0127866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_53#_c_87_n 0.0346763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_M1001_g 0.0415133f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_12 VNB N_A_219_297#_c_165_n 0.00188528f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_13 VNB N_A_219_297#_c_166_n 0.00407348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_219_297#_c_167_n 0.00315488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_219_297#_c_168_n 0.0233712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_219_297#_c_169_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_219_297#_c_170_n 0.0197132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_223_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_256_n 0.0137322f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_20 VNB N_X_c_257_n 0.024426f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_21 VNB N_VGND_c_272_n 6.33456e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_VGND_c_273_n 0.0122945f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_23 VNB N_VGND_c_274_n 0.0164993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_275_n 0.168315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_276_n 0.0174489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_277_n 0.0191933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_278_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_B_N_M1007_g 0.0294136f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_29 VPB B_N 8.85293e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_30 VPB N_B_N_c_57_n 0.0102372f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_31 VPB N_A_27_53#_M1005_g 0.0226524f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_32 VPB N_A_27_53#_c_89_n 0.00457509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_53#_c_85_n 0.00639441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_53#_c_86_n 0.00348764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_53#_c_87_n 0.00826971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_c_130_n 0.043427f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_37 VPB N_A_M1001_g 0.0314341f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_38 VPB A 0.0264491f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_39 VPB N_A_c_133_n 0.0371693f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_40 VPB N_A_219_297#_M1000_g 0.0244633f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_41 VPB N_A_219_297#_c_172_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_219_297#_c_173_n 0.00815415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_219_297#_c_167_n 2.03541e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_219_297#_c_168_n 0.00498459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_224_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_46 VPB N_VPWR_c_225_n 0.0553789f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_VPWR_c_226_n 0.0119713f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_48 VPB N_VPWR_c_227_n 0.0397045f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_49 VPB N_VPWR_c_228_n 0.0176015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_223_n 0.0620391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_230_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_258_n 0.0051537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_X_c_257_n 0.00886361f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_54 VPB X 0.0321952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_B_N_M1003_g N_A_27_53#_c_82_n 0.0125629f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_56 N_B_N_M1003_g N_A_27_53#_c_83_n 0.0129453f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_57 B_N N_A_27_53#_c_83_n 3.15358e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_B_N_M1003_g N_A_27_53#_c_84_n 0.00412847f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_59 B_N N_A_27_53#_c_84_n 0.0254117f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_60 N_B_N_c_57_n N_A_27_53#_c_84_n 0.00729063f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_61 N_B_N_c_57_n N_A_27_53#_c_89_n 0.008428f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B_N_M1003_g N_A_27_53#_c_86_n 0.0100022f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_63 B_N N_A_27_53#_c_86_n 0.0193147f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_64 N_B_N_c_57_n N_A_27_53#_c_87_n 0.00524525f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_65 N_B_N_M1007_g A 2.52857e-19 $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_66 N_B_N_M1007_g N_A_219_297#_c_173_n 0.00135549f $X=0.47 $Y=1.695 $X2=0
+ $Y2=0
cc_67 N_B_N_M1007_g N_VPWR_c_225_n 0.00615653f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_68 B_N N_VPWR_c_225_n 0.020379f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_69 N_B_N_c_57_n N_VPWR_c_225_n 0.0054329f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B_N_M1007_g N_VPWR_c_227_n 0.00317366f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_71 N_B_N_M1007_g N_VPWR_c_223_n 0.00403572f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_72 N_B_N_M1003_g N_VGND_c_275_n 0.0073571f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_73 N_B_N_M1003_g N_VGND_c_276_n 0.00402941f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_74 N_B_N_M1003_g N_VGND_c_277_n 0.00505351f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_75 N_A_27_53#_M1005_g N_A_c_130_n 0.00868417f $X=1.43 $Y=1.695 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_27_53#_M1002_g N_A_M1001_g 0.022046f $X=1.37 $Y=0.475 $X2=0 $Y2=0
cc_77 N_A_27_53#_c_85_n N_A_M1001_g 0.0014977f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_27_53#_c_87_n N_A_M1001_g 0.0652533f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_27_53#_M1005_g A 0.00164982f $X=1.43 $Y=1.695 $X2=0 $Y2=0
cc_80 N_A_27_53#_c_89_n A 0.0122083f $X=0.68 $Y=1.62 $X2=0 $Y2=0
cc_81 N_A_27_53#_M1005_g N_A_219_297#_c_177_n 0.00917186f $X=1.43 $Y=1.695 $X2=0
+ $Y2=0
cc_82 N_A_27_53#_M1002_g N_A_219_297#_c_166_n 0.00310482f $X=1.37 $Y=0.475 $X2=0
+ $Y2=0
cc_83 N_A_27_53#_c_86_n N_A_219_297#_c_166_n 0.00301599f $X=0.72 $Y=0.82 $X2=0
+ $Y2=0
cc_84 N_A_27_53#_c_87_n N_A_219_297#_c_166_n 3.34812e-19 $X=1.43 $Y=1.16 $X2=0
+ $Y2=0
cc_85 N_A_27_53#_M1005_g N_A_219_297#_c_173_n 0.0100132f $X=1.43 $Y=1.695 $X2=0
+ $Y2=0
cc_86 N_A_27_53#_c_89_n N_A_219_297#_c_173_n 0.0253575f $X=0.68 $Y=1.62 $X2=0
+ $Y2=0
cc_87 N_A_27_53#_c_85_n N_A_219_297#_c_173_n 0.0263501f $X=1.22 $Y=1.16 $X2=0
+ $Y2=0
cc_88 N_A_27_53#_c_87_n N_A_219_297#_c_173_n 0.0062777f $X=1.43 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_27_53#_M1002_g N_VGND_c_272_n 5.2524e-19 $X=1.37 $Y=0.475 $X2=0 $Y2=0
cc_90 N_A_27_53#_M1002_g N_VGND_c_273_n 0.00442511f $X=1.37 $Y=0.475 $X2=0 $Y2=0
cc_91 N_A_27_53#_M1002_g N_VGND_c_275_n 0.00779323f $X=1.37 $Y=0.475 $X2=0 $Y2=0
cc_92 N_A_27_53#_c_82_n N_VGND_c_275_n 0.0116656f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_27_53#_c_83_n N_VGND_c_275_n 0.0038498f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_94 N_A_27_53#_c_86_n N_VGND_c_275_n 0.00105248f $X=0.72 $Y=0.82 $X2=0 $Y2=0
cc_95 N_A_27_53#_c_82_n N_VGND_c_276_n 0.0183741f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_27_53#_c_83_n N_VGND_c_276_n 0.00229799f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_97 N_A_27_53#_M1002_g N_VGND_c_277_n 0.00956971f $X=1.37 $Y=0.475 $X2=0 $Y2=0
cc_98 N_A_27_53#_c_85_n N_VGND_c_277_n 0.0188842f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_27_53#_c_86_n N_VGND_c_277_n 0.0214575f $X=0.72 $Y=0.82 $X2=0 $Y2=0
cc_100 N_A_27_53#_c_87_n N_VGND_c_277_n 0.00387909f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_M1001_g N_A_219_297#_M1000_g 0.0251997f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_102 N_A_c_130_n N_A_219_297#_c_177_n 6.94119e-19 $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_103 N_A_M1001_g N_A_219_297#_c_177_n 0.0166311f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_104 A N_A_219_297#_c_177_n 0.0108145f $X=1.07 $Y=2.125 $X2=0 $Y2=0
cc_105 N_A_M1001_g N_A_219_297#_c_165_n 0.0134565f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_106 N_A_c_130_n N_A_219_297#_c_173_n 9.41055e-19 $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_107 N_A_M1001_g N_A_219_297#_c_173_n 0.00122623f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_108 A N_A_219_297#_c_173_n 0.034396f $X=1.07 $Y=2.125 $X2=0 $Y2=0
cc_109 N_A_c_133_n N_A_219_297#_c_173_n 0.00119166f $X=1.175 $Y=2.28 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_A_219_297#_c_168_n 0.0195827f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_111 N_A_M1001_g N_A_219_297#_c_169_n 0.0136533f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_112 N_A_M1001_g N_A_219_297#_c_170_n 0.0172581f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_113 A N_VPWR_c_225_n 0.025857f $X=1.07 $Y=2.125 $X2=0 $Y2=0
cc_114 N_A_c_133_n N_VPWR_c_225_n 0.00100508f $X=1.175 $Y=2.28 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_VPWR_c_226_n 0.00820852f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_116 A N_VPWR_c_226_n 0.0259888f $X=1.07 $Y=2.125 $X2=0 $Y2=0
cc_117 A N_VPWR_c_227_n 0.0587489f $X=1.07 $Y=2.125 $X2=0 $Y2=0
cc_118 N_A_c_133_n N_VPWR_c_227_n 0.0214212f $X=1.175 $Y=2.28 $X2=0 $Y2=0
cc_119 A N_VPWR_c_223_n 0.0432687f $X=1.07 $Y=2.125 $X2=0 $Y2=0
cc_120 N_A_c_133_n N_VPWR_c_223_n 0.0300519f $X=1.175 $Y=2.28 $X2=0 $Y2=0
cc_121 N_A_M1001_g N_VGND_c_272_n 0.00709022f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_122 N_A_M1001_g N_VGND_c_273_n 0.00322006f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_123 N_A_M1001_g N_VGND_c_275_n 0.00390029f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_124 N_A_M1001_g N_VGND_c_277_n 5.59171e-19 $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_125 N_A_219_297#_c_177_n N_VPWR_M1006_d 0.00526233f $X=2.065 $Y=1.58 $X2=0
+ $Y2=0
cc_126 N_A_219_297#_c_173_n N_VPWR_c_225_n 6.48777e-19 $X=1.2 $Y=1.58 $X2=0
+ $Y2=0
cc_127 N_A_219_297#_M1000_g N_VPWR_c_226_n 0.00485906f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_219_297#_c_177_n N_VPWR_c_226_n 0.0190361f $X=2.065 $Y=1.58 $X2=0
+ $Y2=0
cc_129 N_A_219_297#_c_173_n N_VPWR_c_226_n 0.00145048f $X=1.2 $Y=1.58 $X2=0
+ $Y2=0
cc_130 N_A_219_297#_c_168_n N_VPWR_c_226_n 3.85151e-19 $X=2.21 $Y=1.16 $X2=0
+ $Y2=0
cc_131 N_A_219_297#_M1000_g N_VPWR_c_228_n 0.00585385f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_219_297#_M1000_g N_VPWR_c_223_n 0.0128394f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_219_297#_c_177_n A_301_297# 0.0033195f $X=2.065 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_219_297#_c_165_n N_X_c_257_n 0.00357198f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_219_297#_c_172_n N_X_c_257_n 0.00852743f $X=2.15 $Y=1.495 $X2=0 $Y2=0
cc_136 N_A_219_297#_c_167_n N_X_c_257_n 0.0205999f $X=2.21 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_219_297#_c_169_n N_X_c_257_n 0.00848187f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_219_297#_c_170_n N_X_c_257_n 0.0154137f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_219_297#_c_165_n N_VGND_M1001_d 0.00482895f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_140 N_A_219_297#_c_169_n N_VGND_M1001_d 6.98847e-19 $X=2.18 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_219_297#_c_165_n N_VGND_c_272_n 0.020701f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_219_297#_c_168_n N_VGND_c_272_n 4.03696e-19 $X=2.21 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_219_297#_c_170_n N_VGND_c_272_n 0.0132447f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A_219_297#_c_216_p N_VGND_c_273_n 0.00846569f $X=1.58 $Y=0.47 $X2=0
+ $Y2=0
cc_145 N_A_219_297#_c_165_n N_VGND_c_273_n 0.00232396f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_219_297#_c_165_n N_VGND_c_274_n 3.34073e-19 $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_219_297#_c_170_n N_VGND_c_274_n 0.00524631f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_219_297#_c_216_p N_VGND_c_275_n 0.00625722f $X=1.58 $Y=0.47 $X2=0
+ $Y2=0
cc_149 N_A_219_297#_c_165_n N_VGND_c_275_n 0.00637905f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_219_297#_c_170_n N_VGND_c_275_n 0.00951256f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_VPWR_c_223_n N_X_M1000_d 0.0039537f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_152 N_VPWR_c_228_n X 0.0187043f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_223_n X 0.0103212f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_154 N_X_c_256_n N_VGND_c_274_n 0.00876347f $X=2.59 $Y=0.587 $X2=0 $Y2=0
cc_155 N_X_M1004_d N_VGND_c_275_n 0.00411498f $X=2.355 $Y=0.235 $X2=0 $Y2=0
cc_156 N_X_c_256_n N_VGND_c_275_n 0.00924648f $X=2.59 $Y=0.587 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o2bb2ai_2.spice
* Created: Tue Sep  1 19:24:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2bb2ai_2.pex.spice"
.subckt sky130_fd_sc_hd__o2bb2ai_2  VNB VPB A1_N A2_N B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A1_N_M1010_g N_A_113_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_A_113_47#_M1010_s N_A2_N_M1004_g N_A_113_297#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_A_113_47#_M1005_d N_A2_N_M1005_g N_A_113_297#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A1_N_M1011_g N_A_113_47#_M1005_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1012_d N_A_113_297#_M1012_g N_A_471_47#_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.1755 PD=0.92 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1012_d N_A_113_297#_M1015_g N_A_471_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.099125 PD=0.92 PS=0.955 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g N_A_471_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.099125 PD=0.92 PS=0.955 NRD=0 NRS=5.532 M=1 R=4.33333
+ SA=75001.1 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1001 N_A_471_47#_M1001_d N_B2_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 N_A_471_47#_M1001_d N_B2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1009_s N_B1_M1007_g N_A_471_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_113_297#_M1002_d N_A1_N_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.6 A=0.15 P=2.3 MULT=1
MM1014 N_A_113_297#_M1002_d N_A2_N_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1017 N_A_113_297#_M1017_d N_A2_N_M1017_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1013 N_A_113_297#_M1017_d N_A1_N_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.4 PD=1.27 PS=1.8 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75003.3
+ A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1013_s N_A_113_297#_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.4 AS=0.135 PD=1.8 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A_113_297#_M1019_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.135 PD=1.305 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1019_d N_B1_M1000_g N_A_730_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.135 PD=1.305 PS=1.27 NRD=5.8903 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1003 N_A_730_297#_M1000_s N_B2_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.7
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1008 N_A_730_297#_M1008_d N_B2_M1008_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1018_d N_B1_M1018_g N_A_730_297#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_90 VPB 0 3.27631e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__o2bb2ai_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o221ai_1.spice.pex
* Created: Thu Aug 27 14:37:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O221AI_1%C1 1 3 4 6 8 12
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.38
+ $Y=1.16 $X2=0.38 $Y2=1.16
r26 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.23 $Y=1.16 $X2=0.38
+ $Y2=1.16
r27 4 11 38.5363 $w=3.15e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.405 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r29 1 11 38.5363 $w=3.15e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.405 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%B1 3 6 8 11 12 13
r30 11 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=1.16
+ $X2=1.305 $Y2=1.325
r31 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=1.16
+ $X2=1.305 $Y2=0.995
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r33 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.27
+ $Y2=1.16
r34 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.4 $Y=1.985 $X2=1.4
+ $Y2=1.325
r35 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.4 $Y=0.56 $X2=1.4
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%B2 3 7 8 11 13
c37 11 0 8.87346e-20 $X=1.85 $Y=1.16
r38 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=1.325
r39 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=0.995
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.16 $X2=1.85 $Y2=1.16
r41 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.56 $X2=1.82
+ $Y2=0.995
r42 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.79 $Y=1.985
+ $X2=1.79 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%A2 1 3 6 9 11 12 18 20
c46 9 0 8.68947e-20 $X=2.4 $Y=1.445
r47 18 20 14.8143 $w=2.1e-07 $l=2.55e-07 $layer=LI1_cond $X=2.57 $Y=1.615
+ $X2=2.57 $Y2=1.87
r48 12 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.16
+ $X2=2.33 $Y2=1.325
r49 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.16 $X2=2.33 $Y2=1.16
r50 9 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.4 $Y=1.53 $X2=2.57
+ $Y2=1.53
r51 9 11 10.5628 $w=2.08e-07 $l=2e-07 $layer=LI1_cond $X=2.4 $Y=1.445 $X2=2.4
+ $Y2=1.245
r52 6 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.39 $Y=1.985
+ $X2=2.39 $Y2=1.325
r53 1 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=0.995
+ $X2=2.33 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.33 $Y=0.995 $X2=2.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%A1 1 3 6 8 13
c26 8 0 1.83983e-21 $X=2.99 $Y=1.19
r27 10 13 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.935 $Y2=1.16
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.16 $X2=2.935 $Y2=1.16
r29 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.325
+ $X2=2.75 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.325 $X2=2.75
+ $Y2=1.985
r31 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=0.995
+ $X2=2.75 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.995 $X2=2.75
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%Y 1 2 3 10 13 15 17 18 19 22 23 27 28 29
r60 32 34 1.5443 $w=4.74e-07 $l=6e-08 $layer=LI1_cond $X=1.99 $Y=1.6 $X2=1.99
+ $Y2=1.66
r61 29 38 5.40506 $w=4.74e-07 $l=2.1e-07 $layer=LI1_cond $X=1.99 $Y=2.21
+ $X2=1.99 $Y2=2
r62 28 38 3.34599 $w=4.74e-07 $l=1.3e-07 $layer=LI1_cond $X=1.99 $Y=1.87
+ $X2=1.99 $Y2=2
r63 28 34 5.40506 $w=4.74e-07 $l=2.1e-07 $layer=LI1_cond $X=1.99 $Y=1.87
+ $X2=1.99 $Y2=1.66
r64 24 27 5.06322 $w=2.1e-07 $l=1.03e-07 $layer=LI1_cond $X=0.84 $Y=1.6
+ $X2=0.737 $Y2=1.6
r65 23 32 5.52649 $w=2.1e-07 $l=2.55e-07 $layer=LI1_cond $X=1.735 $Y=1.6
+ $X2=1.99 $Y2=1.6
r66 23 24 47.2684 $w=2.08e-07 $l=8.95e-07 $layer=LI1_cond $X=1.735 $Y=1.6
+ $X2=0.84 $Y2=1.6
r67 22 27 1.42948 $w=2.05e-07 $l=1.05e-07 $layer=LI1_cond $X=0.737 $Y=1.495
+ $X2=0.737 $Y2=1.6
r68 21 22 36.2483 $w=2.03e-07 $l=6.7e-07 $layer=LI1_cond $X=0.737 $Y=0.825
+ $X2=0.737 $Y2=1.495
r69 20 26 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.6
+ $X2=0.225 $Y2=1.6
r70 19 27 5.06322 $w=2.1e-07 $l=1.02e-07 $layer=LI1_cond $X=0.635 $Y=1.6
+ $X2=0.737 $Y2=1.6
r71 19 20 14.2597 $w=2.08e-07 $l=2.7e-07 $layer=LI1_cond $X=0.635 $Y=1.6
+ $X2=0.365 $Y2=1.6
r72 17 21 6.85394 $w=1.8e-07 $l=1.39943e-07 $layer=LI1_cond $X=0.635 $Y=0.735
+ $X2=0.737 $Y2=0.825
r73 17 18 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.635 $Y=0.735
+ $X2=0.345 $Y2=0.735
r74 13 26 2.99957 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.225 $Y=1.705
+ $X2=0.225 $Y2=1.6
r75 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=1.705
+ $X2=0.225 $Y2=1.96
r76 10 18 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=0.645
+ $X2=0.345 $Y2=0.735
r77 10 12 2.34615 $w=2.6e-07 $l=5e-08 $layer=LI1_cond $X=0.215 $Y=0.645
+ $X2=0.215 $Y2=0.595
r78 3 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.485 $X2=2 $Y2=2
r79 3 34 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.485 $X2=2 $Y2=1.66
r80 2 26 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r81 2 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
r82 1 12 182 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%VPWR 1 2 7 9 13 15 20 29 37
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 29 32 11.5066 $w=7.88e-07 $l=7.6e-07 $layer=LI1_cond $X=0.945 $Y=1.96
+ $X2=0.945 $Y2=2.72
r45 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 24 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 24 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 23 26 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 21 32 10.1246 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=1.34 $Y=2.72
+ $X2=0.945 $Y2=2.72
r52 21 23 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.34 $Y=2.72 $X2=1.61
+ $Y2=2.72
r53 20 36 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=3.047 $Y2=2.72
r54 20 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 15 32 10.1246 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=0.55 $Y=2.72
+ $X2=0.945 $Y2=2.72
r56 15 17 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=0.23
+ $Y2=2.72
r57 13 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 13 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r59 9 12 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.005 $Y=1.66
+ $X2=3.005 $Y2=2.34
r60 7 36 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.005 $Y=2.635
+ $X2=3.047 $Y2=2.72
r61 7 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.005 $Y=2.635
+ $X2=3.005 $Y2=2.34
r62 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=2.34
r63 2 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.66
r64 1 29 150 $w=1.7e-07 $l=8.13542e-07 $layer=licon1_PDIFF $count=4 $X=0.565
+ $Y=1.485 $X2=1.175 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%A_109_47# 1 2 11
r14 8 11 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.68 $Y=0.39 $X2=1.61
+ $Y2=0.39
r15 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.235 $X2=1.61 $Y2=0.39
r16 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%A_213_123# 1 2 3 10 16 20 23
r43 18 20 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.965 $Y=0.695
+ $X2=2.965 $Y2=0.39
r44 17 23 7.38875 $w=1.75e-07 $l=3.35783e-07 $layer=LI1_cond $X=2.22 $Y=0.78
+ $X2=1.945 $Y2=0.645
r45 16 18 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.795 $Y=0.78
+ $X2=2.965 $Y2=0.695
r46 16 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.795 $Y=0.78
+ $X2=2.22 $Y2=0.78
r47 10 23 7.38875 $w=1.75e-07 $l=9e-08 $layer=LI1_cond $X=1.945 $Y=0.735
+ $X2=1.945 $Y2=0.645
r48 10 12 46.5202 $w=1.78e-07 $l=7.55e-07 $layer=LI1_cond $X=1.945 $Y=0.735
+ $X2=1.19 $Y2=0.735
r49 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.39
r50 2 23 182 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.03 $Y2=0.66
r51 1 12 182 $w=1.7e-07 $l=1.73205e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.615 $X2=1.19 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_1%VGND 1 6 8 10 17 18 21
r40 21 22 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r41 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r42 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r43 15 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.54
+ $Y2=0
r44 15 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.99
+ $Y2=0
r45 10 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.54
+ $Y2=0
r46 10 12 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=2.455 $Y=0 $X2=0.23
+ $Y2=0
r47 8 22 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r48 8 12 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r49 4 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085 $X2=2.54
+ $Y2=0
r50 4 6 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.36
r51 1 6 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.405
+ $Y=0.235 $X2=2.54 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__a221o_4.pxi.spice
* Created: Tue Sep  1 18:52:47 2020
* 
x_PM_SKY130_FD_SC_HD__A221O_4%A_79_21# N_A_79_21#_M1007_d N_A_79_21#_M1009_d
+ N_A_79_21#_M1020_s N_A_79_21#_M1014_s N_A_79_21#_M1002_s N_A_79_21#_c_125_n
+ N_A_79_21#_M1011_g N_A_79_21#_M1003_g N_A_79_21#_c_126_n N_A_79_21#_M1013_g
+ N_A_79_21#_M1005_g N_A_79_21#_c_127_n N_A_79_21#_M1015_g N_A_79_21#_M1016_g
+ N_A_79_21#_c_128_n N_A_79_21#_M1026_g N_A_79_21#_M1025_g N_A_79_21#_c_129_n
+ N_A_79_21#_c_141_n N_A_79_21#_c_142_n N_A_79_21#_c_196_p N_A_79_21#_c_130_n
+ N_A_79_21#_c_166_p N_A_79_21#_c_131_n N_A_79_21#_c_132_n N_A_79_21#_c_174_p
+ N_A_79_21#_c_169_p N_A_79_21#_c_133_n N_A_79_21#_c_134_n N_A_79_21#_c_144_n
+ N_A_79_21#_c_135_n N_A_79_21#_c_136_n PM_SKY130_FD_SC_HD__A221O_4%A_79_21#
x_PM_SKY130_FD_SC_HD__A221O_4%A2 N_A2_c_311_n N_A2_M1019_g N_A2_M1006_g
+ N_A2_c_312_n N_A2_M1024_g N_A2_M1021_g A2 N_A2_c_314_n
+ PM_SKY130_FD_SC_HD__A221O_4%A2
x_PM_SKY130_FD_SC_HD__A221O_4%A1 N_A1_M1001_g N_A1_M1022_g N_A1_c_359_n
+ N_A1_M1007_g N_A1_c_360_n N_A1_M1009_g A1 A1 N_A1_c_362_n N_A1_c_363_n
+ N_A1_c_406_p PM_SKY130_FD_SC_HD__A221O_4%A1
x_PM_SKY130_FD_SC_HD__A221O_4%C1 N_C1_c_418_n N_C1_M1012_g N_C1_M1002_g
+ N_C1_c_419_n N_C1_M1020_g N_C1_M1008_g C1 N_C1_c_420_n N_C1_c_421_n C1
+ PM_SKY130_FD_SC_HD__A221O_4%C1
x_PM_SKY130_FD_SC_HD__A221O_4%B1 N_B1_c_471_n N_B1_M1010_g N_B1_M1017_g
+ N_B1_c_472_n N_B1_M1014_g N_B1_M1023_g N_B1_c_473_n B1 N_B1_c_474_n
+ N_B1_c_475_n PM_SKY130_FD_SC_HD__A221O_4%B1
x_PM_SKY130_FD_SC_HD__A221O_4%B2 N_B2_M1018_g N_B2_c_520_n N_B2_M1000_g
+ N_B2_M1027_g N_B2_c_521_n N_B2_M1004_g B2 N_B2_c_522_n N_B2_c_523_n
+ PM_SKY130_FD_SC_HD__A221O_4%B2
x_PM_SKY130_FD_SC_HD__A221O_4%VPWR N_VPWR_M1003_s N_VPWR_M1005_s N_VPWR_M1025_s
+ N_VPWR_M1021_d N_VPWR_M1022_s N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n
+ N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n
+ N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n
+ N_VPWR_c_577_n VPWR N_VPWR_c_578_n N_VPWR_c_563_n
+ PM_SKY130_FD_SC_HD__A221O_4%VPWR
x_PM_SKY130_FD_SC_HD__A221O_4%X N_X_M1011_s N_X_M1015_s N_X_M1003_d N_X_M1016_d
+ N_X_c_673_n N_X_c_707_n N_X_c_667_n N_X_c_662_n N_X_c_685_n N_X_c_668_n
+ N_X_c_711_n N_X_c_663_n N_X_c_664_n N_X_c_669_n N_X_c_670_n X X X N_X_c_666_n
+ N_X_c_672_n PM_SKY130_FD_SC_HD__A221O_4%X
x_PM_SKY130_FD_SC_HD__A221O_4%A_445_297# N_A_445_297#_M1006_s
+ N_A_445_297#_M1001_d N_A_445_297#_M1017_s N_A_445_297#_M1018_s
+ N_A_445_297#_c_744_n N_A_445_297#_c_745_n N_A_445_297#_c_738_n
+ N_A_445_297#_c_749_n N_A_445_297#_c_739_n N_A_445_297#_c_750_n
+ N_A_445_297#_c_751_n N_A_445_297#_c_740_n N_A_445_297#_c_756_n
+ N_A_445_297#_c_741_n PM_SKY130_FD_SC_HD__A221O_4%A_445_297#
x_PM_SKY130_FD_SC_HD__A221O_4%A_804_297# N_A_804_297#_M1002_d
+ N_A_804_297#_M1008_d N_A_804_297#_M1023_d N_A_804_297#_M1027_d
+ N_A_804_297#_c_810_n N_A_804_297#_c_821_n N_A_804_297#_c_811_n
+ N_A_804_297#_c_844_n PM_SKY130_FD_SC_HD__A221O_4%A_804_297#
x_PM_SKY130_FD_SC_HD__A221O_4%VGND N_VGND_M1011_d N_VGND_M1013_d N_VGND_M1026_d
+ N_VGND_M1024_d N_VGND_M1012_d N_VGND_M1000_d N_VGND_c_845_n N_VGND_c_846_n
+ N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n
+ N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ VGND N_VGND_c_862_n N_VGND_c_863_n PM_SKY130_FD_SC_HD__A221O_4%VGND
x_PM_SKY130_FD_SC_HD__A221O_4%A_445_47# N_A_445_47#_M1019_s N_A_445_47#_M1007_s
+ N_A_445_47#_c_979_n N_A_445_47#_c_972_n N_A_445_47#_c_973_n
+ N_A_445_47#_c_974_n N_A_445_47#_c_975_n N_A_445_47#_c_976_n
+ N_A_445_47#_c_977_n PM_SKY130_FD_SC_HD__A221O_4%A_445_47#
x_PM_SKY130_FD_SC_HD__A221O_4%A_1053_47# N_A_1053_47#_M1010_d
+ N_A_1053_47#_M1000_s N_A_1053_47#_M1004_s N_A_1053_47#_c_1044_n
+ N_A_1053_47#_c_1045_n N_A_1053_47#_c_1046_n N_A_1053_47#_c_1047_n
+ PM_SKY130_FD_SC_HD__A221O_4%A_1053_47#
cc_1 VNB N_A_79_21#_c_125_n 0.0191522f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_126_n 0.0157969f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_127_n 0.0157995f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_128_n 0.0161346f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_129_n 0.00310273f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.18
cc_6 VNB N_A_79_21#_c_130_n 0.00350056f $X=-0.19 $Y=-0.24 $X2=4.055 $Y2=0.39
cc_7 VNB N_A_79_21#_c_131_n 0.00283508f $X=-0.19 $Y=-0.24 $X2=4.18 $Y2=0.725
cc_8 VNB N_A_79_21#_c_132_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=4.815 $Y2=0.815
cc_9 VNB N_A_79_21#_c_133_n 0.00714098f $X=-0.19 $Y=-0.24 $X2=4.98 $Y2=1.455
cc_10 VNB N_A_79_21#_c_134_n 0.00418219f $X=-0.19 $Y=-0.24 $X2=5.82 $Y2=0.38
cc_11 VNB N_A_79_21#_c_135_n 7.47381e-19 $X=-0.19 $Y=-0.24 $X2=4.98 $Y2=0.73
cc_12 VNB N_A_79_21#_c_136_n 0.0677626f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_13 VNB N_A2_c_311_n 0.0154281f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=0.235
cc_14 VNB N_A2_c_312_n 0.0211193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB A2 0.00199071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_314_n 0.0301785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A1_c_359_n 0.0202716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_c_360_n 0.016125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB A1 0.00130173f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_A1_c_362_n 0.0693006f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_21 VNB N_A1_c_363_n 0.00130865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_C1_c_418_n 0.015977f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=0.235
cc_23 VNB N_C1_c_419_n 0.0159693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C1_c_420_n 0.00218913f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_25 VNB N_C1_c_421_n 0.0313814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B1_c_471_n 0.0161181f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=0.235
cc_27 VNB N_B1_c_472_n 0.0214729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_B1_c_473_n 0.0277015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_B1_c_474_n 0.0241668f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_30 VNB N_B1_c_475_n 0.00152344f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_31 VNB N_B2_c_520_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=4.435 $Y2=1.485
cc_32 VNB N_B2_c_521_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_B2_c_522_n 0.0184004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_B2_c_523_n 0.0453669f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_35 VNB N_VPWR_c_563_n 0.326667f $X=-0.19 $Y=-0.24 $X2=5.065 $Y2=0.365
cc_36 VNB N_X_c_662_n 0.00440603f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_37 VNB N_X_c_663_n 9.2445e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_38 VNB N_X_c_664_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_39 VNB X 0.0197123f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_40 VNB N_X_c_666_n 0.00783073f $X=-0.19 $Y=-0.24 $X2=1.68 $Y2=1.16
cc_41 VNB N_VGND_c_845_n 0.0107305f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_42 VNB N_VGND_c_846_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_43 VNB N_VGND_c_847_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_44 VNB N_VGND_c_848_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_849_n 0.00569793f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_46 VNB N_VGND_c_850_n 0.00462966f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_47 VNB N_VGND_c_851_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_48 VNB N_VGND_c_852_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.18
cc_49 VNB N_VGND_c_853_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.18
cc_50 VNB N_VGND_c_854_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_51 VNB N_VGND_c_855_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_856_n 0.0173199f $X=-0.19 $Y=-0.24 $X2=1.68 $Y2=1.16
cc_53 VNB N_VGND_c_857_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=1.68 $Y2=1.16
cc_54 VNB N_VGND_c_858_n 0.0401073f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.455
cc_55 VNB N_VGND_c_859_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=4.405 $Y2=1.54
cc_56 VNB N_VGND_c_860_n 0.0496507f $X=-0.19 $Y=-0.24 $X2=4.055 $Y2=0.39
cc_57 VNB N_VGND_c_861_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=3.3 $Y2=0.39
cc_58 VNB N_VGND_c_862_n 0.0293179f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_59 VNB N_VGND_c_863_n 0.393548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_445_47#_c_972_n 0.00202976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_445_47#_c_973_n 0.00188818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_445_47#_c_974_n 0.0104269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_445_47#_c_975_n 0.00290839f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_64 VNB N_A_445_47#_c_976_n 0.00332212f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_65 VNB N_A_445_47#_c_977_n 0.00305947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1053_47#_c_1044_n 0.0146288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1053_47#_c_1045_n 0.0146572f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_68 VNB N_A_1053_47#_c_1046_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_69 VNB N_A_1053_47#_c_1047_n 5.86661e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VPB N_A_79_21#_M1003_g 0.0219036f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_71 VPB N_A_79_21#_M1005_g 0.0181999f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_72 VPB N_A_79_21#_M1016_g 0.0181974f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_73 VPB N_A_79_21#_M1025_g 0.0187749f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_74 VPB N_A_79_21#_c_141_n 0.00253235f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.455
cc_75 VPB N_A_79_21#_c_142_n 0.0188422f $X=-0.19 $Y=1.305 $X2=4.405 $Y2=1.54
cc_76 VPB N_A_79_21#_c_133_n 0.00281391f $X=-0.19 $Y=1.305 $X2=4.98 $Y2=1.455
cc_77 VPB N_A_79_21#_c_144_n 0.00294106f $X=-0.19 $Y=1.305 $X2=4.57 $Y2=1.62
cc_78 VPB N_A_79_21#_c_136_n 0.0115803f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_79 VPB N_A2_M1006_g 0.0184463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A2_M1021_g 0.0184833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A2_c_314_n 0.00403229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A1_M1001_g 0.0185652f $X=-0.19 $Y=1.305 $X2=4.845 $Y2=0.235
cc_83 VPB N_A1_M1022_g 0.025331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A1_c_362_n 0.0212495f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_85 VPB N_C1_M1002_g 0.0252602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_C1_M1008_g 0.0184521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_C1_c_421_n 0.00409501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_B1_M1017_g 0.0186442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_B1_M1023_g 0.0219398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_B1_c_473_n 0.0037449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_B1_c_474_n 0.00916412f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_92 VPB N_B2_M1018_g 0.0219492f $X=-0.19 $Y=1.305 $X2=4.845 $Y2=0.235
cc_93 VPB N_B2_M1027_g 0.0258456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_B2_c_523_n 0.00977256f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_95 VPB N_VPWR_c_564_n 0.0115433f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_96 VPB N_VPWR_c_565_n 0.00445067f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_97 VPB N_VPWR_c_566_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_567_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_99 VPB N_VPWR_c_568_n 0.00393636f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_100 VPB N_VPWR_c_569_n 0.00456837f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_101 VPB N_VPWR_c_570_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_102 VPB N_VPWR_c_571_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_103 VPB N_VPWR_c_572_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_104 VPB N_VPWR_c_573_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_105 VPB N_VPWR_c_574_n 0.0157745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_575_n 0.00478242f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.18
cc_107 VPB N_VPWR_c_576_n 0.0152829f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_108 VPB N_VPWR_c_577_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_109 VPB N_VPWR_c_578_n 0.0993484f $X=-0.19 $Y=1.305 $X2=4.98 $Y2=1.455
cc_110 VPB N_VPWR_c_563_n 0.069858f $X=-0.19 $Y=1.305 $X2=5.065 $Y2=0.365
cc_111 VPB N_X_c_667_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_112 VPB N_X_c_668_n 0.00226442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_X_c_669_n 0.00100713f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_114 VPB N_X_c_670_n 0.00204609f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_115 VPB X 0.00737886f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_116 VPB N_X_c_672_n 0.00885232f $X=-0.19 $Y=1.305 $X2=1.68 $Y2=1.16
cc_117 VPB N_A_445_297#_c_738_n 0.00222848f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_118 VPB N_A_445_297#_c_739_n 0.00692322f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_119 VPB N_A_445_297#_c_740_n 0.00717103f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_120 VPB N_A_445_297#_c_741_n 0.00208737f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_121 VPB N_A_804_297#_c_810_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_122 VPB N_A_804_297#_c_811_n 0.0039938f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_123 N_A_79_21#_c_128_n N_A2_c_311_n 0.0245549f $X=1.73 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_124 N_A_79_21#_M1025_g N_A2_M1006_g 0.0253675f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_142_n N_A2_M1006_g 0.0162825f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_142_n N_A2_M1021_g 0.0102704f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_129_n A2 0.0115284f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_142_n A2 0.0287857f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_129_n N_A2_c_314_n 0.00191463f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_141_n N_A2_c_314_n 0.00384526f $X=1.9 $Y=1.455 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_142_n N_A2_c_314_n 0.00211509f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_136_n N_A2_c_314_n 0.020495f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_142_n N_A1_M1001_g 0.010346f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_142_n N_A1_M1022_g 0.0124897f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_130_n N_A1_c_359_n 0.00826846f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_130_n N_A1_c_360_n 0.00957565f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_130_n A1 0.00351846f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_131_n A1 4.04651e-19 $X=4.18 $Y=0.725 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_142_n N_A1_c_362_n 0.0187869f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_130_n N_A1_c_362_n 0.00246114f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_142_n N_A1_c_363_n 0.0840565f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_130_n N_A1_c_363_n 0.00124604f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_166_p N_C1_c_418_n 0.00209395f $X=4.18 $Y=0.475 $X2=-0.19
+ $Y2=-0.24
cc_144 N_A_79_21#_c_131_n N_C1_c_418_n 0.0048482f $X=4.18 $Y=0.725 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A_79_21#_c_132_n N_C1_c_418_n 0.00865686f $X=4.815 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_79_21#_c_169_p N_C1_c_418_n 4.58193e-19 $X=4.94 $Y=0.725 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_79_21#_c_142_n N_C1_M1002_g 0.00955985f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_144_n N_C1_M1002_g 0.00512262f $X=4.57 $Y=1.62 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_131_n N_C1_c_419_n 4.58193e-19 $X=4.18 $Y=0.725 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_132_n N_C1_c_419_n 0.00969143f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_174_p N_C1_c_419_n 0.00255288f $X=4.94 $Y=0.475 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_169_p N_C1_c_419_n 0.00376498f $X=4.94 $Y=0.725 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_133_n N_C1_c_419_n 0.00484074f $X=4.98 $Y=1.455 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_135_n N_C1_c_419_n 0.00141025f $X=4.98 $Y=0.73 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_144_n N_C1_M1008_g 0.0115178f $X=4.57 $Y=1.62 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_142_n N_C1_c_420_n 0.0124431f $X=4.405 $Y=1.54 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_131_n N_C1_c_420_n 0.00611226f $X=4.18 $Y=0.725 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_132_n N_C1_c_420_n 0.0300506f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_133_n N_C1_c_420_n 0.016207f $X=4.98 $Y=1.455 $X2=0 $Y2=0
cc_160 N_A_79_21#_c_144_n N_C1_c_420_n 0.0238999f $X=4.57 $Y=1.62 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_132_n N_C1_c_421_n 0.00226432f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_133_n N_C1_c_421_n 0.00526053f $X=4.98 $Y=1.455 $X2=0 $Y2=0
cc_163 N_A_79_21#_c_144_n N_C1_c_421_n 0.00217787f $X=4.57 $Y=1.62 $X2=0 $Y2=0
cc_164 N_A_79_21#_c_135_n N_C1_c_421_n 2.93755e-19 $X=4.98 $Y=0.73 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_133_n N_B1_c_471_n 0.00573857f $X=4.98 $Y=1.455 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_79_21#_c_134_n N_B1_c_471_n 0.0127028f $X=5.82 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_79_21#_c_144_n N_B1_M1017_g 0.00160312f $X=4.57 $Y=1.62 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_134_n N_B1_c_472_n 0.00892725f $X=5.82 $Y=0.38 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_133_n N_B1_c_473_n 0.00432677f $X=4.98 $Y=1.455 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_133_n N_B1_c_475_n 0.0166204f $X=4.98 $Y=1.455 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_134_n N_B2_c_520_n 0.0064046f $X=5.82 $Y=0.38 $X2=0 $Y2=0
cc_172 N_A_79_21#_c_142_n N_VPWR_M1025_s 3.40166e-19 $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_173 N_A_79_21#_c_196_p N_VPWR_M1025_s 0.00156844f $X=1.985 $Y=1.54 $X2=0
+ $Y2=0
cc_174 N_A_79_21#_c_142_n N_VPWR_M1021_d 0.00166235f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_175 N_A_79_21#_c_142_n N_VPWR_M1022_s 0.00276803f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_176 N_A_79_21#_M1003_g N_VPWR_c_565_n 0.00337036f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_79_21#_M1005_g N_VPWR_c_566_n 0.00157837f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_79_21#_M1016_g N_VPWR_c_566_n 0.00157837f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_79_21#_M1025_g N_VPWR_c_567_n 0.00157837f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_79_21#_c_142_n N_VPWR_c_567_n 0.00264836f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_181 N_A_79_21#_c_196_p N_VPWR_c_567_n 0.0108583f $X=1.985 $Y=1.54 $X2=0 $Y2=0
cc_182 N_A_79_21#_M1003_g N_VPWR_c_570_n 0.00585385f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_79_21#_M1005_g N_VPWR_c_570_n 0.00585385f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_79_21#_M1016_g N_VPWR_c_572_n 0.00585385f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_79_21#_M1025_g N_VPWR_c_572_n 0.00585385f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_79_21#_M1002_s N_VPWR_c_563_n 0.00216833f $X=4.435 $Y=1.485 $X2=0
+ $Y2=0
cc_187 N_A_79_21#_M1003_g N_VPWR_c_563_n 0.011391f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_79_21#_M1005_g N_VPWR_c_563_n 0.0104367f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_79_21#_M1016_g N_VPWR_c_563_n 0.0104367f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_79_21#_M1025_g N_VPWR_c_563_n 0.010464f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_125_n N_X_c_673_n 0.0109314f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_126_n N_X_c_673_n 0.00630972f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_127_n N_X_c_673_n 5.22228e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_79_21#_M1005_g N_X_c_667_n 0.0132273f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_79_21#_M1016_g N_X_c_667_n 0.0132131f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_129_n N_X_c_667_n 0.0416643f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_197 N_A_79_21#_c_136_n N_X_c_667_n 0.00211509f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_79_21#_c_126_n N_X_c_662_n 0.00870364f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_79_21#_c_127_n N_X_c_662_n 0.0098365f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_79_21#_c_128_n N_X_c_662_n 0.00255758f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_79_21#_c_129_n N_X_c_662_n 0.0628716f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_202 N_A_79_21#_c_136_n N_X_c_662_n 0.00452472f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_126_n N_X_c_685_n 5.22228e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_79_21#_c_127_n N_X_c_685_n 0.00630972f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_79_21#_c_128_n N_X_c_685_n 0.00630972f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_79_21#_M1025_g N_X_c_668_n 2.57315e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_79_21#_c_129_n N_X_c_668_n 0.0204549f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_196_p N_X_c_668_n 0.00271526f $X=1.985 $Y=1.54 $X2=0 $Y2=0
cc_209 N_A_79_21#_c_136_n N_X_c_668_n 0.00220041f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_79_21#_c_125_n N_X_c_663_n 0.0111076f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_79_21#_c_129_n N_X_c_663_n 0.00134411f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_212 N_A_79_21#_c_125_n N_X_c_664_n 0.00158032f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_79_21#_c_126_n N_X_c_664_n 0.00113286f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_79_21#_c_129_n N_X_c_664_n 0.0266272f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_215 N_A_79_21#_c_136_n N_X_c_664_n 0.00230339f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_79_21#_M1003_g N_X_c_669_n 0.0158771f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_79_21#_c_129_n N_X_c_669_n 0.00413395f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_218 N_A_79_21#_c_129_n N_X_c_670_n 0.0204549f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_136_n N_X_c_670_n 0.00220041f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_79_21#_c_125_n X 0.0206457f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_79_21#_c_129_n X 0.0169898f $X=1.815 $Y=1.18 $X2=0 $Y2=0
cc_222 N_A_79_21#_c_142_n N_A_445_297#_M1006_s 0.00165831f $X=4.405 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_223 N_A_79_21#_c_142_n N_A_445_297#_M1001_d 0.00171146f $X=4.405 $Y=1.54
+ $X2=0 $Y2=0
cc_224 N_A_79_21#_c_142_n N_A_445_297#_c_744_n 0.0315971f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_M1002_s N_A_445_297#_c_745_n 0.0031751f $X=4.435 $Y=1.485
+ $X2=0 $Y2=0
cc_226 N_A_79_21#_c_142_n N_A_445_297#_c_745_n 0.00595197f $X=4.405 $Y=1.54
+ $X2=0 $Y2=0
cc_227 N_A_79_21#_c_144_n N_A_445_297#_c_745_n 0.0312233f $X=4.57 $Y=1.62 $X2=0
+ $Y2=0
cc_228 N_A_79_21#_c_144_n N_A_445_297#_c_738_n 0.0142624f $X=4.57 $Y=1.62 $X2=0
+ $Y2=0
cc_229 N_A_79_21#_c_144_n N_A_445_297#_c_749_n 0.00243741f $X=4.57 $Y=1.62 $X2=0
+ $Y2=0
cc_230 N_A_79_21#_c_142_n N_A_445_297#_c_750_n 0.0126766f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_c_142_n N_A_445_297#_c_751_n 0.0130829f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_c_142_n N_A_445_297#_c_740_n 0.060643f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_c_142_n N_A_804_297#_M1002_d 0.00287043f $X=4.405 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_234 N_A_79_21#_c_144_n N_A_804_297#_M1008_d 0.00346199f $X=4.57 $Y=1.62 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_M1002_s N_A_804_297#_c_811_n 0.00316492f $X=4.435 $Y=1.485
+ $X2=0 $Y2=0
cc_236 N_A_79_21#_c_132_n N_VGND_M1012_d 0.00162089f $X=4.815 $Y=0.815 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_125_n N_VGND_c_846_n 0.00316354f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_79_21#_c_126_n N_VGND_c_847_n 0.00146448f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_79_21#_c_127_n N_VGND_c_847_n 0.00146448f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_c_128_n N_VGND_c_848_n 0.00146448f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_79_21#_c_142_n N_VGND_c_849_n 0.00308977f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_242 N_A_79_21#_c_130_n N_VGND_c_849_n 0.0117888f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_243 N_A_79_21#_c_132_n N_VGND_c_850_n 0.0122559f $X=4.815 $Y=0.815 $X2=0
+ $Y2=0
cc_244 N_A_79_21#_c_125_n N_VGND_c_852_n 0.00424416f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_79_21#_c_126_n N_VGND_c_852_n 0.00423334f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_79_21#_c_127_n N_VGND_c_854_n 0.00423334f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_79_21#_c_128_n N_VGND_c_854_n 0.00541359f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_79_21#_c_130_n N_VGND_c_858_n 0.0418793f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_249 N_A_79_21#_c_166_p N_VGND_c_858_n 0.0114777f $X=4.18 $Y=0.475 $X2=0 $Y2=0
cc_250 N_A_79_21#_c_132_n N_VGND_c_858_n 0.00198695f $X=4.815 $Y=0.815 $X2=0
+ $Y2=0
cc_251 N_A_79_21#_c_132_n N_VGND_c_860_n 0.00198695f $X=4.815 $Y=0.815 $X2=0
+ $Y2=0
cc_252 N_A_79_21#_c_174_p N_VGND_c_860_n 0.015247f $X=4.94 $Y=0.475 $X2=0 $Y2=0
cc_253 N_A_79_21#_c_134_n N_VGND_c_860_n 0.0522924f $X=5.82 $Y=0.38 $X2=0 $Y2=0
cc_254 N_A_79_21#_M1007_d N_VGND_c_863_n 0.00172388f $X=3.175 $Y=0.235 $X2=0
+ $Y2=0
cc_255 N_A_79_21#_M1009_d N_VGND_c_863_n 0.00218529f $X=4.005 $Y=0.235 $X2=0
+ $Y2=0
cc_256 N_A_79_21#_M1020_s N_VGND_c_863_n 0.00215206f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_257 N_A_79_21#_M1014_s N_VGND_c_863_n 0.00209344f $X=5.685 $Y=0.235 $X2=0
+ $Y2=0
cc_258 N_A_79_21#_c_125_n N_VGND_c_863_n 0.00669028f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_79_21#_c_126_n N_VGND_c_863_n 0.0057163f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_79_21#_c_127_n N_VGND_c_863_n 0.0057163f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_79_21#_c_128_n N_VGND_c_863_n 0.00952874f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_79_21#_c_130_n N_VGND_c_863_n 0.0230478f $X=4.055 $Y=0.39 $X2=0 $Y2=0
cc_263 N_A_79_21#_c_166_p N_VGND_c_863_n 0.00913984f $X=4.18 $Y=0.475 $X2=0
+ $Y2=0
cc_264 N_A_79_21#_c_132_n N_VGND_c_863_n 0.00835832f $X=4.815 $Y=0.815 $X2=0
+ $Y2=0
cc_265 N_A_79_21#_c_174_p N_VGND_c_863_n 0.00941474f $X=4.94 $Y=0.475 $X2=0
+ $Y2=0
cc_266 N_A_79_21#_c_134_n N_VGND_c_863_n 0.0329455f $X=5.82 $Y=0.38 $X2=0 $Y2=0
cc_267 N_A_79_21#_c_130_n N_A_445_47#_M1007_s 0.00318958f $X=4.055 $Y=0.39 $X2=0
+ $Y2=0
cc_268 N_A_79_21#_c_128_n N_A_445_47#_c_979_n 5.51569e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_79_21#_M1007_d N_A_445_47#_c_972_n 0.00416469f $X=3.175 $Y=0.235
+ $X2=0 $Y2=0
cc_270 N_A_79_21#_c_130_n N_A_445_47#_c_972_n 0.0148984f $X=4.055 $Y=0.39 $X2=0
+ $Y2=0
cc_271 N_A_79_21#_c_130_n N_A_445_47#_c_973_n 0.0130697f $X=4.055 $Y=0.39 $X2=0
+ $Y2=0
cc_272 N_A_79_21#_c_131_n N_A_445_47#_c_973_n 0.00832371f $X=4.18 $Y=0.725 $X2=0
+ $Y2=0
cc_273 N_A_79_21#_c_142_n N_A_445_47#_c_974_n 0.00579173f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_274 N_A_79_21#_c_130_n N_A_445_47#_c_974_n 0.00208942f $X=4.055 $Y=0.39 $X2=0
+ $Y2=0
cc_275 N_A_79_21#_c_128_n N_A_445_47#_c_975_n 0.00100206f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A_79_21#_c_129_n N_A_445_47#_c_975_n 0.00145773f $X=1.815 $Y=1.18 $X2=0
+ $Y2=0
cc_277 N_A_79_21#_c_142_n N_A_445_47#_c_975_n 0.00475993f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_278 N_A_79_21#_c_128_n N_A_445_47#_c_976_n 0.00132405f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_79_21#_c_129_n N_A_445_47#_c_976_n 0.00899624f $X=1.815 $Y=1.18 $X2=0
+ $Y2=0
cc_280 N_A_79_21#_c_142_n N_A_445_47#_c_976_n 0.00484124f $X=4.405 $Y=1.54 $X2=0
+ $Y2=0
cc_281 N_A_79_21#_M1007_d N_A_445_47#_c_977_n 2.81824e-19 $X=3.175 $Y=0.235
+ $X2=0 $Y2=0
cc_282 N_A_79_21#_c_130_n N_A_445_47#_c_977_n 0.00117584f $X=4.055 $Y=0.39 $X2=0
+ $Y2=0
cc_283 N_A_79_21#_c_131_n N_A_445_47#_c_977_n 8.04547e-19 $X=4.18 $Y=0.725 $X2=0
+ $Y2=0
cc_284 N_A_79_21#_c_134_n N_A_1053_47#_M1010_d 0.00305026f $X=5.82 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_285 N_A_79_21#_M1014_s N_A_1053_47#_c_1044_n 0.0031705f $X=5.685 $Y=0.235
+ $X2=0 $Y2=0
cc_286 N_A_79_21#_c_134_n N_A_1053_47#_c_1044_n 0.0412047f $X=5.82 $Y=0.38 $X2=0
+ $Y2=0
cc_287 N_A_79_21#_c_135_n N_A_1053_47#_c_1044_n 0.00841895f $X=4.98 $Y=0.73
+ $X2=0 $Y2=0
cc_288 N_A2_M1021_g N_A1_M1001_g 0.0445538f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_289 A2 N_A1_c_362_n 7.14059e-19 $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_290 N_A2_c_314_n N_A1_c_362_n 0.0236122f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_291 A2 N_A1_c_363_n 0.0173343f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_292 N_A2_c_314_n N_A1_c_363_n 2.38987e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A2_M1006_g N_VPWR_c_567_n 0.00157837f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A2_M1021_g N_VPWR_c_568_n 0.00157837f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A2_M1006_g N_VPWR_c_574_n 0.00585385f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A2_M1021_g N_VPWR_c_574_n 0.00441875f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A2_M1006_g N_VPWR_c_563_n 0.010464f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A2_M1021_g N_VPWR_c_563_n 0.00588739f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A2_c_311_n N_X_c_685_n 5.22228e-19 $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A2_M1021_g N_A_445_297#_c_744_n 0.0101845f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A2_c_311_n N_VGND_c_848_n 0.00146448f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A2_c_312_n N_VGND_c_849_n 0.00924252f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A2_c_311_n N_VGND_c_856_n 0.00424308f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A2_c_312_n N_VGND_c_856_n 0.00541359f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A2_c_311_n N_VGND_c_863_n 0.00537721f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A2_c_312_n N_VGND_c_863_n 0.00741611f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A2_c_311_n N_A_445_47#_c_979_n 0.0064836f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A2_c_312_n N_A_445_47#_c_979_n 0.00550646f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A2_c_312_n N_A_445_47#_c_972_n 8.90062e-19 $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A2_c_312_n N_A_445_47#_c_974_n 0.00394202f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_311 A2 N_A_445_47#_c_974_n 0.012862f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A2_c_314_n N_A_445_47#_c_974_n 0.00229792f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A2_c_311_n N_A_445_47#_c_975_n 0.00428427f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A2_c_312_n N_A_445_47#_c_975_n 2.36493e-19 $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_c_311_n N_A_445_47#_c_976_n 0.0102373f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A2_c_312_n N_A_445_47#_c_976_n 0.00218533f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_317 A2 N_A_445_47#_c_976_n 0.0168852f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_318 N_A2_c_314_n N_A_445_47#_c_976_n 0.00221535f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A1_c_360_n N_C1_c_418_n 0.0122337f $X=3.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_320 A1 N_C1_c_420_n 0.017972f $X=3.84 $Y=1.105 $X2=0 $Y2=0
cc_321 N_A1_c_362_n N_C1_c_420_n 7.34903e-19 $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_322 A1 N_C1_c_421_n 2.33842e-19 $X=3.84 $Y=1.105 $X2=0 $Y2=0
cc_323 N_A1_c_362_n N_C1_c_421_n 0.0227566f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A1_M1001_g N_VPWR_c_568_n 0.00158508f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A1_M1022_g N_VPWR_c_569_n 0.00338799f $X=3.415 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A1_M1001_g N_VPWR_c_576_n 0.00441875f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A1_M1022_g N_VPWR_c_576_n 0.00441875f $X=3.415 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A1_M1001_g N_VPWR_c_563_n 0.00590064f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A1_M1022_g N_VPWR_c_563_n 0.00719951f $X=3.415 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A1_M1001_g N_A_445_297#_c_744_n 0.0101845f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A1_M1022_g N_A_445_297#_c_740_n 0.0123316f $X=3.415 $Y=1.985 $X2=0
+ $Y2=0
cc_332 N_A1_M1022_g N_A_445_297#_c_756_n 0.00214111f $X=3.415 $Y=1.985 $X2=0
+ $Y2=0
cc_333 N_A1_c_359_n N_VGND_c_849_n 0.00773211f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A1_c_362_n N_VGND_c_849_n 2.20249e-19 $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A1_c_363_n N_VGND_c_849_n 5.53422e-19 $X=3.19 $Y=1.18 $X2=0 $Y2=0
cc_336 N_A1_c_359_n N_VGND_c_858_n 0.00368123f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A1_c_360_n N_VGND_c_858_n 0.00368123f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A1_c_359_n N_VGND_c_863_n 0.00646539f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A1_c_360_n N_VGND_c_863_n 0.00527354f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A1_c_359_n N_A_445_47#_c_972_n 0.0137421f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A1_c_360_n N_A_445_47#_c_972_n 4.69158e-19 $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A1_c_362_n N_A_445_47#_c_972_n 0.00692152f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A1_c_406_p N_A_445_47#_c_972_n 0.0249475f $X=3.71 $Y=1.18 $X2=0 $Y2=0
cc_344 N_A1_c_360_n N_A_445_47#_c_973_n 0.00372211f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_345 A1 N_A_445_47#_c_973_n 0.0130337f $X=3.84 $Y=1.105 $X2=0 $Y2=0
cc_346 N_A1_c_362_n N_A_445_47#_c_973_n 0.00225807f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A1_c_406_p N_A_445_47#_c_973_n 0.0062631f $X=3.71 $Y=1.18 $X2=0 $Y2=0
cc_348 N_A1_c_362_n N_A_445_47#_c_974_n 0.0129453f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A1_c_363_n N_A_445_47#_c_974_n 0.0129381f $X=3.19 $Y=1.18 $X2=0 $Y2=0
cc_350 N_A1_c_406_p N_A_445_47#_c_974_n 0.00326261f $X=3.71 $Y=1.18 $X2=0 $Y2=0
cc_351 N_A1_c_359_n N_A_445_47#_c_977_n 0.00267467f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A1_c_360_n N_A_445_47#_c_977_n 9.56291e-19 $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_353 N_A1_c_362_n N_A_445_47#_c_977_n 0.00305448f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A1_c_406_p N_A_445_47#_c_977_n 0.00753862f $X=3.71 $Y=1.18 $X2=0 $Y2=0
cc_355 N_C1_c_419_n N_B1_c_471_n 0.00912669f $X=4.77 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_356 N_C1_M1008_g N_B1_M1017_g 0.0222405f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_357 N_C1_c_421_n N_B1_c_473_n 0.0362035f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_358 N_C1_M1002_g N_VPWR_c_569_n 0.00214231f $X=4.36 $Y=1.985 $X2=0 $Y2=0
cc_359 N_C1_M1002_g N_VPWR_c_578_n 0.00357877f $X=4.36 $Y=1.985 $X2=0 $Y2=0
cc_360 N_C1_M1008_g N_VPWR_c_578_n 0.00357877f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_361 N_C1_M1002_g N_VPWR_c_563_n 0.00655123f $X=4.36 $Y=1.985 $X2=0 $Y2=0
cc_362 N_C1_M1008_g N_VPWR_c_563_n 0.00525237f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_363 N_C1_M1002_g N_A_445_297#_c_745_n 0.0124134f $X=4.36 $Y=1.985 $X2=0 $Y2=0
cc_364 N_C1_M1008_g N_A_445_297#_c_745_n 0.0106545f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_365 N_C1_M1008_g N_A_445_297#_c_749_n 0.00107149f $X=4.78 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_C1_M1002_g N_A_804_297#_c_811_n 0.00970685f $X=4.36 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_C1_M1008_g N_A_804_297#_c_811_n 0.00970685f $X=4.78 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_C1_c_418_n N_VGND_c_850_n 0.00268723f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_369 N_C1_c_419_n N_VGND_c_850_n 0.00268723f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_370 N_C1_c_418_n N_VGND_c_858_n 0.00423866f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_371 N_C1_c_419_n N_VGND_c_860_n 0.00421816f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_372 N_C1_c_418_n N_VGND_c_863_n 0.0057566f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_373 N_C1_c_419_n N_VGND_c_863_n 0.00575258f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_374 N_B1_M1023_g N_B2_M1018_g 0.0096257f $X=5.62 $Y=1.985 $X2=0 $Y2=0
cc_375 N_B1_c_474_n N_B2_c_522_n 9.15201e-19 $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_376 N_B1_c_475_n N_B2_c_522_n 0.0144818f $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_377 N_B1_c_474_n N_B2_c_523_n 0.0157691f $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_378 N_B1_c_475_n N_B2_c_523_n 2.34902e-19 $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_379 N_B1_M1017_g N_VPWR_c_578_n 0.00357877f $X=5.2 $Y=1.985 $X2=0 $Y2=0
cc_380 N_B1_M1023_g N_VPWR_c_578_n 0.00357877f $X=5.62 $Y=1.985 $X2=0 $Y2=0
cc_381 N_B1_M1017_g N_VPWR_c_563_n 0.00525237f $X=5.2 $Y=1.985 $X2=0 $Y2=0
cc_382 N_B1_M1023_g N_VPWR_c_563_n 0.00597864f $X=5.62 $Y=1.985 $X2=0 $Y2=0
cc_383 N_B1_M1017_g N_A_445_297#_c_745_n 0.0113842f $X=5.2 $Y=1.985 $X2=0 $Y2=0
cc_384 N_B1_M1023_g N_A_445_297#_c_745_n 0.00228614f $X=5.62 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_B1_c_475_n N_A_445_297#_c_745_n 2.34443e-19 $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_386 N_B1_M1017_g N_A_445_297#_c_738_n 0.00258632f $X=5.2 $Y=1.985 $X2=0 $Y2=0
cc_387 N_B1_M1023_g N_A_445_297#_c_738_n 0.00123487f $X=5.62 $Y=1.985 $X2=0
+ $Y2=0
cc_388 N_B1_c_473_n N_A_445_297#_c_738_n 0.0022284f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_389 N_B1_c_475_n N_A_445_297#_c_738_n 0.0264095f $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_390 N_B1_M1017_g N_A_445_297#_c_749_n 0.0044999f $X=5.2 $Y=1.985 $X2=0 $Y2=0
cc_391 N_B1_M1023_g N_A_445_297#_c_749_n 0.0082924f $X=5.62 $Y=1.985 $X2=0 $Y2=0
cc_392 N_B1_M1023_g N_A_445_297#_c_739_n 0.0101816f $X=5.62 $Y=1.985 $X2=0 $Y2=0
cc_393 N_B1_c_474_n N_A_445_297#_c_739_n 0.00796921f $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_394 N_B1_c_475_n N_A_445_297#_c_739_n 0.0328967f $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_395 N_B1_M1017_g N_A_804_297#_c_811_n 0.00970559f $X=5.2 $Y=1.985 $X2=0 $Y2=0
cc_396 N_B1_M1023_g N_A_804_297#_c_811_n 0.0113267f $X=5.62 $Y=1.985 $X2=0 $Y2=0
cc_397 N_B1_c_471_n N_VGND_c_860_n 0.00357877f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_398 N_B1_c_472_n N_VGND_c_860_n 0.00357877f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_399 N_B1_c_471_n N_VGND_c_863_n 0.00525237f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_400 N_B1_c_472_n N_VGND_c_863_n 0.00655123f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_401 N_B1_c_471_n N_A_1053_47#_c_1044_n 0.00372684f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_402 N_B1_c_472_n N_A_1053_47#_c_1044_n 0.0141922f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_403 N_B1_c_473_n N_A_1053_47#_c_1044_n 0.0110255f $X=5.695 $Y=1.16 $X2=0
+ $Y2=0
cc_404 N_B1_c_475_n N_A_1053_47#_c_1044_n 0.0593719f $X=5.87 $Y=1.16 $X2=0 $Y2=0
cc_405 N_B2_M1018_g N_VPWR_c_578_n 0.00357877f $X=6.46 $Y=1.985 $X2=0 $Y2=0
cc_406 N_B2_M1027_g N_VPWR_c_578_n 0.00357877f $X=6.88 $Y=1.985 $X2=0 $Y2=0
cc_407 N_B2_M1018_g N_VPWR_c_563_n 0.00597864f $X=6.46 $Y=1.985 $X2=0 $Y2=0
cc_408 N_B2_M1027_g N_VPWR_c_563_n 0.00655123f $X=6.88 $Y=1.985 $X2=0 $Y2=0
cc_409 N_B2_M1018_g N_A_445_297#_c_739_n 0.0124772f $X=6.46 $Y=1.985 $X2=0 $Y2=0
cc_410 N_B2_c_522_n N_A_445_297#_c_739_n 0.0204068f $X=6.845 $Y=1.16 $X2=0 $Y2=0
cc_411 N_B2_c_523_n N_A_445_297#_c_739_n 0.00105696f $X=6.97 $Y=1.16 $X2=0 $Y2=0
cc_412 N_B2_M1027_g N_A_445_297#_c_741_n 0.00101193f $X=6.88 $Y=1.985 $X2=0
+ $Y2=0
cc_413 N_B2_c_522_n N_A_445_297#_c_741_n 0.020533f $X=6.845 $Y=1.16 $X2=0 $Y2=0
cc_414 N_B2_c_523_n N_A_445_297#_c_741_n 0.00256468f $X=6.97 $Y=1.16 $X2=0 $Y2=0
cc_415 N_B2_M1018_g N_A_804_297#_c_810_n 0.00984328f $X=6.46 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_B2_M1027_g N_A_804_297#_c_810_n 0.0121747f $X=6.88 $Y=1.985 $X2=0 $Y2=0
cc_417 N_B2_c_522_n N_A_804_297#_c_821_n 0.00859468f $X=6.845 $Y=1.16 $X2=0
+ $Y2=0
cc_418 N_B2_c_523_n N_A_804_297#_c_821_n 0.00138343f $X=6.97 $Y=1.16 $X2=0 $Y2=0
cc_419 N_B2_c_520_n N_VGND_c_851_n 0.00268723f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_420 N_B2_c_521_n N_VGND_c_851_n 0.00268723f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_421 N_B2_c_520_n N_VGND_c_860_n 0.00435595f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_422 N_B2_c_521_n N_VGND_c_862_n 0.00423334f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_423 N_B2_c_520_n N_VGND_c_863_n 0.00726879f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_424 N_B2_c_521_n N_VGND_c_863_n 0.00704237f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_425 N_B2_c_522_n N_A_1053_47#_c_1044_n 0.0542204f $X=6.845 $Y=1.16 $X2=0
+ $Y2=0
cc_426 N_B2_c_523_n N_A_1053_47#_c_1044_n 0.00374513f $X=6.97 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_B2_c_520_n N_A_1053_47#_c_1045_n 0.00869873f $X=6.55 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_B2_c_521_n N_A_1053_47#_c_1045_n 0.00999285f $X=6.97 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_B2_c_522_n N_A_1053_47#_c_1045_n 0.0223991f $X=6.845 $Y=1.16 $X2=0
+ $Y2=0
cc_430 N_B2_c_523_n N_A_1053_47#_c_1045_n 0.00260689f $X=6.97 $Y=1.16 $X2=0
+ $Y2=0
cc_431 N_B2_c_520_n N_A_1053_47#_c_1046_n 7.04871e-19 $X=6.55 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_B2_c_521_n N_A_1053_47#_c_1046_n 0.00640821f $X=6.97 $Y=0.995 $X2=0
+ $Y2=0
cc_433 N_B2_c_520_n N_A_1053_47#_c_1047_n 0.00339214f $X=6.55 $Y=0.995 $X2=0
+ $Y2=0
cc_434 N_B2_c_521_n N_A_1053_47#_c_1047_n 2.31028e-19 $X=6.97 $Y=0.995 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_563_n N_X_M1003_d 0.00284632f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_436 N_VPWR_c_563_n N_X_M1016_d 0.00284632f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_437 N_VPWR_c_570_n N_X_c_707_n 0.0142343f $X=0.975 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_c_563_n N_X_c_707_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_439 N_VPWR_M1005_s N_X_c_667_n 0.00165831f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_440 N_VPWR_c_566_n N_X_c_667_n 0.0126919f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_441 N_VPWR_c_572_n N_X_c_711_n 0.0142343f $X=1.815 $Y=2.72 $X2=0 $Y2=0
cc_442 N_VPWR_c_563_n N_X_c_711_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_443 N_VPWR_c_565_n N_X_c_669_n 0.00102118f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_444 N_VPWR_M1003_s N_X_c_672_n 0.00343744f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_445 N_VPWR_c_565_n N_X_c_672_n 0.0152373f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_446 N_VPWR_c_563_n N_A_445_297#_M1006_s 0.00253991f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_447 N_VPWR_c_563_n N_A_445_297#_M1001_d 0.00227365f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_563_n N_A_445_297#_M1017_s 0.00216833f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_563_n N_A_445_297#_M1018_s 0.0021603f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_450 N_VPWR_M1021_d N_A_445_297#_c_744_n 0.00325422f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_568_n N_A_445_297#_c_744_n 0.0123012f $X=2.78 $Y=2.3 $X2=0 $Y2=0
cc_452 N_VPWR_c_574_n N_A_445_297#_c_744_n 0.00201582f $X=2.655 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_576_n N_A_445_297#_c_744_n 0.00201582f $X=3.5 $Y=2.72 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_563_n N_A_445_297#_c_744_n 0.00800071f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_574_n N_A_445_297#_c_750_n 0.0142224f $X=2.655 $Y=2.72 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_563_n N_A_445_297#_c_750_n 0.00954719f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_576_n N_A_445_297#_c_751_n 0.0145736f $X=3.5 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_563_n N_A_445_297#_c_751_n 0.00973967f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_459 N_VPWR_M1022_s N_A_445_297#_c_740_n 0.0047504f $X=3.49 $Y=1.485 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_569_n N_A_445_297#_c_740_n 0.0159284f $X=3.625 $Y=2.3 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_576_n N_A_445_297#_c_740_n 0.00201582f $X=3.5 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_578_n N_A_445_297#_c_740_n 0.00272871f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_563_n N_A_445_297#_c_740_n 0.0096447f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_563_n N_A_804_297#_M1002_d 0.00213443f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_465 N_VPWR_c_563_n N_A_804_297#_M1008_d 0.00215227f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_563_n N_A_804_297#_M1023_d 0.0055807f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_563_n N_A_804_297#_M1027_d 0.00217519f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_578_n N_A_804_297#_c_810_n 0.0162911f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_563_n N_A_804_297#_c_810_n 0.00962794f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_569_n N_A_804_297#_c_811_n 0.0195142f $X=3.625 $Y=2.3 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_578_n N_A_804_297#_c_811_n 0.178343f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_472 N_VPWR_c_563_n N_A_804_297#_c_811_n 0.109864f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_473 N_X_c_666_n N_VGND_M1011_d 0.0031268f $X=0.21 $Y=0.905 $X2=-0.19
+ $Y2=-0.24
cc_474 N_X_c_662_n N_VGND_M1013_d 0.00162089f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_475 N_X_c_666_n N_VGND_c_845_n 0.00130186f $X=0.21 $Y=0.905 $X2=0 $Y2=0
cc_476 N_X_c_663_n N_VGND_c_846_n 9.38992e-19 $X=0.515 $Y=0.82 $X2=0 $Y2=0
cc_477 N_X_c_666_n N_VGND_c_846_n 0.0122878f $X=0.21 $Y=0.905 $X2=0 $Y2=0
cc_478 N_X_c_662_n N_VGND_c_847_n 0.0122559f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_479 N_X_c_673_n N_VGND_c_852_n 0.0188551f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_480 N_X_c_662_n N_VGND_c_852_n 0.00198695f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_481 N_X_c_663_n N_VGND_c_852_n 0.00193763f $X=0.515 $Y=0.82 $X2=0 $Y2=0
cc_482 N_X_c_662_n N_VGND_c_854_n 0.00198695f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_483 N_X_c_685_n N_VGND_c_854_n 0.0188551f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_484 N_X_M1011_s N_VGND_c_863_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_485 N_X_M1015_s N_VGND_c_863_n 0.00215201f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_486 N_X_c_673_n N_VGND_c_863_n 0.0122069f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_487 N_X_c_662_n N_VGND_c_863_n 0.00835832f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_488 N_X_c_685_n N_VGND_c_863_n 0.0122069f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_489 N_X_c_663_n N_VGND_c_863_n 0.00388553f $X=0.515 $Y=0.82 $X2=0 $Y2=0
cc_490 N_X_c_666_n N_VGND_c_863_n 0.00292923f $X=0.21 $Y=0.905 $X2=0 $Y2=0
cc_491 N_X_c_662_n N_A_445_47#_c_979_n 3.09105e-19 $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_492 N_X_c_685_n N_A_445_47#_c_979_n 0.00518536f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_493 N_X_c_662_n N_A_445_47#_c_975_n 0.00106395f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_494 N_X_c_662_n N_A_445_47#_c_976_n 0.00697112f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_495 N_A_445_297#_c_740_n N_A_804_297#_M1002_d 0.00120897f $X=4.06 $Y=1.92
+ $X2=-0.19 $Y2=1.305
cc_496 N_A_445_297#_c_756_n N_A_804_297#_M1002_d 0.00571063f $X=4.23 $Y=1.92
+ $X2=-0.19 $Y2=1.305
cc_497 N_A_445_297#_c_745_n N_A_804_297#_M1008_d 0.00351203f $X=5.245 $Y=1.96
+ $X2=0 $Y2=0
cc_498 N_A_445_297#_c_739_n N_A_804_297#_M1023_d 0.00867684f $X=6.555 $Y=1.54
+ $X2=0 $Y2=0
cc_499 N_A_445_297#_M1018_s N_A_804_297#_c_810_n 0.00312348f $X=6.535 $Y=1.485
+ $X2=0 $Y2=0
cc_500 N_A_445_297#_c_739_n N_A_804_297#_c_810_n 0.00320918f $X=6.555 $Y=1.54
+ $X2=0 $Y2=0
cc_501 N_A_445_297#_c_741_n N_A_804_297#_c_810_n 0.0118729f $X=6.67 $Y=1.62
+ $X2=0 $Y2=0
cc_502 N_A_445_297#_M1017_s N_A_804_297#_c_811_n 0.00316082f $X=5.275 $Y=1.485
+ $X2=0 $Y2=0
cc_503 N_A_445_297#_c_745_n N_A_804_297#_c_811_n 0.0166283f $X=5.245 $Y=1.96
+ $X2=0 $Y2=0
cc_504 N_A_445_297#_c_739_n N_A_804_297#_c_811_n 0.00297464f $X=6.555 $Y=1.54
+ $X2=0 $Y2=0
cc_505 N_A_445_297#_c_740_n N_A_804_297#_c_811_n 0.0064354f $X=4.06 $Y=1.92
+ $X2=0 $Y2=0
cc_506 N_A_445_297#_c_756_n N_A_804_297#_c_811_n 0.0626083f $X=4.23 $Y=1.92
+ $X2=0 $Y2=0
cc_507 N_A_445_297#_c_739_n N_A_804_297#_c_844_n 0.0465891f $X=6.555 $Y=1.54
+ $X2=0 $Y2=0
cc_508 N_A_445_297#_c_739_n N_A_1053_47#_c_1044_n 0.00813617f $X=6.555 $Y=1.54
+ $X2=0 $Y2=0
cc_509 N_VGND_c_863_n N_A_445_47#_M1019_s 0.00177024f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_510 N_VGND_c_863_n N_A_445_47#_M1007_s 0.00212583f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_856_n N_A_445_47#_c_979_n 0.0188551f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_863_n N_A_445_47#_c_979_n 0.00578691f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_849_n N_A_445_47#_c_972_n 0.0060966f $X=2.78 $Y=0.73 $X2=0 $Y2=0
cc_514 N_VGND_M1024_d N_A_445_47#_c_974_n 0.00126326f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_515 N_VGND_c_849_n N_A_445_47#_c_974_n 0.0116865f $X=2.78 $Y=0.73 $X2=0 $Y2=0
cc_516 N_VGND_c_863_n N_A_445_47#_c_974_n 0.0528913f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_M1026_d N_A_445_47#_c_975_n 5.72321e-19 $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_518 N_VGND_c_848_n N_A_445_47#_c_975_n 4.77004e-19 $X=1.94 $Y=0.39 $X2=0
+ $Y2=0
cc_519 N_VGND_c_863_n N_A_445_47#_c_975_n 0.0139713f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_M1026_d N_A_445_47#_c_976_n 0.00143564f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_521 N_VGND_c_848_n N_A_445_47#_c_976_n 0.0111567f $X=1.94 $Y=0.39 $X2=0 $Y2=0
cc_522 N_VGND_c_849_n N_A_445_47#_c_976_n 0.00789021f $X=2.78 $Y=0.73 $X2=0
+ $Y2=0
cc_523 N_VGND_c_856_n N_A_445_47#_c_976_n 0.00200982f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_863_n N_A_445_47#_c_976_n 0.00149178f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_849_n N_A_445_47#_c_977_n 2.40232e-19 $X=2.78 $Y=0.73 $X2=0
+ $Y2=0
cc_526 N_VGND_c_863_n N_A_445_47#_c_977_n 0.0143563f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_863_n N_A_1053_47#_M1010_d 0.00216833f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_528 N_VGND_c_863_n N_A_1053_47#_M1000_s 0.00308734f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_863_n N_A_1053_47#_M1004_s 0.00209319f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_860_n N_A_1053_47#_c_1044_n 0.00884209f $X=6.675 $Y=0 $X2=0
+ $Y2=0
cc_531 N_VGND_c_863_n N_A_1053_47#_c_1044_n 0.0161857f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_M1000_d N_A_1053_47#_c_1045_n 0.00162089f $X=6.625 $Y=0.235 $X2=0
+ $Y2=0
cc_533 N_VGND_c_851_n N_A_1053_47#_c_1045_n 0.0122559f $X=6.76 $Y=0.39 $X2=0
+ $Y2=0
cc_534 N_VGND_c_860_n N_A_1053_47#_c_1045_n 0.00198695f $X=6.675 $Y=0 $X2=0
+ $Y2=0
cc_535 N_VGND_c_862_n N_A_1053_47#_c_1045_n 0.00198695f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_863_n N_A_1053_47#_c_1045_n 0.00835832f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_862_n N_A_1053_47#_c_1046_n 0.0209752f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_863_n N_A_1053_47#_c_1046_n 0.0124119f $X=7.59 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkdlybuf4s50_2.spice
* Created: Thu Aug 27 14:12:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s50_2.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s50_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819196 AS=0.1134 PD=0.792897 PS=1.38 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_283_47#_M1002_d N_A_27_47#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.5
+ W=0.65 AD=0.17225 AS=0.12678 PD=1.83 PS=1.2271 NRD=0 NRS=4.608 M=1 R=1.3
+ SA=250000 SB=250000 A=0.325 P=2.3 MULT=1
MM1000 N_VGND_M1000_d N_A_283_47#_M1000_g N_A_390_47#_M1000_s VNB NSHORT L=0.5
+ W=0.65 AD=0.119126 AS=0.169 PD=1.19065 PS=1.82 NRD=0 NRS=0 M=1 R=1.3 SA=250000
+ SB=250001 A=0.325 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_390_47#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.0769738 PD=0.695 PS=0.769346 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1001_d N_A_390_47#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.1638 PD=0.695 PS=1.62 NRD=0 NRS=35.712 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.186923 AS=0.27 PD=1.49451 PS=2.54 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1008 N_A_283_47#_M1008_d N_A_27_47#_M1008_g N_VPWR_M1006_d VPB PHIGHVT L=0.5
+ W=0.82 AD=0.2173 AS=0.153277 PD=2.17 PS=1.22549 NRD=0 NRS=2.3837 M=1 R=1.64
+ SA=250001 SB=250000 A=0.41 P=2.64 MULT=1
MM1007 N_VPWR_M1007_d N_A_283_47#_M1007_g N_A_390_47#_M1007_s VPB PHIGHVT L=0.5
+ W=0.82 AD=0.142193 AS=0.2132 PD=1.19846 PS=2.16 NRD=0 NRS=0 M=1 R=1.64
+ SA=250000 SB=250001 A=0.41 P=2.64 MULT=1
MM1004 N_VPWR_M1007_d N_A_390_47#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.173407 AS=0.1375 PD=1.46154 PS=1.275 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.9 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_390_47#_M1009_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.39 AS=0.1375 PD=2.78 PS=1.275 NRD=24.6053 NRS=0 M=1 R=6.66667 SA=75001.3
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__clkdlybuf4s50_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__dfsbp_1.pxi.spice
* Created: Thu Aug 27 14:15:01 2020
* 
x_PM_SKY130_FD_SC_HD__DFSBP_1%CLK N_CLK_c_235_n N_CLK_c_230_n N_CLK_M1032_g
+ N_CLK_c_236_n N_CLK_M1018_g N_CLK_c_231_n N_CLK_c_237_n CLK CLK N_CLK_c_233_n
+ N_CLK_c_234_n PM_SKY130_FD_SC_HD__DFSBP_1%CLK
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_27_47# N_A_27_47#_M1032_s N_A_27_47#_M1018_s
+ N_A_27_47#_M1022_g N_A_27_47#_M1000_g N_A_27_47#_c_275_n N_A_27_47#_M1030_g
+ N_A_27_47#_M1033_g N_A_27_47#_M1005_g N_A_27_47#_M1012_g N_A_27_47#_c_530_p
+ N_A_27_47#_c_276_n N_A_27_47#_c_277_n N_A_27_47#_c_291_n N_A_27_47#_c_403_p
+ N_A_27_47#_c_278_n N_A_27_47#_c_279_n N_A_27_47#_c_280_n N_A_27_47#_c_281_n
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_c_295_n N_A_27_47#_c_284_n
+ N_A_27_47#_c_285_n N_A_27_47#_c_296_n N_A_27_47#_c_297_n N_A_27_47#_c_298_n
+ N_A_27_47#_c_299_n N_A_27_47#_c_300_n N_A_27_47#_c_286_n N_A_27_47#_c_302_n
+ N_A_27_47#_c_303_n N_A_27_47#_c_304_n N_A_27_47#_c_305_n N_A_27_47#_c_287_n
+ PM_SKY130_FD_SC_HD__DFSBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DFSBP_1%D N_D_M1009_g N_D_M1027_g D D N_D_c_548_n
+ N_D_c_549_n PM_SKY130_FD_SC_HD__DFSBP_1%D
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_193_47# N_A_193_47#_M1022_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1010_g N_A_193_47#_c_586_n N_A_193_47#_c_587_n
+ N_A_193_47#_M1020_g N_A_193_47#_c_589_n N_A_193_47#_M1011_g
+ N_A_193_47#_c_591_n N_A_193_47#_M1028_g N_A_193_47#_c_592_n
+ N_A_193_47#_c_593_n N_A_193_47#_c_594_n N_A_193_47#_c_595_n
+ N_A_193_47#_c_596_n N_A_193_47#_c_597_n N_A_193_47#_c_598_n
+ N_A_193_47#_c_599_n N_A_193_47#_c_600_n N_A_193_47#_c_601_n
+ N_A_193_47#_c_602_n N_A_193_47#_c_603_n PM_SKY130_FD_SC_HD__DFSBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_652_21# N_A_652_21#_M1006_d N_A_652_21#_M1029_d
+ N_A_652_21#_M1025_g N_A_652_21#_M1008_g N_A_652_21#_c_788_n
+ N_A_652_21#_c_872_p N_A_652_21#_c_789_n N_A_652_21#_c_783_n
+ N_A_652_21#_c_784_n N_A_652_21#_c_791_n N_A_652_21#_c_792_n
+ N_A_652_21#_c_793_n N_A_652_21#_c_785_n PM_SKY130_FD_SC_HD__DFSBP_1%A_652_21#
x_PM_SKY130_FD_SC_HD__DFSBP_1%SET_B N_SET_B_c_897_n N_SET_B_M1029_g
+ N_SET_B_M1004_g N_SET_B_M1021_g N_SET_B_M1001_g N_SET_B_c_901_n
+ N_SET_B_c_912_n N_SET_B_c_902_n N_SET_B_c_903_n SET_B N_SET_B_c_905_n
+ N_SET_B_c_906_n N_SET_B_c_907_n N_SET_B_c_908_n
+ PM_SKY130_FD_SC_HD__DFSBP_1%SET_B
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_476_47# N_A_476_47#_M1030_d N_A_476_47#_M1010_d
+ N_A_476_47#_c_1032_n N_A_476_47#_M1006_g N_A_476_47#_c_1033_n
+ N_A_476_47#_M1023_g N_A_476_47#_c_1034_n N_A_476_47#_M1016_g
+ N_A_476_47#_c_1035_n N_A_476_47#_M1024_g N_A_476_47#_c_1036_n
+ N_A_476_47#_c_1059_n N_A_476_47#_c_1064_n N_A_476_47#_c_1044_n
+ N_A_476_47#_c_1037_n N_A_476_47#_c_1038_n N_A_476_47#_c_1039_n
+ N_A_476_47#_c_1040_n N_A_476_47#_c_1041_n
+ PM_SKY130_FD_SC_HD__DFSBP_1%A_476_47#
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_1178_261# N_A_1178_261#_M1017_d
+ N_A_1178_261#_M1026_d N_A_1178_261#_c_1193_n N_A_1178_261#_M1013_g
+ N_A_1178_261#_M1014_g N_A_1178_261#_c_1190_n N_A_1178_261#_c_1196_n
+ N_A_1178_261#_c_1247_p N_A_1178_261#_c_1191_n N_A_1178_261#_c_1192_n
+ N_A_1178_261#_c_1198_n N_A_1178_261#_c_1199_n
+ PM_SKY130_FD_SC_HD__DFSBP_1%A_1178_261#
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_1028_413# N_A_1028_413#_M1011_d
+ N_A_1028_413#_M1005_d N_A_1028_413#_M1001_s N_A_1028_413#_M1017_g
+ N_A_1028_413#_M1026_g N_A_1028_413#_c_1266_n N_A_1028_413#_c_1267_n
+ N_A_1028_413#_M1007_g N_A_1028_413#_M1019_g N_A_1028_413#_c_1270_n
+ N_A_1028_413#_c_1271_n N_A_1028_413#_c_1272_n N_A_1028_413#_c_1273_n
+ N_A_1028_413#_M1003_g N_A_1028_413#_c_1286_n N_A_1028_413#_M1002_g
+ N_A_1028_413#_c_1274_n N_A_1028_413#_c_1275_n N_A_1028_413#_c_1276_n
+ N_A_1028_413#_c_1287_n N_A_1028_413#_c_1295_n N_A_1028_413#_c_1288_n
+ N_A_1028_413#_c_1303_n N_A_1028_413#_c_1277_n N_A_1028_413#_c_1278_n
+ N_A_1028_413#_c_1290_n N_A_1028_413#_c_1279_n N_A_1028_413#_c_1291_n
+ N_A_1028_413#_c_1292_n N_A_1028_413#_c_1375_n N_A_1028_413#_c_1280_n
+ N_A_1028_413#_c_1281_n PM_SKY130_FD_SC_HD__DFSBP_1%A_1028_413#
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_1786_47# N_A_1786_47#_M1003_s
+ N_A_1786_47#_M1002_s N_A_1786_47#_M1015_g N_A_1786_47#_M1031_g
+ N_A_1786_47#_c_1454_n N_A_1786_47#_c_1460_n N_A_1786_47#_c_1455_n
+ N_A_1786_47#_c_1456_n N_A_1786_47#_c_1457_n N_A_1786_47#_c_1458_n
+ PM_SKY130_FD_SC_HD__DFSBP_1%A_1786_47#
x_PM_SKY130_FD_SC_HD__DFSBP_1%VPWR N_VPWR_M1018_d N_VPWR_M1027_s N_VPWR_M1008_d
+ N_VPWR_M1023_d N_VPWR_M1013_d N_VPWR_M1001_d N_VPWR_M1019_s N_VPWR_M1002_d
+ N_VPWR_c_1508_n N_VPWR_c_1509_n N_VPWR_c_1510_n N_VPWR_c_1511_n
+ N_VPWR_c_1512_n N_VPWR_c_1513_n N_VPWR_c_1514_n N_VPWR_c_1515_n
+ N_VPWR_c_1516_n N_VPWR_c_1517_n VPWR VPWR N_VPWR_c_1518_n N_VPWR_c_1519_n
+ N_VPWR_c_1520_n N_VPWR_c_1521_n N_VPWR_c_1522_n N_VPWR_c_1523_n
+ N_VPWR_c_1507_n N_VPWR_c_1525_n N_VPWR_c_1526_n N_VPWR_c_1527_n
+ N_VPWR_c_1528_n N_VPWR_c_1529_n N_VPWR_c_1530_n N_VPWR_c_1531_n
+ PM_SKY130_FD_SC_HD__DFSBP_1%VPWR
x_PM_SKY130_FD_SC_HD__DFSBP_1%A_381_47# N_A_381_47#_M1009_d N_A_381_47#_M1027_d
+ N_A_381_47#_c_1687_n N_A_381_47#_c_1692_n N_A_381_47#_c_1688_n
+ N_A_381_47#_c_1694_n N_A_381_47#_c_1690_n N_A_381_47#_c_1696_n
+ N_A_381_47#_c_1697_n PM_SKY130_FD_SC_HD__DFSBP_1%A_381_47#
x_PM_SKY130_FD_SC_HD__DFSBP_1%Q_N N_Q_N_M1007_d N_Q_N_M1019_d Q_N Q_N Q_N Q_N
+ Q_N Q_N N_Q_N_c_1753_n PM_SKY130_FD_SC_HD__DFSBP_1%Q_N
x_PM_SKY130_FD_SC_HD__DFSBP_1%Q N_Q_M1015_d N_Q_M1031_d N_Q_c_1775_n
+ N_Q_c_1778_n N_Q_c_1776_n Q Q Q PM_SKY130_FD_SC_HD__DFSBP_1%Q
x_PM_SKY130_FD_SC_HD__DFSBP_1%VGND N_VGND_M1032_d N_VGND_M1009_s N_VGND_M1025_d
+ N_VGND_M1024_s N_VGND_M1021_d N_VGND_M1007_s N_VGND_M1003_d N_VGND_c_1791_n
+ N_VGND_c_1792_n N_VGND_c_1793_n N_VGND_c_1794_n N_VGND_c_1795_n
+ N_VGND_c_1796_n N_VGND_c_1797_n N_VGND_c_1798_n N_VGND_c_1799_n VGND VGND
+ N_VGND_c_1800_n N_VGND_c_1801_n N_VGND_c_1802_n N_VGND_c_1803_n
+ N_VGND_c_1804_n N_VGND_c_1805_n N_VGND_c_1806_n N_VGND_c_1807_n
+ N_VGND_c_1808_n N_VGND_c_1809_n N_VGND_c_1810_n N_VGND_c_1811_n
+ N_VGND_c_1812_n PM_SKY130_FD_SC_HD__DFSBP_1%VGND
cc_1 VNB N_CLK_c_230_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_231_n 0.0229857f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK 0.0187424f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_c_233_n 0.01953f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_CLK_c_234_n 0.0141141f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1022_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_275_n 0.0180457f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_8 VNB N_A_27_47#_c_276_n 0.00174761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_277_n 0.00643757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_278_n 0.00246672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_279_n 0.00445416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_280_n 0.0327378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_281_n 0.0065365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_282_n 0.00811013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_283_n 0.00157243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_284_n 0.00506957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_285_n 0.0254426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_286_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_287_n 0.0159476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_M1009_g 0.0205663f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_21 VNB N_D_c_548_n 0.0258802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_D_c_549_n 0.00442451f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_23 VNB N_A_193_47#_c_586_n 0.0132632f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_24 VNB N_A_193_47#_c_587_n 0.00435992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_M1020_g 0.0199482f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_26 VNB N_A_193_47#_c_589_n 0.00803437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_M1011_g 0.0339128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_591_n 0.0101365f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_29 VNB N_A_193_47#_c_592_n 0.0177609f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_30 VNB N_A_193_47#_c_593_n 0.0194566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_594_n 0.00568843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_595_n 0.00105673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_596_n 0.0167211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_597_n 0.00113053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_598_n 0.00189817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_599_n 0.00500582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_600_n 0.00145876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_601_n 0.00222242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_602_n 0.0246637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_603_n 0.0161628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_652_21#_M1025_g 0.0422386f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_42 VNB N_A_652_21#_c_783_n 0.00136482f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_652_21#_c_784_n 0.00320601f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_44 VNB N_A_652_21#_c_785_n 0.00519354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_SET_B_c_897_n 0.0308821f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_46 VNB N_SET_B_M1029_g 0.00706345f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_47 VNB N_SET_B_M1004_g 0.0179723f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_48 VNB N_SET_B_M1021_g 0.0183761f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_49 VNB N_SET_B_c_901_n 0.0075909f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_50 VNB N_SET_B_c_902_n 0.0252701f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_51 VNB N_SET_B_c_903_n 0.00436858f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_52 VNB SET_B 0.00646661f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_53 VNB N_SET_B_c_905_n 0.0135879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_906_n 0.00185354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_907_n 3.85333e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_SET_B_c_908_n 0.00287603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_476_47#_c_1032_n 0.017726f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_58 VNB N_A_476_47#_c_1033_n 0.0138425f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_59 VNB N_A_476_47#_c_1034_n 0.0551178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_476_47#_c_1035_n 0.0177765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_476_47#_c_1036_n 0.00507008f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_62 VNB N_A_476_47#_c_1037_n 0.00430167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_476_47#_c_1038_n 0.00446117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_476_47#_c_1039_n 0.00393532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_476_47#_c_1040_n 0.00107462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_476_47#_c_1041_n 0.0145904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1178_261#_M1014_g 0.0370862f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_68 VNB N_A_1178_261#_c_1190_n 0.00831243f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_69 VNB N_A_1178_261#_c_1191_n 0.00592339f $X=-0.19 $Y=-0.24 $X2=0.265
+ $Y2=1.53
cc_70 VNB N_A_1178_261#_c_1192_n 0.0048553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1028_413#_M1017_g 0.0277072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1028_413#_c_1266_n 0.063811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1028_413#_c_1267_n 0.0154019f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_74 VNB N_A_1028_413#_M1007_g 0.0249669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1028_413#_M1019_g 5.92051e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_76 VNB N_A_1028_413#_c_1270_n 0.054487f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_77 VNB N_A_1028_413#_c_1271_n 0.0081567f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_78 VNB N_A_1028_413#_c_1272_n 4.83176e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1028_413#_c_1273_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1028_413#_c_1274_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1028_413#_c_1275_n 0.0181388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1028_413#_c_1276_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1028_413#_c_1277_n 0.00479234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1028_413#_c_1278_n 0.00125329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1028_413#_c_1279_n 0.00897687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1028_413#_c_1280_n 8.45714e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1028_413#_c_1281_n 0.00455313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1786_47#_c_1454_n 0.00773792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1786_47#_c_1455_n 0.00613607f $X=-0.19 $Y=-0.24 $X2=0.245
+ $Y2=1.235
cc_90 VNB N_A_1786_47#_c_1456_n 0.0266366f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_91 VNB N_A_1786_47#_c_1457_n 3.01905e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_92 VNB N_A_1786_47#_c_1458_n 0.0203853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VPWR_c_1507_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_381_47#_c_1687_n 0.00882912f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_95 VNB N_A_381_47#_c_1688_n 0.00229945f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_96 VNB N_Q_N_c_1753_n 0.00680658f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_97 VNB N_Q_c_1775_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_98 VNB N_Q_c_1776_n 0.0230748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB Q 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_100 VNB N_VGND_c_1791_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_101 VNB N_VGND_c_1792_n 0.00492922f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_102 VNB N_VGND_c_1793_n 0.00404464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1794_n 0.0101869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1795_n 0.0183409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1796_n 0.00706267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1797_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1798_n 0.033128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1799_n 0.00324376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1800_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1801_n 0.0164349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1802_n 0.0451324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1803_n 0.0192996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1804_n 0.0304243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1805_n 0.522696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1806_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1807_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1808_n 0.0056662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1809_n 0.00651127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1810_n 0.0402451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1811_n 0.0122102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1812_n 0.00345893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VPB N_CLK_c_235_n 0.0118724f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_123 VPB N_CLK_c_236_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_124 VPB N_CLK_c_237_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_125 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_126 VPB N_CLK_c_233_n 0.0100888f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_127 VPB N_A_27_47#_M1000_g 0.0364742f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_128 VPB N_A_27_47#_M1033_g 0.021588f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_129 VPB N_A_27_47#_M1005_g 0.0202815f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_130 VPB N_A_27_47#_c_291_n 0.00196457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_278_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_279_n 0.00245013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_281_n 0.00551288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_295_n 0.00355155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_296_n 0.0141666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_297_n 0.00111704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_298_n 0.0113093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_299_n 0.0015212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_300_n 0.0036941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_286_n 0.0115872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_302_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_303_n 0.00564526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_304_n 0.0280489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_305_n 0.00604462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_D_M1027_g 0.0293669f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_146 VPB N_D_c_548_n 0.00538482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_D_c_549_n 0.00459652f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_148 VPB N_A_193_47#_M1010_g 0.0465266f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_149 VPB N_A_193_47#_c_586_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_150 VPB N_A_193_47#_c_587_n 0.00328709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_193_47#_c_591_n 0.0110014f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_152 VPB N_A_193_47#_M1028_g 0.0394336f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_153 VPB N_A_193_47#_c_592_n 0.0120454f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_154 VPB N_A_193_47#_c_601_n 0.00234279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_193_47#_c_603_n 0.0183573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_652_21#_M1025_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_157 VPB N_A_652_21#_M1008_g 0.0208799f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_158 VPB N_A_652_21#_c_788_n 0.00189033f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_159 VPB N_A_652_21#_c_789_n 0.00247793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_652_21#_c_784_n 0.00270641f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_161 VPB N_A_652_21#_c_791_n 0.00460198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_652_21#_c_792_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_163 VPB N_A_652_21#_c_793_n 0.00112185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_SET_B_M1029_g 0.0474843f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_165 VPB N_SET_B_M1001_g 0.0382448f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_166 VPB N_SET_B_c_901_n 0.0122147f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_167 VPB N_SET_B_c_912_n 0.00986298f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_168 VPB N_A_476_47#_M1023_g 0.0334449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_476_47#_M1016_g 0.0319182f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_170 VPB N_A_476_47#_c_1044_n 0.0121124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_476_47#_c_1038_n 0.00542515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_476_47#_c_1039_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_476_47#_c_1040_n 0.00262972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_476_47#_c_1041_n 0.030786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1178_261#_c_1193_n 0.0156579f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_176 VPB N_A_1178_261#_M1013_g 0.0268643f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=0.805
cc_177 VPB N_A_1178_261#_c_1190_n 0.02817f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_178 VPB N_A_1178_261#_c_1196_n 0.0179597f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_179 VPB N_A_1178_261#_c_1191_n 0.00603546f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.53
cc_180 VPB N_A_1178_261#_c_1198_n 0.0176834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_1178_261#_c_1199_n 0.0088754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1028_413#_M1026_g 0.0263696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1028_413#_c_1267_n 0.0117326f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_184 VPB N_A_1028_413#_M1019_g 0.0277449f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_185 VPB N_A_1028_413#_c_1272_n 0.0181611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1028_413#_c_1286_n 0.0183825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1028_413#_c_1287_n 0.0184988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1028_413#_c_1288_n 0.00417505f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1028_413#_c_1277_n 0.00164622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1028_413#_c_1290_n 0.0147146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1028_413#_c_1291_n 0.0037282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1028_413#_c_1292_n 2.84285e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1028_413#_c_1280_n 0.00129905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1028_413#_c_1281_n 0.00450937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_1786_47#_M1031_g 0.0234933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1786_47#_c_1460_n 0.0131569f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_197 VPB N_A_1786_47#_c_1455_n 0.00640788f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_198 VPB N_A_1786_47#_c_1456_n 0.00684089f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_199 VPB N_VPWR_c_1508_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_200 VPB N_VPWR_c_1509_n 0.00578936f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_201 VPB N_VPWR_c_1510_n 0.0114969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1511_n 3.97306e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1512_n 0.00366994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1513_n 0.0192032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1514_n 0.0067824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1515_n 0.00472845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1516_n 0.0331155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1517_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1518_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1519_n 0.0163072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1520_n 0.0416374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1521_n 0.0310195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1522_n 0.01851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1523_n 0.0304243f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1507_n 0.0922733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1525_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1526_n 0.00507833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1527_n 0.0091704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1528_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1529_n 0.0112536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1530_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1531_n 0.00343303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_381_47#_c_1687_n 0.00799292f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_224 VPB N_A_381_47#_c_1690_n 0.00185519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_Q_N_c_1753_n 0.0101709f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_226 VPB N_Q_c_1778_n 0.00617439f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_227 VPB N_Q_c_1776_n 0.00721226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB Q 0.0341455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 N_CLK_c_230_n N_A_27_47#_M1022_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_230 CLK N_A_27_47#_M1022_g 3.09846e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_231 N_CLK_c_234_n N_A_27_47#_M1022_g 0.00508029f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_232 N_CLK_c_237_n N_A_27_47#_M1000_g 0.0276478f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_233 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_234 N_CLK_c_233_n N_A_27_47#_M1000_g 0.00530924f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_235 N_CLK_c_230_n N_A_27_47#_c_276_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_236 N_CLK_c_231_n N_A_27_47#_c_276_n 0.00787672f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_237 CLK N_A_27_47#_c_276_n 0.00736322f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_238 N_CLK_c_231_n N_A_27_47#_c_277_n 0.0059979f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_239 CLK N_A_27_47#_c_277_n 0.014414f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_240 N_CLK_c_233_n N_A_27_47#_c_277_n 3.2891e-19 $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_241 N_CLK_c_236_n N_A_27_47#_c_291_n 0.0128144f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_237_n N_A_27_47#_c_291_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_243 CLK N_A_27_47#_c_291_n 0.00728212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_244 N_CLK_c_231_n N_A_27_47#_c_278_n 0.00189711f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_245 N_CLK_c_237_n N_A_27_47#_c_278_n 0.00440146f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_246 CLK N_A_27_47#_c_278_n 0.0517133f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_247 N_CLK_c_233_n N_A_27_47#_c_278_n 9.99252e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_248 N_CLK_c_234_n N_A_27_47#_c_278_n 0.00246929f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_249 N_CLK_c_236_n N_A_27_47#_c_295_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_250 N_CLK_c_237_n N_A_27_47#_c_295_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_251 CLK N_A_27_47#_c_295_n 0.0153363f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_252 N_CLK_c_233_n N_A_27_47#_c_295_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_253 N_CLK_c_236_n N_A_27_47#_c_297_n 0.00100532f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_254 CLK N_A_27_47#_c_286_n 0.00161876f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_255 N_CLK_c_233_n N_A_27_47#_c_286_n 0.0169694f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_256 N_CLK_c_236_n N_VPWR_c_1508_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_257 N_CLK_c_236_n N_VPWR_c_1518_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_258 N_CLK_c_236_n N_VPWR_c_1507_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_259 N_CLK_c_230_n N_VGND_c_1791_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_260 N_CLK_c_230_n N_VGND_c_1800_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_261 N_CLK_c_231_n N_VGND_c_1800_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_262 N_CLK_c_230_n N_VGND_c_1805_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_275_n N_D_M1009_g 0.0210908f $X=2.305 $Y=0.705 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_279_n N_D_M1009_g 0.00120175f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_303_n N_D_M1027_g 7.92917e-19 $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_279_n N_D_c_548_n 0.00106119f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_280_n N_D_c_548_n 0.00155965f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_279_n N_D_c_549_n 0.0453933f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_280_n N_D_c_549_n 2.37218e-19 $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_296_n N_D_c_549_n 0.00575757f $X=2.385 $Y=1.87 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_303_n N_D_c_549_n 0.00408526f $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_296_n N_A_193_47#_M1000_d 6.81311e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1033_g N_A_193_47#_M1010_g 0.0191849f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_279_n N_A_193_47#_M1010_g 0.0053439f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_296_n N_A_193_47#_M1010_g 0.00702647f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_299_n N_A_193_47#_M1010_g 5.22576e-19 $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_302_n N_A_193_47#_M1010_g 0.0174486f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_303_n N_A_193_47#_M1010_g 0.010416f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_279_n N_A_193_47#_c_586_n 0.0101526f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_298_n N_A_193_47#_c_586_n 3.63007e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_302_n N_A_193_47#_c_586_n 0.0212215f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_303_n N_A_193_47#_c_586_n 0.00655916f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_279_n N_A_193_47#_c_587_n 0.00204176f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_280_n N_A_193_47#_c_587_n 0.0232669f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_275_n N_A_193_47#_M1020_g 0.0128045f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_279_n N_A_193_47#_M1020_g 4.48322e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_280_n N_A_193_47#_M1020_g 0.0214244f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_281_n N_A_193_47#_M1011_g 0.00410946f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_282_n N_A_193_47#_M1011_g 0.0119245f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_284_n N_A_193_47#_M1011_g 0.00270619f $X=5.985 $Y=0.81 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_285_n N_A_193_47#_M1011_g 0.020941f $X=5.985 $Y=0.93 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_287_n N_A_193_47#_M1011_g 0.0125268f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1005_g N_A_193_47#_M1028_g 0.0175915f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_281_n N_A_193_47#_M1028_g 0.00220834f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_295 N_A_27_47#_c_300_n N_A_193_47#_M1028_g 0.00434444f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_304_n N_A_193_47#_M1028_g 0.0159793f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_305_n N_A_193_47#_M1028_g 0.00188266f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_281_n N_A_193_47#_c_592_n 0.00357994f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_299 N_A_27_47#_c_282_n N_A_193_47#_c_592_n 0.00341997f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_300_n N_A_193_47#_c_592_n 2.28797e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_304_n N_A_193_47#_c_592_n 0.00943741f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_305_n N_A_193_47#_c_592_n 9.97637e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_279_n N_A_193_47#_c_593_n 0.0173405f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_280_n N_A_193_47#_c_593_n 0.0059767f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1022_g N_A_193_47#_c_594_n 0.00656242f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_276_n N_A_193_47#_c_594_n 0.00216565f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_278_n N_A_193_47#_c_594_n 0.00510004f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_279_n N_A_193_47#_c_595_n 0.00886175f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_281_n N_A_193_47#_c_596_n 0.0120133f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_282_n N_A_193_47#_c_596_n 0.00159218f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_300_n N_A_193_47#_c_596_n 0.00185678f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_304_n N_A_193_47#_c_596_n 8.62653e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_305_n N_A_193_47#_c_596_n 0.00270002f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_298_n N_A_193_47#_c_597_n 0.0947033f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_279_n N_A_193_47#_c_598_n 5.02791e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_275_n N_A_193_47#_c_599_n 5.21885e-19 $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_c_279_n N_A_193_47#_c_599_n 0.0209059f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_280_n N_A_193_47#_c_599_n 0.00155193f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_302_n N_A_193_47#_c_599_n 3.45191e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_303_n N_A_193_47#_c_599_n 0.00332918f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_281_n N_A_193_47#_c_600_n 0.00256294f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_282_n N_A_193_47#_c_600_n 0.00147046f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_300_n N_A_193_47#_c_600_n 0.0122409f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_305_n N_A_193_47#_c_600_n 0.00173324f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_281_n N_A_193_47#_c_601_n 0.0285015f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_282_n N_A_193_47#_c_601_n 0.0123872f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_300_n N_A_193_47#_c_601_n 0.0012049f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_304_n N_A_193_47#_c_601_n 4.94166e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_305_n N_A_193_47#_c_601_n 0.0107523f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_279_n N_A_193_47#_c_602_n 0.00673428f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_M1022_g N_A_193_47#_c_603_n 0.0272829f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_276_n N_A_193_47#_c_603_n 0.0118856f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_403_p N_A_193_47#_c_603_n 0.00826606f $X=0.725 $Y=1.795
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_278_n N_A_193_47#_c_603_n 0.0701054f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_296_n N_A_193_47#_c_603_n 0.0247331f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_297_n N_A_193_47#_c_603_n 0.00247964f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_279_n N_A_652_21#_M1025_g 5.35023e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_298_n N_A_652_21#_M1008_g 0.00197541f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_298_n N_A_652_21#_c_788_n 0.0147195f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1005_g N_A_652_21#_c_789_n 6.75516e-19 $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_298_n N_A_652_21#_c_789_n 0.0219758f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_300_n N_A_652_21#_c_789_n 9.37384e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_305_n N_A_652_21#_c_789_n 0.00836434f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_281_n N_A_652_21#_c_784_n 0.0382594f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_298_n N_A_652_21#_c_784_n 0.00690195f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_304_n N_A_652_21#_c_784_n 2.34093e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_305_n N_A_652_21#_c_784_n 0.0123795f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_298_n N_A_652_21#_c_791_n 0.0157473f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_M1033_g N_A_652_21#_c_792_n 0.0161874f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_298_n N_A_652_21#_c_792_n 0.00193898f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_302_n N_A_652_21#_c_792_n 0.00927772f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_298_n N_A_652_21#_c_793_n 0.00782494f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_281_n N_A_652_21#_c_785_n 0.0122166f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_283_n N_A_652_21#_c_785_n 0.0108313f $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_298_n N_SET_B_M1029_g 0.00205491f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_281_n N_SET_B_c_905_n 0.00401475f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_282_n N_SET_B_c_905_n 0.0293235f $X=5.82 $Y=0.81 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_283_n N_SET_B_c_905_n 0.00586008f $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_284_n N_SET_B_c_905_n 0.0167082f $X=5.985 $Y=0.81 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_281_n N_A_476_47#_c_1033_n 3.00397e-19 $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_298_n N_A_476_47#_M1023_g 0.00187886f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_281_n N_A_476_47#_c_1034_n 0.0046475f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_282_n N_A_476_47#_c_1034_n 0.00749989f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_283_n N_A_476_47#_c_1034_n 0.00616785f $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_304_n N_A_476_47#_c_1034_n 0.00246296f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_366 N_A_27_47#_c_298_n N_A_476_47#_M1016_g 0.00301713f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_304_n N_A_476_47#_M1016_g 0.0626933f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_305_n N_A_476_47#_M1016_g 0.00173271f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_282_n N_A_476_47#_c_1035_n 0.00413822f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1033_g N_A_476_47#_c_1059_n 0.0090453f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_298_n N_A_476_47#_c_1059_n 0.00517144f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_299_n N_A_476_47#_c_1059_n 0.00306479f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_302_n N_A_476_47#_c_1059_n 0.00186639f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_303_n N_A_476_47#_c_1059_n 0.015267f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_279_n N_A_476_47#_c_1064_n 0.00676006f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_280_n N_A_476_47#_c_1064_n 9.25786e-19 $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_M1033_g N_A_476_47#_c_1044_n 0.00650943f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_279_n N_A_476_47#_c_1044_n 0.00666284f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_298_n N_A_476_47#_c_1044_n 0.013911f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_299_n N_A_476_47#_c_1044_n 0.00145075f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_302_n N_A_476_47#_c_1044_n 0.00203066f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_303_n N_A_476_47#_c_1044_n 0.0283088f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_298_n N_A_476_47#_c_1038_n 0.00472657f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_279_n N_A_476_47#_c_1039_n 0.007273f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_298_n N_A_476_47#_c_1039_n 0.00456576f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_298_n N_A_476_47#_c_1040_n 0.00248872f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_281_n N_A_476_47#_c_1041_n 0.00636379f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_298_n N_A_476_47#_c_1041_n 0.00148193f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_284_n N_A_1178_261#_M1014_g 8.41348e-19 $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_287_n N_A_1178_261#_M1014_g 0.0627906f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_284_n N_A_1178_261#_c_1190_n 3.96308e-19 $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_285_n N_A_1178_261#_c_1190_n 0.0149285f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_M1005_g N_A_1028_413#_c_1295_n 0.00494425f $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_300_n N_A_1028_413#_c_1295_n 0.00403604f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_304_n N_A_1028_413#_c_1295_n 9.00165e-19 $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_305_n N_A_1028_413#_c_1295_n 0.0148431f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_281_n N_A_1028_413#_c_1288_n 0.00537753f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_300_n N_A_1028_413#_c_1288_n 0.00765291f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_304_n N_A_1028_413#_c_1288_n 4.06473e-19 $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_305_n N_A_1028_413#_c_1288_n 0.0190128f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_282_n N_A_1028_413#_c_1303_n 0.00680222f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_284_n N_A_1028_413#_c_1303_n 0.0126727f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_285_n N_A_1028_413#_c_1303_n 5.72459e-19 $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_287_n N_A_1028_413#_c_1303_n 0.00790984f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_282_n N_A_1028_413#_c_1277_n 0.00194166f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_284_n N_A_1028_413#_c_1277_n 0.0183126f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_285_n N_A_1028_413#_c_1277_n 0.00247612f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_282_n N_A_1028_413#_c_1278_n 0.00583458f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_284_n N_A_1028_413#_c_1279_n 0.0218685f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_285_n N_A_1028_413#_c_1279_n 0.00156489f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_287_n N_A_1028_413#_c_1279_n 0.00248854f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_M1005_g N_A_1028_413#_c_1292_n 9.72583e-19 $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_403_p N_VPWR_M1018_d 6.91013e-19 $X=0.725 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_414 N_A_27_47#_c_297_n N_VPWR_M1018_d 0.00172249f $X=0.875 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_415 N_A_27_47#_M1000_g N_VPWR_c_1508_n 0.00827983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_291_n N_VPWR_c_1508_n 0.0029318f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_417 N_A_27_47#_c_403_p N_VPWR_c_1508_n 0.0133497f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_295_n N_VPWR_c_1508_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_419 N_A_27_47#_c_297_n N_VPWR_c_1508_n 0.00318756f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1000_g N_VPWR_c_1509_n 0.00190407f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_296_n N_VPWR_c_1509_n 0.00166908f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1005_g N_VPWR_c_1511_n 0.0019199f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_298_n N_VPWR_c_1511_n 0.001212f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_424 N_A_27_47#_c_291_n N_VPWR_c_1518_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_425 N_A_27_47#_c_295_n N_VPWR_c_1518_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_426 N_A_27_47#_M1000_g N_VPWR_c_1519_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_M1033_g N_VPWR_c_1520_n 0.00367119f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_M1005_g N_VPWR_c_1521_n 0.00427125f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_305_n N_VPWR_c_1521_n 0.00292005f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_M1000_g N_VPWR_c_1507_n 0.00533769f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_M1033_g N_VPWR_c_1507_n 0.00563088f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1005_g N_VPWR_c_1507_n 0.00577339f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_291_n N_VPWR_c_1507_n 0.00406578f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_295_n N_VPWR_c_1507_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_296_n N_VPWR_c_1507_n 0.0707422f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_297_n N_VPWR_c_1507_n 0.0146019f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_298_n N_VPWR_c_1507_n 0.112045f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_438 N_A_27_47#_c_299_n N_VPWR_c_1507_n 0.0160044f $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_300_n N_VPWR_c_1507_n 0.016077f $X=5.29 $Y=1.87 $X2=0 $Y2=0
cc_440 N_A_27_47#_c_303_n N_VPWR_c_1507_n 2.46058e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_c_305_n N_VPWR_c_1507_n 0.00223302f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_298_n N_VPWR_c_1527_n 0.0014214f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_296_n N_A_381_47#_M1027_d 8.84929e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_275_n N_A_381_47#_c_1692_n 0.00223782f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_279_n N_A_381_47#_c_1692_n 0.00713576f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_296_n N_A_381_47#_c_1694_n 0.019313f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_296_n N_A_381_47#_c_1690_n 0.0157335f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_275_n N_A_381_47#_c_1696_n 0.00399753f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_449 N_A_27_47#_c_296_n N_A_381_47#_c_1697_n 0.0109514f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_299_n N_A_381_47#_c_1697_n 0.00146426f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_451 N_A_27_47#_c_303_n N_A_381_47#_c_1697_n 0.00827001f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_276_n N_VGND_M1032_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_453 N_A_27_47#_M1022_g N_VGND_c_1791_n 0.0078844f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_276_n N_VGND_c_1791_n 0.0170164f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_455 N_A_27_47#_c_286_n N_VGND_c_1791_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_M1022_g N_VGND_c_1792_n 0.00296522f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_275_n N_VGND_c_1792_n 0.00120909f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_282_n N_VGND_c_1794_n 3.70426e-19 $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_283_n N_VGND_c_1794_n 0.0129707f $X=5.07 $Y=0.81 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_530_p N_VGND_c_1800_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_276_n N_VGND_c_1800_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_M1022_g N_VGND_c_1801_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_275_n N_VGND_c_1802_n 0.00556304f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_279_n N_VGND_c_1802_n 0.00113905f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_280_n N_VGND_c_1802_n 2.48118e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_M1032_s N_VGND_c_1805_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_M1022_g N_VGND_c_1805_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_275_n N_VGND_c_1805_n 0.00678262f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_c_530_p N_VGND_c_1805_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_276_n N_VGND_c_1805_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_279_n N_VGND_c_1805_n 0.00122477f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_282_n N_VGND_c_1805_n 0.00610914f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_283_n N_VGND_c_1805_n 4.92512e-19 $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_287_n N_VGND_c_1805_n 0.00522127f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_282_n N_VGND_c_1810_n 0.00797153f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_287_n N_VGND_c_1810_n 0.00368123f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_477 N_D_M1027_g N_A_193_47#_c_587_n 0.0303627f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_478 N_D_c_548_n N_A_193_47#_c_587_n 0.00467503f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_479 N_D_c_549_n N_A_193_47#_c_587_n 0.00330794f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_480 N_D_M1009_g N_A_193_47#_c_593_n 0.00395556f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_481 N_D_c_548_n N_A_193_47#_c_593_n 8.88354e-19 $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_482 N_D_c_549_n N_A_193_47#_c_593_n 0.0127149f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_483 N_D_M1009_g N_A_193_47#_c_603_n 0.00372305f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_484 N_D_M1027_g N_A_193_47#_c_603_n 0.00471318f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_485 N_D_M1027_g N_VPWR_c_1509_n 0.0116766f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_486 N_D_M1027_g N_VPWR_c_1520_n 0.0035268f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_487 N_D_M1027_g N_VPWR_c_1507_n 0.00402871f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_488 N_D_M1009_g N_A_381_47#_c_1687_n 0.00557005f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_489 N_D_M1027_g N_A_381_47#_c_1687_n 0.0115166f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_490 N_D_c_548_n N_A_381_47#_c_1687_n 0.00753248f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_491 N_D_c_549_n N_A_381_47#_c_1687_n 0.0473419f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_492 N_D_M1009_g N_A_381_47#_c_1692_n 0.0126635f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_493 N_D_c_548_n N_A_381_47#_c_1692_n 0.0014463f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_494 N_D_c_549_n N_A_381_47#_c_1692_n 0.0217898f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_495 N_D_M1027_g N_A_381_47#_c_1694_n 0.011823f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_496 N_D_c_549_n N_A_381_47#_c_1694_n 0.0109323f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_497 N_D_c_549_n N_A_381_47#_c_1697_n 0.0137404f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_498 N_D_M1009_g N_VGND_c_1792_n 0.00942273f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_499 N_D_M1009_g N_VGND_c_1802_n 0.00339367f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_500 N_D_M1009_g N_VGND_c_1805_n 0.00393034f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_501 N_A_193_47#_M1020_g N_A_652_21#_M1025_g 0.024565f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_502 N_A_193_47#_c_589_n N_A_652_21#_M1025_g 0.0114519f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_503 N_A_193_47#_c_596_n N_A_652_21#_M1025_g 9.99732e-19 $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_504 N_A_193_47#_c_598_n N_A_652_21#_M1025_g 0.00631121f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_505 N_A_193_47#_c_599_n N_A_652_21#_M1025_g 0.00191013f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_506 N_A_193_47#_c_602_n N_A_652_21#_M1025_g 0.0200607f $X=2.915 $Y=0.93 $X2=0
+ $Y2=0
cc_507 N_A_193_47#_c_596_n N_A_652_21#_c_788_n 5.47854e-19 $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_508 N_A_193_47#_c_596_n N_A_652_21#_c_789_n 0.00115455f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_509 N_A_193_47#_c_596_n N_A_652_21#_c_784_n 0.0142042f $X=5.185 $Y=1.19 $X2=0
+ $Y2=0
cc_510 N_A_193_47#_c_596_n N_A_652_21#_c_791_n 8.37667e-19 $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_511 N_A_193_47#_c_596_n N_A_652_21#_c_785_n 0.00655125f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_512 N_A_193_47#_c_596_n N_SET_B_c_897_n 0.00381498f $X=5.185 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_513 N_A_193_47#_c_596_n N_SET_B_M1029_g 0.00121673f $X=5.185 $Y=1.19 $X2=0
+ $Y2=0
cc_514 N_A_193_47#_c_596_n SET_B 0.00570533f $X=5.185 $Y=1.19 $X2=0 $Y2=0
cc_515 N_A_193_47#_M1011_g N_SET_B_c_905_n 0.00480049f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_516 N_A_193_47#_c_591_n N_SET_B_c_905_n 3.54642e-19 $X=5.605 $Y=1.455 $X2=0
+ $Y2=0
cc_517 N_A_193_47#_c_592_n N_SET_B_c_905_n 3.96195e-19 $X=5.47 $Y=1.26 $X2=0
+ $Y2=0
cc_518 N_A_193_47#_c_596_n N_SET_B_c_905_n 0.0895102f $X=5.185 $Y=1.19 $X2=0
+ $Y2=0
cc_519 N_A_193_47#_c_600_n N_SET_B_c_905_n 0.02693f $X=5.33 $Y=1.19 $X2=0 $Y2=0
cc_520 N_A_193_47#_c_601_n N_SET_B_c_905_n 0.00112669f $X=5.33 $Y=1.19 $X2=0
+ $Y2=0
cc_521 N_A_193_47#_c_596_n N_SET_B_c_906_n 0.0263312f $X=5.185 $Y=1.19 $X2=0
+ $Y2=0
cc_522 N_A_193_47#_c_596_n N_A_476_47#_c_1033_n 0.00253485f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_523 N_A_193_47#_c_592_n N_A_476_47#_c_1034_n 0.00775418f $X=5.47 $Y=1.26
+ $X2=0 $Y2=0
cc_524 N_A_193_47#_c_596_n N_A_476_47#_c_1034_n 0.001113f $X=5.185 $Y=1.19 $X2=0
+ $Y2=0
cc_525 N_A_193_47#_c_601_n N_A_476_47#_c_1034_n 2.11256e-19 $X=5.33 $Y=1.19
+ $X2=0 $Y2=0
cc_526 N_A_193_47#_M1011_g N_A_476_47#_c_1035_n 0.0518139f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_527 N_A_193_47#_M1010_g N_A_476_47#_c_1059_n 0.00278769f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_528 N_A_193_47#_M1020_g N_A_476_47#_c_1064_n 0.008828f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_529 N_A_193_47#_c_593_n N_A_476_47#_c_1064_n 0.00573977f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_530 N_A_193_47#_c_598_n N_A_476_47#_c_1064_n 0.00194059f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_531 N_A_193_47#_c_599_n N_A_476_47#_c_1064_n 0.0194974f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_532 N_A_193_47#_c_602_n N_A_476_47#_c_1064_n 5.24271e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_533 N_A_193_47#_M1010_g N_A_476_47#_c_1044_n 8.73767e-19 $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_534 N_A_193_47#_c_597_n N_A_476_47#_c_1044_n 3.07745e-19 $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_535 N_A_193_47#_M1020_g N_A_476_47#_c_1037_n 0.00118778f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_536 N_A_193_47#_c_589_n N_A_476_47#_c_1037_n 7.74259e-19 $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_c_596_n N_A_476_47#_c_1037_n 0.0146154f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_538 N_A_193_47#_c_598_n N_A_476_47#_c_1037_n 0.0134967f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_539 N_A_193_47#_c_599_n N_A_476_47#_c_1037_n 0.0244992f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_540 N_A_193_47#_c_602_n N_A_476_47#_c_1037_n 7.73887e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_541 N_A_193_47#_c_596_n N_A_476_47#_c_1038_n 0.0232188f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_542 N_A_193_47#_c_589_n N_A_476_47#_c_1039_n 0.00262762f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_c_596_n N_A_476_47#_c_1039_n 0.0121342f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_544 N_A_193_47#_c_597_n N_A_476_47#_c_1039_n 0.00535278f $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_599_n N_A_476_47#_c_1039_n 0.00527199f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_602_n N_A_476_47#_c_1039_n 5.70501e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_c_596_n N_A_476_47#_c_1040_n 0.00996075f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_c_591_n N_A_476_47#_c_1041_n 5.77474e-19 $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_592_n N_A_476_47#_c_1041_n 0.0044662f $X=5.47 $Y=1.26 $X2=0
+ $Y2=0
cc_550 N_A_193_47#_c_596_n N_A_476_47#_c_1041_n 0.00413707f $X=5.185 $Y=1.19
+ $X2=0 $Y2=0
cc_551 N_A_193_47#_M1011_g N_A_1178_261#_M1014_g 0.00242755f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_552 N_A_193_47#_c_591_n N_A_1178_261#_c_1190_n 0.0407002f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_553 N_A_193_47#_M1028_g N_A_1178_261#_c_1196_n 0.0407002f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_554 N_A_193_47#_M1028_g N_A_1028_413#_c_1295_n 0.00929093f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_555 N_A_193_47#_c_591_n N_A_1028_413#_c_1288_n 0.00100314f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_556 N_A_193_47#_M1028_g N_A_1028_413#_c_1288_n 0.00996215f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_557 N_A_193_47#_c_601_n N_A_1028_413#_c_1288_n 0.00496129f $X=5.33 $Y=1.19
+ $X2=0 $Y2=0
cc_558 N_A_193_47#_c_591_n N_A_1028_413#_c_1278_n 0.0075541f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_559 N_A_193_47#_c_600_n N_A_1028_413#_c_1278_n 0.00200974f $X=5.33 $Y=1.19
+ $X2=0 $Y2=0
cc_560 N_A_193_47#_c_601_n N_A_1028_413#_c_1278_n 0.0123133f $X=5.33 $Y=1.19
+ $X2=0 $Y2=0
cc_561 N_A_193_47#_M1028_g N_A_1028_413#_c_1290_n 2.12512e-19 $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_562 N_A_193_47#_M1011_g N_A_1028_413#_c_1279_n 0.00203086f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_563 N_A_193_47#_M1028_g N_A_1028_413#_c_1292_n 0.0109424f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_564 N_A_193_47#_c_603_n N_VPWR_c_1508_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_565 N_A_193_47#_M1010_g N_VPWR_c_1509_n 0.00113058f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_566 N_A_193_47#_c_603_n N_VPWR_c_1509_n 0.0226552f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_567 N_A_193_47#_c_603_n N_VPWR_c_1519_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_568 N_A_193_47#_M1010_g N_VPWR_c_1520_n 0.00541732f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_569 N_A_193_47#_M1028_g N_VPWR_c_1521_n 0.00369452f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_570 N_A_193_47#_M1010_g N_VPWR_c_1507_n 0.00628966f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_571 N_A_193_47#_M1028_g N_VPWR_c_1507_n 0.00544637f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_572 N_A_193_47#_c_603_n N_VPWR_c_1507_n 0.00409094f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_573 N_A_193_47#_M1028_g N_VPWR_c_1529_n 0.00192611f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_574 N_A_193_47#_c_593_n N_A_381_47#_M1009_d 4.25819e-19 $X=2.845 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_575 N_A_193_47#_c_593_n N_A_381_47#_c_1687_n 0.0148354f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_576 N_A_193_47#_c_594_n N_A_381_47#_c_1687_n 0.00135406f $X=1.295 $Y=0.85
+ $X2=0 $Y2=0
cc_577 N_A_193_47#_c_603_n N_A_381_47#_c_1687_n 0.0675361f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_578 N_A_193_47#_c_593_n N_A_381_47#_c_1692_n 0.0198802f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_579 N_A_193_47#_c_599_n N_A_381_47#_c_1692_n 0.00201969f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_580 N_A_193_47#_c_593_n N_A_381_47#_c_1688_n 0.00435863f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_581 N_A_193_47#_c_594_n N_A_381_47#_c_1688_n 0.00140429f $X=1.295 $Y=0.85
+ $X2=0 $Y2=0
cc_582 N_A_193_47#_c_603_n N_A_381_47#_c_1688_n 0.0138352f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_583 N_A_193_47#_c_603_n N_A_381_47#_c_1690_n 0.011423f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_584 N_A_193_47#_M1010_g N_A_381_47#_c_1697_n 0.0102511f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_585 N_A_193_47#_c_593_n N_VGND_c_1792_n 0.0012296f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_586 N_A_193_47#_c_603_n N_VGND_c_1792_n 0.00823827f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_587 N_A_193_47#_c_603_n N_VGND_c_1801_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_588 N_A_193_47#_M1020_g N_VGND_c_1802_n 0.00359964f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_589 N_A_193_47#_M1022_d N_VGND_c_1805_n 0.00324958f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_590 N_A_193_47#_M1020_g N_VGND_c_1805_n 0.0056346f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_591 N_A_193_47#_M1011_g N_VGND_c_1805_n 0.00571363f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_592 N_A_193_47#_c_593_n N_VGND_c_1805_n 0.072327f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_593 N_A_193_47#_c_594_n N_VGND_c_1805_n 0.0151383f $X=1.295 $Y=0.85 $X2=0
+ $Y2=0
cc_594 N_A_193_47#_c_598_n N_VGND_c_1805_n 0.0151785f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_595 N_A_193_47#_c_603_n N_VGND_c_1805_n 0.00372614f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_596 N_A_193_47#_M1011_g N_VGND_c_1810_n 0.00437852f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_597 N_A_193_47#_c_599_n A_586_47# 0.00109469f $X=2.99 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_598 N_A_652_21#_M1025_g N_SET_B_c_897_n 0.0189903f $X=3.335 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_599 N_A_652_21#_c_784_n N_SET_B_c_897_n 7.60504e-19 $X=4.625 $Y=1.835
+ $X2=-0.19 $Y2=-0.24
cc_600 N_A_652_21#_M1025_g N_SET_B_M1029_g 0.0137896f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_601 N_A_652_21#_M1008_g N_SET_B_M1029_g 0.0113783f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_602 N_A_652_21#_c_788_n N_SET_B_M1029_g 0.0139954f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_603 N_A_652_21#_c_791_n N_SET_B_M1029_g 0.00563707f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_604 N_A_652_21#_c_792_n N_SET_B_M1029_g 0.0201938f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_605 N_A_652_21#_M1025_g N_SET_B_M1004_g 0.0141659f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_606 N_A_652_21#_c_783_n N_SET_B_M1004_g 0.00124922f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_607 N_A_652_21#_c_785_n N_SET_B_M1004_g 3.79232e-19 $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_608 N_A_652_21#_M1025_g SET_B 0.00110794f $X=3.335 $Y=0.445 $X2=0 $Y2=0
cc_609 N_A_652_21#_c_785_n SET_B 0.0144281f $X=4.625 $Y=0.895 $X2=0 $Y2=0
cc_610 N_A_652_21#_c_783_n N_SET_B_c_905_n 9.52814e-19 $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_611 N_A_652_21#_c_785_n N_SET_B_c_905_n 0.019808f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_612 N_A_652_21#_c_785_n N_SET_B_c_906_n 0.00250762f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_613 N_A_652_21#_c_783_n N_A_476_47#_c_1032_n 0.00809901f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_614 N_A_652_21#_c_785_n N_A_476_47#_c_1032_n 4.65467e-19 $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_615 N_A_652_21#_c_784_n N_A_476_47#_c_1033_n 0.00246574f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_616 N_A_652_21#_c_785_n N_A_476_47#_c_1033_n 0.0035345f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_617 N_A_652_21#_c_789_n N_A_476_47#_M1023_g 0.0138123f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_618 N_A_652_21#_c_784_n N_A_476_47#_M1023_g 0.00531645f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_619 N_A_652_21#_c_783_n N_A_476_47#_c_1034_n 0.00253676f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_620 N_A_652_21#_c_784_n N_A_476_47#_c_1034_n 2.06235e-19 $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_621 N_A_652_21#_c_785_n N_A_476_47#_c_1034_n 0.0150104f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_622 N_A_652_21#_c_789_n N_A_476_47#_M1016_g 0.00849064f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_623 N_A_652_21#_c_784_n N_A_476_47#_M1016_g 0.00519116f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_624 N_A_652_21#_c_783_n N_A_476_47#_c_1035_n 0.00422581f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_625 N_A_652_21#_c_785_n N_A_476_47#_c_1036_n 0.00182302f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_626 N_A_652_21#_M1008_g N_A_476_47#_c_1059_n 0.00202046f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_627 N_A_652_21#_M1025_g N_A_476_47#_c_1064_n 0.00854236f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_628 N_A_652_21#_M1025_g N_A_476_47#_c_1044_n 0.015293f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_629 N_A_652_21#_c_791_n N_A_476_47#_c_1044_n 0.0366983f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_630 N_A_652_21#_M1025_g N_A_476_47#_c_1037_n 0.0188229f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_631 N_A_652_21#_c_788_n N_A_476_47#_c_1038_n 0.00881126f $X=3.99 $Y=1.96
+ $X2=0 $Y2=0
cc_632 N_A_652_21#_c_793_n N_A_476_47#_c_1038_n 0.00337624f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_633 N_A_652_21#_M1025_g N_A_476_47#_c_1039_n 0.0109017f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_634 N_A_652_21#_c_791_n N_A_476_47#_c_1039_n 0.0171213f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_635 N_A_652_21#_c_792_n N_A_476_47#_c_1039_n 0.0011995f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_636 N_A_652_21#_c_789_n N_A_476_47#_c_1040_n 0.0079382f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_637 N_A_652_21#_c_784_n N_A_476_47#_c_1040_n 0.0229291f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_638 N_A_652_21#_c_793_n N_A_476_47#_c_1040_n 0.00169427f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_639 N_A_652_21#_c_785_n N_A_476_47#_c_1040_n 0.0037745f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_640 N_A_652_21#_c_789_n N_A_476_47#_c_1041_n 0.0029883f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_641 N_A_652_21#_c_784_n N_A_476_47#_c_1041_n 0.0132275f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_642 N_A_652_21#_c_785_n N_A_476_47#_c_1041_n 0.00437877f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_643 N_A_652_21#_c_788_n N_VPWR_M1008_d 0.00131929f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_644 N_A_652_21#_c_791_n N_VPWR_M1008_d 0.00154452f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_645 N_A_652_21#_c_789_n N_VPWR_M1023_d 0.00161389f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_646 N_A_652_21#_c_788_n N_VPWR_c_1510_n 0.00266175f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_647 N_A_652_21#_c_872_p N_VPWR_c_1510_n 0.0070924f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_648 N_A_652_21#_c_789_n N_VPWR_c_1510_n 0.00248431f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_649 N_A_652_21#_c_789_n N_VPWR_c_1511_n 0.0155298f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_650 N_A_652_21#_M1008_g N_VPWR_c_1520_n 0.00532975f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_651 N_A_652_21#_c_791_n N_VPWR_c_1520_n 0.00105935f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_652 N_A_652_21#_c_789_n N_VPWR_c_1521_n 8.80252e-19 $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_653 N_A_652_21#_M1029_d N_VPWR_c_1507_n 0.00202389f $X=3.94 $Y=2.065 $X2=0
+ $Y2=0
cc_654 N_A_652_21#_M1008_g N_VPWR_c_1507_n 0.0066225f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_655 N_A_652_21#_c_788_n N_VPWR_c_1507_n 0.00255051f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_656 N_A_652_21#_c_872_p N_VPWR_c_1507_n 0.00288476f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_657 N_A_652_21#_c_789_n N_VPWR_c_1507_n 0.0034475f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_658 N_A_652_21#_c_791_n N_VPWR_c_1507_n 0.00138626f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_659 N_A_652_21#_M1008_g N_VPWR_c_1527_n 0.00326498f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_660 N_A_652_21#_c_788_n N_VPWR_c_1527_n 0.0101842f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_661 N_A_652_21#_c_791_n N_VPWR_c_1527_n 0.0109284f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_662 N_A_652_21#_c_792_n N_VPWR_c_1527_n 6.81742e-19 $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_663 N_A_652_21#_M1025_g N_VGND_c_1793_n 0.0040279f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_664 N_A_652_21#_c_783_n N_VGND_c_1794_n 0.0192612f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_665 N_A_652_21#_M1025_g N_VGND_c_1802_n 0.0035977f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_666 N_A_652_21#_c_783_n N_VGND_c_1803_n 0.0118981f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_667 N_A_652_21#_c_785_n N_VGND_c_1803_n 0.00244068f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_668 N_A_652_21#_M1006_d N_VGND_c_1805_n 0.00186029f $X=4.34 $Y=0.235 $X2=0
+ $Y2=0
cc_669 N_A_652_21#_M1025_g N_VGND_c_1805_n 0.00580574f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_670 N_A_652_21#_c_783_n N_VGND_c_1805_n 0.00426169f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_671 N_A_652_21#_c_785_n N_VGND_c_1805_n 0.00183644f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_672 N_SET_B_M1004_g N_A_476_47#_c_1032_n 0.0270653f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_897_n N_A_476_47#_c_1033_n 0.0146844f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_905_n N_A_476_47#_c_1033_n 8.12862e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_906_n N_A_476_47#_c_1033_n 7.28461e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_676 N_SET_B_M1029_g N_A_476_47#_M1023_g 0.0336841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_905_n N_A_476_47#_c_1034_n 0.00272702f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_897_n N_A_476_47#_c_1036_n 0.0270653f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_679 SET_B N_A_476_47#_c_1036_n 0.0021684f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_680 N_SET_B_c_905_n N_A_476_47#_c_1036_n 0.00277782f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_906_n N_A_476_47#_c_1036_n 7.28461e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_897_n N_A_476_47#_c_1037_n 0.00218199f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_683 N_SET_B_M1029_g N_A_476_47#_c_1037_n 6.04572e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_684 N_SET_B_M1004_g N_A_476_47#_c_1037_n 0.00184201f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_685 SET_B N_A_476_47#_c_1037_n 0.0243988f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_686 N_SET_B_c_906_n N_A_476_47#_c_1037_n 0.00116251f $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_897_n N_A_476_47#_c_1038_n 0.00307815f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_688 N_SET_B_M1029_g N_A_476_47#_c_1038_n 0.0103672f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_689 SET_B N_A_476_47#_c_1038_n 0.0263655f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_690 N_SET_B_c_905_n N_A_476_47#_c_1038_n 3.66303e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_906_n N_A_476_47#_c_1038_n 5.23607e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_692 N_SET_B_M1029_g N_A_476_47#_c_1039_n 5.20457e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_693 N_SET_B_M1029_g N_A_476_47#_c_1040_n 0.00354841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_905_n N_A_476_47#_c_1040_n 0.00236582f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_695 N_SET_B_M1029_g N_A_476_47#_c_1041_n 0.0205296f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_901_n N_A_1178_261#_c_1193_n 0.00246223f $X=6.895 $Y=1.535
+ $X2=0 $Y2=0
cc_697 N_SET_B_M1021_g N_A_1178_261#_M1014_g 0.0658096f $X=6.765 $Y=0.445 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_901_n N_A_1178_261#_M1014_g 0.0116464f $X=6.895 $Y=1.535 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_903_n N_A_1178_261#_M1014_g 0.00104156f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_700 N_SET_B_M1001_g N_A_1178_261#_c_1196_n 0.00297289f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_701 N_SET_B_c_912_n N_A_1178_261#_c_1196_n 0.00246223f $X=6.895 $Y=1.685
+ $X2=0 $Y2=0
cc_702 N_SET_B_c_902_n N_A_1178_261#_c_1191_n 3.84308e-19 $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_903_n N_A_1178_261#_c_1191_n 0.00169497f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_907_n N_A_1178_261#_c_1191_n 0.00146176f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_908_n N_A_1178_261#_c_1191_n 0.0115867f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_706 N_SET_B_M1001_g N_A_1178_261#_c_1198_n 0.00934654f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_707 N_SET_B_c_912_n N_A_1178_261#_c_1198_n 0.00775501f $X=6.895 $Y=1.685
+ $X2=0 $Y2=0
cc_708 N_SET_B_M1021_g N_A_1028_413#_M1017_g 0.0164357f $X=6.765 $Y=0.445 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_902_n N_A_1028_413#_M1017_g 0.00975744f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_903_n N_A_1028_413#_M1017_g 5.97128e-19 $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_711 N_SET_B_c_908_n N_A_1028_413#_M1017_g 0.00790355f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_901_n N_A_1028_413#_M1026_g 0.00412516f $X=6.895 $Y=1.535 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_912_n N_A_1028_413#_M1026_g 0.0260901f $X=6.895 $Y=1.685 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_902_n N_A_1028_413#_c_1267_n 0.0216918f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_908_n N_A_1028_413#_c_1267_n 0.00349124f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_905_n N_A_1028_413#_c_1303_n 0.00655755f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_905_n N_A_1028_413#_c_1277_n 0.0101452f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_905_n N_A_1028_413#_c_1278_n 0.00400606f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_719 N_SET_B_M1001_g N_A_1028_413#_c_1290_n 0.00433068f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_720 N_SET_B_M1021_g N_A_1028_413#_c_1279_n 0.00258467f $X=6.765 $Y=0.445
+ $X2=0 $Y2=0
cc_721 N_SET_B_c_901_n N_A_1028_413#_c_1279_n 0.00102632f $X=6.895 $Y=1.535
+ $X2=0 $Y2=0
cc_722 N_SET_B_c_902_n N_A_1028_413#_c_1279_n 0.00158445f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_903_n N_A_1028_413#_c_1279_n 0.0254752f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_905_n N_A_1028_413#_c_1279_n 0.0180658f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_907_n N_A_1028_413#_c_1279_n 3.39847e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_901_n N_A_1028_413#_c_1280_n 6.19496e-19 $X=6.895 $Y=1.535
+ $X2=0 $Y2=0
cc_727 N_SET_B_c_907_n N_A_1028_413#_c_1280_n 8.97025e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_908_n N_A_1028_413#_c_1280_n 0.0128812f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_901_n N_A_1028_413#_c_1281_n 0.0101835f $X=6.895 $Y=1.535 $X2=0
+ $Y2=0
cc_730 N_SET_B_c_912_n N_A_1028_413#_c_1281_n 5.5231e-19 $X=6.895 $Y=1.685 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_902_n N_A_1028_413#_c_1281_n 0.00347344f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_903_n N_A_1028_413#_c_1281_n 0.0229264f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_905_n N_A_1028_413#_c_1281_n 0.00838415f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_734 N_SET_B_c_907_n N_A_1028_413#_c_1281_n 0.00102488f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_908_n N_A_1028_413#_c_1281_n 0.00830557f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_SET_B_M1029_g N_VPWR_c_1510_n 0.00368415f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_737 N_SET_B_M1029_g N_VPWR_c_1511_n 7.26951e-19 $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_738 N_SET_B_M1001_g N_VPWR_c_1512_n 0.00327827f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_739 N_SET_B_M1001_g N_VPWR_c_1522_n 0.00585385f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_740 N_SET_B_M1029_g N_VPWR_c_1507_n 0.00406312f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_741 N_SET_B_M1001_g N_VPWR_c_1507_n 0.0121898f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_742 N_SET_B_M1029_g N_VPWR_c_1527_n 0.00699603f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_743 N_SET_B_M1001_g N_VPWR_c_1529_n 0.00306241f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_744 N_SET_B_c_907_n N_VGND_M1021_d 0.00132095f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_745 N_SET_B_c_908_n N_VGND_M1021_d 9.16065e-19 $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_746 N_SET_B_c_897_n N_VGND_c_1793_n 0.00103531f $X=3.865 $Y=1.145 $X2=0 $Y2=0
cc_747 N_SET_B_M1004_g N_VGND_c_1793_n 0.0134999f $X=3.905 $Y=0.445 $X2=0 $Y2=0
cc_748 SET_B N_VGND_c_1793_n 0.0213368f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_749 N_SET_B_c_906_n N_VGND_c_1793_n 0.00267196f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_750 N_SET_B_c_905_n N_VGND_c_1794_n 0.00622223f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_751 N_SET_B_c_903_n N_VGND_c_1805_n 0.00105154f $X=6.99 $Y=0.9 $X2=0 $Y2=0
cc_752 SET_B N_VGND_c_1805_n 9.94995e-19 $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_753 N_SET_B_c_905_n N_VGND_c_1805_n 0.134825f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_754 N_SET_B_c_906_n N_VGND_c_1805_n 0.0146581f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_755 N_SET_B_c_907_n N_VGND_c_1805_n 0.0145559f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_756 N_SET_B_M1021_g N_VGND_c_1811_n 0.0199195f $X=6.765 $Y=0.445 $X2=0 $Y2=0
cc_757 N_SET_B_c_902_n N_VGND_c_1811_n 6.12458e-19 $X=6.825 $Y=0.98 $X2=0 $Y2=0
cc_758 N_SET_B_c_903_n N_VGND_c_1811_n 0.0401429f $X=6.99 $Y=0.9 $X2=0 $Y2=0
cc_759 N_SET_B_c_905_n N_VGND_c_1811_n 0.00146726f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_760 N_SET_B_c_907_n N_VGND_c_1811_n 0.00339972f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_761 N_A_476_47#_M1016_g N_A_1028_413#_c_1295_n 8.83644e-19 $X=4.705 $Y=2.275
+ $X2=0 $Y2=0
cc_762 N_A_476_47#_M1023_g N_VPWR_c_1510_n 0.00339367f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_763 N_A_476_47#_M1023_g N_VPWR_c_1511_n 0.00730335f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_764 N_A_476_47#_M1016_g N_VPWR_c_1511_n 0.00909428f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_765 N_A_476_47#_c_1059_n N_VPWR_c_1520_n 0.0377433f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_766 N_A_476_47#_M1016_g N_VPWR_c_1521_n 0.00414121f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_767 N_A_476_47#_M1010_d N_VPWR_c_1507_n 0.00172638f $X=2.39 $Y=2.065 $X2=0
+ $Y2=0
cc_768 N_A_476_47#_M1023_g N_VPWR_c_1507_n 0.00379591f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_769 N_A_476_47#_M1016_g N_VPWR_c_1507_n 0.00402125f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_770 N_A_476_47#_c_1059_n N_VPWR_c_1507_n 0.0132505f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_771 N_A_476_47#_M1023_g N_VPWR_c_1527_n 7.14614e-19 $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_772 N_A_476_47#_c_1059_n N_A_381_47#_c_1697_n 0.0102747f $X=3.02 $Y=2.335
+ $X2=0 $Y2=0
cc_773 N_A_476_47#_c_1059_n A_562_413# 0.00859792f $X=3.02 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_774 N_A_476_47#_c_1044_n A_562_413# 0.00578953f $X=3.105 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_775 N_A_476_47#_c_1032_n N_VGND_c_1793_n 0.00301834f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_776 N_A_476_47#_c_1032_n N_VGND_c_1794_n 0.00375773f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_777 N_A_476_47#_c_1034_n N_VGND_c_1794_n 0.00746256f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_778 N_A_476_47#_c_1035_n N_VGND_c_1794_n 0.00458594f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_779 N_A_476_47#_c_1064_n N_VGND_c_1802_n 0.055608f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_780 N_A_476_47#_c_1032_n N_VGND_c_1803_n 0.00541969f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_781 N_A_476_47#_c_1034_n N_VGND_c_1803_n 0.00110285f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_782 N_A_476_47#_M1030_d N_VGND_c_1805_n 0.00275359f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_783 N_A_476_47#_c_1032_n N_VGND_c_1805_n 0.00742824f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_784 N_A_476_47#_c_1034_n N_VGND_c_1805_n 3.98471e-19 $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_785 N_A_476_47#_c_1035_n N_VGND_c_1805_n 0.00674913f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_786 N_A_476_47#_c_1064_n N_VGND_c_1805_n 0.0223868f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_787 N_A_476_47#_c_1035_n N_VGND_c_1810_n 0.00437852f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_788 N_A_476_47#_c_1064_n A_586_47# 0.00628999f $X=3.27 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_789 N_A_1178_261#_c_1191_n N_A_1028_413#_M1017_g 0.00743522f $X=7.735
+ $Y=1.575 $X2=0 $Y2=0
cc_790 N_A_1178_261#_c_1198_n N_A_1028_413#_M1026_g 0.0144868f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_791 N_A_1178_261#_c_1191_n N_A_1028_413#_c_1266_n 0.0241648f $X=7.735
+ $Y=1.575 $X2=0 $Y2=0
cc_792 N_A_1178_261#_c_1192_n N_A_1028_413#_c_1266_n 0.00356732f $X=7.735
+ $Y=0.515 $X2=0 $Y2=0
cc_793 N_A_1178_261#_c_1199_n N_A_1028_413#_c_1266_n 0.00367651f $X=7.735
+ $Y=1.67 $X2=0 $Y2=0
cc_794 N_A_1178_261#_c_1191_n N_A_1028_413#_c_1267_n 0.00666201f $X=7.735
+ $Y=1.575 $X2=0 $Y2=0
cc_795 N_A_1178_261#_c_1198_n N_A_1028_413#_c_1267_n 0.0032134f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_796 N_A_1178_261#_c_1191_n N_A_1028_413#_M1007_g 0.00237066f $X=7.735
+ $Y=1.575 $X2=0 $Y2=0
cc_797 N_A_1178_261#_c_1191_n N_A_1028_413#_M1019_g 0.00326859f $X=7.735
+ $Y=1.575 $X2=0 $Y2=0
cc_798 N_A_1178_261#_c_1190_n N_A_1028_413#_c_1288_n 0.00412466f $X=6.405
+ $Y=1.38 $X2=0 $Y2=0
cc_799 N_A_1178_261#_c_1198_n N_A_1028_413#_c_1288_n 0.0133831f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_800 N_A_1178_261#_M1014_g N_A_1028_413#_c_1303_n 0.00576956f $X=6.405
+ $Y=0.445 $X2=0 $Y2=0
cc_801 N_A_1178_261#_c_1190_n N_A_1028_413#_c_1277_n 0.0144229f $X=6.405 $Y=1.38
+ $X2=0 $Y2=0
cc_802 N_A_1178_261#_c_1198_n N_A_1028_413#_c_1277_n 0.026737f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_803 N_A_1178_261#_M1013_g N_A_1028_413#_c_1290_n 0.0121476f $X=5.965 $Y=2.275
+ $X2=0 $Y2=0
cc_804 N_A_1178_261#_c_1196_n N_A_1028_413#_c_1290_n 0.00514123f $X=6.095
+ $Y=1.66 $X2=0 $Y2=0
cc_805 N_A_1178_261#_c_1198_n N_A_1028_413#_c_1290_n 0.0639862f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_806 N_A_1178_261#_M1014_g N_A_1028_413#_c_1279_n 0.0142383f $X=6.405 $Y=0.445
+ $X2=0 $Y2=0
cc_807 N_A_1178_261#_M1013_g N_A_1028_413#_c_1291_n 0.00296198f $X=5.965
+ $Y=2.275 $X2=0 $Y2=0
cc_808 N_A_1178_261#_M1013_g N_A_1028_413#_c_1292_n 0.00455504f $X=5.965
+ $Y=2.275 $X2=0 $Y2=0
cc_809 N_A_1178_261#_c_1196_n N_A_1028_413#_c_1292_n 0.00412466f $X=6.095
+ $Y=1.66 $X2=0 $Y2=0
cc_810 N_A_1178_261#_M1014_g N_A_1028_413#_c_1375_n 0.00331097f $X=6.405
+ $Y=0.445 $X2=0 $Y2=0
cc_811 N_A_1178_261#_c_1190_n N_A_1028_413#_c_1375_n 0.00412185f $X=6.405
+ $Y=1.38 $X2=0 $Y2=0
cc_812 N_A_1178_261#_c_1198_n N_A_1028_413#_c_1375_n 0.0136304f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_813 N_A_1178_261#_c_1191_n N_A_1028_413#_c_1280_n 0.0181507f $X=7.735
+ $Y=1.575 $X2=0 $Y2=0
cc_814 N_A_1178_261#_c_1198_n N_A_1028_413#_c_1281_n 0.0708842f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_815 N_A_1178_261#_c_1198_n N_VPWR_M1001_d 0.00225674f $X=7.51 $Y=1.67 $X2=0
+ $Y2=0
cc_816 N_A_1178_261#_c_1198_n N_VPWR_c_1512_n 0.0195228f $X=7.51 $Y=1.67 $X2=0
+ $Y2=0
cc_817 N_A_1178_261#_c_1247_p N_VPWR_c_1513_n 0.00727431f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_818 N_A_1178_261#_c_1247_p N_VPWR_c_1514_n 0.0267353f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_819 N_A_1178_261#_c_1191_n N_VPWR_c_1514_n 0.00657492f $X=7.735 $Y=1.575
+ $X2=0 $Y2=0
cc_820 N_A_1178_261#_c_1199_n N_VPWR_c_1514_n 0.0143842f $X=7.735 $Y=1.67 $X2=0
+ $Y2=0
cc_821 N_A_1178_261#_M1013_g N_VPWR_c_1521_n 0.00113358f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_822 N_A_1178_261#_M1026_d N_VPWR_c_1507_n 0.00535012f $X=7.46 $Y=1.645 $X2=0
+ $Y2=0
cc_823 N_A_1178_261#_M1013_g N_VPWR_c_1507_n 0.00171818f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_824 N_A_1178_261#_c_1247_p N_VPWR_c_1507_n 0.00614354f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_825 N_A_1178_261#_M1013_g N_VPWR_c_1529_n 0.0139543f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_826 N_A_1178_261#_c_1191_n N_Q_N_c_1753_n 0.0171749f $X=7.735 $Y=1.575 $X2=0
+ $Y2=0
cc_827 N_A_1178_261#_c_1192_n N_VGND_c_1795_n 0.0131701f $X=7.735 $Y=0.515 $X2=0
+ $Y2=0
cc_828 N_A_1178_261#_c_1191_n N_VGND_c_1796_n 0.0155836f $X=7.735 $Y=1.575 $X2=0
+ $Y2=0
cc_829 N_A_1178_261#_c_1192_n N_VGND_c_1796_n 0.0237335f $X=7.735 $Y=0.515 $X2=0
+ $Y2=0
cc_830 N_A_1178_261#_M1017_d N_VGND_c_1805_n 0.00391384f $X=7.46 $Y=0.235 $X2=0
+ $Y2=0
cc_831 N_A_1178_261#_M1014_g N_VGND_c_1805_n 0.00495706f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_832 N_A_1178_261#_c_1192_n N_VGND_c_1805_n 0.0114301f $X=7.735 $Y=0.515 $X2=0
+ $Y2=0
cc_833 N_A_1178_261#_M1014_g N_VGND_c_1810_n 0.00367922f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_834 N_A_1178_261#_M1014_g N_VGND_c_1811_n 0.00248483f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_835 N_A_1028_413#_c_1272_n N_A_1786_47#_M1031_g 0.0064039f $X=9.135 $Y=1.62
+ $X2=0 $Y2=0
cc_836 N_A_1028_413#_c_1287_n N_A_1786_47#_M1031_g 0.0128064f $X=9.265 $Y=1.695
+ $X2=0 $Y2=0
cc_837 N_A_1028_413#_M1007_g N_A_1786_47#_c_1454_n 0.00124425f $X=8.325 $Y=0.56
+ $X2=0 $Y2=0
cc_838 N_A_1028_413#_c_1271_n N_A_1786_47#_c_1454_n 0.00392984f $X=9.135
+ $Y=1.025 $X2=0 $Y2=0
cc_839 N_A_1028_413#_c_1273_n N_A_1786_47#_c_1454_n 0.00968345f $X=9.265 $Y=0.73
+ $X2=0 $Y2=0
cc_840 N_A_1028_413#_c_1275_n N_A_1786_47#_c_1454_n 0.0100252f $X=9.265 $Y=0.805
+ $X2=0 $Y2=0
cc_841 N_A_1028_413#_M1019_g N_A_1786_47#_c_1460_n 0.00191035f $X=8.325 $Y=1.985
+ $X2=0 $Y2=0
cc_842 N_A_1028_413#_c_1272_n N_A_1786_47#_c_1460_n 0.0101898f $X=9.135 $Y=1.62
+ $X2=0 $Y2=0
cc_843 N_A_1028_413#_c_1286_n N_A_1786_47#_c_1460_n 0.010339f $X=9.265 $Y=1.77
+ $X2=0 $Y2=0
cc_844 N_A_1028_413#_c_1287_n N_A_1786_47#_c_1460_n 0.0102457f $X=9.265 $Y=1.695
+ $X2=0 $Y2=0
cc_845 N_A_1028_413#_c_1275_n N_A_1786_47#_c_1455_n 0.00562989f $X=9.265
+ $Y=0.805 $X2=0 $Y2=0
cc_846 N_A_1028_413#_c_1287_n N_A_1786_47#_c_1455_n 0.0046403f $X=9.265 $Y=1.695
+ $X2=0 $Y2=0
cc_847 N_A_1028_413#_c_1271_n N_A_1786_47#_c_1456_n 0.0131369f $X=9.135 $Y=1.025
+ $X2=0 $Y2=0
cc_848 N_A_1028_413#_c_1270_n N_A_1786_47#_c_1457_n 0.0123611f $X=9.06 $Y=1.16
+ $X2=0 $Y2=0
cc_849 N_A_1028_413#_c_1271_n N_A_1786_47#_c_1457_n 0.00118555f $X=9.135
+ $Y=1.025 $X2=0 $Y2=0
cc_850 N_A_1028_413#_c_1272_n N_A_1786_47#_c_1457_n 0.00118555f $X=9.135 $Y=1.62
+ $X2=0 $Y2=0
cc_851 N_A_1028_413#_c_1276_n N_A_1786_47#_c_1457_n 0.00732445f $X=9.135 $Y=1.16
+ $X2=0 $Y2=0
cc_852 N_A_1028_413#_c_1271_n N_A_1786_47#_c_1458_n 0.00248624f $X=9.135
+ $Y=1.025 $X2=0 $Y2=0
cc_853 N_A_1028_413#_c_1273_n N_A_1786_47#_c_1458_n 0.0162698f $X=9.265 $Y=0.73
+ $X2=0 $Y2=0
cc_854 N_A_1028_413#_c_1290_n N_VPWR_M1013_d 0.00216018f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_855 N_A_1028_413#_c_1295_n N_VPWR_c_1511_n 0.00559306f $X=5.59 $Y=2.29 $X2=0
+ $Y2=0
cc_856 N_A_1028_413#_M1026_g N_VPWR_c_1512_n 0.0165029f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_857 N_A_1028_413#_c_1290_n N_VPWR_c_1512_n 0.00850121f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_858 N_A_1028_413#_M1026_g N_VPWR_c_1513_n 0.0046653f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_859 N_A_1028_413#_M1026_g N_VPWR_c_1514_n 0.00576686f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_860 N_A_1028_413#_c_1266_n N_VPWR_c_1514_n 0.00383624f $X=8.25 $Y=1.16 $X2=0
+ $Y2=0
cc_861 N_A_1028_413#_M1019_g N_VPWR_c_1514_n 0.00450985f $X=8.325 $Y=1.985 $X2=0
+ $Y2=0
cc_862 N_A_1028_413#_c_1286_n N_VPWR_c_1515_n 0.00496692f $X=9.265 $Y=1.77 $X2=0
+ $Y2=0
cc_863 N_A_1028_413#_M1019_g N_VPWR_c_1516_n 0.00541359f $X=8.325 $Y=1.985 $X2=0
+ $Y2=0
cc_864 N_A_1028_413#_c_1286_n N_VPWR_c_1516_n 0.00541359f $X=9.265 $Y=1.77 $X2=0
+ $Y2=0
cc_865 N_A_1028_413#_c_1295_n N_VPWR_c_1521_n 0.0210044f $X=5.59 $Y=2.29 $X2=0
+ $Y2=0
cc_866 N_A_1028_413#_c_1290_n N_VPWR_c_1521_n 0.00249003f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_867 N_A_1028_413#_c_1292_n N_VPWR_c_1521_n 0.00729403f $X=5.675 $Y=2 $X2=0
+ $Y2=0
cc_868 N_A_1028_413#_c_1290_n N_VPWR_c_1522_n 0.0036467f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_869 N_A_1028_413#_c_1291_n N_VPWR_c_1522_n 0.0101929f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_870 N_A_1028_413#_M1005_d N_VPWR_c_1507_n 0.0026466f $X=5.14 $Y=2.065 $X2=0
+ $Y2=0
cc_871 N_A_1028_413#_M1001_s N_VPWR_c_1507_n 0.00394021f $X=6.57 $Y=2.065 $X2=0
+ $Y2=0
cc_872 N_A_1028_413#_M1026_g N_VPWR_c_1507_n 0.00934473f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_873 N_A_1028_413#_M1019_g N_VPWR_c_1507_n 0.0121537f $X=8.325 $Y=1.985 $X2=0
+ $Y2=0
cc_874 N_A_1028_413#_c_1286_n N_VPWR_c_1507_n 0.011107f $X=9.265 $Y=1.77 $X2=0
+ $Y2=0
cc_875 N_A_1028_413#_c_1295_n N_VPWR_c_1507_n 0.0105058f $X=5.59 $Y=2.29 $X2=0
+ $Y2=0
cc_876 N_A_1028_413#_c_1290_n N_VPWR_c_1507_n 0.012123f $X=6.54 $Y=2 $X2=0 $Y2=0
cc_877 N_A_1028_413#_c_1291_n N_VPWR_c_1507_n 0.0086238f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_878 N_A_1028_413#_c_1292_n N_VPWR_c_1507_n 0.00588869f $X=5.675 $Y=2 $X2=0
+ $Y2=0
cc_879 N_A_1028_413#_c_1290_n N_VPWR_c_1529_n 0.0263196f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_880 N_A_1028_413#_c_1291_n N_VPWR_c_1529_n 0.00885365f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_881 N_A_1028_413#_c_1292_n N_VPWR_c_1529_n 0.0120166f $X=5.675 $Y=2 $X2=0
+ $Y2=0
cc_882 N_A_1028_413#_c_1290_n A_1136_413# 0.00131812f $X=6.54 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_883 N_A_1028_413#_c_1292_n A_1136_413# 0.00354334f $X=5.675 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_884 N_A_1028_413#_M1007_g N_Q_N_c_1753_n 0.0120523f $X=8.325 $Y=0.56 $X2=0
+ $Y2=0
cc_885 N_A_1028_413#_M1019_g N_Q_N_c_1753_n 0.0178678f $X=8.325 $Y=1.985 $X2=0
+ $Y2=0
cc_886 N_A_1028_413#_c_1270_n N_Q_N_c_1753_n 0.0218272f $X=9.06 $Y=1.16 $X2=0
+ $Y2=0
cc_887 N_A_1028_413#_c_1272_n N_Q_N_c_1753_n 0.00144713f $X=9.135 $Y=1.62 $X2=0
+ $Y2=0
cc_888 N_A_1028_413#_c_1273_n N_Q_N_c_1753_n 0.00106211f $X=9.265 $Y=0.73 $X2=0
+ $Y2=0
cc_889 N_A_1028_413#_c_1286_n N_Q_N_c_1753_n 0.00126529f $X=9.265 $Y=1.77 $X2=0
+ $Y2=0
cc_890 N_A_1028_413#_c_1274_n N_Q_N_c_1753_n 0.00792324f $X=8.325 $Y=1.16 $X2=0
+ $Y2=0
cc_891 N_A_1028_413#_c_1275_n N_Q_N_c_1753_n 8.98323e-19 $X=9.265 $Y=0.805 $X2=0
+ $Y2=0
cc_892 N_A_1028_413#_M1017_g N_VGND_c_1795_n 0.00505556f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_893 N_A_1028_413#_M1017_g N_VGND_c_1796_n 0.00472587f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_894 N_A_1028_413#_c_1266_n N_VGND_c_1796_n 0.00418302f $X=8.25 $Y=1.16 $X2=0
+ $Y2=0
cc_895 N_A_1028_413#_M1007_g N_VGND_c_1796_n 0.00484144f $X=8.325 $Y=0.56 $X2=0
+ $Y2=0
cc_896 N_A_1028_413#_c_1273_n N_VGND_c_1797_n 0.00392236f $X=9.265 $Y=0.73 $X2=0
+ $Y2=0
cc_897 N_A_1028_413#_M1007_g N_VGND_c_1798_n 0.00541359f $X=8.325 $Y=0.56 $X2=0
+ $Y2=0
cc_898 N_A_1028_413#_c_1273_n N_VGND_c_1798_n 0.00541359f $X=9.265 $Y=0.73 $X2=0
+ $Y2=0
cc_899 N_A_1028_413#_c_1275_n N_VGND_c_1798_n 2.96334e-19 $X=9.265 $Y=0.805
+ $X2=0 $Y2=0
cc_900 N_A_1028_413#_M1011_d N_VGND_c_1805_n 0.00218745f $X=5.64 $Y=0.235 $X2=0
+ $Y2=0
cc_901 N_A_1028_413#_M1017_g N_VGND_c_1805_n 0.00991048f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_902 N_A_1028_413#_M1007_g N_VGND_c_1805_n 0.0121537f $X=8.325 $Y=0.56 $X2=0
+ $Y2=0
cc_903 N_A_1028_413#_c_1273_n N_VGND_c_1805_n 0.0111969f $X=9.265 $Y=0.73 $X2=0
+ $Y2=0
cc_904 N_A_1028_413#_c_1303_n N_VGND_c_1805_n 0.0135115f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_905 N_A_1028_413#_c_1303_n N_VGND_c_1810_n 0.0361566f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_906 N_A_1028_413#_M1017_g N_VGND_c_1811_n 0.0188993f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_907 N_A_1028_413#_c_1280_n N_VGND_c_1811_n 2.67651e-19 $X=7.305 $Y=1.26 $X2=0
+ $Y2=0
cc_908 N_A_1028_413#_c_1303_n A_1224_47# 0.00244121f $X=6.32 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_909 N_A_1786_47#_M1031_g N_VPWR_c_1515_n 0.00276849f $X=9.74 $Y=1.985 $X2=0
+ $Y2=0
cc_910 N_A_1786_47#_c_1460_n N_VPWR_c_1515_n 0.0380859f $X=9.055 $Y=2 $X2=0
+ $Y2=0
cc_911 N_A_1786_47#_c_1455_n N_VPWR_c_1515_n 0.00618937f $X=9.655 $Y=1.16 $X2=0
+ $Y2=0
cc_912 N_A_1786_47#_c_1456_n N_VPWR_c_1515_n 0.00173485f $X=9.655 $Y=1.16 $X2=0
+ $Y2=0
cc_913 N_A_1786_47#_c_1460_n N_VPWR_c_1516_n 0.0210382f $X=9.055 $Y=2 $X2=0
+ $Y2=0
cc_914 N_A_1786_47#_M1031_g N_VPWR_c_1523_n 0.00585385f $X=9.74 $Y=1.985 $X2=0
+ $Y2=0
cc_915 N_A_1786_47#_M1002_s N_VPWR_c_1507_n 0.00209319f $X=8.93 $Y=1.845 $X2=0
+ $Y2=0
cc_916 N_A_1786_47#_M1031_g N_VPWR_c_1507_n 0.0121467f $X=9.74 $Y=1.985 $X2=0
+ $Y2=0
cc_917 N_A_1786_47#_c_1460_n N_VPWR_c_1507_n 0.0124268f $X=9.055 $Y=2 $X2=0
+ $Y2=0
cc_918 N_A_1786_47#_c_1454_n N_Q_N_c_1753_n 0.0569423f $X=9.055 $Y=0.51 $X2=0
+ $Y2=0
cc_919 N_A_1786_47#_c_1460_n N_Q_N_c_1753_n 0.0877426f $X=9.055 $Y=2 $X2=0 $Y2=0
cc_920 N_A_1786_47#_c_1457_n N_Q_N_c_1753_n 0.0246108f $X=9.055 $Y=1.16 $X2=0
+ $Y2=0
cc_921 N_A_1786_47#_M1031_g N_Q_c_1778_n 0.00595806f $X=9.74 $Y=1.985 $X2=0
+ $Y2=0
cc_922 N_A_1786_47#_c_1460_n N_Q_c_1778_n 0.00599032f $X=9.055 $Y=2 $X2=0 $Y2=0
cc_923 N_A_1786_47#_c_1455_n N_Q_c_1776_n 0.0266603f $X=9.655 $Y=1.16 $X2=0
+ $Y2=0
cc_924 N_A_1786_47#_c_1458_n N_Q_c_1776_n 0.0189779f $X=9.667 $Y=0.995 $X2=0
+ $Y2=0
cc_925 N_A_1786_47#_c_1454_n N_VGND_c_1797_n 0.019638f $X=9.055 $Y=0.51 $X2=0
+ $Y2=0
cc_926 N_A_1786_47#_c_1455_n N_VGND_c_1797_n 0.00720145f $X=9.655 $Y=1.16 $X2=0
+ $Y2=0
cc_927 N_A_1786_47#_c_1456_n N_VGND_c_1797_n 0.00185111f $X=9.655 $Y=1.16 $X2=0
+ $Y2=0
cc_928 N_A_1786_47#_c_1458_n N_VGND_c_1797_n 0.00281691f $X=9.667 $Y=0.995 $X2=0
+ $Y2=0
cc_929 N_A_1786_47#_c_1454_n N_VGND_c_1798_n 0.0210709f $X=9.055 $Y=0.51 $X2=0
+ $Y2=0
cc_930 N_A_1786_47#_c_1458_n N_VGND_c_1804_n 0.00585385f $X=9.667 $Y=0.995 $X2=0
+ $Y2=0
cc_931 N_A_1786_47#_M1003_s N_VGND_c_1805_n 0.00210122f $X=8.93 $Y=0.235 $X2=0
+ $Y2=0
cc_932 N_A_1786_47#_c_1454_n N_VGND_c_1805_n 0.0124992f $X=9.055 $Y=0.51 $X2=0
+ $Y2=0
cc_933 N_A_1786_47#_c_1458_n N_VGND_c_1805_n 0.0121467f $X=9.667 $Y=0.995 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1507_n N_A_381_47#_M1027_d 0.00325229f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_935 N_VPWR_M1027_s N_A_381_47#_c_1687_n 0.00237137f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_936 N_VPWR_M1027_s N_A_381_47#_c_1694_n 0.00471078f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1509_n N_A_381_47#_c_1694_n 0.00880041f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1520_n N_A_381_47#_c_1694_n 0.0018545f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_939 N_VPWR_c_1507_n N_A_381_47#_c_1694_n 0.00198108f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_940 N_VPWR_M1027_s N_A_381_47#_c_1690_n 0.00187968f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1509_n N_A_381_47#_c_1690_n 0.0114817f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1519_n N_A_381_47#_c_1690_n 3.86777e-19 $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1507_n N_A_381_47#_c_1690_n 7.1462e-19 $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1520_n N_A_381_47#_c_1697_n 0.0115924f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1507_n N_A_381_47#_c_1697_n 0.00307944f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_946 N_VPWR_c_1507_n A_562_413# 0.00355877f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_947 N_VPWR_c_1507_n A_956_413# 0.00259672f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_948 N_VPWR_c_1507_n A_1136_413# 0.00216227f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_949 N_VPWR_c_1507_n N_Q_N_M1019_d 0.00209319f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_950 N_VPWR_c_1514_n N_Q_N_c_1753_n 0.0371113f $X=8.115 $Y=1.66 $X2=0 $Y2=0
cc_951 N_VPWR_c_1516_n N_Q_N_c_1753_n 0.0210382f $X=9.445 $Y=2.72 $X2=0 $Y2=0
cc_952 N_VPWR_c_1507_n N_Q_N_c_1753_n 0.0124268f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_953 N_VPWR_c_1507_n N_Q_M1031_d 0.00387172f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_954 N_VPWR_c_1523_n Q 0.018001f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_955 N_VPWR_c_1507_n Q 0.00993603f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_956 N_VPWR_c_1514_n N_VGND_c_1796_n 0.00705082f $X=8.115 $Y=1.66 $X2=0 $Y2=0
cc_957 N_A_381_47#_c_1687_n N_VGND_M1009_s 0.00105184f $X=1.515 $Y=1.795 $X2=0
+ $Y2=0
cc_958 N_A_381_47#_c_1692_n N_VGND_M1009_s 0.00264874f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_959 N_A_381_47#_c_1688_n N_VGND_M1009_s 0.0019591f $X=1.6 $Y=0.73 $X2=0 $Y2=0
cc_960 N_A_381_47#_c_1692_n N_VGND_c_1792_n 0.00883988f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_961 N_A_381_47#_c_1688_n N_VGND_c_1792_n 0.0114461f $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_962 N_A_381_47#_c_1688_n N_VGND_c_1801_n 4.97798e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_963 N_A_381_47#_c_1692_n N_VGND_c_1802_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_964 N_A_381_47#_c_1696_n N_VGND_c_1802_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_965 N_A_381_47#_M1009_d N_VGND_c_1805_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_966 N_A_381_47#_c_1692_n N_VGND_c_1805_n 0.00232804f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_967 N_A_381_47#_c_1688_n N_VGND_c_1805_n 8.52239e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_968 N_A_381_47#_c_1696_n N_VGND_c_1805_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_969 N_Q_N_c_1753_n N_VGND_c_1796_n 0.0251106f $X=8.535 $Y=0.4 $X2=0 $Y2=0
cc_970 N_Q_N_c_1753_n N_VGND_c_1798_n 0.0210382f $X=8.535 $Y=0.4 $X2=0 $Y2=0
cc_971 N_Q_N_M1007_d N_VGND_c_1805_n 0.00209319f $X=8.4 $Y=0.235 $X2=0 $Y2=0
cc_972 N_Q_N_c_1753_n N_VGND_c_1805_n 0.0124268f $X=8.535 $Y=0.4 $X2=0 $Y2=0
cc_973 Q N_VGND_c_1804_n 0.0179668f $X=9.865 $Y=0.425 $X2=0 $Y2=0
cc_974 N_Q_M1015_d N_VGND_c_1805_n 0.00387172f $X=9.815 $Y=0.235 $X2=0 $Y2=0
cc_975 Q N_VGND_c_1805_n 0.00992828f $X=9.865 $Y=0.425 $X2=0 $Y2=0
cc_976 N_VGND_c_1805_n A_586_47# 0.00231384f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_977 N_VGND_c_1805_n A_796_47# 0.00240916f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_978 N_VGND_c_1805_n A_1056_47# 0.00198596f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_979 N_VGND_c_1805_n A_1224_47# 0.00140476f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_980 N_VGND_c_1805_n A_1296_47# 0.00259801f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24

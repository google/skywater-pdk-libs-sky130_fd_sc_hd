# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__and3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 0.635000 1.020000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 2.125000 1.345000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.145000 0.305000 1.365000 0.790000 ;
        RECT 1.145000 0.790000 1.475000 1.215000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.765000 2.215000 2.465000 ;
        RECT 1.955000 0.255000 2.215000 0.735000 ;
        RECT 2.045000 0.735000 2.215000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.300000 0.085000 ;
        RECT 1.535000  0.085000 1.785000 0.625000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.300000 2.805000 ;
        RECT 0.085000 1.980000 0.700000 2.080000 ;
        RECT 0.085000 2.080000 0.690000 2.635000 ;
        RECT 0.515000 1.710000 0.845000 1.955000 ;
        RECT 0.515000 1.955000 0.700000 1.980000 ;
        RECT 1.515000 2.090000 1.770000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.295000 0.975000 0.465000 ;
      RECT 0.085000 1.190000 0.975000 1.260000 ;
      RECT 0.085000 1.260000 0.980000 1.285000 ;
      RECT 0.085000 1.285000 0.990000 1.300000 ;
      RECT 0.085000 1.300000 0.995000 1.315000 ;
      RECT 0.085000 1.315000 1.005000 1.320000 ;
      RECT 0.085000 1.320000 1.010000 1.330000 ;
      RECT 0.085000 1.330000 1.015000 1.340000 ;
      RECT 0.085000 1.340000 1.025000 1.345000 ;
      RECT 0.085000 1.345000 1.035000 1.355000 ;
      RECT 0.085000 1.355000 1.045000 1.360000 ;
      RECT 0.085000 1.360000 0.345000 1.810000 ;
      RECT 0.710000 1.360000 1.045000 1.365000 ;
      RECT 0.710000 1.365000 1.060000 1.370000 ;
      RECT 0.710000 1.370000 1.075000 1.380000 ;
      RECT 0.710000 1.380000 1.100000 1.385000 ;
      RECT 0.710000 1.385000 1.875000 1.390000 ;
      RECT 0.740000 1.390000 1.875000 1.425000 ;
      RECT 0.775000 1.425000 1.875000 1.450000 ;
      RECT 0.805000 0.465000 0.975000 1.190000 ;
      RECT 0.805000 1.450000 1.875000 1.480000 ;
      RECT 0.825000 1.480000 1.875000 1.510000 ;
      RECT 0.845000 1.510000 1.875000 1.540000 ;
      RECT 0.915000 1.540000 1.875000 1.550000 ;
      RECT 0.940000 1.550000 1.875000 1.560000 ;
      RECT 0.960000 1.560000 1.875000 1.575000 ;
      RECT 0.980000 1.575000 1.875000 1.590000 ;
      RECT 0.985000 1.590000 1.770000 1.600000 ;
      RECT 1.000000 1.600000 1.770000 1.635000 ;
      RECT 1.015000 1.635000 1.770000 1.885000 ;
      RECT 1.645000 0.990000 1.875000 1.385000 ;
  END
END sky130_fd_sc_hd__and3_1

* File: sky130_fd_sc_hd__ebufn_2.pxi.spice
* Created: Tue Sep  1 19:07:13 2020
* 
x_PM_SKY130_FD_SC_HD__EBUFN_2%A N_A_M1009_g N_A_M1006_g A A N_A_c_79_n
+ PM_SKY130_FD_SC_HD__EBUFN_2%A
x_PM_SKY130_FD_SC_HD__EBUFN_2%TE_B N_TE_B_M1008_g N_TE_B_M1010_g N_TE_B_c_113_n
+ N_TE_B_c_114_n N_TE_B_M1001_g N_TE_B_c_115_n N_TE_B_c_116_n N_TE_B_M1011_g
+ N_TE_B_c_117_n TE_B N_TE_B_c_111_n PM_SKY130_FD_SC_HD__EBUFN_2%TE_B
x_PM_SKY130_FD_SC_HD__EBUFN_2%A_214_47# N_A_214_47#_M1008_d N_A_214_47#_M1010_d
+ N_A_214_47#_c_170_n N_A_214_47#_M1005_g N_A_214_47#_c_171_n
+ N_A_214_47#_c_172_n N_A_214_47#_M1007_g N_A_214_47#_c_173_n
+ N_A_214_47#_c_180_n N_A_214_47#_c_174_n N_A_214_47#_c_175_n
+ N_A_214_47#_c_176_n N_A_214_47#_c_182_n N_A_214_47#_c_177_n
+ N_A_214_47#_c_178_n N_A_214_47#_c_179_n PM_SKY130_FD_SC_HD__EBUFN_2%A_214_47#
x_PM_SKY130_FD_SC_HD__EBUFN_2%A_27_47# N_A_27_47#_M1009_s N_A_27_47#_M1006_s
+ N_A_27_47#_M1003_g N_A_27_47#_M1000_g N_A_27_47#_M1004_g N_A_27_47#_M1002_g
+ N_A_27_47#_c_260_n N_A_27_47#_c_261_n N_A_27_47#_c_252_n N_A_27_47#_c_253_n
+ N_A_27_47#_c_254_n N_A_27_47#_c_255_n N_A_27_47#_c_264_n N_A_27_47#_c_256_n
+ N_A_27_47#_c_257_n PM_SKY130_FD_SC_HD__EBUFN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__EBUFN_2%VPWR N_VPWR_M1006_d N_VPWR_M1001_d N_VPWR_c_330_n
+ N_VPWR_c_331_n VPWR N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n
+ N_VPWR_c_329_n N_VPWR_c_336_n N_VPWR_c_337_n PM_SKY130_FD_SC_HD__EBUFN_2%VPWR
x_PM_SKY130_FD_SC_HD__EBUFN_2%A_320_309# N_A_320_309#_M1001_s
+ N_A_320_309#_M1011_s N_A_320_309#_M1002_d N_A_320_309#_c_387_n
+ N_A_320_309#_c_379_n N_A_320_309#_c_380_n N_A_320_309#_c_381_n
+ N_A_320_309#_c_383_n N_A_320_309#_c_406_n
+ PM_SKY130_FD_SC_HD__EBUFN_2%A_320_309#
x_PM_SKY130_FD_SC_HD__EBUFN_2%Z N_Z_M1003_d N_Z_M1000_s N_Z_c_433_n N_Z_c_420_n
+ N_Z_c_421_n N_Z_c_422_n Z Z Z Z Z Z Z Z N_Z_c_419_n
+ PM_SKY130_FD_SC_HD__EBUFN_2%Z
x_PM_SKY130_FD_SC_HD__EBUFN_2%VGND N_VGND_M1009_d N_VGND_M1005_d N_VGND_c_474_n
+ N_VGND_c_475_n VGND N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n PM_SKY130_FD_SC_HD__EBUFN_2%VGND
x_PM_SKY130_FD_SC_HD__EBUFN_2%A_392_47# N_A_392_47#_M1005_s N_A_392_47#_M1007_s
+ N_A_392_47#_M1004_s N_A_392_47#_c_527_n N_A_392_47#_c_532_n
+ N_A_392_47#_c_528_n N_A_392_47#_c_561_n N_A_392_47#_c_529_n
+ PM_SKY130_FD_SC_HD__EBUFN_2%A_392_47#
cc_1 VNB N_A_M1009_g 0.0325187f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.00512854f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_3 VNB N_A_c_79_n 0.0269023f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_4 VNB N_TE_B_M1008_g 0.0379714f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB TE_B 0.00432929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_TE_B_c_111_n 0.0286654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_214_47#_c_170_n 0.0175424f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_8 VNB N_A_214_47#_c_171_n 0.0125703f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_9 VNB N_A_214_47#_c_172_n 0.00844702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_214_47#_c_173_n 0.0124642f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_11 VNB N_A_214_47#_c_174_n 0.0122986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_214_47#_c_175_n 0.00135223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_214_47#_c_176_n 0.0187671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_214_47#_c_177_n 0.0025313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_214_47#_c_178_n 0.0337826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_214_47#_c_179_n 0.015062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_M1003_g 0.0184978f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_18 VNB N_A_27_47#_M1000_g 6.84067e-19 $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.16
cc_19 VNB N_A_27_47#_M1004_g 0.0208147f $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.325
cc_20 VNB N_A_27_47#_M1002_g 4.53022e-19 $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_21 VNB N_A_27_47#_c_252_n 0.0131055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_253_n 0.0135755f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_254_n 0.0113244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_255_n 0.0284854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_256_n 8.30803e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_257_n 0.0322743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_329_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB Z 0.0215341f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_29 VNB N_Z_c_419_n 0.0098129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_474_n 0.00279657f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_31 VNB N_VGND_c_475_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.16
cc_32 VNB N_VGND_c_476_n 0.0151734f $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.325
cc_33 VNB N_VGND_c_477_n 0.0362594f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.53
cc_34 VNB N_VGND_c_478_n 0.0362003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_479_n 0.22969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_480_n 0.00517167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_481_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_392_47#_c_527_n 0.00498807f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_39 VNB N_A_392_47#_c_528_n 0.00265725f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_40 VNB N_A_392_47#_c_529_n 0.00871563f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_41 VPB N_A_M1006_g 0.042548f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_42 VPB A 0.00563944f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_43 VPB N_A_c_79_n 0.00605063f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_44 VPB N_TE_B_M1010_g 0.0357236f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_45 VPB N_TE_B_c_113_n 0.0398485f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_46 VPB N_TE_B_c_114_n 0.0167451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_TE_B_c_115_n 0.0252744f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_48 VPB N_TE_B_c_116_n 0.0172196f $X=-0.19 $Y=1.305 $X2=0.552 $Y2=0.995
cc_49 VPB N_TE_B_c_117_n 0.00612638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_TE_B_c_111_n 0.0137819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_214_47#_c_180_n 0.0106505f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_52 VPB N_A_214_47#_c_175_n 6.99428e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_214_47#_c_182_n 0.0128368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_M1000_g 0.0267161f $X=-0.19 $Y=1.305 $X2=0.552 $Y2=1.16
cc_55 VPB N_A_27_47#_M1002_g 0.0230799f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_56 VPB N_A_27_47#_c_260_n 0.00528662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_261_n 0.0189425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_254_n 0.00161002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_255_n 0.0275234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_264_n 0.00188398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_330_n 0.00364243f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_62 VPB N_VPWR_c_331_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.552 $Y2=1.16
cc_63 VPB N_VPWR_c_332_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0.552 $Y2=1.325
cc_64 VPB N_VPWR_c_333_n 0.0251591f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.53
cc_65 VPB N_VPWR_c_334_n 0.0434782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_329_n 0.0529156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_336_n 0.00585573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_337_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_320_309#_c_379_n 0.00130839f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_70 VPB N_A_320_309#_c_380_n 0.00759475f $X=-0.19 $Y=1.305 $X2=0.552 $Y2=0.995
cc_71 VPB N_A_320_309#_c_381_n 0.0194249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_Z_c_420_n 0.00110732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_Z_c_421_n 0.00568641f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_74 VPB N_Z_c_422_n 0.0017893f $X=-0.19 $Y=1.305 $X2=0.552 $Y2=0.995
cc_75 VPB Z 0.00693953f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_76 VPB Z 0.0082414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 N_A_M1009_g N_TE_B_M1008_g 0.0210944f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_78 A N_TE_B_M1008_g 0.00773576f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_c_79_n N_TE_B_M1008_g 0.0212945f $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_M1009_g TE_B 2.00312e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_81 A TE_B 0.038411f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A_c_79_n TE_B 3.65211e-19 $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_TE_B_c_111_n 0.0188416f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_84 A N_A_214_47#_c_175_n 0.00474768f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_85 A N_A_214_47#_c_182_n 0.0121505f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_86 A N_A_27_47#_c_253_n 0.0194626f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_87 N_A_c_79_n N_A_27_47#_c_253_n 0.00964443f $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_88 A N_A_27_47#_c_254_n 0.00274795f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_c_79_n N_A_27_47#_c_254_n 0.00262964f $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_M1009_g N_A_27_47#_c_255_n 0.032091f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_91 A N_A_27_47#_c_255_n 0.0671931f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_VPWR_c_330_n 0.0132729f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_93 A N_VPWR_c_330_n 0.0208956f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_94 N_A_c_79_n N_VPWR_c_330_n 5.35719e-19 $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_M1006_g N_VPWR_c_332_n 0.0046653f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_96 N_A_M1006_g N_VPWR_c_329_n 0.00895857f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_97 N_A_M1009_g N_VGND_c_474_n 0.0112241f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_98 A N_VGND_c_474_n 0.0200531f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_99 N_A_c_79_n N_VGND_c_474_n 6.62542e-19 $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_M1009_g N_VGND_c_476_n 0.0046653f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_M1009_g N_VGND_c_479_n 0.00818925f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_102 A N_VGND_c_479_n 0.00190664f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_103 N_TE_B_c_115_n N_A_214_47#_c_171_n 2.6249e-19 $X=2.28 $Y=1.395 $X2=0
+ $Y2=0
cc_104 N_TE_B_c_115_n N_A_214_47#_c_172_n 0.0133877f $X=2.28 $Y=1.395 $X2=0
+ $Y2=0
cc_105 N_TE_B_M1008_g N_A_214_47#_c_173_n 0.00516105f $X=0.995 $Y=0.445 $X2=0
+ $Y2=0
cc_106 TE_B N_A_214_47#_c_173_n 0.0181259f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_107 N_TE_B_c_111_n N_A_214_47#_c_173_n 7.72975e-19 $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_TE_B_M1010_g N_A_214_47#_c_180_n 0.00773658f $X=0.995 $Y=2.165 $X2=0
+ $Y2=0
cc_109 N_TE_B_c_114_n N_A_214_47#_c_180_n 0.0059364f $X=1.935 $Y=1.47 $X2=0
+ $Y2=0
cc_110 N_TE_B_c_111_n N_A_214_47#_c_180_n 8.62733e-19 $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_TE_B_M1008_g N_A_214_47#_c_174_n 0.00550308f $X=0.995 $Y=0.445 $X2=0
+ $Y2=0
cc_112 TE_B N_A_214_47#_c_174_n 0.021343f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_113 N_TE_B_c_113_n N_A_214_47#_c_175_n 0.0201809f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_114 N_TE_B_c_111_n N_A_214_47#_c_175_n 0.00128122f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_TE_B_c_113_n N_A_214_47#_c_176_n 0.0165609f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_116 N_TE_B_M1010_g N_A_214_47#_c_182_n 0.0094476f $X=0.995 $Y=2.165 $X2=0
+ $Y2=0
cc_117 N_TE_B_c_113_n N_A_214_47#_c_182_n 0.0138273f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_118 N_TE_B_c_114_n N_A_214_47#_c_182_n 0.00614532f $X=1.935 $Y=1.47 $X2=0
+ $Y2=0
cc_119 TE_B N_A_214_47#_c_182_n 0.0112925f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_120 N_TE_B_c_111_n N_A_214_47#_c_182_n 0.00524648f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_121 TE_B N_A_214_47#_c_177_n 0.0190634f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_122 N_TE_B_c_111_n N_A_214_47#_c_177_n 0.00499695f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_123 N_TE_B_c_113_n N_A_27_47#_c_253_n 0.00385524f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_124 TE_B N_A_27_47#_c_253_n 0.0244937f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_125 N_TE_B_c_111_n N_A_27_47#_c_253_n 0.00469111f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_126 N_TE_B_M1010_g N_VPWR_c_330_n 0.013653f $X=0.995 $Y=2.165 $X2=0 $Y2=0
cc_127 N_TE_B_c_114_n N_VPWR_c_331_n 0.00812695f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_128 N_TE_B_c_116_n N_VPWR_c_331_n 0.00815483f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_129 N_TE_B_M1010_g N_VPWR_c_333_n 0.0046653f $X=0.995 $Y=2.165 $X2=0 $Y2=0
cc_130 N_TE_B_c_114_n N_VPWR_c_333_n 0.00337001f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_131 N_TE_B_c_116_n N_VPWR_c_334_n 0.00337001f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_132 N_TE_B_M1010_g N_VPWR_c_329_n 0.00934473f $X=0.995 $Y=2.165 $X2=0 $Y2=0
cc_133 N_TE_B_c_114_n N_VPWR_c_329_n 0.00523175f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_134 N_TE_B_c_116_n N_VPWR_c_329_n 0.00523175f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_135 N_TE_B_c_113_n N_A_320_309#_c_379_n 0.00118255f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_136 N_TE_B_c_114_n N_A_320_309#_c_383_n 0.0132889f $X=1.935 $Y=1.47 $X2=0
+ $Y2=0
cc_137 N_TE_B_c_115_n N_A_320_309#_c_383_n 3.36696e-19 $X=2.28 $Y=1.395 $X2=0
+ $Y2=0
cc_138 N_TE_B_c_116_n N_A_320_309#_c_383_n 0.0133852f $X=2.355 $Y=1.47 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_114_n N_Z_c_421_n 0.00956756f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_140 N_TE_B_c_115_n N_Z_c_421_n 0.00662881f $X=2.28 $Y=1.395 $X2=0 $Y2=0
cc_141 N_TE_B_c_116_n N_Z_c_421_n 0.0166982f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_142 N_TE_B_c_117_n N_Z_c_421_n 0.00144299f $X=1.935 $Y=1.395 $X2=0 $Y2=0
cc_143 N_TE_B_M1008_g N_VGND_c_474_n 0.00630084f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_144 N_TE_B_M1008_g N_VGND_c_477_n 0.00509549f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_145 N_TE_B_M1008_g N_VGND_c_479_n 0.00841714f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_146 TE_B N_VGND_c_479_n 0.0027627f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_147 N_A_214_47#_c_178_n N_A_27_47#_M1003_g 0.0231998f $X=2.8 $Y=1.035 $X2=0
+ $Y2=0
cc_148 N_A_214_47#_c_179_n N_A_27_47#_M1003_g 0.0147131f $X=2.8 $Y=0.96 $X2=0
+ $Y2=0
cc_149 N_A_214_47#_c_173_n N_A_27_47#_c_253_n 0.00692194f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_150 N_A_214_47#_c_176_n N_A_27_47#_c_253_n 0.056439f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_214_47#_c_182_n N_A_27_47#_c_253_n 0.00995529f $X=1.592 $Y=1.605
+ $X2=0 $Y2=0
cc_152 N_A_214_47#_c_177_n N_A_27_47#_c_253_n 0.0243818f $X=1.592 $Y=1.15 $X2=0
+ $Y2=0
cc_153 N_A_214_47#_c_178_n N_A_27_47#_c_253_n 6.94548e-19 $X=2.8 $Y=1.035 $X2=0
+ $Y2=0
cc_154 N_A_214_47#_c_176_n N_A_27_47#_c_264_n 3.80502e-19 $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_214_47#_c_176_n N_A_27_47#_c_256_n 0.0106399f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_214_47#_c_178_n N_A_27_47#_c_256_n 3.94165e-19 $X=2.8 $Y=1.035 $X2=0
+ $Y2=0
cc_157 N_A_214_47#_c_176_n N_A_27_47#_c_257_n 0.00100223f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_214_47#_c_180_n N_VPWR_c_333_n 0.0201949f $X=1.205 $Y=2.22 $X2=0
+ $Y2=0
cc_159 N_A_214_47#_M1010_d N_VPWR_c_329_n 0.00387172f $X=1.07 $Y=1.845 $X2=0
+ $Y2=0
cc_160 N_A_214_47#_c_180_n N_VPWR_c_329_n 0.0110999f $X=1.205 $Y=2.22 $X2=0
+ $Y2=0
cc_161 N_A_214_47#_c_182_n N_A_320_309#_M1001_s 0.00410412f $X=1.592 $Y=1.605
+ $X2=-0.19 $Y2=-0.24
cc_162 N_A_214_47#_c_180_n N_A_320_309#_c_387_n 0.0259828f $X=1.205 $Y=2.22
+ $X2=0 $Y2=0
cc_163 N_A_214_47#_c_180_n N_A_320_309#_c_379_n 0.0134641f $X=1.205 $Y=2.22
+ $X2=0 $Y2=0
cc_164 N_A_214_47#_c_176_n N_A_320_309#_c_379_n 0.00217928f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_214_47#_c_182_n N_A_320_309#_c_379_n 0.011254f $X=1.592 $Y=1.605
+ $X2=0 $Y2=0
cc_166 N_A_214_47#_c_176_n N_A_320_309#_c_383_n 0.00193213f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_214_47#_c_171_n N_Z_c_421_n 0.00101771f $X=2.635 $Y=1.035 $X2=0 $Y2=0
cc_168 N_A_214_47#_c_176_n N_Z_c_421_n 0.0750347f $X=2.8 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_214_47#_c_182_n N_Z_c_421_n 0.0276028f $X=1.592 $Y=1.605 $X2=0 $Y2=0
cc_170 N_A_214_47#_c_178_n N_Z_c_421_n 0.00832899f $X=2.8 $Y=1.035 $X2=0 $Y2=0
cc_171 N_A_214_47#_c_173_n N_VGND_c_474_n 0.0279767f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_172 N_A_214_47#_c_170_n N_VGND_c_475_n 0.00856801f $X=2.295 $Y=0.96 $X2=0
+ $Y2=0
cc_173 N_A_214_47#_c_179_n N_VGND_c_475_n 0.00829743f $X=2.8 $Y=0.96 $X2=0 $Y2=0
cc_174 N_A_214_47#_c_170_n N_VGND_c_477_n 0.00341689f $X=2.295 $Y=0.96 $X2=0
+ $Y2=0
cc_175 N_A_214_47#_c_173_n N_VGND_c_477_n 0.0468578f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_176 N_A_214_47#_c_179_n N_VGND_c_478_n 0.00341689f $X=2.8 $Y=0.96 $X2=0 $Y2=0
cc_177 N_A_214_47#_M1008_d N_VGND_c_479_n 0.00210147f $X=1.07 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_214_47#_c_170_n N_VGND_c_479_n 0.00540327f $X=2.295 $Y=0.96 $X2=0
+ $Y2=0
cc_179 N_A_214_47#_c_173_n N_VGND_c_479_n 0.0268076f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_180 N_A_214_47#_c_179_n N_VGND_c_479_n 0.004321f $X=2.8 $Y=0.96 $X2=0 $Y2=0
cc_181 N_A_214_47#_c_173_n N_A_392_47#_c_527_n 0.029754f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_182 N_A_214_47#_c_174_n N_A_392_47#_c_527_n 0.00477906f $X=1.59 $Y=1.025
+ $X2=0 $Y2=0
cc_183 N_A_214_47#_c_170_n N_A_392_47#_c_532_n 0.0121972f $X=2.295 $Y=0.96 $X2=0
+ $Y2=0
cc_184 N_A_214_47#_c_171_n N_A_392_47#_c_532_n 0.00186586f $X=2.635 $Y=1.035
+ $X2=0 $Y2=0
cc_185 N_A_214_47#_c_176_n N_A_392_47#_c_532_n 0.046904f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_186 N_A_214_47#_c_178_n N_A_392_47#_c_532_n 0.0031161f $X=2.8 $Y=1.035 $X2=0
+ $Y2=0
cc_187 N_A_214_47#_c_179_n N_A_392_47#_c_532_n 0.0115842f $X=2.8 $Y=0.96 $X2=0
+ $Y2=0
cc_188 N_A_214_47#_c_174_n N_A_392_47#_c_528_n 0.0174868f $X=1.59 $Y=1.025 $X2=0
+ $Y2=0
cc_189 N_A_214_47#_c_176_n N_A_392_47#_c_528_n 0.02076f $X=2.8 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_253_n N_VPWR_c_330_n 0.00680952f $X=3.32 $Y=1.19 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_261_n N_VPWR_c_332_n 0.0179925f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_192 N_A_27_47#_M1000_g N_VPWR_c_334_n 0.00357877f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1002_g N_VPWR_c_334_n 0.00357877f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1006_s N_VPWR_c_329_n 0.00387172f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1000_g N_VPWR_c_329_n 0.00664112f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1002_g N_VPWR_c_329_n 0.00617937f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_261_n N_VPWR_c_329_n 0.0099338f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_198 N_A_27_47#_M1000_g N_A_320_309#_c_380_n 0.0130654f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_M1002_g N_A_320_309#_c_380_n 0.00941684f $X=3.67 $Y=1.985
+ $X2=0 $Y2=0
cc_200 N_A_27_47#_M1003_g N_Z_c_433_n 0.00304334f $X=3.25 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_27_47#_M1004_g N_Z_c_433_n 0.0127197f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_264_n N_Z_c_433_n 0.00194826f $X=3.465 $Y=1.19 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_256_n N_Z_c_433_n 0.0207501f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_257_n N_Z_c_433_n 6.48684e-19 $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_27_47#_M1002_g N_Z_c_420_n 0.0118398f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_256_n N_Z_c_420_n 0.00201091f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_27_47#_M1000_g N_Z_c_421_n 0.0162143f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_253_n N_Z_c_421_n 0.0187092f $X=3.32 $Y=1.19 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_256_n N_Z_c_421_n 0.00324626f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1000_g N_Z_c_422_n 0.00173244f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_27_47#_M1002_g N_Z_c_422_n 0.00800327f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_264_n N_Z_c_422_n 0.00843249f $X=3.465 $Y=1.19 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_256_n N_Z_c_422_n 0.0233644f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_257_n N_Z_c_422_n 0.00163105f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_27_47#_M1000_g Z 0.00990987f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_27_47#_M1002_g Z 0.00529685f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1004_g Z 0.0203863f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_264_n Z 0.00264045f $X=3.465 $Y=1.19 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_256_n Z 0.0181927f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_253_n N_VGND_c_474_n 0.00373214f $X=3.32 $Y=1.19 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1003_g N_VGND_c_475_n 0.0011614f $X=3.25 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_252_n N_VGND_c_476_n 0.0154629f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A_27_47#_M1003_g N_VGND_c_478_n 0.00362032f $X=3.25 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1004_g N_VGND_c_478_n 0.00362032f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1009_s N_VGND_c_479_n 0.00388065f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_M1003_g N_VGND_c_479_n 0.00556431f $X=3.25 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1004_g N_VGND_c_479_n 0.00618478f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_252_n N_VGND_c_479_n 0.00979848f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_253_n N_A_392_47#_c_532_n 0.00958353f $X=3.32 $Y=1.19 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_253_n N_A_392_47#_c_528_n 0.00183114f $X=3.32 $Y=1.19 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1003_g N_A_392_47#_c_529_n 0.0122643f $X=3.25 $Y=0.56 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1004_g N_A_392_47#_c_529_n 0.00828053f $X=3.67 $Y=0.56 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_256_n N_A_392_47#_c_529_n 0.00129798f $X=3.46 $Y=1.16 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_329_n N_A_320_309#_M1001_s 0.00224186f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_235 N_VPWR_c_329_n N_A_320_309#_M1011_s 0.00620436f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_329_n N_A_320_309#_M1002_d 0.00209324f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_333_n N_A_320_309#_c_387_n 0.0141623f $X=1.98 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_329_n N_A_320_309#_c_387_n 0.00795901f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_334_n N_A_320_309#_c_380_n 0.0180525f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_329_n N_A_320_309#_c_380_n 0.010004f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_241 N_VPWR_M1001_d N_A_320_309#_c_383_n 0.00313513f $X=2.01 $Y=1.545 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_331_n N_A_320_309#_c_383_n 0.0158599f $X=2.145 $Y=2.36 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_333_n N_A_320_309#_c_383_n 0.00256355f $X=1.98 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_334_n N_A_320_309#_c_383_n 0.00256355f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_329_n N_A_320_309#_c_383_n 0.0100471f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_334_n N_A_320_309#_c_406_n 0.0796448f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_329_n N_A_320_309#_c_406_n 0.0481784f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_329_n N_Z_M1000_s 0.00216833f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_M1001_d N_Z_c_421_n 0.00169505f $X=2.01 $Y=1.545 $X2=0 $Y2=0
cc_250 N_A_320_309#_c_380_n N_Z_M1000_s 0.00312348f $X=3.795 $Y=2.38 $X2=0 $Y2=0
cc_251 N_A_320_309#_M1002_d N_Z_c_420_n 2.34277e-19 $X=3.745 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_320_309#_c_380_n N_Z_c_420_n 0.00257436f $X=3.795 $Y=2.38 $X2=0 $Y2=0
cc_253 N_A_320_309#_c_381_n N_Z_c_420_n 0.00183942f $X=3.88 $Y=1.96 $X2=0 $Y2=0
cc_254 N_A_320_309#_M1011_s N_Z_c_421_n 0.0128017f $X=2.43 $Y=1.545 $X2=0 $Y2=0
cc_255 N_A_320_309#_c_380_n N_Z_c_421_n 0.0033549f $X=3.795 $Y=2.38 $X2=0 $Y2=0
cc_256 N_A_320_309#_c_383_n N_Z_c_421_n 0.0824067f $X=2.48 $Y=2.2 $X2=0 $Y2=0
cc_257 N_A_320_309#_c_380_n Z 0.015949f $X=3.795 $Y=2.38 $X2=0 $Y2=0
cc_258 N_A_320_309#_M1002_d Z 0.00261185f $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_259 N_A_320_309#_c_381_n Z 0.0207974f $X=3.88 $Y=1.96 $X2=0 $Y2=0
cc_260 N_Z_M1003_d N_VGND_c_479_n 0.00217706f $X=3.325 $Y=0.235 $X2=0 $Y2=0
cc_261 N_Z_c_419_n N_VGND_c_479_n 7.23694e-19 $X=3.94 $Y=0.855 $X2=0 $Y2=0
cc_262 N_Z_c_433_n N_A_392_47#_M1004_s 6.34565e-19 $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_263 Z N_A_392_47#_M1004_s 4.61372e-19 $X=3.84 $Y=0.765 $X2=0 $Y2=0
cc_264 N_Z_c_419_n N_A_392_47#_M1004_s 0.00289486f $X=3.94 $Y=0.855 $X2=0 $Y2=0
cc_265 N_Z_c_421_n N_A_392_47#_c_532_n 0.00220399f $X=3.295 $Y=1.605 $X2=0 $Y2=0
cc_266 N_Z_M1003_d N_A_392_47#_c_529_n 0.00309251f $X=3.325 $Y=0.235 $X2=0 $Y2=0
cc_267 N_Z_c_433_n N_A_392_47#_c_529_n 0.0241481f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_268 N_Z_c_419_n N_A_392_47#_c_529_n 0.0175569f $X=3.94 $Y=0.855 $X2=0 $Y2=0
cc_269 N_VGND_c_479_n N_A_392_47#_M1005_s 0.00229009f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_270 N_VGND_c_479_n N_A_392_47#_M1007_s 0.00329894f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_271 N_VGND_c_479_n N_A_392_47#_M1004_s 0.00210181f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_477_n N_A_392_47#_c_527_n 0.0185481f $X=2.34 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_c_479_n N_A_392_47#_c_527_n 0.0102875f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_M1005_d N_A_392_47#_c_532_n 0.00293186f $X=2.37 $Y=0.235 $X2=0
+ $Y2=0
cc_275 N_VGND_c_475_n N_A_392_47#_c_532_n 0.0162338f $X=2.505 $Y=0.36 $X2=0
+ $Y2=0
cc_276 N_VGND_c_477_n N_A_392_47#_c_532_n 0.00234306f $X=2.34 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_478_n N_A_392_47#_c_532_n 0.00234306f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_479_n N_A_392_47#_c_532_n 0.00978207f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_478_n N_A_392_47#_c_561_n 0.0171369f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_479_n N_A_392_47#_c_561_n 0.0108223f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_478_n N_A_392_47#_c_529_n 0.0463624f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_479_n N_A_392_47#_c_529_n 0.0326703f $X=3.91 $Y=0 $X2=0 $Y2=0

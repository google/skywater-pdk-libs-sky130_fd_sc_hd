* NGSPICE file created from sky130_fd_sc_hd__a31oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=2.1125e+11p ps=1.95e+06u
M1001 Y B1 a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=5.95e+11p ps=5.19e+06u
M1002 VPWR A2 a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.65e+11p pd=5.13e+06u as=0p ps=0u
M1003 a_181_47# A2 a_109_47# VNB nshort w=650000u l=150000u
+  ad=2.3725e+11p pd=2.03e+06u as=1.365e+11p ps=1.72e+06u
M1004 Y A1 a_181_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_109_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_109_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_109_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


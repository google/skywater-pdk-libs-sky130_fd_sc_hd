* NGSPICE file created from sky130_fd_sc_hd__a2111oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=9.1325e+11p pd=6.71e+06u as=6.3375e+11p ps=4.55e+06u
M1001 a_316_297# C1 a_217_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.7e+11p pd=2.74e+06u as=3.45e+11p ps=2.69e+06u
M1002 a_568_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1003 Y D1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_420_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=8.7e+11p pd=5.74e+06u as=2.75e+11p ps=2.55e+06u
M1006 a_217_297# D1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=7.55e+11p ps=3.51e+06u
M1007 VPWR A1 a_420_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_420_297# B1 a_316_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_568_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


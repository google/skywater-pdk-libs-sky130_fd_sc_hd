* File: sky130_fd_sc_hd__clkdlybuf4s50_1.spice.SKY130_FD_SC_HD__CLKDLYBUF4S50_1.pxi
* Created: Thu Aug 27 14:12:01 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A N_A_M1002_g N_A_M1003_g A N_A_c_60_n
+ N_A_c_61_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_27_47# N_A_27_47#_M1002_s
+ N_A_27_47#_M1003_s N_A_27_47#_M1001_g N_A_27_47#_M1005_g N_A_27_47#_c_90_n
+ N_A_27_47#_c_96_n N_A_27_47#_c_91_n N_A_27_47#_c_92_n N_A_27_47#_c_97_n
+ N_A_27_47#_c_98_n N_A_27_47#_c_93_n N_A_27_47#_c_94_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_283_47# N_A_283_47#_M1001_d
+ N_A_283_47#_M1005_d N_A_283_47#_M1006_g N_A_283_47#_M1004_g
+ N_A_283_47#_c_159_n N_A_283_47#_c_160_n N_A_283_47#_c_161_n
+ N_A_283_47#_c_165_n N_A_283_47#_c_162_n N_A_283_47#_c_163_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_283_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_390_47# N_A_390_47#_M1006_s
+ N_A_390_47#_M1004_s N_A_390_47#_M1000_g N_A_390_47#_M1007_g
+ N_A_390_47#_c_220_n N_A_390_47#_c_216_n N_A_390_47#_c_212_n
+ N_A_390_47#_c_236_n N_A_390_47#_c_213_n N_A_390_47#_c_214_n
+ N_A_390_47#_c_219_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_390_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%VPWR N_VPWR_M1003_d N_VPWR_M1004_d
+ N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n VPWR
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_269_n N_VPWR_c_277_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%X N_X_M1000_d N_X_M1007_d X X X X X X
+ N_X_c_312_n X PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%VGND N_VGND_M1002_d N_VGND_M1006_d
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n VGND
+ N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%VGND
cc_1 VNB N_A_M1002_g 0.0386267f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.445
cc_2 VNB N_A_c_60_n 0.0308097f $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.16
cc_3 VNB N_A_c_61_n 0.0104592f $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.16
cc_4 VNB N_A_27_47#_M1001_g 0.0440303f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_M1005_g 8.8112e-19 $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.16
cc_6 VNB N_A_27_47#_c_90_n 0.0193392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_91_n 0.00311413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_92_n 0.0100727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_93_n 0.00273063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_94_n 0.0323829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_283_47#_M1006_g 0.0444279f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_A_283_47#_M1004_g 8.32628e-19 $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.16
cc_13 VNB N_A_283_47#_c_159_n 0.032249f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.31
cc_14 VNB N_A_283_47#_c_160_n 0.0172639f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.182
cc_15 VNB N_A_283_47#_c_161_n 0.0101161f $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.182
cc_16 VNB N_A_283_47#_c_162_n 0.00644785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_283_47#_c_163_n 0.0011734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_390_47#_M1000_g 0.0343963f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_19 VNB N_A_390_47#_c_212_n 0.00149056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_390_47#_c_213_n 0.00294554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_390_47#_c_214_n 0.0232901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_269_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB X 0.0348518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_312_n 0.0157672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_325_n 0.00557099f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB N_VGND_c_326_n 0.00283171f $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.16
cc_27 VNB N_VGND_c_327_n 0.0477363f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.182
cc_28 VNB N_VGND_c_328_n 0.00510866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_329_n 0.0169264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_330_n 0.0193417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_331_n 0.209423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_332_n 0.00631673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A_M1003_g 0.0278439f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_34 VPB N_A_c_60_n 0.00527711f $X=-0.19 $Y=1.305 $X2=0.37 $Y2=1.16
cc_35 VPB N_A_27_47#_M1005_g 0.0657215f $X=-0.19 $Y=1.305 $X2=0.37 $Y2=1.16
cc_36 VPB N_A_27_47#_c_96_n 0.0331199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_c_97_n 0.00200795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_98_n 0.009619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_93_n 0.00213103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_283_47#_M1004_g 0.0674932f $X=-0.19 $Y=1.305 $X2=0.37 $Y2=1.16
cc_41 VPB N_A_283_47#_c_165_n 0.013976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_283_47#_c_162_n 0.0114214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_390_47#_M1007_g 0.0229339f $X=-0.19 $Y=1.305 $X2=0.37 $Y2=1.16
cc_44 VPB N_A_390_47#_c_216_n 3.5835e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_390_47#_c_213_n 0.00333787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_390_47#_c_214_n 0.00527602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_390_47#_c_219_n 0.00360956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_270_n 0.00284395f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_49 VPB N_VPWR_c_271_n 0.00283171f $X=-0.19 $Y=1.305 $X2=0.37 $Y2=1.16
cc_50 VPB N_VPWR_c_272_n 0.0479842f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.182
cc_51 VPB N_VPWR_c_273_n 0.00510842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_274_n 0.0178855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_275_n 0.0193417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_269_n 0.0535145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_277_n 0.00516427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB X 0.0177313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB X 0.0313376f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_58 N_A_M1002_g N_A_27_47#_M1001_g 0.0185951f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_59 N_A_c_60_n N_A_27_47#_M1005_g 0.0294785f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_A_27_47#_c_90_n 0.00815405f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_A_27_47#_c_96_n 0.013155f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_A_27_47#_c_91_n 0.0102842f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_63 N_A_c_61_n N_A_27_47#_c_91_n 0.00824931f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_A_27_47#_c_92_n 0.00376316f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_65 N_A_c_60_n N_A_27_47#_c_92_n 0.00488555f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_61_n N_A_27_47#_c_92_n 0.0273569f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_A_27_47#_c_97_n 0.0117678f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_c_61_n N_A_27_47#_c_97_n 0.00721391f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_A_27_47#_c_98_n 0.00423547f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A_c_60_n N_A_27_47#_c_98_n 0.00466819f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_61_n N_A_27_47#_c_98_n 0.0286225f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_A_27_47#_c_93_n 0.00764772f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A_c_61_n N_A_27_47#_c_93_n 0.0177763f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_c_60_n N_A_27_47#_c_94_n 0.0135475f $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_c_61_n N_A_27_47#_c_94_n 2.14536e-19 $X=0.37 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_VPWR_c_270_n 0.00669214f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_VPWR_c_274_n 0.0054895f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1003_g N_VPWR_c_269_n 0.0109548f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_VGND_c_325_n 0.00315263f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_M1002_g N_VGND_c_329_n 0.00435288f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A_M1002_g N_VGND_c_331_n 0.00710212f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_94_n N_A_283_47#_c_159_n 0.00537157f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_83 N_A_27_47#_M1001_g N_A_283_47#_c_161_n 0.0308531f $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_84 N_A_27_47#_c_93_n N_A_283_47#_c_161_n 0.0161564f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_85 N_A_27_47#_c_94_n N_A_283_47#_c_161_n 0.00154027f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_86 N_A_27_47#_M1005_g N_A_283_47#_c_165_n 0.042907f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_87 N_A_27_47#_c_93_n N_A_283_47#_c_165_n 0.0145167f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_88 N_A_27_47#_M1005_g N_A_283_47#_c_163_n 0.00111405f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_89 N_A_27_47#_c_93_n N_A_283_47#_c_163_n 0.0150997f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_c_94_n N_A_283_47#_c_163_n 0.00872239f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_M1001_g N_A_390_47#_c_220_n 0.00100752f $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_M1005_g N_A_390_47#_c_216_n 0.00157375f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_M1001_g N_A_390_47#_c_212_n 6.91146e-19 $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_M1005_g N_A_390_47#_c_219_n 6.83015e-19 $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_97_n N_VPWR_M1003_d 9.77978e-19 $X=0.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_27_47#_c_93_n N_VPWR_M1003_d 0.00110662f $X=0.97 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_27_47#_M1005_g N_VPWR_c_270_n 0.0228238f $X=1.165 $Y=2.075 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_97_n N_VPWR_c_270_n 0.00752987f $X=0.705 $Y=1.545 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_93_n N_VPWR_c_270_n 0.0177016f $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_94_n N_VPWR_c_270_n 3.36728e-19 $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_27_47#_M1005_g N_VPWR_c_272_n 0.0183935f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_96_n N_VPWR_c_274_n 0.0221174f $X=0.265 $Y=1.965 $X2=0 $Y2=0
cc_103 N_A_27_47#_M1003_s N_VPWR_c_269_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_M1005_g N_VPWR_c_269_n 0.0304754f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_96_n N_VPWR_c_269_n 0.0130273f $X=0.265 $Y=1.965 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_91_n N_VGND_M1002_d 4.05015e-19 $X=0.705 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_27_47#_c_93_n N_VGND_M1002_d 0.001654f $X=0.97 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_27_47#_M1001_g N_VGND_c_325_n 0.00345654f $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_91_n N_VGND_c_325_n 0.00824264f $X=0.705 $Y=0.82 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_93_n N_VGND_c_325_n 0.013265f $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_94_n N_VGND_c_325_n 3.60019e-19 $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_27_47#_M1001_g N_VGND_c_327_n 0.017623f $X=1.165 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_93_n N_VGND_c_327_n 0.00201552f $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_90_n N_VGND_c_329_n 0.0210314f $X=0.265 $Y=0.435 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_91_n N_VGND_c_329_n 0.0022703f $X=0.705 $Y=0.82 $X2=0 $Y2=0
cc_116 N_A_27_47#_M1002_s N_VGND_c_331_n 0.00217517f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_M1001_g N_VGND_c_331_n 0.0280953f $X=1.165 $Y=0.56 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_90_n N_VGND_c_331_n 0.0125034f $X=0.265 $Y=0.435 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_91_n N_VGND_c_331_n 0.00415859f $X=0.705 $Y=0.82 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_93_n N_VGND_c_331_n 0.00408646f $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_283_47#_M1006_g N_A_390_47#_M1000_g 0.0204037f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_122 N_A_283_47#_M1004_g N_A_390_47#_M1007_g 0.0232662f $X=2.465 $Y=2.075
+ $X2=0 $Y2=0
cc_123 N_A_283_47#_M1006_g N_A_390_47#_c_220_n 0.0169044f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_124 N_A_283_47#_c_161_n N_A_390_47#_c_220_n 0.0281823f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_125 N_A_283_47#_M1004_g N_A_390_47#_c_216_n 0.0262639f $X=2.465 $Y=2.075
+ $X2=0 $Y2=0
cc_126 N_A_283_47#_c_165_n N_A_390_47#_c_216_n 0.0475123f $X=1.555 $Y=1.965
+ $X2=0 $Y2=0
cc_127 N_A_283_47#_M1006_g N_A_390_47#_c_212_n 0.0341515f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_128 N_A_283_47#_M1004_g N_A_390_47#_c_212_n 0.00107104f $X=2.465 $Y=2.075
+ $X2=0 $Y2=0
cc_129 N_A_283_47#_c_159_n N_A_390_47#_c_212_n 0.00528171f $X=2.215 $Y=1.16
+ $X2=0 $Y2=0
cc_130 N_A_283_47#_c_160_n N_A_390_47#_c_212_n 0.00980465f $X=2.465 $Y=1.16
+ $X2=0 $Y2=0
cc_131 N_A_283_47#_c_161_n N_A_390_47#_c_212_n 0.0108095f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_132 N_A_283_47#_c_162_n N_A_390_47#_c_212_n 0.0413587f $X=2.075 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_283_47#_M1004_g N_A_390_47#_c_236_n 0.0124362f $X=2.465 $Y=2.075
+ $X2=0 $Y2=0
cc_134 N_A_283_47#_M1006_g N_A_390_47#_c_213_n 0.00641624f $X=2.465 $Y=0.56
+ $X2=0 $Y2=0
cc_135 N_A_283_47#_M1004_g N_A_390_47#_c_213_n 0.00649821f $X=2.465 $Y=2.075
+ $X2=0 $Y2=0
cc_136 N_A_283_47#_c_160_n N_A_390_47#_c_213_n 0.00605761f $X=2.465 $Y=1.16
+ $X2=0 $Y2=0
cc_137 N_A_283_47#_M1006_g N_A_390_47#_c_214_n 0.0196666f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_138 N_A_283_47#_M1004_g N_A_390_47#_c_219_n 0.0324943f $X=2.465 $Y=2.075
+ $X2=0 $Y2=0
cc_139 N_A_283_47#_c_159_n N_A_390_47#_c_219_n 0.00147245f $X=2.215 $Y=1.16
+ $X2=0 $Y2=0
cc_140 N_A_283_47#_c_165_n N_A_390_47#_c_219_n 0.010964f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_141 N_A_283_47#_c_162_n N_A_390_47#_c_219_n 0.0188032f $X=2.075 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_283_47#_c_165_n N_VPWR_c_270_n 0.0227813f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_143 N_A_283_47#_M1004_g N_VPWR_c_271_n 0.0231578f $X=2.465 $Y=2.075 $X2=0
+ $Y2=0
cc_144 N_A_283_47#_M1004_g N_VPWR_c_272_n 0.0181551f $X=2.465 $Y=2.075 $X2=0
+ $Y2=0
cc_145 N_A_283_47#_c_165_n N_VPWR_c_272_n 0.0224476f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_146 N_A_283_47#_M1005_d N_VPWR_c_269_n 0.00213418f $X=1.415 $Y=1.665 $X2=0
+ $Y2=0
cc_147 N_A_283_47#_M1004_g N_VPWR_c_269_n 0.030231f $X=2.465 $Y=2.075 $X2=0
+ $Y2=0
cc_148 N_A_283_47#_c_165_n N_VPWR_c_269_n 0.0131742f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_149 N_A_283_47#_c_161_n N_VGND_c_325_n 0.0115672f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_150 N_A_283_47#_M1006_g N_VGND_c_326_n 0.0156639f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_151 N_A_283_47#_M1006_g N_VGND_c_327_n 0.0148233f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_152 N_A_283_47#_c_161_n N_VGND_c_327_n 0.0224545f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_153 N_A_283_47#_M1001_d N_VGND_c_331_n 0.00209319f $X=1.415 $Y=0.235 $X2=0
+ $Y2=0
cc_154 N_A_283_47#_M1006_g N_VGND_c_331_n 0.0196071f $X=2.465 $Y=0.56 $X2=0
+ $Y2=0
cc_155 N_A_283_47#_c_161_n N_VGND_c_331_n 0.0131742f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_156 N_A_390_47#_M1007_g N_VPWR_c_271_n 0.00313672f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_390_47#_c_216_n N_VPWR_c_271_n 0.0210376f $X=2.075 $Y=1.96 $X2=0
+ $Y2=0
cc_158 N_A_390_47#_c_213_n N_VPWR_c_271_n 0.0105408f $X=3.075 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_390_47#_c_214_n N_VPWR_c_271_n 0.00131009f $X=3.075 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A_390_47#_c_216_n N_VPWR_c_272_n 0.0153696f $X=2.075 $Y=1.96 $X2=0
+ $Y2=0
cc_161 N_A_390_47#_M1007_g N_VPWR_c_275_n 0.00585385f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_390_47#_M1004_s N_VPWR_c_269_n 0.00355752f $X=1.95 $Y=1.665 $X2=0
+ $Y2=0
cc_163 N_A_390_47#_M1007_g N_VPWR_c_269_n 0.0116522f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_390_47#_c_216_n N_VPWR_c_269_n 0.00936871f $X=2.075 $Y=1.96 $X2=0
+ $Y2=0
cc_165 N_A_390_47#_M1000_g X 0.0110953f $X=3.115 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_390_47#_M1007_g X 0.0114596f $X=3.115 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_390_47#_c_213_n X 0.0269587f $X=3.075 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_390_47#_c_214_n X 0.00750121f $X=3.075 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_390_47#_M1000_g N_VGND_c_326_n 0.0031594f $X=3.115 $Y=0.445 $X2=0
+ $Y2=0
cc_170 N_A_390_47#_c_220_n N_VGND_c_326_n 0.0115206f $X=2.075 $Y=0.435 $X2=0
+ $Y2=0
cc_171 N_A_390_47#_c_213_n N_VGND_c_326_n 0.0127813f $X=3.075 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_390_47#_c_214_n N_VGND_c_326_n 0.00144312f $X=3.075 $Y=1.16 $X2=0
+ $Y2=0
cc_173 N_A_390_47#_c_220_n N_VGND_c_327_n 0.0153182f $X=2.075 $Y=0.435 $X2=0
+ $Y2=0
cc_174 N_A_390_47#_c_212_n N_VGND_c_327_n 0.00474075f $X=2.495 $Y=1.325 $X2=0
+ $Y2=0
cc_175 N_A_390_47#_M1000_g N_VGND_c_330_n 0.00585385f $X=3.115 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A_390_47#_M1006_s N_VGND_c_331_n 0.00355752f $X=1.95 $Y=0.235 $X2=0
+ $Y2=0
cc_177 N_A_390_47#_M1000_g N_VGND_c_331_n 0.0117573f $X=3.115 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_390_47#_c_220_n N_VGND_c_331_n 0.00935558f $X=2.075 $Y=0.435 $X2=0
+ $Y2=0
cc_179 N_A_390_47#_c_212_n N_VGND_c_331_n 0.0075282f $X=2.495 $Y=1.325 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_269_n N_X_M1007_d 0.002872f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_181 N_VPWR_c_275_n X 0.0264556f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_182 N_VPWR_c_269_n X 0.0155202f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_183 N_X_c_312_n N_VGND_c_330_n 0.0261793f $X=3.345 $Y=0.435 $X2=0 $Y2=0
cc_184 N_X_M1000_d N_VGND_c_331_n 0.002872f $X=3.19 $Y=0.235 $X2=0 $Y2=0
cc_185 N_X_c_312_n N_VGND_c_331_n 0.0154359f $X=3.345 $Y=0.435 $X2=0 $Y2=0

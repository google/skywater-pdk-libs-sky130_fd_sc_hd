* File: sky130_fd_sc_hd__a21oi_4.pxi.spice
* Created: Tue Sep  1 18:52:30 2020
* 
x_PM_SKY130_FD_SC_HD__A21OI_4%B1 N_B1_c_89_n N_B1_M1008_g N_B1_M1006_g
+ N_B1_c_90_n N_B1_M1013_g N_B1_M1011_g N_B1_c_91_n N_B1_M1014_g N_B1_M1012_g
+ N_B1_c_92_n N_B1_M1023_g N_B1_M1022_g N_B1_c_93_n B1 N_B1_c_100_n N_B1_c_94_n
+ PM_SKY130_FD_SC_HD__A21OI_4%B1
x_PM_SKY130_FD_SC_HD__A21OI_4%A2 N_A2_M1001_g N_A2_M1000_g N_A2_c_162_n
+ N_A2_M1005_g N_A2_M1010_g N_A2_c_163_n N_A2_M1017_g N_A2_M1016_g N_A2_c_164_n
+ N_A2_M1021_g N_A2_M1020_g N_A2_c_165_n N_A2_c_166_n N_A2_c_185_n N_A2_c_167_n
+ N_A2_c_178_n A2 N_A2_c_168_n N_A2_c_169_n N_A2_c_170_n
+ PM_SKY130_FD_SC_HD__A21OI_4%A2
x_PM_SKY130_FD_SC_HD__A21OI_4%A1 N_A1_c_290_n N_A1_M1003_g N_A1_M1002_g
+ N_A1_c_292_n N_A1_M1004_g N_A1_M1007_g N_A1_c_294_n N_A1_M1018_g N_A1_M1009_g
+ N_A1_c_296_n N_A1_M1019_g N_A1_M1015_g A1 PM_SKY130_FD_SC_HD__A21OI_4%A1
x_PM_SKY130_FD_SC_HD__A21OI_4%A_28_297# N_A_28_297#_M1006_d N_A_28_297#_M1011_d
+ N_A_28_297#_M1022_d N_A_28_297#_M1002_s N_A_28_297#_M1009_s
+ N_A_28_297#_M1010_s N_A_28_297#_M1020_s N_A_28_297#_c_421_p
+ N_A_28_297#_c_364_n N_A_28_297#_c_366_n N_A_28_297#_c_377_n
+ N_A_28_297#_c_368_n N_A_28_297#_c_413_p N_A_28_297#_c_381_n
+ N_A_28_297#_c_416_p N_A_28_297#_c_382_n N_A_28_297#_c_419_p
+ N_A_28_297#_c_384_n N_A_28_297#_c_362_n N_A_28_297#_c_363_n
+ N_A_28_297#_c_390_n N_A_28_297#_c_391_n N_A_28_297#_c_392_n
+ PM_SKY130_FD_SC_HD__A21OI_4%A_28_297#
x_PM_SKY130_FD_SC_HD__A21OI_4%Y N_Y_M1008_d N_Y_M1014_d N_Y_M1003_s N_Y_M1018_s
+ N_Y_M1006_s N_Y_M1012_s N_Y_c_450_n N_Y_c_502_p N_Y_c_445_n N_Y_c_460_n
+ N_Y_c_446_n N_Y_c_447_n N_Y_c_463_n N_Y_c_448_n Y N_Y_c_465_n
+ PM_SKY130_FD_SC_HD__A21OI_4%Y
x_PM_SKY130_FD_SC_HD__A21OI_4%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_M1015_d
+ N_VPWR_M1016_d N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n N_VPWR_c_524_n
+ N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n
+ N_VPWR_c_530_n VPWR N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_520_n
+ N_VPWR_c_534_n PM_SKY130_FD_SC_HD__A21OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A21OI_4%VGND N_VGND_M1008_s N_VGND_M1013_s N_VGND_M1023_s
+ N_VGND_M1005_d N_VGND_M1021_d N_VGND_c_623_n N_VGND_c_624_n N_VGND_c_625_n
+ N_VGND_c_626_n N_VGND_c_627_n N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n
+ N_VGND_c_631_n N_VGND_c_632_n VGND N_VGND_c_633_n N_VGND_c_634_n
+ N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n
+ PM_SKY130_FD_SC_HD__A21OI_4%VGND
x_PM_SKY130_FD_SC_HD__A21OI_4%A_462_47# N_A_462_47#_M1000_s N_A_462_47#_M1004_d
+ N_A_462_47#_M1019_d N_A_462_47#_M1017_s N_A_462_47#_c_718_n
+ N_A_462_47#_c_719_n N_A_462_47#_c_720_n N_A_462_47#_c_716_n
+ N_A_462_47#_c_717_n N_A_462_47#_c_731_n PM_SKY130_FD_SC_HD__A21OI_4%A_462_47#
cc_1 VNB N_B1_c_89_n 0.0212151f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_B1_c_90_n 0.0160046f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_B1_c_91_n 0.0159819f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_4 VNB N_B1_c_92_n 0.0154089f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.995
cc_5 VNB N_B1_c_93_n 0.0126238f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.205
cc_6 VNB N_B1_c_94_n 0.0830682f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_7 VNB N_A2_c_162_n 0.016129f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_8 VNB N_A2_c_163_n 0.0159999f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_9 VNB N_A2_c_164_n 0.0219817f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.995
cc_10 VNB N_A2_c_165_n 0.00159939f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_11 VNB N_A2_c_166_n 0.0238251f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_12 VNB N_A2_c_167_n 0.00235101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_168_n 0.016777f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=1.16
cc_14 VNB N_A2_c_169_n 0.061598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_170_n 0.00961897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_290_n 0.0160486f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_17 VNB N_A1_M1002_g 3.5465e-19 $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_18 VNB N_A1_c_292_n 0.0158334f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_19 VNB N_A1_M1007_g 3.82449e-19 $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_20 VNB N_A1_c_294_n 0.0158329f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_21 VNB N_A1_M1009_g 3.82449e-19 $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.985
cc_22 VNB N_A1_c_296_n 0.0879521f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.995
cc_23 VNB N_A1_M1015_g 4.33197e-19 $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.985
cc_24 VNB A1 0.00170867f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.225
cc_25 VNB N_Y_c_445_n 0.0042958f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.985
cc_26 VNB N_Y_c_446_n 4.56702e-19 $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.225
cc_27 VNB N_Y_c_447_n 0.00972875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_448_n 0.00656144f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=1.16
cc_29 VNB N_VPWR_c_520_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_623_n 0.0103023f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.56
cc_31 VNB N_VGND_c_624_n 0.025217f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.325
cc_32 VNB N_VGND_c_625_n 3.12649e-19 $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.995
cc_33 VNB N_VGND_c_626_n 0.00252906f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.985
cc_34 VNB N_VGND_c_627_n 0.00421457f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.205
cc_35 VNB N_VGND_c_628_n 0.0359713f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.205
cc_36 VNB N_VGND_c_629_n 0.0547347f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_37 VNB N_VGND_c_630_n 0.00362081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_631_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_39 VNB N_VGND_c_632_n 0.00499771f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=1.16
cc_40 VNB N_VGND_c_633_n 0.0125022f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.16
cc_41 VNB N_VGND_c_634_n 0.0120227f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=1.225
cc_42 VNB N_VGND_c_635_n 0.0134401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_636_n 0.304744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_637_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_638_n 0.0042586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_462_47#_c_716_n 0.00452179f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.56
cc_47 VNB N_A_462_47#_c_717_n 0.003364f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.56
cc_48 VPB N_B1_M1006_g 0.0241139f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_49 VPB N_B1_M1011_g 0.0180113f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_50 VPB N_B1_M1012_g 0.0179965f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_51 VPB N_B1_M1022_g 0.0177211f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_52 VPB N_B1_c_93_n 0.0114231f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.205
cc_53 VPB N_B1_c_100_n 0.00683265f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=1.16
cc_54 VPB N_B1_c_94_n 0.021017f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.16
cc_55 VPB N_A2_M1001_g 0.0176318f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_56 VPB N_A2_M1010_g 0.0171445f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_57 VPB N_A2_M1016_g 0.017124f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_58 VPB N_A2_M1020_g 0.0222503f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_59 VPB N_A2_c_165_n 0.00276621f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_60 VPB N_A2_c_166_n 0.00631169f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_61 VPB N_A2_c_167_n 0.00197902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A2_c_178_n 0.0136346f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_63 VPB N_A2_c_169_n 0.0123305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A2_c_170_n 0.00733094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A1_M1002_g 0.0196283f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_66 VPB N_A1_M1007_g 0.0193016f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_67 VPB N_A1_M1009_g 0.0193016f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_68 VPB N_A1_M1015_g 0.0196386f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_69 VPB A1 0.00799673f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.225
cc_70 VPB N_A_28_297#_c_362_n 0.0112688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_28_297#_c_363_n 0.0137952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_Y_c_445_n 0.00238794f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_73 VPB N_VPWR_c_521_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=1.335 $Y2=0.995
cc_74 VPB N_VPWR_c_522_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_75 VPB N_VPWR_c_523_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=1.765 $Y2=0.56
cc_76 VPB N_VPWR_c_524_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_77 VPB N_VPWR_c_525_n 0.0113516f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.205
cc_78 VPB N_VPWR_c_526_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_79 VPB N_VPWR_c_527_n 0.0113516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_528_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.205
cc_81 VPB N_VPWR_c_529_n 0.0113994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_530_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_83 VPB N_VPWR_c_531_n 0.0542572f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_84 VPB N_VPWR_c_532_n 0.0228555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_520_n 0.0568425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_534_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 N_B1_M1022_g N_A2_M1001_g 0.0357673f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_88 N_B1_M1022_g N_A2_c_165_n 5.08272e-19 $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B1_c_94_n N_A2_c_165_n 2.96609e-19 $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B1_c_94_n N_A2_c_166_n 0.0207157f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B1_M1022_g N_A2_c_185_n 8.40721e-19 $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B1_c_92_n N_A2_c_168_n 0.0218566f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_93 N_B1_c_93_n N_A_28_297#_c_364_n 0.00879422f $X=0.4 $Y=1.205 $X2=0 $Y2=0
cc_94 N_B1_c_94_n N_A_28_297#_c_364_n 0.00104676f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B1_M1006_g N_A_28_297#_c_366_n 0.0146159f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_96 N_B1_M1011_g N_A_28_297#_c_366_n 0.00863478f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B1_M1011_g N_A_28_297#_c_368_n 0.00128732f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B1_M1012_g N_A_28_297#_c_368_n 0.0100298f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_99 N_B1_M1022_g N_A_28_297#_c_368_n 0.0166494f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B1_c_90_n N_Y_c_450_n 0.0122034f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_c_91_n N_Y_c_450_n 0.0115395f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_100_n N_Y_c_450_n 0.0418688f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B1_c_94_n N_Y_c_450_n 0.00237219f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B1_c_91_n N_Y_c_445_n 0.00220255f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B1_M1012_g N_Y_c_445_n 0.0040742f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B1_c_92_n N_Y_c_445_n 0.0024509f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_M1022_g N_Y_c_445_n 0.0190092f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B1_c_100_n N_Y_c_445_n 0.030578f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B1_c_94_n N_Y_c_445_n 0.0141892f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B1_c_91_n N_Y_c_460_n 7.42475e-19 $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B1_c_92_n N_Y_c_460_n 0.00899399f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B1_c_94_n N_Y_c_460_n 0.00454735f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B1_c_100_n N_Y_c_463_n 0.0143498f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_c_94_n N_Y_c_463_n 0.00241784f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B1_M1011_g N_Y_c_465_n 0.0166049f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_M1012_g N_Y_c_465_n 0.0170404f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B1_c_100_n N_Y_c_465_n 0.060644f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_118 N_B1_c_94_n N_Y_c_465_n 0.00499462f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_M1022_g N_VPWR_c_521_n 0.00101195f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_M1006_g N_VPWR_c_531_n 0.00357877f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B1_M1011_g N_VPWR_c_531_n 0.00357842f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1012_g N_VPWR_c_531_n 0.00357668f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1022_g N_VPWR_c_531_n 0.00357668f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_M1006_g N_VPWR_c_520_n 0.00621154f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_125 N_B1_M1011_g N_VPWR_c_520_n 0.00527891f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_M1012_g N_VPWR_c_520_n 0.00527877f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B1_M1022_g N_VPWR_c_520_n 0.00537502f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B1_c_89_n N_VGND_c_624_n 0.0118723f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B1_c_90_n N_VGND_c_624_n 8.28108e-19 $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_93_n N_VGND_c_624_n 0.0216211f $X=0.4 $Y=1.205 $X2=0 $Y2=0
cc_131 N_B1_c_100_n N_VGND_c_624_n 0.00145496f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B1_c_94_n N_VGND_c_624_n 0.00650316f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_133 N_B1_c_89_n N_VGND_c_625_n 7.79461e-19 $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B1_c_90_n N_VGND_c_625_n 0.00709932f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B1_c_91_n N_VGND_c_625_n 0.00630134f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B1_c_92_n N_VGND_c_625_n 5.06577e-19 $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_91_n N_VGND_c_626_n 5.08148e-19 $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_92_n N_VGND_c_626_n 0.00574609f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_89_n N_VGND_c_633_n 0.00486043f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_90_n N_VGND_c_633_n 0.00351072f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_c_91_n N_VGND_c_634_n 0.00351072f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_92_n N_VGND_c_634_n 0.00418359f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B1_c_89_n N_VGND_c_636_n 0.00830219f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B1_c_90_n N_VGND_c_636_n 0.00411677f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B1_c_91_n N_VGND_c_636_n 0.0040731f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B1_c_92_n N_VGND_c_636_n 0.0048233f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A2_c_168_n N_A1_c_290_n 0.0245688f $X=2.215 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A2_M1001_g N_A1_M1002_g 0.0419819f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A2_c_165_n N_A1_M1002_g 0.00392475f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_178_n N_A1_M1002_g 0.0125777f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_151 N_A2_c_178_n N_A1_M1007_g 0.0125621f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_152 N_A2_c_178_n N_A1_M1009_g 0.0125621f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_153 N_A2_c_162_n N_A1_c_296_n 0.0240403f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A2_c_165_n N_A1_c_296_n 7.52702e-19 $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_166_n N_A1_c_296_n 0.0223423f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_c_167_n N_A1_c_296_n 0.00648306f $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_157 N_A2_c_178_n N_A1_c_296_n 0.00207346f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_158 N_A2_c_169_n N_A1_c_296_n 0.0240403f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_M1010_g N_A1_M1015_g 0.0240403f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A2_c_178_n N_A1_M1015_g 0.0134561f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_161 N_A2_c_165_n A1 0.0215566f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A2_c_166_n A1 8.88438e-19 $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A2_c_167_n A1 0.0167772f $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_164 N_A2_c_178_n A1 0.109007f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_165 N_A2_c_169_n A1 3.1221e-19 $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A2_c_185_n N_A_28_297#_M1022_d 0.00239676f $X=2.395 $Y=1.592 $X2=0
+ $Y2=0
cc_167 N_A2_c_178_n N_A_28_297#_M1002_s 0.00177993f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_168 N_A2_c_178_n N_A_28_297#_M1009_s 0.00177993f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_169 N_A2_c_167_n N_A_28_297#_M1010_s 2.54531e-19 $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_170 N_A2_c_170_n N_A_28_297#_M1010_s 0.00157145f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A2_c_170_n N_A_28_297#_M1020_s 0.0109084f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_M1001_g N_A_28_297#_c_377_n 0.0135032f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_c_185_n N_A_28_297#_c_377_n 0.0147522f $X=2.395 $Y=1.592 $X2=0 $Y2=0
cc_174 N_A2_c_178_n N_A_28_297#_c_377_n 0.02103f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_175 N_A2_c_185_n N_A_28_297#_c_368_n 0.00381962f $X=2.395 $Y=1.592 $X2=0
+ $Y2=0
cc_176 N_A2_c_178_n N_A_28_297#_c_381_n 0.0337896f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_177 N_A2_M1010_g N_A_28_297#_c_382_n 0.0137977f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_c_178_n N_A_28_297#_c_382_n 0.0348689f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_179 N_A2_M1016_g N_A_28_297#_c_384_n 0.0138609f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A2_M1020_g N_A_28_297#_c_384_n 0.01108f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A2_c_169_n N_A_28_297#_c_384_n 3.267e-19 $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A2_c_170_n N_A_28_297#_c_384_n 0.03668f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A2_c_169_n N_A_28_297#_c_362_n 2.48761e-19 $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A2_c_170_n N_A_28_297#_c_362_n 0.00821211f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A2_c_178_n N_A_28_297#_c_390_n 0.01361f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_186 N_A2_c_178_n N_A_28_297#_c_391_n 0.01361f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_187 N_A2_c_167_n N_A_28_297#_c_392_n 0.0146138f $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_188 N_A2_c_169_n N_A_28_297#_c_392_n 3.5494e-19 $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_M1001_g N_Y_c_445_n 0.0014992f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A2_c_165_n N_Y_c_445_n 0.0331237f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A2_c_166_n N_Y_c_445_n 0.0030176f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A2_c_185_n N_Y_c_445_n 0.00488434f $X=2.395 $Y=1.592 $X2=0 $Y2=0
cc_193 N_A2_c_168_n N_Y_c_445_n 0.00201402f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_166_n N_Y_c_446_n 0.00171462f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A2_c_168_n N_Y_c_446_n 0.00464606f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_178_n N_Y_c_447_n 0.00563538f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_197 N_A2_c_165_n N_Y_c_448_n 0.0270822f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A2_c_166_n N_Y_c_448_n 0.00274735f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A2_c_168_n N_Y_c_448_n 0.00906787f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_185_n N_VPWR_M1001_d 4.097e-19 $X=2.395 $Y=1.592 $X2=-0.19
+ $Y2=-0.24
cc_201 N_A2_c_178_n N_VPWR_M1001_d 0.00147256f $X=4.225 $Y=1.39 $X2=-0.19
+ $Y2=-0.24
cc_202 N_A2_c_178_n N_VPWR_M1007_d 0.00178427f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_203 N_A2_c_167_n N_VPWR_M1015_d 3.10624e-19 $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_204 N_A2_c_178_n N_VPWR_M1015_d 0.00147256f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_205 N_A2_c_170_n N_VPWR_M1016_d 0.00184156f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A2_M1001_g N_VPWR_c_521_n 0.00685925f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A2_M1010_g N_VPWR_c_523_n 0.00621909f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_M1016_g N_VPWR_c_523_n 4.98572e-19 $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_M1010_g N_VPWR_c_524_n 5.01519e-19 $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1016_g N_VPWR_c_524_n 0.0062985f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A2_M1020_g N_VPWR_c_524_n 0.00788945f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A2_M1010_g N_VPWR_c_529_n 0.00351072f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A2_M1016_g N_VPWR_c_529_n 0.00351072f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A2_M1001_g N_VPWR_c_531_n 0.00379212f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A2_M1020_g N_VPWR_c_532_n 0.00351072f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A2_M1001_g N_VPWR_c_520_n 0.00445145f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A2_M1010_g N_VPWR_c_520_n 0.0040731f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A2_M1016_g N_VPWR_c_520_n 0.0040731f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A2_M1020_g N_VPWR_c_520_n 0.00517613f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A2_c_168_n N_VGND_c_626_n 0.00293166f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A2_c_162_n N_VGND_c_627_n 0.00275982f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_163_n N_VGND_c_627_n 0.00151324f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_164_n N_VGND_c_628_n 0.00325061f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_169_n N_VGND_c_628_n 0.00183945f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A2_c_170_n N_VGND_c_628_n 0.00793512f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A2_c_162_n N_VGND_c_629_n 0.00425616f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A2_c_168_n N_VGND_c_629_n 0.00420889f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_163_n N_VGND_c_631_n 0.00427134f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A2_c_164_n N_VGND_c_631_n 0.0054895f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A2_c_162_n N_VGND_c_636_n 0.00583934f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A2_c_163_n N_VGND_c_636_n 0.00580493f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A2_c_164_n N_VGND_c_636_n 0.0108297f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A2_c_168_n N_VGND_c_636_n 0.00587292f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_168_n N_A_462_47#_c_718_n 0.0030746f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_162_n N_A_462_47#_c_719_n 0.00274319f $X=4.385 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A2_c_162_n N_A_462_47#_c_720_n 0.00354489f $X=4.385 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A2_c_163_n N_A_462_47#_c_720_n 4.5244e-19 $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A2_c_162_n N_A_462_47#_c_716_n 0.00883987f $X=4.385 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A2_c_163_n N_A_462_47#_c_716_n 0.00975354f $X=4.815 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A2_c_164_n N_A_462_47#_c_716_n 0.00312188f $X=5.245 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A2_c_167_n N_A_462_47#_c_716_n 0.040856f $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_242 N_A2_c_169_n N_A_462_47#_c_716_n 0.00502404f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A2_c_170_n N_A_462_47#_c_716_n 0.0287976f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A2_c_162_n N_A_462_47#_c_717_n 9.23859e-19 $X=4.385 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A2_c_167_n N_A_462_47#_c_717_n 0.00994332f $X=4.54 $Y=1.39 $X2=0 $Y2=0
cc_246 N_A2_c_178_n N_A_462_47#_c_717_n 0.00548957f $X=4.225 $Y=1.39 $X2=0 $Y2=0
cc_247 N_A2_c_162_n N_A_462_47#_c_731_n 5.22552e-19 $X=4.385 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A2_c_163_n N_A_462_47#_c_731_n 0.00627823f $X=4.815 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A2_c_164_n N_A_462_47#_c_731_n 0.00529965f $X=5.245 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A1_M1002_g N_A_28_297#_c_377_n 0.0110962f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A1_M1007_g N_A_28_297#_c_381_n 0.01108f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A1_M1009_g N_A_28_297#_c_381_n 0.01108f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A1_M1015_g N_A_28_297#_c_382_n 0.0110168f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A1_c_290_n N_Y_c_447_n 0.00981933f $X=2.665 $Y=0.99 $X2=0 $Y2=0
cc_255 N_A1_c_292_n N_Y_c_447_n 0.00987975f $X=3.095 $Y=0.99 $X2=0 $Y2=0
cc_256 N_A1_c_294_n N_Y_c_447_n 0.00987975f $X=3.525 $Y=0.99 $X2=0 $Y2=0
cc_257 N_A1_c_296_n N_Y_c_447_n 0.0102606f $X=3.955 $Y=0.99 $X2=0 $Y2=0
cc_258 A1 N_Y_c_447_n 0.0987456f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_259 N_A1_M1002_g N_VPWR_c_521_n 0.00626401f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A1_M1007_g N_VPWR_c_521_n 4.98572e-19 $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A1_M1002_g N_VPWR_c_522_n 4.98572e-19 $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A1_M1007_g N_VPWR_c_522_n 0.00625485f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_M1009_g N_VPWR_c_522_n 0.00625485f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A1_M1015_g N_VPWR_c_522_n 4.98572e-19 $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A1_M1009_g N_VPWR_c_523_n 4.98572e-19 $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A1_M1015_g N_VPWR_c_523_n 0.00621909f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A1_M1002_g N_VPWR_c_525_n 0.00351072f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A1_M1007_g N_VPWR_c_525_n 0.00351072f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A1_M1009_g N_VPWR_c_527_n 0.00351072f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A1_M1015_g N_VPWR_c_527_n 0.00351072f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A1_M1002_g N_VPWR_c_520_n 0.0040731f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A1_M1007_g N_VPWR_c_520_n 0.0040731f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A1_M1009_g N_VPWR_c_520_n 0.0040731f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A1_M1015_g N_VPWR_c_520_n 0.0040731f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A1_c_290_n N_VGND_c_629_n 0.00357877f $X=2.665 $Y=0.99 $X2=0 $Y2=0
cc_276 N_A1_c_292_n N_VGND_c_629_n 0.00357877f $X=3.095 $Y=0.99 $X2=0 $Y2=0
cc_277 N_A1_c_294_n N_VGND_c_629_n 0.00357877f $X=3.525 $Y=0.99 $X2=0 $Y2=0
cc_278 N_A1_c_296_n N_VGND_c_629_n 0.00357877f $X=3.955 $Y=0.99 $X2=0 $Y2=0
cc_279 N_A1_c_290_n N_VGND_c_636_n 0.00530427f $X=2.665 $Y=0.99 $X2=0 $Y2=0
cc_280 N_A1_c_292_n N_VGND_c_636_n 0.00527894f $X=3.095 $Y=0.99 $X2=0 $Y2=0
cc_281 N_A1_c_294_n N_VGND_c_636_n 0.00527894f $X=3.525 $Y=0.99 $X2=0 $Y2=0
cc_282 N_A1_c_296_n N_VGND_c_636_n 0.00530427f $X=3.955 $Y=0.99 $X2=0 $Y2=0
cc_283 N_A1_c_290_n N_A_462_47#_c_718_n 0.00979905f $X=2.665 $Y=0.99 $X2=0 $Y2=0
cc_284 N_A1_c_292_n N_A_462_47#_c_718_n 0.00979905f $X=3.095 $Y=0.99 $X2=0 $Y2=0
cc_285 N_A1_c_294_n N_A_462_47#_c_718_n 0.00979905f $X=3.525 $Y=0.99 $X2=0 $Y2=0
cc_286 N_A1_c_296_n N_A_462_47#_c_718_n 0.0119595f $X=3.955 $Y=0.99 $X2=0 $Y2=0
cc_287 A1 N_A_462_47#_c_718_n 0.00255981f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_288 N_A1_c_296_n N_A_462_47#_c_717_n 4.2252e-19 $X=3.955 $Y=0.99 $X2=0 $Y2=0
cc_289 N_A_28_297#_c_366_n N_Y_M1006_s 0.00341119f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_290 N_A_28_297#_c_368_n N_Y_M1012_s 0.00335313f $X=2.115 $Y=1.99 $X2=0 $Y2=0
cc_291 N_A_28_297#_c_368_n N_Y_c_445_n 0.023777f $X=2.115 $Y=1.99 $X2=0 $Y2=0
cc_292 N_A_28_297#_M1011_d N_Y_c_465_n 0.00338071f $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_293 N_A_28_297#_c_366_n N_Y_c_465_n 0.0206064f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_294 N_A_28_297#_c_368_n N_Y_c_465_n 0.0357328f $X=2.115 $Y=1.99 $X2=0 $Y2=0
cc_295 N_A_28_297#_c_377_n N_VPWR_M1001_d 0.00367764f $X=2.785 $Y=1.99 $X2=-0.19
+ $Y2=1.305
cc_296 N_A_28_297#_c_381_n N_VPWR_M1007_d 0.00339518f $X=3.645 $Y=1.99 $X2=0
+ $Y2=0
cc_297 N_A_28_297#_c_382_n N_VPWR_M1015_d 0.00349236f $X=4.505 $Y=1.99 $X2=0
+ $Y2=0
cc_298 N_A_28_297#_c_384_n N_VPWR_M1016_d 0.00338714f $X=5.365 $Y=1.99 $X2=0
+ $Y2=0
cc_299 N_A_28_297#_c_377_n N_VPWR_c_521_n 0.0162775f $X=2.785 $Y=1.99 $X2=0
+ $Y2=0
cc_300 N_A_28_297#_c_381_n N_VPWR_c_522_n 0.0162283f $X=3.645 $Y=1.99 $X2=0
+ $Y2=0
cc_301 N_A_28_297#_c_382_n N_VPWR_c_523_n 0.0162283f $X=4.505 $Y=1.99 $X2=0
+ $Y2=0
cc_302 N_A_28_297#_c_384_n N_VPWR_c_524_n 0.0162283f $X=5.365 $Y=1.99 $X2=0
+ $Y2=0
cc_303 N_A_28_297#_c_377_n N_VPWR_c_525_n 0.00263122f $X=2.785 $Y=1.99 $X2=0
+ $Y2=0
cc_304 N_A_28_297#_c_413_p N_VPWR_c_525_n 0.0123333f $X=2.88 $Y=2.3 $X2=0 $Y2=0
cc_305 N_A_28_297#_c_381_n N_VPWR_c_525_n 0.00263122f $X=3.645 $Y=1.99 $X2=0
+ $Y2=0
cc_306 N_A_28_297#_c_381_n N_VPWR_c_527_n 0.00263122f $X=3.645 $Y=1.99 $X2=0
+ $Y2=0
cc_307 N_A_28_297#_c_416_p N_VPWR_c_527_n 0.0123333f $X=3.74 $Y=2.3 $X2=0 $Y2=0
cc_308 N_A_28_297#_c_382_n N_VPWR_c_527_n 0.00263122f $X=4.505 $Y=1.99 $X2=0
+ $Y2=0
cc_309 N_A_28_297#_c_382_n N_VPWR_c_529_n 0.00263838f $X=4.505 $Y=1.99 $X2=0
+ $Y2=0
cc_310 N_A_28_297#_c_419_p N_VPWR_c_529_n 0.0119785f $X=4.6 $Y=2.3 $X2=0 $Y2=0
cc_311 N_A_28_297#_c_384_n N_VPWR_c_529_n 0.00274153f $X=5.365 $Y=1.99 $X2=0
+ $Y2=0
cc_312 N_A_28_297#_c_421_p N_VPWR_c_531_n 0.0125853f $X=0.277 $Y=2.215 $X2=0
+ $Y2=0
cc_313 N_A_28_297#_c_366_n N_VPWR_c_531_n 0.0330048f $X=0.955 $Y=2.34 $X2=0
+ $Y2=0
cc_314 N_A_28_297#_c_377_n N_VPWR_c_531_n 0.00270999f $X=2.785 $Y=1.99 $X2=0
+ $Y2=0
cc_315 N_A_28_297#_c_368_n N_VPWR_c_531_n 0.0668997f $X=2.115 $Y=1.99 $X2=0
+ $Y2=0
cc_316 N_A_28_297#_c_384_n N_VPWR_c_532_n 0.00263122f $X=5.365 $Y=1.99 $X2=0
+ $Y2=0
cc_317 N_A_28_297#_c_363_n N_VPWR_c_532_n 0.0176323f $X=5.46 $Y=2.3 $X2=0 $Y2=0
cc_318 N_A_28_297#_M1006_d N_VPWR_c_520_n 0.00348184f $X=0.14 $Y=1.485 $X2=0
+ $Y2=0
cc_319 N_A_28_297#_M1011_d N_VPWR_c_520_n 0.00223231f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_320 N_A_28_297#_M1022_d N_VPWR_c_520_n 0.00258751f $X=1.84 $Y=1.485 $X2=0
+ $Y2=0
cc_321 N_A_28_297#_M1002_s N_VPWR_c_520_n 0.00251209f $X=2.74 $Y=1.485 $X2=0
+ $Y2=0
cc_322 N_A_28_297#_M1009_s N_VPWR_c_520_n 0.00251209f $X=3.6 $Y=1.485 $X2=0
+ $Y2=0
cc_323 N_A_28_297#_M1010_s N_VPWR_c_520_n 0.00254571f $X=4.46 $Y=1.485 $X2=0
+ $Y2=0
cc_324 N_A_28_297#_M1020_s N_VPWR_c_520_n 0.00227407f $X=5.32 $Y=1.485 $X2=0
+ $Y2=0
cc_325 N_A_28_297#_c_421_p N_VPWR_c_520_n 0.00750689f $X=0.277 $Y=2.215 $X2=0
+ $Y2=0
cc_326 N_A_28_297#_c_366_n N_VPWR_c_520_n 0.0204525f $X=0.955 $Y=2.34 $X2=0
+ $Y2=0
cc_327 N_A_28_297#_c_377_n N_VPWR_c_520_n 0.0100933f $X=2.785 $Y=1.99 $X2=0
+ $Y2=0
cc_328 N_A_28_297#_c_368_n N_VPWR_c_520_n 0.0420965f $X=2.115 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_28_297#_c_413_p N_VPWR_c_520_n 0.00721345f $X=2.88 $Y=2.3 $X2=0 $Y2=0
cc_330 N_A_28_297#_c_381_n N_VPWR_c_520_n 0.0101289f $X=3.645 $Y=1.99 $X2=0
+ $Y2=0
cc_331 N_A_28_297#_c_416_p N_VPWR_c_520_n 0.00721345f $X=3.74 $Y=2.3 $X2=0 $Y2=0
cc_332 N_A_28_297#_c_382_n N_VPWR_c_520_n 0.0101396f $X=4.505 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_28_297#_c_419_p N_VPWR_c_520_n 0.00682467f $X=4.6 $Y=2.3 $X2=0 $Y2=0
cc_334 N_A_28_297#_c_384_n N_VPWR_c_520_n 0.0104307f $X=5.365 $Y=1.99 $X2=0
+ $Y2=0
cc_335 N_A_28_297#_c_363_n N_VPWR_c_520_n 0.00989931f $X=5.46 $Y=2.3 $X2=0 $Y2=0
cc_336 N_Y_M1006_s N_VPWR_c_520_n 0.00224864f $X=0.55 $Y=1.485 $X2=0 $Y2=0
cc_337 N_Y_M1012_s N_VPWR_c_520_n 0.00224837f $X=1.41 $Y=1.485 $X2=0 $Y2=0
cc_338 N_Y_c_450_n N_VGND_M1013_s 0.00325948f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_339 N_Y_c_448_n N_VGND_M1023_s 0.00213857f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_340 N_Y_c_450_n N_VGND_c_625_n 0.0163189f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_341 N_Y_c_460_n N_VGND_c_626_n 2.80485e-19 $X=1.88 $Y=0.795 $X2=0 $Y2=0
cc_342 N_Y_c_448_n N_VGND_c_626_n 0.0161669f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_343 N_Y_c_448_n N_VGND_c_629_n 0.00202288f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_344 N_Y_c_450_n N_VGND_c_633_n 0.00264265f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_345 N_Y_c_463_n N_VGND_c_633_n 0.00699602f $X=0.69 $Y=0.535 $X2=0 $Y2=0
cc_346 N_Y_c_450_n N_VGND_c_634_n 0.00264265f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_347 N_Y_c_502_p N_VGND_c_634_n 0.0123798f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_348 N_Y_c_460_n N_VGND_c_634_n 0.00264231f $X=1.88 $Y=0.795 $X2=0 $Y2=0
cc_349 N_Y_M1008_d N_VGND_c_636_n 0.00408233f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_350 N_Y_M1014_d N_VGND_c_636_n 0.00256266f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_351 N_Y_M1003_s N_VGND_c_636_n 0.00224864f $X=2.74 $Y=0.235 $X2=0 $Y2=0
cc_352 N_Y_M1018_s N_VGND_c_636_n 0.00224864f $X=3.6 $Y=0.235 $X2=0 $Y2=0
cc_353 N_Y_c_450_n N_VGND_c_636_n 0.0102198f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_354 N_Y_c_502_p N_VGND_c_636_n 0.00722448f $X=1.55 $Y=0.42 $X2=0 $Y2=0
cc_355 N_Y_c_460_n N_VGND_c_636_n 0.00490637f $X=1.88 $Y=0.795 $X2=0 $Y2=0
cc_356 N_Y_c_446_n N_VGND_c_636_n 0.00313233f $X=2.385 $Y=0.785 $X2=0 $Y2=0
cc_357 N_Y_c_463_n N_VGND_c_636_n 0.00672198f $X=0.69 $Y=0.535 $X2=0 $Y2=0
cc_358 N_Y_c_448_n N_VGND_c_636_n 0.00467993f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_359 N_Y_c_447_n N_A_462_47#_M1000_s 0.00152947f $X=3.74 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_360 N_Y_c_447_n N_A_462_47#_M1004_d 0.00172716f $X=3.74 $Y=0.76 $X2=0 $Y2=0
cc_361 N_Y_M1003_s N_A_462_47#_c_718_n 0.00324321f $X=2.74 $Y=0.235 $X2=0 $Y2=0
cc_362 N_Y_M1018_s N_A_462_47#_c_718_n 0.00324321f $X=3.6 $Y=0.235 $X2=0 $Y2=0
cc_363 N_Y_c_446_n N_A_462_47#_c_718_n 0.0821126f $X=2.385 $Y=0.785 $X2=0 $Y2=0
cc_364 N_Y_c_447_n N_A_462_47#_c_717_n 0.00710427f $X=3.74 $Y=0.76 $X2=0 $Y2=0
cc_365 N_VGND_c_636_n N_A_462_47#_M1000_s 0.00223258f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_366 N_VGND_c_636_n N_A_462_47#_M1004_d 0.00223258f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_636_n N_A_462_47#_M1019_d 0.00223235f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_636_n N_A_462_47#_M1017_s 0.00223231f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_629_n N_A_462_47#_c_718_n 0.100183f $X=4.505 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_636_n N_A_462_47#_c_718_n 0.064026f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_629_n N_A_462_47#_c_719_n 0.0157493f $X=4.505 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_636_n N_A_462_47#_c_719_n 0.00981451f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_M1005_d N_A_462_47#_c_716_n 0.00172391f $X=4.46 $Y=0.235 $X2=0
+ $Y2=0
cc_374 N_VGND_c_627_n N_A_462_47#_c_716_n 0.0130261f $X=4.6 $Y=0.4 $X2=0 $Y2=0
cc_375 N_VGND_c_629_n N_A_462_47#_c_716_n 0.00196536f $X=4.505 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_c_631_n N_A_462_47#_c_716_n 0.00196536f $X=5.365 $Y=0 $X2=0 $Y2=0
cc_377 N_VGND_c_636_n N_A_462_47#_c_716_n 0.00828266f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_631_n N_A_462_47#_c_731_n 0.0188765f $X=5.365 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_636_n N_A_462_47#_c_731_n 0.0122527f $X=5.75 $Y=0 $X2=0 $Y2=0

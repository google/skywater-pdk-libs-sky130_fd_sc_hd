* NGSPICE file created from sky130_fd_sc_hd__sdfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1781_295# a_1597_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.65815e+12p ps=1.79e+07u
M1001 a_193_369# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=2.4568e+12p ps=2.316e+07u
M1002 a_1350_47# a_1006_47# a_1132_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u
M1003 VGND CLK a_652_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1004 a_181_47# D a_193_369# VPB phighvt w=640000u l=150000u
+  ad=3.204e+11p pd=3.3e+06u as=0p ps=0u
M1005 VPWR a_1597_329# a_2501_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1006 VPWR a_2501_47# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 a_1006_47# a_818_47# a_181_47# VPB phighvt w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1008 a_1132_21# a_1006_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.428e+11p pd=1.52e+06u as=0p ps=0u
M1009 VPWR a_1781_295# a_1723_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1010 VPWR CLK a_652_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1011 VGND a_1597_329# a_2501_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1012 VPWR a_1597_329# Q_N VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1013 a_1597_329# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=4.158e+11p pd=4e+06u as=0p ps=0u
M1014 VGND SET_B a_1885_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1015 a_1525_329# a_1006_47# VPWR VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1016 a_181_47# SCE a_109_47# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=8.82e+10p ps=1.26e+06u
M1017 Q a_2501_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1813_47# a_652_47# a_1597_329# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.44e+11p ps=2.18e+06u
M1019 a_1090_47# a_818_47# a_1006_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.134e+11p ps=1.38e+06u
M1020 a_1885_47# a_1781_295# a_1813_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1597_329# a_652_47# a_1525_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1132_21# a_1090_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1517_47# a_1006_47# VGND VNB nshort w=640000u l=150000u
+  ad=4.672e+11p pd=2.74e+06u as=0p ps=0u
M1024 VGND SCE a_328_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1025 VPWR SCD a_27_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.29225e+11p ps=3.6e+06u
M1026 a_1781_295# a_1597_329# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1027 a_265_47# D a_181_47# VNB nshort w=420000u l=150000u
+  ad=1.323e+11p pd=1.47e+06u as=0p ps=0u
M1028 Q_N a_1597_329# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR SCE a_328_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.62825e+11p ps=1.8e+06u
M1030 a_1006_47# a_652_47# a_181_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_818_47# a_652_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1032 a_27_369# a_328_21# a_181_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR SET_B a_1132_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1102_413# a_652_47# a_1006_47# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1035 VGND a_1597_329# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1036 VGND a_328_21# a_265_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SET_B a_1350_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q_N a_1597_329# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1723_413# a_818_47# a_1597_329# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_2501_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1041 a_109_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 Q a_2501_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1597_329# a_818_47# a_1517_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_1132_21# a_1102_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_818_47# a_652_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__o311ai_2.spice
* Created: Thu Aug 27 14:39:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o311ai_2.pex.spice"
.subckt sky130_fd_sc_hd__o311ai_2  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_A_55_47#_M1003_d N_A1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_55_47#_M1016_d N_A1_M1016_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_55_47#_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1009_d N_A2_M1018_g N_A_55_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1013 N_A_55_47#_M1018_s N_A3_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.23075 PD=0.92 PS=1.36 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.9
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1014 N_A_55_47#_M1014_d N_A3_M1014_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.23075 PD=0.92 PS=1.36 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_A_55_47#_M1014_d N_B1_M1005_g N_A_729_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_55_47#_M1008_d N_B1_M1008_g N_A_729_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g N_A_729_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_Y_M1017_d N_C1_M1017_g N_A_729_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_51_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1002_d N_A1_M1019_g N_A_51_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1006 N_A_51_297#_M1019_s N_A2_M1006_g N_A_301_297#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_51_297#_M1010_d N_A2_M1010_g N_A_301_297#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A3_M1000_g N_A_301_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A3_M1001_g N_A_301_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1011 N_Y_M1001_d N_B1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.305 PD=1.27 PS=1.61 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001.9 A=0.15
+ P=2.3 MULT=1
MM1015 N_Y_M1015_d N_B1_M1015_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.205
+ AS=0.305 PD=1.41 PS=1.61 NRD=12.7853 NRS=0 M=1 R=6.66667 SA=75001.8 SB=75001.2
+ A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1015_d N_C1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.205
+ AS=0.135 PD=1.41 PS=1.27 NRD=12.7853 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1012_d N_C1_M1012_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_53 VNB 0 1.40125e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__o311ai_2.pxi.spice"
*
.ends
*
*

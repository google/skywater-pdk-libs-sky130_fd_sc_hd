* File: sky130_fd_sc_hd__clkbuf_8.pxi.spice
* Created: Thu Aug 27 14:11:08 2020
* 
x_PM_SKY130_FD_SC_HD__CLKBUF_8%A N_A_M1004_g N_A_c_87_n N_A_M1007_g N_A_M1012_g
+ N_A_c_88_n N_A_M1018_g A A N_A_c_86_n PM_SKY130_FD_SC_HD__CLKBUF_8%A
x_PM_SKY130_FD_SC_HD__CLKBUF_8%A_110_47# N_A_110_47#_M1004_d N_A_110_47#_M1007_d
+ N_A_110_47#_M1001_g N_A_110_47#_M1000_g N_A_110_47#_M1006_g
+ N_A_110_47#_M1002_g N_A_110_47#_M1008_g N_A_110_47#_M1003_g
+ N_A_110_47#_M1010_g N_A_110_47#_M1005_g N_A_110_47#_M1014_g
+ N_A_110_47#_M1009_g N_A_110_47#_M1016_g N_A_110_47#_M1011_g
+ N_A_110_47#_M1017_g N_A_110_47#_M1013_g N_A_110_47#_c_129_n
+ N_A_110_47#_M1019_g N_A_110_47#_M1015_g N_A_110_47#_c_131_n
+ N_A_110_47#_c_142_n N_A_110_47#_c_132_n N_A_110_47#_c_155_n
+ PM_SKY130_FD_SC_HD__CLKBUF_8%A_110_47#
x_PM_SKY130_FD_SC_HD__CLKBUF_8%VPWR N_VPWR_M1007_s N_VPWR_M1018_s N_VPWR_M1002_s
+ N_VPWR_M1005_s N_VPWR_M1011_s N_VPWR_M1015_s N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n
+ N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n
+ N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n VPWR N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_268_n N_VPWR_c_287_n PM_SKY130_FD_SC_HD__CLKBUF_8%VPWR
x_PM_SKY130_FD_SC_HD__CLKBUF_8%X N_X_M1001_s N_X_M1008_s N_X_M1014_s N_X_M1017_s
+ N_X_M1000_d N_X_M1003_d N_X_M1009_d N_X_M1013_d N_X_c_346_n N_X_c_347_n
+ N_X_c_348_n N_X_c_370_n N_X_c_349_n N_X_c_350_n N_X_c_380_n N_X_c_351_n
+ N_X_c_352_n N_X_c_389_n N_X_c_353_n N_X_c_394_n N_X_c_354_n N_X_c_398_n
+ N_X_c_355_n N_X_c_402_n X X X PM_SKY130_FD_SC_HD__CLKBUF_8%X
x_PM_SKY130_FD_SC_HD__CLKBUF_8%VGND N_VGND_M1004_s N_VGND_M1012_s N_VGND_M1006_d
+ N_VGND_M1010_d N_VGND_M1016_d N_VGND_M1019_d N_VGND_c_463_n N_VGND_c_464_n
+ N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n
+ N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n VGND N_VGND_c_478_n
+ N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n PM_SKY130_FD_SC_HD__CLKBUF_8%VGND
cc_1 VNB N_A_M1004_g 0.0280927f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_M1012_g 0.0234436f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_3 VNB A 0.0260861f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_A_c_86_n 0.0669956f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.155
cc_5 VNB N_A_110_47#_M1001_g 0.0260664f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_6 VNB N_A_110_47#_M1006_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_110_47#_M1008_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_110_47#_M1010_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_110_47#_M1014_g 0.0241252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_110_47#_M1016_g 0.0241164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_110_47#_M1017_g 0.023767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_110_47#_c_129_n 0.151577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_110_47#_M1019_g 0.0320587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_110_47#_c_131_n 0.00445674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_c_132_n 0.00442652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_268_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_346_n 0.00160391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_347_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_348_n 0.00419804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_349_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_350_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_351_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_352_n 0.00400554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_353_n 0.0013724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_354_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_355_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB X 0.0301966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_463_n 0.0112866f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.155
cc_29 VNB N_VGND_c_464_n 0.00454665f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_30 VNB N_VGND_c_465_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_466_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.16
cc_32 VNB N_VGND_c_467_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_468_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_469_n 0.0177301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_470_n 0.0160902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_471_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_472_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_473_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_474_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_475_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_476_n 0.0154599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_477_n 0.00574315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_478_n 0.0166984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_479_n 0.0126445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_480_n 0.266016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_481_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VPB N_A_c_87_n 0.0192408f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.41
cc_48 VPB N_A_c_88_n 0.0145802f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.41
cc_49 VPB A 0.00123221f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_50 VPB N_A_c_86_n 0.0273976f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.155
cc_51 VPB N_A_110_47#_M1000_g 0.0190615f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_52 VPB N_A_110_47#_M1002_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_53 VPB N_A_110_47#_M1003_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.16
cc_54 VPB N_A_110_47#_M1005_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_110_47#_M1009_g 0.0187459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_110_47#_M1011_g 0.0187139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_110_47#_M1013_g 0.0173762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_110_47#_c_129_n 0.0250755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_110_47#_M1015_g 0.0224494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_110_47#_c_142_n 0.00140018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_110_47#_c_132_n 0.00331269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_269_n 0.0108797f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.155
cc_63 VPB N_VPWR_c_270_n 0.0416587f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_64 VPB N_VPWR_c_271_n 0.00400996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_272_n 0.00400996f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.16
cc_66 VPB N_VPWR_c_273_n 0.00400996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_274_n 0.00400996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_275_n 0.0272286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_276_n 0.016626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_277_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_278_n 0.016626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_279_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_280_n 0.016626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_281_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_282_n 0.016626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_283_n 0.00564836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_284_n 0.0167191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_285_n 0.0127268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_268_n 0.0532032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_287_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB X 0.010431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB X 0.0107432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 N_A_M1012_g N_A_110_47#_M1001_g 0.0204718f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_c_88_n N_A_110_47#_M1000_g 0.0204718f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_86_n N_A_110_47#_c_129_n 0.0204718f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_A_110_47#_c_131_n 0.0030957f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_M1012_g N_A_110_47#_c_131_n 0.00356184f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_88 A N_A_110_47#_c_131_n 0.0277994f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_c_86_n N_A_110_47#_c_131_n 0.0116674f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_90 N_A_c_87_n N_A_110_47#_c_142_n 0.00287039f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_88_n N_A_110_47#_c_142_n 0.00291483f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_86_n N_A_110_47#_c_142_n 0.00945812f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_93 N_A_c_86_n N_A_110_47#_c_132_n 0.0213857f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_94 A N_A_110_47#_c_155_n 0.0198893f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_95 N_A_c_86_n N_A_110_47#_c_155_n 0.00950927f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_96 N_A_c_87_n N_VPWR_c_270_n 0.00763298f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_97 A N_VPWR_c_270_n 0.0206626f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A_c_86_n N_VPWR_c_270_n 0.00767867f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_99 N_A_c_88_n N_VPWR_c_271_n 0.00258231f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_87_n N_VPWR_c_284_n 0.00585385f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_88_n N_VPWR_c_284_n 0.00585385f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_87_n N_VPWR_c_268_n 0.0116115f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_88_n N_VPWR_c_268_n 0.0106694f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_104 A N_VGND_c_463_n 0.00101698f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A_M1004_g N_VGND_c_464_n 0.00339198f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_106 A N_VGND_c_464_n 0.0191362f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_107 N_A_c_86_n N_VGND_c_464_n 0.00113059f $X=0.905 $Y=1.155 $X2=0 $Y2=0
cc_108 N_A_M1012_g N_VGND_c_465_n 0.00168046f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_M1004_g N_VGND_c_478_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_M1012_g N_VGND_c_478_n 0.00585385f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_M1004_g N_VGND_c_480_n 0.011499f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_M1012_g N_VGND_c_480_n 0.0106694f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_113 A N_VGND_c_480_n 0.00301823f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_114 N_A_110_47#_M1000_g N_VPWR_c_271_n 0.00258231f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_110_47#_c_132_n N_VPWR_c_271_n 0.0158218f $X=3.245 $Y=1.16 $X2=0
+ $Y2=0
cc_116 N_A_110_47#_M1002_g N_VPWR_c_272_n 0.00248982f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_110_47#_M1003_g N_VPWR_c_272_n 0.00248982f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_110_47#_M1005_g N_VPWR_c_273_n 0.00248982f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_110_47#_M1009_g N_VPWR_c_273_n 0.00248982f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_110_47#_M1011_g N_VPWR_c_274_n 0.00248982f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_110_47#_M1013_g N_VPWR_c_274_n 0.00248982f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_110_47#_M1015_g N_VPWR_c_275_n 0.00723036f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_110_47#_M1000_g N_VPWR_c_276_n 0.00585385f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_110_47#_M1002_g N_VPWR_c_276_n 0.00585385f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_110_47#_M1003_g N_VPWR_c_278_n 0.00585385f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_110_47#_M1005_g N_VPWR_c_278_n 0.00585385f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_110_47#_M1009_g N_VPWR_c_280_n 0.00585385f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_110_47#_M1011_g N_VPWR_c_280_n 0.00585385f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_110_47#_M1013_g N_VPWR_c_282_n 0.00585385f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_110_47#_M1015_g N_VPWR_c_282_n 0.00585385f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_110_47#_c_142_n N_VPWR_c_284_n 0.0141362f $X=0.69 $Y=1.69 $X2=0 $Y2=0
cc_132 N_A_110_47#_M1007_d N_VPWR_c_268_n 0.00336062f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_133 N_A_110_47#_M1000_g N_VPWR_c_268_n 0.0106694f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_110_47#_M1002_g N_VPWR_c_268_n 0.010643f $X=1.765 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_110_47#_M1003_g N_VPWR_c_268_n 0.010643f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_110_47#_M1005_g N_VPWR_c_268_n 0.010643f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_110_47#_M1009_g N_VPWR_c_268_n 0.010643f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_110_47#_M1011_g N_VPWR_c_268_n 0.010643f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_110_47#_M1013_g N_VPWR_c_268_n 0.010643f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_110_47#_M1015_g N_VPWR_c_268_n 0.0117793f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_110_47#_c_142_n N_VPWR_c_268_n 0.00952853f $X=0.69 $Y=1.69 $X2=0
+ $Y2=0
cc_142 N_A_110_47#_M1001_g N_X_c_346_n 0.00120255f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_110_47#_M1006_g N_X_c_346_n 0.00120255f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_110_47#_c_131_n N_X_c_346_n 0.00257148f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_110_47#_M1006_g N_X_c_347_n 0.0119364f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_110_47#_M1008_g N_X_c_347_n 0.0122327f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_110_47#_c_129_n N_X_c_347_n 0.00267078f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_148 N_A_110_47#_c_132_n N_X_c_347_n 0.0429599f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_110_47#_M1001_g N_X_c_348_n 0.00289158f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_110_47#_c_129_n N_X_c_348_n 0.00277135f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_151 N_A_110_47#_c_131_n N_X_c_348_n 0.00599637f $X=0.69 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A_110_47#_c_132_n N_X_c_348_n 0.0213686f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_110_47#_M1002_g N_X_c_370_n 0.0151109f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_110_47#_M1003_g N_X_c_370_n 0.015045f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_110_47#_c_129_n N_X_c_370_n 0.00232005f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_156 N_A_110_47#_c_132_n N_X_c_370_n 0.0385727f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_110_47#_M1008_g N_X_c_349_n 0.00120255f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_110_47#_M1010_g N_X_c_349_n 0.00120255f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_110_47#_M1010_g N_X_c_350_n 0.0122792f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_110_47#_M1014_g N_X_c_350_n 0.0122792f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_110_47#_c_129_n N_X_c_350_n 0.00267078f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_162 N_A_110_47#_c_132_n N_X_c_350_n 0.0429599f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_110_47#_M1005_g N_X_c_380_n 0.0151109f $X=2.625 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_110_47#_M1009_g N_X_c_380_n 0.0151109f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_110_47#_c_129_n N_X_c_380_n 0.00232005f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_166 N_A_110_47#_c_132_n N_X_c_380_n 0.0385727f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_110_47#_M1014_g N_X_c_351_n 0.00120255f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_110_47#_M1016_g N_X_c_351_n 0.00120255f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_110_47#_M1016_g N_X_c_352_n 0.0122792f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_170 N_A_110_47#_c_129_n N_X_c_352_n 0.00320502f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_171 N_A_110_47#_c_132_n N_X_c_352_n 0.0133842f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_110_47#_M1011_g N_X_c_389_n 0.0151109f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_110_47#_c_129_n N_X_c_389_n 0.00278134f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_174 N_A_110_47#_c_132_n N_X_c_389_n 0.0121568f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_110_47#_M1017_g N_X_c_353_n 0.00120255f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A_110_47#_M1019_g N_X_c_353_n 0.00221636f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A_110_47#_c_129_n N_X_c_394_n 0.00238948f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_178 N_A_110_47#_c_132_n N_X_c_394_n 0.0168441f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_110_47#_c_129_n N_X_c_354_n 0.00277135f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_180 N_A_110_47#_c_132_n N_X_c_354_n 0.0213686f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_110_47#_c_129_n N_X_c_398_n 0.00238948f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_182 N_A_110_47#_c_132_n N_X_c_398_n 0.0168441f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_110_47#_c_129_n N_X_c_355_n 0.00277135f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_184 N_A_110_47#_c_132_n N_X_c_355_n 0.0213686f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_110_47#_c_129_n N_X_c_402_n 0.00238948f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_186 N_A_110_47#_c_132_n N_X_c_402_n 0.0168441f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_110_47#_M1016_g X 0.00116814f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_110_47#_M1011_g X 0.00448672f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_110_47#_M1017_g X 0.0116551f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_110_47#_M1013_g X 0.0053012f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_110_47#_c_129_n X 0.0458412f $X=4.345 $Y=0.95 $X2=0 $Y2=0
cc_192 N_A_110_47#_M1019_g X 0.0136957f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_110_47#_M1015_g X 0.00773738f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_110_47#_c_132_n X 0.0208936f $X=3.245 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_110_47#_M1013_g X 0.0139693f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_110_47#_M1015_g X 0.0159698f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_110_47#_M1001_g N_VGND_c_465_n 0.00168046f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_198 N_A_110_47#_c_132_n N_VGND_c_465_n 0.00869033f $X=3.245 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_110_47#_M1006_g N_VGND_c_466_n 0.00161372f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_A_110_47#_M1008_g N_VGND_c_466_n 0.00161372f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_110_47#_M1010_g N_VGND_c_467_n 0.00161372f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_110_47#_M1014_g N_VGND_c_467_n 0.00161372f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_110_47#_M1016_g N_VGND_c_468_n 0.00161372f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_110_47#_M1017_g N_VGND_c_468_n 0.00161372f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_110_47#_M1019_g N_VGND_c_469_n 0.00341923f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_110_47#_M1001_g N_VGND_c_470_n 0.00585385f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_110_47#_M1006_g N_VGND_c_470_n 0.00439206f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_110_47#_M1008_g N_VGND_c_472_n 0.00439206f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_110_47#_M1010_g N_VGND_c_472_n 0.00439206f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_210 N_A_110_47#_M1014_g N_VGND_c_474_n 0.00439206f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_110_47#_M1016_g N_VGND_c_474_n 0.00439206f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_212 N_A_110_47#_M1017_g N_VGND_c_476_n 0.00439071f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_213 N_A_110_47#_M1019_g N_VGND_c_476_n 0.00439071f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_214 N_A_110_47#_c_131_n N_VGND_c_478_n 0.0137163f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_110_47#_M1004_d N_VGND_c_480_n 0.00336236f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_A_110_47#_M1001_g N_VGND_c_480_n 0.0106694f $X=1.335 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_110_47#_M1006_g N_VGND_c_480_n 0.00590932f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_110_47#_M1008_g N_VGND_c_480_n 0.00590932f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_A_110_47#_M1010_g N_VGND_c_480_n 0.00590932f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_110_47#_M1014_g N_VGND_c_480_n 0.00590932f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_110_47#_M1016_g N_VGND_c_480_n 0.00590932f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A_110_47#_M1017_g N_VGND_c_480_n 0.00590684f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_110_47#_M1019_g N_VGND_c_480_n 0.00700101f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_110_47#_c_131_n N_VGND_c_480_n 0.00950576f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_268_n N_X_M1000_d 0.00301352f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_c_268_n N_X_M1003_d 0.00301352f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_c_268_n N_X_M1009_d 0.00301352f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_268_n N_X_M1013_d 0.00301352f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_M1002_s N_X_c_370_n 0.00334014f $X=1.84 $Y=1.485 $X2=0 $Y2=0
cc_230 N_VPWR_c_272_n N_X_c_370_n 0.0138265f $X=1.98 $Y=2.22 $X2=0 $Y2=0
cc_231 N_VPWR_M1005_s N_X_c_380_n 0.00334014f $X=2.7 $Y=1.485 $X2=0 $Y2=0
cc_232 N_VPWR_c_273_n N_X_c_380_n 0.0138265f $X=2.84 $Y=2.22 $X2=0 $Y2=0
cc_233 N_VPWR_M1011_s N_X_c_389_n 0.00362232f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_234 N_VPWR_c_274_n N_X_c_389_n 0.0118724f $X=3.7 $Y=2.22 $X2=0 $Y2=0
cc_235 N_VPWR_c_276_n N_X_c_394_n 0.0144808f $X=1.85 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_c_268_n N_X_c_394_n 0.00991274f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_278_n N_X_c_398_n 0.0144808f $X=2.71 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_c_268_n N_X_c_398_n 0.00991274f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_239 N_VPWR_c_280_n N_X_c_402_n 0.0144808f $X=3.57 $Y=2.72 $X2=0 $Y2=0
cc_240 N_VPWR_c_268_n N_X_c_402_n 0.00991274f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_241 N_VPWR_M1011_s X 2.43457e-19 $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_242 N_VPWR_M1015_s X 0.00343092f $X=4.42 $Y=1.485 $X2=0 $Y2=0
cc_243 N_VPWR_c_274_n X 0.00202864f $X=3.7 $Y=2.22 $X2=0 $Y2=0
cc_244 N_VPWR_c_275_n X 0.0224079f $X=4.56 $Y=2.22 $X2=0 $Y2=0
cc_245 N_VPWR_c_282_n X 0.0144808f $X=4.43 $Y=2.72 $X2=0 $Y2=0
cc_246 N_VPWR_c_268_n X 0.00991274f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_247 N_X_c_347_n N_VGND_c_466_n 0.0164628f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_248 N_X_c_350_n N_VGND_c_467_n 0.0164628f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_249 N_X_c_352_n N_VGND_c_468_n 0.0129787f $X=3.76 $Y=0.82 $X2=0 $Y2=0
cc_250 X N_VGND_c_468_n 0.00403581f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_251 X N_VGND_c_469_n 0.0243348f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_252 N_X_c_346_n N_VGND_c_470_n 0.0128416f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_253 N_X_c_347_n N_VGND_c_470_n 0.00224999f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_254 N_X_c_347_n N_VGND_c_472_n 0.00224999f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_255 N_X_c_349_n N_VGND_c_472_n 0.0128416f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_256 N_X_c_350_n N_VGND_c_472_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_257 N_X_c_350_n N_VGND_c_474_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_258 N_X_c_351_n N_VGND_c_474_n 0.0128416f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_259 N_X_c_352_n N_VGND_c_474_n 0.00224999f $X=3.76 $Y=0.82 $X2=0 $Y2=0
cc_260 N_X_c_353_n N_VGND_c_476_n 0.0129027f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_261 X N_VGND_c_476_n 0.00498855f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_262 N_X_M1001_s N_VGND_c_480_n 0.00268444f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_263 N_X_M1008_s N_VGND_c_480_n 0.00234574f $X=2.27 $Y=0.235 $X2=0 $Y2=0
cc_264 N_X_M1014_s N_VGND_c_480_n 0.00234574f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_265 N_X_M1017_s N_VGND_c_480_n 0.00234544f $X=3.99 $Y=0.235 $X2=0 $Y2=0
cc_266 N_X_c_346_n N_VGND_c_480_n 0.00979224f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_267 N_X_c_347_n N_VGND_c_480_n 0.00829353f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_268 N_X_c_349_n N_VGND_c_480_n 0.00979224f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_269 N_X_c_350_n N_VGND_c_480_n 0.00829353f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_270 N_X_c_351_n N_VGND_c_480_n 0.00979224f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_271 N_X_c_352_n N_VGND_c_480_n 0.00436967f $X=3.76 $Y=0.82 $X2=0 $Y2=0
cc_272 N_X_c_353_n N_VGND_c_480_n 0.00981584f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_273 X N_VGND_c_480_n 0.00944699f $X=3.825 $Y=0.765 $X2=0 $Y2=0

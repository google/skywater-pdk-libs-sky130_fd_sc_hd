* File: sky130_fd_sc_hd__o22ai_2.spice
* Created: Thu Aug 27 14:37:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o22ai_2.pex.spice"
.subckt sky130_fd_sc_hd__o22ai_2  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_A_27_47#_M1004_d N_B1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1007_d N_B1_M1007_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g N_A_27_47#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1002_d N_B2_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.26975 PD=0.92 PS=1.48 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.26975 PD=0.92 PS=1.48 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1008_d N_A2_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 N_A_27_47#_M1014_s N_A1_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_A_27_47#_M1011_d N_A1_M1011_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1001_d N_B1_M1015_g N_A_27_297#_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1010 N_A_27_297#_M1015_s N_B2_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_A_27_297#_M1012_d N_B2_M1012_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_475_297#_M1000_d N_A2_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1003 N_A_475_297#_M1003_d N_A2_M1003_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1005 N_A_475_297#_M1003_d N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_A_475_297#_M1013_d N_A1_M1013_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__o22ai_2.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
M1000 a_147_105# SHORT VGND VNB nshort w=360000u l=150000u
+  ad=7.56e+10p pd=1.14e+06u as=9.36e+10p ps=1.24e+06u
M1001 a_291_105# SHORT a_219_105# VNB nshort w=360000u l=150000u
+  ad=7.56e+10p pd=1.14e+06u as=7.56e+10p ps=1.14e+06u
M1002 VPWR SHORT a_363_105# VNB nshort w=360000u l=150000u
+  ad=9.36e+10p pd=1.24e+06u as=7.56e+10p ps=1.14e+06u
M1003 a_363_105# SHORT a_291_105# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_219_105# SHORT a_147_105# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__and4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.450000 1.675000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.420000 1.800000 1.695000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 0.420000 2.295000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 0.665000 2.825000 1.695000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 0.295000 3.590000 0.340000 ;
        RECT 3.255000 0.340000 3.595000 0.805000 ;
        RECT 3.335000 1.495000 3.595000 2.465000 ;
        RECT 3.425000 0.805000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 2.755000  0.085000 3.085000 0.465000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.515000 2.195000 0.845000 2.635000 ;
        RECT 1.555000 2.225000 2.225000 2.635000 ;
        RECT 2.810000 2.225000 3.140000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.170000 0.255000 0.345000 0.655000 ;
      RECT 0.170000 0.655000 0.800000 0.825000 ;
      RECT 0.170000 1.845000 0.800000 2.015000 ;
      RECT 0.170000 2.015000 0.345000 2.465000 ;
      RECT 0.630000 0.825000 0.800000 0.995000 ;
      RECT 0.630000 0.995000 0.980000 1.325000 ;
      RECT 0.630000 1.325000 0.800000 1.845000 ;
      RECT 1.090000 0.255000 1.320000 0.585000 ;
      RECT 1.150000 0.585000 1.320000 1.875000 ;
      RECT 1.150000 1.875000 3.165000 2.045000 ;
      RECT 1.150000 2.045000 1.320000 2.465000 ;
      RECT 2.440000 2.045000 2.610000 2.465000 ;
      RECT 2.995000 0.995000 3.255000 1.325000 ;
      RECT 2.995000 1.325000 3.165000 1.875000 ;
  END
END sky130_fd_sc_hd__and4b_1

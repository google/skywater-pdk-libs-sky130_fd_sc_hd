* File: sky130_fd_sc_hd__o211ai_2.pex.spice
* Created: Tue Sep  1 19:20:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O211AI_2%C1 1 3 6 8 10 13 15 19 22
c41 8 0 3.31329e-20 $X=0.925 $Y=0.995
r42 21 22 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.925 $Y2=1.16
r43 18 21 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.495 $Y2=1.16
r44 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r45 15 19 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.53
+ $X2=0.23 $Y2=1.16
r46 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.325
+ $X2=0.925 $Y2=1.16
r47 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.325
+ $X2=0.925 $Y2=1.985
r48 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=0.995
+ $X2=0.925 $Y2=1.16
r49 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.925 $Y=0.995
+ $X2=0.925 $Y2=0.56
r50 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r51 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.985
r52 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=1.16
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%B1 1 3 6 8 10 13 15 25
c47 1 0 1.03048e-19 $X=1.355 $Y=0.995
r48 23 25 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.685 $Y=1.16
+ $X2=1.785 $Y2=1.16
r49 21 23 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.355 $Y=1.16
+ $X2=1.685 $Y2=1.16
r50 18 21 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.355 $Y2=1.16
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=1.16 $X2=1.345 $Y2=1.16
r52 15 19 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=1.61 $Y=1.22
+ $X2=1.345 $Y2=1.22
r53 15 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.685
+ $Y=1.16 $X2=1.685 $Y2=1.16
r54 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.16
r55 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.985
r56 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=0.995
+ $X2=1.785 $Y2=1.16
r57 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.785 $Y=0.995
+ $X2=1.785 $Y2=0.56
r58 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.325
+ $X2=1.355 $Y2=1.16
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.355 $Y=1.325
+ $X2=1.355 $Y2=1.985
r60 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=0.995
+ $X2=1.355 $Y2=1.16
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.355 $Y=0.995
+ $X2=1.355 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%A2 1 3 6 8 10 13 15 21 22
r43 20 22 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.17 $Y=1.16
+ $X2=3.205 $Y2=1.16
r44 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.17
+ $Y=1.16 $X2=3.17 $Y2=1.16
r45 17 20 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=2.775 $Y=1.16
+ $X2=3.17 $Y2=1.16
r46 15 21 26.3416 $w=2.78e-07 $l=6.4e-07 $layer=LI1_cond $X=2.53 $Y=1.215
+ $X2=3.17 $Y2=1.215
r47 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.325
+ $X2=3.205 $Y2=1.16
r48 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.205 $Y=1.325
+ $X2=3.205 $Y2=1.985
r49 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=0.995
+ $X2=3.205 $Y2=1.16
r50 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.205 $Y=0.995
+ $X2=3.205 $Y2=0.56
r51 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.325
+ $X2=2.775 $Y2=1.16
r52 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.775 $Y=1.325
+ $X2=2.775 $Y2=1.985
r53 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=0.995
+ $X2=2.775 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.775 $Y=0.995
+ $X2=2.775 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%A1 1 3 6 8 10 13 15 22 26
c39 26 0 1.55445e-19 $X=4.37 $Y=0.85
c40 6 0 8.33406e-20 $X=3.635 $Y=1.985
r41 21 26 13.3902 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.01 $Y=1.075
+ $X2=4.37 $Y2=1.075
r42 20 22 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.01 $Y=1.16
+ $X2=4.065 $Y2=1.16
r43 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.01
+ $Y=1.16 $X2=4.01 $Y2=1.16
r44 17 20 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.635 $Y=1.16
+ $X2=4.01 $Y2=1.16
r45 15 26 4.5877 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=4.37 $Y=0.85 $X2=4.37
+ $Y2=1.075
r46 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=1.325
+ $X2=4.065 $Y2=1.16
r47 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.065 $Y=1.325
+ $X2=4.065 $Y2=1.985
r48 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=0.995
+ $X2=4.065 $Y2=1.16
r49 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.065 $Y=0.995
+ $X2=4.065 $Y2=0.56
r50 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=1.325
+ $X2=3.635 $Y2=1.16
r51 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.635 $Y=1.325
+ $X2=3.635 $Y2=1.985
r52 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=0.995
+ $X2=3.635 $Y2=1.16
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.635 $Y=0.995
+ $X2=3.635 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%VPWR 1 2 3 4 13 15 19 23 27 29 31 36 41 51
+ 52 58 61 64
r69 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r71 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 52 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r74 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.85 $Y2=2.72
r75 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r78 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r79 45 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r82 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.165 $Y=2.72 $X2=2
+ $Y2=2.72
r83 42 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.53 $Y2=2.72
r84 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.85 $Y2=2.72
r85 41 47 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 40 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r89 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.14 $Y2=2.72
r90 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.61 $Y2=2.72
r91 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=2.72 $X2=2
+ $Y2=2.72
r92 36 39 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 35 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 32 55 4.09637 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.187 $Y2=2.72
r96 32 34 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.69 $Y2=2.72
r97 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.14 $Y2=2.72
r98 31 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.69 $Y2=2.72
r99 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r100 29 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r101 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.72
r102 25 27 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=1.95
r103 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=2.635 $X2=2
+ $Y2=2.72
r104 21 23 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2 $Y=2.635 $X2=2
+ $Y2=2
r105 17 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.72
r106 17 19 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2
r107 13 55 3.11585 $w=2.6e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.187 $Y2=2.72
r108 13 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2.34
r109 4 27 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=3.71
+ $Y=1.485 $X2=3.85 $Y2=1.95
r110 3 23 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.485 $X2=2 $Y2=2
r111 2 19 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.485 $X2=1.14 $Y2=2
r112 1 15 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%Y 1 2 3 4 15 17 21 23 28 29 31 32 35
c49 31 0 8.33406e-20 $X=2.99 $Y=1.7
r50 32 35 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.71 $Y=0.85 $X2=0.71
+ $Y2=0.76
r51 27 32 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.71 $Y=1.54
+ $X2=0.71 $Y2=0.85
r52 27 28 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.54
+ $X2=0.71 $Y2=1.625
r53 24 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.665 $Y=1.625
+ $X2=1.57 $Y2=1.625
r54 23 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=1.625
+ $X2=2.99 $Y2=1.625
r55 23 24 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.825 $Y=1.625
+ $X2=1.665 $Y2=1.625
r56 19 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=1.71
+ $X2=1.57 $Y2=1.625
r57 19 21 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.57 $Y=1.71
+ $X2=1.57 $Y2=1.845
r58 18 28 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.625
+ $X2=0.71 $Y2=1.625
r59 17 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.475 $Y=1.625
+ $X2=1.57 $Y2=1.625
r60 17 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.475 $Y=1.625
+ $X2=0.875 $Y2=1.625
r61 13 28 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.675 $Y=1.71
+ $X2=0.71 $Y2=1.625
r62 13 15 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=0.675 $Y=1.71
+ $X2=0.675 $Y2=1.82
r63 4 31 300 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=1.485 $X2=2.99 $Y2=1.7
r64 3 21 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=1.485 $X2=1.57 $Y2=1.845
r65 2 15 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.485 $X2=0.71 $Y2=1.82
r66 1 35 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%A_487_297# 1 2 3 10 16 20 23
r26 23 25 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=2.525 $Y=2.3 $X2=2.525
+ $Y2=2.38
r27 18 20 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=4.315 $Y=1.695
+ $X2=4.315 $Y2=1.96
r28 16 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.185 $Y=1.61
+ $X2=4.315 $Y2=1.695
r29 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.185 $Y=1.61
+ $X2=3.515 $Y2=1.61
r30 13 15 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=3.42 $Y=2.295
+ $X2=3.42 $Y2=1.825
r31 12 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.42 $Y=1.695
+ $X2=3.515 $Y2=1.61
r32 12 15 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=3.42 $Y=1.695
+ $X2=3.42 $Y2=1.825
r33 11 25 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.525 $Y2=2.38
r34 10 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.325 $Y=2.38
+ $X2=3.42 $Y2=2.295
r35 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.325 $Y=2.38
+ $X2=2.655 $Y2=2.38
r36 3 20 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=4.14
+ $Y=1.485 $X2=4.28 $Y2=1.96
r37 2 15 300 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=1.485 $X2=3.42 $Y2=1.825
r38 1 23 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.485 $X2=2.56 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%A_27_47# 1 2 3 10 16 20 23
c28 16 0 1.36181e-19 $X=1.14 $Y=0.705
r29 18 23 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=1.235 $Y=0.36 $X2=1.14
+ $Y2=0.36
r30 18 20 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=1.235 $Y=0.36 $X2=2
+ $Y2=0.36
r31 14 23 1.5279 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=1.14 $Y=0.465
+ $X2=1.14 $Y2=0.36
r32 14 16 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=1.14 $Y=0.465
+ $X2=1.14 $Y2=0.705
r33 10 23 4.9491 $w=2e-07 $l=9.98749e-08 $layer=LI1_cond $X=1.045 $Y=0.35
+ $X2=1.14 $Y2=0.36
r34 10 12 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=1.045 $Y=0.35
+ $X2=0.28 $Y2=0.35
r35 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2 $Y2=0.36
r36 2 23 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.36
r37 2 16 182 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.705
r38 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%A_286_47# 1 2 3 10 17
r29 17 19 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=3.85 $Y=0.68 $X2=3.85
+ $Y2=0.74
r30 12 15 74.9957 $w=2.08e-07 $l=1.42e-06 $layer=LI1_cond $X=1.57 $Y=0.74
+ $X2=2.99 $Y2=0.74
r31 10 19 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=3.755 $Y=0.74
+ $X2=3.85 $Y2=0.74
r32 10 15 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=3.755 $Y=0.74
+ $X2=2.99 $Y2=0.74
r33 3 17 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.235 $X2=3.85 $Y2=0.68
r34 2 15 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.235 $X2=2.99 $Y2=0.74
r35 1 12 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_2%VGND 1 2 3 12 16 18 20 22 24 32 37 43 46 50
c62 18 0 1.55445e-19 $X=4.28 $Y=0.085
r63 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r64 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r65 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r66 41 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r67 41 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r68 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r69 38 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r70 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.91
+ $Y2=0
r71 37 49 4.65202 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.357
+ $Y2=0
r72 37 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=3.91
+ $Y2=0
r73 36 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r74 36 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r75 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r76 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.56
+ $Y2=0
r77 33 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.99
+ $Y2=0
r78 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r79 32 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r80 31 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r81 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r82 26 30 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r83 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.56
+ $Y2=0
r84 24 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.07
+ $Y2=0
r85 22 31 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r86 22 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r87 18 49 3.11416 $w=3.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.357 $Y2=0
r88 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0.36
r89 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r90 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.36
r91 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r92 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.36
r93 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.14
+ $Y=0.235 $X2=4.28 $Y2=0.36
r94 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.235 $X2=3.42 $Y2=0.36
r95 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.56 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__nand4bb_1.spice
* Created: Thu Aug 27 14:30:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4bb_1.pex.spice"
.subckt sky130_fd_sc_hd__nand4bb_1  VNB VPB B_N D C A_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_B_N_M1011_g N_A_27_93#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0940093 AS=0.1092 PD=0.820374 PS=1.36 NRD=48.228 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1005 A_218_47# N_D_M1005_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65 AD=0.12675
+ AS=0.145491 PD=1.04 PS=1.26963 NRD=25.836 NRS=10.152 M=1 R=4.33333 SA=75000.6
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1009 A_326_47# N_C_M1009_g A_218_47# VNB NSHORT L=0.15 W=0.65 AD=0.11375
+ AS=0.12675 PD=1 PS=1.04 NRD=22.152 NRS=25.836 M=1 R=4.33333 SA=75001.1
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 A_426_47# N_A_27_93#_M1007_g A_326_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.11375 PD=1 PS=1 NRD=22.152 NRS=22.152 M=1 R=4.33333 SA=75001.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A_496_21#_M1006_g A_426_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.11375 PD=1.82 PS=1 NRD=0 NRS=22.152 M=1 R=4.33333 SA=75002.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_496_21#_M1001_d N_A_N_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1827 AS=0.1092 PD=1.71 PS=1.36 NRD=25.704 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B_N_M1003_g N_A_27_93#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.103965 AS=0.1092 PD=0.825211 PS=1.36 NRD=35.1645 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_D_M1008_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.247535 PD=1.39 PS=1.96479 NRD=10.8153 NRS=7.8603 M=1 R=6.66667 SA=75000.4
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_Y_M1008_d VPB PHIGHVT L=0.15 W=1 AD=0.175
+ AS=0.195 PD=1.35 PS=1.39 NRD=6.8753 NRS=10.8153 M=1 R=6.66667 SA=75001
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_A_27_93#_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=6.8753 NRS=6.8753 M=1 R=6.66667
+ SA=75001.5 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_496_21#_M1004_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.175 PD=2.52 PS=1.35 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75002
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1010 N_A_496_21#_M1010_d N_A_N_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1827 AS=0.1092 PD=1.71 PS=1.36 NRD=42.1974 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.4 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__nand4bb_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__probe_p_8.pex.spice
* Created: Tue Sep  1 19:29:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__PROBE_P_8%A 3 7 11 15 17 19 23 25 26 27
c77 27 0 1.27947e-19 $X=1.155 $Y=1.19
r78 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.16 $X2=0.985 $Y2=1.16
r79 32 34 28.8152 $w=2.76e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.16
+ $X2=0.47 $Y2=1.16
r80 27 38 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=0.985 $Y2=1.175
r81 26 38 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.985 $Y2=1.175
r82 25 26 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r83 25 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r84 17 37 56.7572 $w=2.76e-07 $l=3.25e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=0.985 $Y2=1.16
r85 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r86 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r87 9 37 16.5906 $w=2.76e-07 $l=9.5e-08 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.985 $Y2=1.16
r88 9 34 73.3478 $w=2.76e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.47 $Y2=1.16
r89 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r90 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r91 5 34 17.0164 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r92 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r93 1 34 17.0164 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r94 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__PROBE_P_8%A_27_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 85 87 88 89 90 93 99 101 104 106 112 116 118 119
+ 130
c296 130 0 1.27947e-19 $X=4.67 $Y=1.16
c297 67 0 1.42997e-20 $X=4.25 $Y=1.985
c298 43 0 1.88697e-19 $X=2.99 $Y=1.985
c299 39 0 1.3987e-19 $X=2.99 $Y=0.56
r300 129 130 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.67 $Y2=1.16
r301 126 127 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.83 $Y2=1.16
r302 125 126 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.41 $Y2=1.16
r303 124 125 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r304 123 124 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r305 113 129 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=3.88 $Y=1.16
+ $X2=4.25 $Y2=1.16
r306 113 127 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=3.88 $Y=1.16
+ $X2=3.83 $Y2=1.16
r307 112 113 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r308 110 123 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=2.15 $Y2=1.16
r309 110 120 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=1.73 $Y2=1.16
r310 109 112 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.84 $Y=1.16
+ $X2=3.88 $Y2=1.16
r311 109 110 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.84
+ $Y=1.16 $X2=1.84 $Y2=1.16
r312 107 119 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.507 $Y2=1.16
r313 107 109 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.84 $Y2=1.16
r314 106 116 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.445
+ $X2=1.507 $Y2=1.53
r315 105 119 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.16
r316 105 106 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.445
r317 104 119 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.075
+ $X2=1.507 $Y2=1.16
r318 103 104 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.507 $Y=0.905
+ $X2=1.507 $Y2=1.075
r319 102 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.82
+ $X2=1.1 $Y2=0.82
r320 101 103 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.42 $Y=0.82
+ $X2=1.507 $Y2=0.905
r321 101 102 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.42 $Y=0.82
+ $X2=1.185 $Y2=0.82
r322 97 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.82
r323 97 99 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.56
r324 93 95 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.1 $Y=1.63 $X2=1.1
+ $Y2=2.31
r325 91 116 26.5529 $w=1.68e-07 $l=4.07e-07 $layer=LI1_cond $X=1.1 $Y=1.53
+ $X2=1.507 $Y2=1.53
r326 91 93 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.1 $Y=1.615
+ $X2=1.1 $Y2=1.63
r327 89 91 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.53
+ $X2=1.1 $Y2=1.53
r328 89 90 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=1.53
+ $X2=0.425 $Y2=1.53
r329 87 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.82
+ $X2=1.1 $Y2=0.82
r330 87 88 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.82
+ $X2=0.345 $Y2=0.82
r331 83 88 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.345 $Y2=0.82
r332 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.56
r333 79 81 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r334 77 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r335 77 79 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r336 73 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.16
r337 73 75 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.985
r338 69 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=1.16
r339 69 71 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=0.56
r340 65 129 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.16
r341 65 67 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.985
r342 61 129 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=1.16
r343 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
r344 57 127 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.16
r345 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.985
r346 53 127 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.16
r347 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
r348 49 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r349 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r350 45 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r351 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r352 41 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r353 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r354 37 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r355 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r356 33 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r357 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r358 29 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r359 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r360 25 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r361 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r362 21 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r363 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r364 17 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r365 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r366 13 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r367 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r368 4 95 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.31
r369 4 93 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.63
r370 3 81 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r371 3 79 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r372 2 99 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.56
r373 1 85 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__PROBE_P_8%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 43 48
+ 49 51 52 54 55 56 57 58 60 76 83 84 87 90
c118 43 0 2.19555e-19 $X=4.88 $Y=1.66
c119 39 0 1.93771e-19 $X=4.04 $Y=2
r120 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r122 84 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r124 81 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=4.88 $Y2=2.72
r125 81 83 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=5.29 $Y2=2.72
r126 80 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r127 80 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r128 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r129 77 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.72
+ $X2=4.04 $Y2=2.72
r130 77 79 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.72
+ $X2=4.37 $Y2=2.72
r131 76 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.88 $Y2=2.72
r132 76 79 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 75 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r134 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r135 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r136 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r137 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r138 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 60 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 58 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r141 56 74 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.99 $Y2=2.72
r142 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.2 $Y2=2.72
r143 54 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r144 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.36 $Y2=2.72
r145 53 74 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.99 $Y2=2.72
r146 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.36 $Y2=2.72
r147 51 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.52 $Y2=2.72
r149 50 71 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=2.07 $Y2=2.72
r150 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.52 $Y2=2.72
r151 48 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r153 47 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=1.15 $Y2=2.72
r154 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r155 43 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.88 $Y=1.66
+ $X2=4.88 $Y2=2.34
r156 41 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2.72
r157 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2.34
r158 37 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.635
+ $X2=4.04 $Y2=2.72
r159 37 39 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.04 $Y=2.635
+ $X2=4.04 $Y2=2
r160 36 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.72
+ $X2=3.2 $Y2=2.72
r161 35 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.72
+ $X2=4.04 $Y2=2.72
r162 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=2.72
+ $X2=3.365 $Y2=2.72
r163 31 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635 $X2=3.2
+ $Y2=2.72
r164 31 33 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2
r165 27 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r166 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2
r167 23 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r168 23 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2
r169 19 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r170 19 21 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2
r171 6 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2.34
r172 6 43 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.66
r173 5 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=2
r174 4 33 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2
r175 3 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2
r176 2 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
r177 1 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__PROBE_P_8%noxref_6 1 2 3 4 5 6 7 8 27 31 33 34 35 36
+ 39 43 45 47 51 55 57 59 62 65 69 71 72 73 74 75 76 80 82 83 85 87 88 91 93 100
c262 100 0 1.3987e-19 $X=3.945 $Y=1.19
c263 88 0 3.16339e-19 $X=3.56 $Y=1.27
c264 87 0 9.69875e-20 $X=3.56 $Y=1.27
c265 85 0 1.88697e-19 $X=3.975 $Y=1.19
c266 83 0 1.42997e-20 $X=4.765 $Y=1.19
r267 99 100 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=3.945 $Y=1.19
+ $X2=3.945 $Y2=1.19
r268 91 100 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=3.985 $Y=1.19
+ $X2=3.985 $Y2=1.19
r269 88 93 0.00650012 $w=3.02e-06 $l=6.75e-07 $layer=MET5_cond $X=2.76 $Y=1.27
+ $X2=2.76 $Y2=1.945
r270 87 91 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=3.985 $Y=1.19
+ $X2=3.985 $Y2=1.19
r271 87 88 0.19 $w=8e-07 $l=1.6e-06 $layer=via4_notcap2m $count=2 $X=3.56
+ $Y=1.27 $X2=3.56 $Y2=1.27
r272 85 99 0.0170272 $w=2.6e-07 $l=3e-08 $layer=MET1_cond $X=3.975 $Y=1.19
+ $X2=3.945 $Y2=1.19
r273 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.765 $Y=1.19
+ $X2=4.765 $Y2=1.19
r274 80 85 0.0749482 $w=2.6e-07 $l=1.3e-07 $layer=MET1_cond $X=4.105 $Y=1.19
+ $X2=3.975 $Y2=1.19
r275 80 82 0.423459 $w=2.3e-07 $l=6.6e-07 $layer=MET1_cond $X=4.105 $Y=1.19
+ $X2=4.765 $Y2=1.19
r276 77 83 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=4.545 $Y=1.185
+ $X2=4.765 $Y2=1.185
r277 76 77 0.597719 $w=2.6e-07 $l=1.28e-07 $layer=LI1_cond $X=4.417 $Y=1.185
+ $X2=4.545 $Y2=1.185
r278 69 79 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.46 $Y=1.755
+ $X2=4.46 $Y2=1.615
r279 63 75 4.27425 $w=2.12e-07 $l=1.04307e-07 $layer=LI1_cond $X=4.46 $Y=0.735
+ $X2=4.417 $Y2=0.82
r280 63 65 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.46 $Y=0.735
+ $X2=4.46 $Y2=0.56
r281 62 76 5.8752 $w=2.53e-07 $l=1.3e-07 $layer=LI1_cond $X=4.417 $Y=1.055
+ $X2=4.417 $Y2=1.185
r282 61 75 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=4.417 $Y=0.905
+ $X2=4.417 $Y2=0.82
r283 61 62 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=4.417 $Y=0.905
+ $X2=4.417 $Y2=1.055
r284 60 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=1.53
+ $X2=3.62 $Y2=1.53
r285 59 79 5.12497 $w=2.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.417 $Y=1.53
+ $X2=4.417 $Y2=1.615
r286 59 76 15.5919 $w=2.53e-07 $l=3.45e-07 $layer=LI1_cond $X=4.417 $Y=1.53
+ $X2=4.417 $Y2=1.185
r287 59 60 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.29 $Y=1.53
+ $X2=3.705 $Y2=1.53
r288 58 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0.82
+ $X2=3.62 $Y2=0.82
r289 57 75 2.15711 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.29 $Y=0.82
+ $X2=4.417 $Y2=0.82
r290 57 58 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.29 $Y=0.82
+ $X2=3.705 $Y2=0.82
r291 53 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.615
+ $X2=3.62 $Y2=1.53
r292 53 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.62 $Y=1.615
+ $X2=3.62 $Y2=1.755
r293 49 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.82
r294 49 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.56
r295 48 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.53
+ $X2=2.78 $Y2=1.53
r296 47 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=1.53
+ $X2=3.62 $Y2=1.53
r297 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=1.53
+ $X2=2.865 $Y2=1.53
r298 46 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=2.78 $Y2=0.82
r299 45 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.82
+ $X2=3.62 $Y2=0.82
r300 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=0.82
+ $X2=2.865 $Y2=0.82
r301 41 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=1.615
+ $X2=2.78 $Y2=1.53
r302 41 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=1.615
+ $X2=2.78 $Y2=1.755
r303 37 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.82
r304 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.56
r305 35 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=1.53
+ $X2=2.78 $Y2=1.53
r306 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=1.53
+ $X2=2.025 $Y2=1.53
r307 33 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.82
+ $X2=2.78 $Y2=0.82
r308 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=0.82
+ $X2=2.025 $Y2=0.82
r309 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=2.025 $Y2=1.53
r310 29 31 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=1.94 $Y2=1.755
r311 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=2.025 $Y2=0.82
r312 25 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.56
r313 8 69 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=1.755
r314 7 55 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.755
r315 6 43 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.755
r316 5 31 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.755
r317 4 65 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.56
r318 3 51 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.56
r319 2 39 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.56
r320 1 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__PROBE_P_8%VGND 1 2 3 4 5 6 21 25 29 33 35 39 43 46
+ 47 49 50 51 52 53 55 57 62 74 81 82 85 88 91
r134 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r135 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r136 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r137 82 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r138 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r139 79 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=4.88
+ $Y2=0
r140 79 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.29
+ $Y2=0
r141 78 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r142 78 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r143 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r144 75 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0 $X2=4.04
+ $Y2=0
r145 75 77 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0
+ $X2=4.37 $Y2=0
r146 74 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.88
+ $Y2=0
r147 74 77 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.37
+ $Y2=0
r148 73 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r149 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r150 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r151 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r152 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r153 67 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r154 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r155 64 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r156 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r157 57 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r158 55 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r159 55 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r160 53 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=0
+ $X2=0.515 $Y2=0
r161 53 62 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r162 51 72 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.99
+ $Y2=0
r163 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.2
+ $Y2=0
r164 49 69 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=0
+ $X2=2.07 $Y2=0
r165 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.36
+ $Y2=0
r166 48 72 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=2.99 $Y2=0
r167 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.36
+ $Y2=0
r168 46 66 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.15 $Y2=0
r169 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r170 45 69 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=0
+ $X2=2.07 $Y2=0
r171 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r172 41 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r173 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.38
r174 37 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r175 37 39 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.4
r176 36 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.2
+ $Y2=0
r177 35 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.04
+ $Y2=0
r178 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=0
+ $X2=3.365 $Y2=0
r179 31 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.085 $X2=3.2
+ $Y2=0
r180 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0.4
r181 27 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r182 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.4
r183 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r184 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r185 19 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r186 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r187 6 43 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.38
r188 5 39 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.4
r189 4 33 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.4
r190 3 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.4
r191 2 25 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r192 1 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__PROBE_P_8%X 1 3
r23 1 3 0.00103039 $w=3.02e-06 $l=1.07e-07 $layer=MET5_cond $X=2.76 $Y=2.057
+ $X2=2.76 $Y2=1.95
.ends


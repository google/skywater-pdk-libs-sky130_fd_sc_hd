* File: sky130_fd_sc_hd__clkinv_16.spice.pex
* Created: Thu Aug 27 14:12:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINV_16%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55
+ 59 63 67 71 73 74 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 153 157 161 163 165 170 171 172 174 212 213
r306 211 213 16.8304 $w=3.6e-07 $l=1.05e-07 $layer=POLY_cond $X=10.46 $Y=1.17
+ $X2=10.565 $Y2=1.17
r307 211 212 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.46
+ $Y=1.16 $X2=10.46 $Y2=1.16
r308 209 211 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=10.135 $Y=1.17
+ $X2=10.46 $Y2=1.17
r309 208 209 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=9.705 $Y=1.17
+ $X2=10.135 $Y2=1.17
r310 207 208 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=9.275 $Y=1.17
+ $X2=9.705 $Y2=1.17
r311 205 207 28.0507 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=9.1 $Y=1.17
+ $X2=9.275 $Y2=1.17
r312 205 206 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.1
+ $Y=1.16 $X2=9.1 $Y2=1.16
r313 203 205 40.8738 $w=3.6e-07 $l=2.55e-07 $layer=POLY_cond $X=8.845 $Y=1.17
+ $X2=9.1 $Y2=1.17
r314 202 203 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=8.415 $Y=1.17
+ $X2=8.845 $Y2=1.17
r315 201 202 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=7.985 $Y=1.17
+ $X2=8.415 $Y2=1.17
r316 200 201 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=7.555 $Y=1.17
+ $X2=7.985 $Y2=1.17
r317 199 200 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=7.125 $Y=1.17
+ $X2=7.555 $Y2=1.17
r318 198 199 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=6.695 $Y=1.17
+ $X2=7.125 $Y2=1.17
r319 197 198 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=6.265 $Y=1.17
+ $X2=6.695 $Y2=1.17
r320 196 197 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=5.835 $Y=1.17
+ $X2=6.265 $Y2=1.17
r321 195 196 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=5.405 $Y=1.17
+ $X2=5.835 $Y2=1.17
r322 193 194 74.5346 $w=3.6e-07 $l=4.65e-07 $layer=POLY_cond $X=4.355 $Y=1.17
+ $X2=4.82 $Y2=1.17
r323 192 193 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=3.925 $Y=1.17
+ $X2=4.355 $Y2=1.17
r324 191 192 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=3.495 $Y=1.17
+ $X2=3.925 $Y2=1.17
r325 190 191 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=3.065 $Y=1.17
+ $X2=3.495 $Y2=1.17
r326 189 190 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=2.635 $Y=1.17
+ $X2=3.065 $Y2=1.17
r327 188 189 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=2.205 $Y=1.17
+ $X2=2.635 $Y2=1.17
r328 186 188 40.8738 $w=3.6e-07 $l=2.55e-07 $layer=POLY_cond $X=1.95 $Y=1.17
+ $X2=2.205 $Y2=1.17
r329 184 186 28.0507 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=1.775 $Y=1.17
+ $X2=1.95 $Y2=1.17
r330 183 184 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=1.345 $Y=1.17
+ $X2=1.775 $Y2=1.17
r331 182 183 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=0.915 $Y=1.17
+ $X2=1.345 $Y2=1.17
r332 180 182 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=0.59 $Y=1.17
+ $X2=0.915 $Y2=1.17
r333 180 181 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r334 177 180 16.8304 $w=3.6e-07 $l=1.05e-07 $layer=POLY_cond $X=0.485 $Y=1.17
+ $X2=0.59 $Y2=1.17
r335 175 212 17.2866 $w=3.78e-07 $l=5.7e-07 $layer=LI1_cond $X=9.89 $Y=1.085
+ $X2=10.46 $Y2=1.085
r336 175 206 23.9587 $w=3.78e-07 $l=7.9e-07 $layer=LI1_cond $X=9.89 $Y=1.085
+ $X2=9.1 $Y2=1.085
r337 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=1.19
+ $X2=9.89 $Y2=1.19
r338 172 174 0.314386 $w=2.3e-07 $l=4.9e-07 $layer=MET1_cond $X=9.4 $Y=1.19
+ $X2=9.89 $Y2=1.19
r339 170 172 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.285 $Y=1.19
+ $X2=9.4 $Y2=1.19
r340 170 171 8.74998 $w=1.4e-07 $l=7.07e-06 $layer=MET1_cond $X=9.285 $Y=1.19
+ $X2=2.215 $Y2=1.19
r341 165 171 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=2.1 $Y=1.19
+ $X2=2.215 $Y2=1.19
r342 165 167 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=2.1 $Y=1.19
+ $X2=2.07 $Y2=1.19
r343 163 181 41.2453 $w=3.78e-07 $l=1.36e-06 $layer=LI1_cond $X=1.95 $Y=1.085
+ $X2=0.59 $Y2=1.085
r344 163 186 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r345 163 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.19
r346 159 213 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=10.565 $Y=1.35
+ $X2=10.565 $Y2=1.17
r347 159 161 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.565 $Y=1.35
+ $X2=10.565 $Y2=1.985
r348 155 209 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=10.135 $Y=1.35
+ $X2=10.135 $Y2=1.17
r349 155 157 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.135 $Y=1.35
+ $X2=10.135 $Y2=1.985
r350 151 208 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=9.705 $Y=1.35
+ $X2=9.705 $Y2=1.17
r351 151 153 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.705 $Y=1.35
+ $X2=9.705 $Y2=1.985
r352 147 207 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=9.275 $Y=1.35
+ $X2=9.275 $Y2=1.17
r353 147 149 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.275 $Y=1.35
+ $X2=9.275 $Y2=1.985
r354 143 203 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.845 $Y=1.35
+ $X2=8.845 $Y2=1.17
r355 143 145 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.845 $Y=1.35
+ $X2=8.845 $Y2=1.985
r356 139 203 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.845 $Y=0.99
+ $X2=8.845 $Y2=1.17
r357 139 141 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=8.845 $Y=0.99
+ $X2=8.845 $Y2=0.445
r358 135 202 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.415 $Y=1.35
+ $X2=8.415 $Y2=1.17
r359 135 137 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.415 $Y=1.35
+ $X2=8.415 $Y2=1.985
r360 131 202 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.415 $Y=0.99
+ $X2=8.415 $Y2=1.17
r361 131 133 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=8.415 $Y=0.99
+ $X2=8.415 $Y2=0.445
r362 127 201 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.985 $Y=1.35
+ $X2=7.985 $Y2=1.17
r363 127 129 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.985 $Y=1.35
+ $X2=7.985 $Y2=1.985
r364 123 201 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.985 $Y=0.99
+ $X2=7.985 $Y2=1.17
r365 123 125 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.985 $Y=0.99
+ $X2=7.985 $Y2=0.445
r366 119 200 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=1.17
r367 119 121 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=1.985
r368 115 200 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.555 $Y=0.99
+ $X2=7.555 $Y2=1.17
r369 115 117 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.555 $Y=0.99
+ $X2=7.555 $Y2=0.445
r370 111 199 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=1.17
r371 111 113 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=1.985
r372 107 199 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.125 $Y=0.99
+ $X2=7.125 $Y2=1.17
r373 107 109 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.125 $Y=0.99
+ $X2=7.125 $Y2=0.445
r374 103 198 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.17
r375 103 105 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.985
r376 99 198 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.695 $Y=0.99
+ $X2=6.695 $Y2=1.17
r377 99 101 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.695 $Y=0.99
+ $X2=6.695 $Y2=0.445
r378 95 197 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.17
r379 95 97 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.985
r380 91 197 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.265 $Y=0.99
+ $X2=6.265 $Y2=1.17
r381 91 93 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.265 $Y=0.99
+ $X2=6.265 $Y2=0.445
r382 87 196 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.17
r383 87 89 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.985
r384 83 196 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.835 $Y=0.99
+ $X2=5.835 $Y2=1.17
r385 83 85 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.835 $Y=0.99
+ $X2=5.835 $Y2=0.445
r386 79 195 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.17
r387 79 81 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.985
r388 75 195 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.405 $Y=0.99
+ $X2=5.405 $Y2=1.17
r389 75 77 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.405 $Y=0.99
+ $X2=5.405 $Y2=0.445
r390 74 194 12.0217 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=4.895 $Y=1.17
+ $X2=4.82 $Y2=1.17
r391 73 195 12.0217 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.17
+ $X2=5.405 $Y2=1.17
r392 73 74 69.7259 $w=3.6e-07 $l=4.35e-07 $layer=POLY_cond $X=5.33 $Y=1.17
+ $X2=4.895 $Y2=1.17
r393 69 194 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.82 $Y=1.35
+ $X2=4.82 $Y2=1.17
r394 69 71 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.82 $Y=1.35
+ $X2=4.82 $Y2=1.985
r395 65 194 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.82 $Y=0.99
+ $X2=4.82 $Y2=1.17
r396 65 67 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.82 $Y=0.99
+ $X2=4.82 $Y2=0.445
r397 61 193 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.355 $Y2=1.17
r398 61 63 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.355 $Y2=1.985
r399 57 193 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.355 $Y=0.99
+ $X2=4.355 $Y2=1.17
r400 57 59 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.355 $Y=0.99
+ $X2=4.355 $Y2=0.445
r401 53 192 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=1.17
r402 53 55 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=1.985
r403 49 192 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.925 $Y=0.99
+ $X2=3.925 $Y2=1.17
r404 49 51 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.925 $Y=0.99
+ $X2=3.925 $Y2=0.445
r405 45 191 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=1.17
r406 45 47 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=1.985
r407 41 191 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.495 $Y=0.99
+ $X2=3.495 $Y2=1.17
r408 41 43 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.495 $Y=0.99
+ $X2=3.495 $Y2=0.445
r409 37 190 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=1.17
r410 37 39 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=1.985
r411 33 190 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.065 $Y=0.99
+ $X2=3.065 $Y2=1.17
r412 33 35 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.065 $Y=0.99
+ $X2=3.065 $Y2=0.445
r413 29 189 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=1.17
r414 29 31 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=1.985
r415 25 189 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.635 $Y=0.99
+ $X2=2.635 $Y2=1.17
r416 25 27 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.635 $Y=0.99
+ $X2=2.635 $Y2=0.445
r417 21 188 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=1.17
r418 21 23 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=1.985
r419 17 188 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.205 $Y=0.99
+ $X2=2.205 $Y2=1.17
r420 17 19 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.205 $Y=0.99
+ $X2=2.205 $Y2=0.445
r421 13 184 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.775 $Y=1.35
+ $X2=1.775 $Y2=1.17
r422 13 15 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.775 $Y=1.35
+ $X2=1.775 $Y2=1.985
r423 9 183 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.345 $Y=1.35
+ $X2=1.345 $Y2=1.17
r424 9 11 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.345 $Y=1.35
+ $X2=1.345 $Y2=1.985
r425 5 182 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.915 $Y=1.35
+ $X2=0.915 $Y2=1.17
r426 5 7 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.915 $Y=1.35
+ $X2=0.915 $Y2=1.985
r427 1 177 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.485 $Y=1.35
+ $X2=0.485 $Y2=1.17
r428 1 3 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.485 $Y=1.35
+ $X2=0.485 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42
+ 48 52 56 60 64 68 73 76 80 84 86 90 94 96 98 101 102 104 105 107 108 110 111
+ 114 115 117 118 120 121 122 123 124 126 156 161 170 173 176 180
r172 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r173 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r174 173 174 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r175 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r176 165 180 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r177 165 177 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.89 $Y2=2.72
r178 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r179 162 176 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.05 $Y=2.72
+ $X2=9.922 $Y2=2.72
r180 162 164 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.05 $Y=2.72
+ $X2=10.35 $Y2=2.72
r181 161 179 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=10.65 $Y=2.72
+ $X2=10.845 $Y2=2.72
r182 161 164 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.65 $Y=2.72
+ $X2=10.35 $Y2=2.72
r183 160 177 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r184 160 174 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r185 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r186 157 173 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.19 $Y=2.72
+ $X2=9.062 $Y2=2.72
r187 157 159 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.19 $Y=2.72
+ $X2=9.43 $Y2=2.72
r188 156 176 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=9.922 $Y2=2.72
r189 156 159 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=9.43 $Y2=2.72
r190 155 174 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r191 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r192 152 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r193 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r194 149 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r195 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r196 146 149 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r197 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r198 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r199 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r200 140 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r201 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r202 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r203 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r204 134 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r205 134 171 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r206 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r207 131 170 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.26 $Y=2.72
+ $X2=1.13 $Y2=2.72
r208 131 133 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.26 $Y=2.72
+ $X2=1.61 $Y2=2.72
r209 130 171 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r210 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r211 127 167 4.10994 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r212 127 129 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.69 $Y2=2.72
r213 126 170 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=1.13
+ $Y2=2.72
r214 126 129 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1 $Y=2.72
+ $X2=0.69 $Y2=2.72
r215 124 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r216 124 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r217 122 154 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.075 $Y=2.72
+ $X2=8.05 $Y2=2.72
r218 122 123 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.075 $Y=2.72
+ $X2=8.202 $Y2=2.72
r219 120 151 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=2.72
+ $X2=7.13 $Y2=2.72
r220 120 121 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.215 $Y=2.72
+ $X2=7.342 $Y2=2.72
r221 119 154 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.47 $Y=2.72
+ $X2=8.05 $Y2=2.72
r222 119 121 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.47 $Y=2.72
+ $X2=7.342 $Y2=2.72
r223 117 148 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.355 $Y=2.72
+ $X2=6.21 $Y2=2.72
r224 117 118 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=6.355 $Y=2.72
+ $X2=6.482 $Y2=2.72
r225 116 151 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.61 $Y=2.72
+ $X2=7.13 $Y2=2.72
r226 116 118 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=6.61 $Y=2.72
+ $X2=6.482 $Y2=2.72
r227 114 145 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.29 $Y2=2.72
r228 114 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.62 $Y2=2.72
r229 113 148 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r230 113 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=5.62 $Y2=2.72
r231 110 142 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.465 $Y=2.72
+ $X2=4.37 $Y2=2.72
r232 110 111 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.465 $Y=2.72
+ $X2=4.592 $Y2=2.72
r233 109 145 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=5.29 $Y2=2.72
r234 109 111 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.592 $Y2=2.72
r235 107 139 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.45 $Y2=2.72
r236 107 108 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.712 $Y2=2.72
r237 106 142 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.84 $Y=2.72
+ $X2=4.37 $Y2=2.72
r238 106 108 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.84 $Y=2.72
+ $X2=3.712 $Y2=2.72
r239 104 136 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.72 $Y=2.72
+ $X2=2.53 $Y2=2.72
r240 104 105 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.72 $Y=2.72
+ $X2=2.85 $Y2=2.72
r241 103 139 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=3.45 $Y2=2.72
r242 103 105 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=2.85 $Y2=2.72
r243 101 133 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=1.61 $Y2=2.72
r244 101 102 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=1.992 $Y2=2.72
r245 100 136 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.12 $Y=2.72
+ $X2=2.53 $Y2=2.72
r246 100 102 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.12 $Y=2.72
+ $X2=1.992 $Y2=2.72
r247 96 179 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=10.78 $Y=2.635
+ $X2=10.845 $Y2=2.72
r248 96 98 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=10.78 $Y=2.635
+ $X2=10.78 $Y2=2
r249 92 176 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.922 $Y=2.635
+ $X2=9.922 $Y2=2.72
r250 92 94 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=9.922 $Y=2.635
+ $X2=9.922 $Y2=2
r251 88 173 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.062 $Y=2.635
+ $X2=9.062 $Y2=2.72
r252 88 90 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=9.062 $Y=2.635
+ $X2=9.062 $Y2=2
r253 87 123 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.33 $Y=2.72
+ $X2=8.202 $Y2=2.72
r254 86 173 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.935 $Y=2.72
+ $X2=9.062 $Y2=2.72
r255 86 87 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.935 $Y=2.72
+ $X2=8.33 $Y2=2.72
r256 82 123 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.202 $Y=2.635
+ $X2=8.202 $Y2=2.72
r257 82 84 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=8.202 $Y=2.635
+ $X2=8.202 $Y2=2
r258 78 121 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.342 $Y=2.635
+ $X2=7.342 $Y2=2.72
r259 78 80 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=7.342 $Y=2.635
+ $X2=7.342 $Y2=2
r260 74 118 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=6.482 $Y=2.635
+ $X2=6.482 $Y2=2.72
r261 74 76 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=6.482 $Y=2.635
+ $X2=6.482 $Y2=2
r262 71 115 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.62 $Y=2.635
+ $X2=5.62 $Y2=2.72
r263 71 73 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.62 $Y=2.635
+ $X2=5.62 $Y2=2.34
r264 70 112 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.62 $Y=2.25
+ $X2=5.62 $Y2=2.12
r265 70 73 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=5.62 $Y=2.25 $X2=5.62
+ $Y2=2.34
r266 68 112 5.42326 $w=2.53e-07 $l=1.2e-07 $layer=LI1_cond $X=5.617 $Y=2
+ $X2=5.617 $Y2=2.12
r267 62 111 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.592 $Y=2.635
+ $X2=4.592 $Y2=2.72
r268 62 64 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=4.592 $Y=2.635
+ $X2=4.592 $Y2=2
r269 58 108 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.712 $Y=2.635
+ $X2=3.712 $Y2=2.72
r270 58 60 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=3.712 $Y=2.635
+ $X2=3.712 $Y2=2
r271 54 105 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=2.635
+ $X2=2.85 $Y2=2.72
r272 54 56 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=2.85 $Y=2.635
+ $X2=2.85 $Y2=2
r273 50 102 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.992 $Y=2.635
+ $X2=1.992 $Y2=2.72
r274 50 52 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=1.992 $Y=2.635
+ $X2=1.992 $Y2=2
r275 46 170 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2.72
r276 46 48 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2
r277 42 45 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=0.272 $Y=1.66
+ $X2=0.272 $Y2=2.34
r278 40 167 3.13813 $w=2.65e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.272 $Y=2.635
+ $X2=0.202 $Y2=2.72
r279 40 45 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.272 $Y=2.635
+ $X2=0.272 $Y2=2.34
r280 13 98 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=10.64
+ $Y=1.485 $X2=10.775 $Y2=2
r281 12 94 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=9.78
+ $Y=1.485 $X2=9.92 $Y2=2
r282 11 90 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=8.92
+ $Y=1.485 $X2=9.06 $Y2=2
r283 10 84 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=8.06
+ $Y=1.485 $X2=8.2 $Y2=2
r284 9 80 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=7.2
+ $Y=1.485 $X2=7.34 $Y2=2
r285 8 76 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=6.34
+ $Y=1.485 $X2=6.48 $Y2=2
r286 7 73 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.48
+ $Y=1.485 $X2=5.615 $Y2=2.34
r287 7 68 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=5.48
+ $Y=1.485 $X2=5.615 $Y2=2
r288 6 64 300 $w=1.7e-07 $l=5.89597e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.485 $X2=4.59 $Y2=2
r289 5 60 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=3.57
+ $Y=1.485 $X2=3.71 $Y2=2
r290 4 56 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=1.485 $X2=2.85 $Y2=2
r291 3 52 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1.85
+ $Y=1.485 $X2=1.99 $Y2=2
r292 2 48 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=0.99
+ $Y=1.485 $X2=1.13 $Y2=2
r293 1 45 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.34
r294 1 42 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 61 63 65 69 73 77 81 85 89 93 97 103 107 111 115 119 123 127 131
+ 135 142 144 146 148 149 151 153 155 157 159 161 162 167
r232 165 167 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=5.28 $Y=1.54
+ $X2=5.29 $Y2=1.54
r233 162 165 4.25218 $w=2.5e-07 $l=1.88e-07 $layer=LI1_cond $X=5.092 $Y=1.54
+ $X2=5.28 $Y2=1.54
r234 162 167 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=5.327 $Y=1.54
+ $X2=5.29 $Y2=1.54
r235 149 162 27.5664 $w=2.48e-07 $l=5.98e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=5.327 $Y2=1.54
r236 149 151 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=6.05 $Y2=1.54
r237 136 159 5.7647 $w=2.1e-07 $l=1.2e-07 $layer=LI1_cond $X=9.605 $Y=1.56
+ $X2=9.485 $Y2=1.56
r238 135 161 3.77708 $w=2.1e-07 $l=1.27e-07 $layer=LI1_cond $X=10.225 $Y=1.56
+ $X2=10.352 $Y2=1.56
r239 135 136 32.7446 $w=2.08e-07 $l=6.2e-07 $layer=LI1_cond $X=10.225 $Y=1.56
+ $X2=9.605 $Y2=1.56
r240 132 157 3.30809 $w=2.1e-07 $l=1.34629e-07 $layer=LI1_cond $X=8.755 $Y=1.56
+ $X2=8.63 $Y2=1.54
r241 131 159 5.7647 $w=2.1e-07 $l=1.2e-07 $layer=LI1_cond $X=9.365 $Y=1.56
+ $X2=9.485 $Y2=1.56
r242 131 132 32.2164 $w=2.08e-07 $l=6.1e-07 $layer=LI1_cond $X=9.365 $Y=1.56
+ $X2=8.755 $Y2=1.56
r243 125 157 2.79962 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.63 $Y=1.415
+ $X2=8.63 $Y2=1.54
r244 125 127 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=8.63 $Y=1.415
+ $X2=8.63 $Y2=0.445
r245 124 155 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.895 $Y=1.54
+ $X2=7.77 $Y2=1.54
r246 123 157 3.30809 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.505 $Y=1.54
+ $X2=8.63 $Y2=1.54
r247 123 124 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=8.505 $Y=1.54
+ $X2=7.895 $Y2=1.54
r248 117 155 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.77 $Y=1.415
+ $X2=7.77 $Y2=1.54
r249 117 119 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=7.77 $Y=1.415
+ $X2=7.77 $Y2=0.445
r250 116 153 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.035 $Y=1.54
+ $X2=6.91 $Y2=1.54
r251 115 155 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.645 $Y=1.54
+ $X2=7.77 $Y2=1.54
r252 115 116 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.645 $Y=1.54
+ $X2=7.035 $Y2=1.54
r253 109 153 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.91 $Y=1.415
+ $X2=6.91 $Y2=1.54
r254 109 111 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=6.91 $Y=1.415
+ $X2=6.91 $Y2=0.445
r255 108 151 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.175 $Y=1.54
+ $X2=6.05 $Y2=1.54
r256 107 153 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=6.91 $Y2=1.54
r257 107 108 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=6.175 $Y2=1.54
r258 101 151 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.05 $Y=1.415
+ $X2=6.05 $Y2=1.54
r259 101 103 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=6.05 $Y=1.415
+ $X2=6.05 $Y2=0.445
r260 95 162 1.99954 $w=3.5e-07 $l=1.30863e-07 $layer=LI1_cond $X=5.08 $Y=1.415
+ $X2=5.092 $Y2=1.54
r261 95 97 31.9391 $w=3.48e-07 $l=9.7e-07 $layer=LI1_cond $X=5.08 $Y=1.415
+ $X2=5.08 $Y2=0.445
r262 94 148 5.856 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.255 $Y=1.54
+ $X2=4.135 $Y2=1.54
r263 93 162 4.25218 $w=2.5e-07 $l=1.87e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=5.092 $Y2=1.54
r264 93 94 29.9635 $w=2.48e-07 $l=6.5e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=4.255 $Y2=1.54
r265 87 148 6.35417 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=4.135 $Y=1.415
+ $X2=4.135 $Y2=1.54
r266 87 89 46.5779 $w=2.38e-07 $l=9.7e-07 $layer=LI1_cond $X=4.135 $Y=1.415
+ $X2=4.135 $Y2=0.445
r267 86 146 6.1976 $w=2.5e-07 $l=1.28e-07 $layer=LI1_cond $X=3.41 $Y=1.54
+ $X2=3.282 $Y2=1.54
r268 85 148 5.856 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.015 $Y=1.54
+ $X2=4.135 $Y2=1.54
r269 85 86 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=4.015 $Y=1.54
+ $X2=3.41 $Y2=1.54
r270 79 146 5.98039 $w=2.55e-07 $l=1.25e-07 $layer=LI1_cond $X=3.282 $Y=1.415
+ $X2=3.282 $Y2=1.54
r271 79 81 43.838 $w=2.53e-07 $l=9.7e-07 $layer=LI1_cond $X=3.282 $Y=1.415
+ $X2=3.282 $Y2=0.445
r272 78 144 2.98324 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=2.55 $Y=1.54
+ $X2=2.437 $Y2=1.54
r273 77 146 6.1976 $w=2.5e-07 $l=1.27e-07 $layer=LI1_cond $X=3.155 $Y=1.54
+ $X2=3.282 $Y2=1.54
r274 77 78 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=3.155 $Y=1.54
+ $X2=2.55 $Y2=1.54
r275 71 144 3.11731 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=2.437 $Y=1.415
+ $X2=2.437 $Y2=1.54
r276 71 73 49.6831 $w=2.23e-07 $l=9.7e-07 $layer=LI1_cond $X=2.437 $Y=1.415
+ $X2=2.437 $Y2=0.445
r277 70 142 6.05271 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=1.69 $Y=1.56
+ $X2=1.562 $Y2=1.56
r278 69 144 2.98324 $w=2.1e-07 $l=1.21589e-07 $layer=LI1_cond $X=2.325 $Y=1.56
+ $X2=2.437 $Y2=1.54
r279 69 70 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=2.325 $Y=1.56
+ $X2=1.69 $Y2=1.56
r280 66 140 3.79048 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=0.83 $Y=1.56
+ $X2=0.702 $Y2=1.56
r281 65 142 6.05271 $w=2.1e-07 $l=1.27e-07 $layer=LI1_cond $X=1.435 $Y=1.56
+ $X2=1.562 $Y2=1.56
r282 65 66 31.9524 $w=2.08e-07 $l=6.05e-07 $layer=LI1_cond $X=1.435 $Y=1.56
+ $X2=0.83 $Y2=1.56
r283 61 140 3.10938 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=0.702 $Y=1.665
+ $X2=0.702 $Y2=1.56
r284 61 63 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.702 $Y=1.665
+ $X2=0.702 $Y2=2.3
r285 20 161 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=10.21
+ $Y=1.485 $X2=10.35 $Y2=1.62
r286 19 159 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=9.35
+ $Y=1.485 $X2=9.49 $Y2=1.62
r287 18 157 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=1.485 $X2=8.63 $Y2=1.62
r288 17 155 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=7.63
+ $Y=1.485 $X2=7.77 $Y2=1.62
r289 16 153 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=6.77
+ $Y=1.485 $X2=6.91 $Y2=1.62
r290 15 151 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.485 $X2=6.05 $Y2=1.62
r291 14 162 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.485 $X2=5.165 $Y2=1.62
r292 13 148 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=4
+ $Y=1.485 $X2=4.14 $Y2=1.62
r293 12 146 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=3.14
+ $Y=1.485 $X2=3.28 $Y2=1.62
r294 11 144 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=2.28
+ $Y=1.485 $X2=2.42 $Y2=1.62
r295 10 142 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=1.42
+ $Y=1.485 $X2=1.56 $Y2=1.62
r296 9 140 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.7 $Y2=1.62
r297 9 63 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.7 $Y2=2.3
r298 8 127 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.49
+ $Y=0.235 $X2=8.63 $Y2=0.445
r299 7 119 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.63
+ $Y=0.235 $X2=7.77 $Y2=0.445
r300 6 111 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.235 $X2=6.91 $Y2=0.445
r301 5 103 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.235 $X2=6.05 $Y2=0.445
r302 4 97 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=4.895
+ $Y=0.235 $X2=5.065 $Y2=0.445
r303 3 89 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.235 $X2=4.14 $Y2=0.445
r304 2 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.14
+ $Y=0.235 $X2=3.28 $Y2=0.445
r305 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.42 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_16%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 58 60 64 67 68 70 71 73 74 76 77 79 80 82 83 85 86 87 88 89 124 125 128
r121 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r122 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r123 122 125 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r124 122 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r125 121 124 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r126 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r127 119 128 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.062 $Y2=0
r128 119 121 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.43 $Y2=0
r129 118 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r130 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r131 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r132 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r133 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r134 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r135 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r136 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r137 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r138 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r139 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r140 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r141 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r142 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r143 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r144 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r145 92 96 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r146 89 97 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.61 $Y2=0
r147 89 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r148 87 117 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.05
+ $Y2=0
r149 87 88 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.202
+ $Y2=0
r150 85 114 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.21 $Y=0 $X2=7.13
+ $Y2=0
r151 85 86 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.21 $Y=0 $X2=7.342
+ $Y2=0
r152 84 117 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=8.05 $Y2=0
r153 84 86 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.342 $Y2=0
r154 82 111 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.35 $Y=0 $X2=6.21
+ $Y2=0
r155 82 83 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=6.35 $Y=0 $X2=6.462
+ $Y2=0
r156 81 114 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=7.13 $Y2=0
r157 81 83 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.462 $Y2=0
r158 79 108 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.49 $Y=0 $X2=5.29
+ $Y2=0
r159 79 80 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.49 $Y=0 $X2=5.622
+ $Y2=0
r160 78 111 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=6.21 $Y2=0
r161 78 80 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.622 $Y2=0
r162 76 105 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.37 $Y2=0
r163 76 77 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.597 $Y2=0
r164 75 108 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=5.29
+ $Y2=0
r165 75 77 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.597
+ $Y2=0
r166 73 102 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.45
+ $Y2=0
r167 73 74 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.712
+ $Y2=0
r168 72 105 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.845 $Y=0
+ $X2=4.37 $Y2=0
r169 72 74 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.845 $Y=0
+ $X2=3.712 $Y2=0
r170 70 99 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.53
+ $Y2=0
r171 70 71 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.852
+ $Y2=0
r172 69 102 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=3.45 $Y2=0
r173 69 71 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=2.852 $Y2=0
r174 67 96 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r175 67 68 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.99
+ $Y2=0
r176 66 99 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=0
+ $X2=2.53 $Y2=0
r177 66 68 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.99
+ $Y2=0
r178 62 128 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=9.062 $Y=0.085
+ $X2=9.062 $Y2=0
r179 62 64 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=9.062 $Y=0.085
+ $X2=9.062 $Y2=0.445
r180 61 88 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.335 $Y=0
+ $X2=8.202 $Y2=0
r181 60 128 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.93 $Y=0
+ $X2=9.062 $Y2=0
r182 60 61 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=8.93 $Y=0
+ $X2=8.335 $Y2=0
r183 56 88 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=8.202 $Y=0.085
+ $X2=8.202 $Y2=0
r184 56 58 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=8.202 $Y=0.085
+ $X2=8.202 $Y2=0.445
r185 52 86 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.342 $Y=0.085
+ $X2=7.342 $Y2=0
r186 52 54 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=7.342 $Y=0.085
+ $X2=7.342 $Y2=0.445
r187 48 83 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=6.462 $Y=0.085
+ $X2=6.462 $Y2=0
r188 48 50 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=6.462 $Y=0.085
+ $X2=6.462 $Y2=0.445
r189 44 80 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.622 $Y=0.085
+ $X2=5.622 $Y2=0
r190 44 46 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=5.622 $Y=0.085
+ $X2=5.622 $Y2=0.445
r191 40 77 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.597 $Y=0.085
+ $X2=4.597 $Y2=0
r192 40 42 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=4.597 $Y=0.085
+ $X2=4.597 $Y2=0.445
r193 36 74 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.712 $Y=0.085
+ $X2=3.712 $Y2=0
r194 36 38 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=3.712 $Y=0.085
+ $X2=3.712 $Y2=0.445
r195 32 71 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.852 $Y=0.085
+ $X2=2.852 $Y2=0
r196 32 34 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=2.852 $Y=0.085
+ $X2=2.852 $Y2=0.445
r197 28 68 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r198 28 30 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.445
r199 9 64 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.92
+ $Y=0.235 $X2=9.06 $Y2=0.445
r200 8 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.06
+ $Y=0.235 $X2=8.2 $Y2=0.445
r201 7 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.235 $X2=7.34 $Y2=0.445
r202 6 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.48 $Y2=0.445
r203 5 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.235 $X2=5.62 $Y2=0.445
r204 4 42 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.235 $X2=4.595 $Y2=0.445
r205 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.445
r206 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.85 $Y2=0.445
r207 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.235 $X2=1.99 $Y2=0.445
.ends


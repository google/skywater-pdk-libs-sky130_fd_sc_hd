* File: sky130_fd_sc_hd__a211oi_1.spice.SKY130_FD_SC_HD__A211OI_1.pxi
* Created: Thu Aug 27 13:59:42 2020
* 
x_PM_SKY130_FD_SC_HD__A211OI_1%A2 N_A2_c_45_n N_A2_M1002_g N_A2_M1007_g A2 A2
+ N_A2_c_47_n PM_SKY130_FD_SC_HD__A211OI_1%A2
x_PM_SKY130_FD_SC_HD__A211OI_1%A1 N_A1_M1003_g N_A1_M1000_g A1 A1 A1 A1
+ N_A1_c_74_n N_A1_c_75_n PM_SKY130_FD_SC_HD__A211OI_1%A1
x_PM_SKY130_FD_SC_HD__A211OI_1%B1 N_B1_M1004_g N_B1_M1005_g B1 B1 B1 B1
+ N_B1_c_108_n N_B1_c_109_n N_B1_c_110_n PM_SKY130_FD_SC_HD__A211OI_1%B1
x_PM_SKY130_FD_SC_HD__A211OI_1%C1 N_C1_c_143_n N_C1_M1001_g N_C1_M1006_g C1 C1
+ N_C1_c_145_n PM_SKY130_FD_SC_HD__A211OI_1%C1
x_PM_SKY130_FD_SC_HD__A211OI_1%A_56_297# N_A_56_297#_M1007_s N_A_56_297#_M1000_d
+ N_A_56_297#_c_173_n N_A_56_297#_c_175_n N_A_56_297#_c_174_n
+ N_A_56_297#_c_183_p PM_SKY130_FD_SC_HD__A211OI_1%A_56_297#
x_PM_SKY130_FD_SC_HD__A211OI_1%VPWR N_VPWR_M1007_d N_VPWR_c_190_n VPWR
+ N_VPWR_c_191_n N_VPWR_c_189_n N_VPWR_c_193_n PM_SKY130_FD_SC_HD__A211OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A211OI_1%Y N_Y_M1003_d N_Y_M1001_d N_Y_M1006_d N_Y_c_247_p
+ N_Y_c_226_n N_Y_c_225_n N_Y_c_250_p Y Y Y Y Y N_Y_c_221_n Y N_Y_c_224_n
+ PM_SKY130_FD_SC_HD__A211OI_1%Y
x_PM_SKY130_FD_SC_HD__A211OI_1%VGND N_VGND_M1002_s N_VGND_M1004_d N_VGND_c_256_n
+ N_VGND_c_257_n N_VGND_c_258_n VGND N_VGND_c_259_n N_VGND_c_260_n
+ N_VGND_c_261_n N_VGND_c_262_n PM_SKY130_FD_SC_HD__A211OI_1%VGND
cc_1 VNB N_A2_c_45_n 0.0188907f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=0.995
cc_2 VNB A2 0.0212651f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A2_c_47_n 0.0397136f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_4 VNB A1 0.00152833f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_5 VNB A1 0.00505989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A1_c_74_n 0.0212992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A1_c_75_n 0.0166487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B1_c_108_n 0.0204722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_109_n 0.00377768f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=0.85
cc_10 VNB N_B1_c_110_n 0.0167957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_C1_c_143_n 0.0202298f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=0.995
cc_12 VNB C1 0.00209371f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_13 VNB N_C1_c_145_n 0.0341016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_189_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=0.85
cc_15 VNB N_Y_c_221_n 0.02141f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB Y 0.0259888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_256_n 0.0114263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_257_n 0.020468f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_VGND_c_258_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_20 VNB N_VGND_c_259_n 0.0297299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_260_n 0.0246591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_261_n 0.165263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_262_n 0.00436092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_A2_M1007_g 0.0261857f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.985
cc_25 VPB A2 0.00869346f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_26 VPB N_A2_c_47_n 0.0107745f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_27 VPB N_A1_M1000_g 0.0191391f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.985
cc_28 VPB A1 0.00286938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A1_c_74_n 0.00391271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_B1_M1005_g 0.0187934f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.985
cc_31 VPB B1 9.54222e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_B1_c_108_n 0.00496919f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_C1_M1006_g 0.0237272f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.985
cc_34 VPB C1 0.00159926f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_35 VPB N_C1_c_145_n 0.00947836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_56_297#_c_173_n 0.0272566f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_37 VPB N_A_56_297#_c_174_n 0.00856363f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_38 VPB N_VPWR_c_190_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_39 VPB N_VPWR_c_191_n 0.0466323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_189_n 0.0535122f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=0.85
cc_41 VPB N_VPWR_c_193_n 0.0244979f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_42 VPB Y 0.0257493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_Y_c_224_n 0.0466322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 N_A2_M1007_g N_A1_M1000_g 0.0291506f $X=0.62 $Y=1.985 $X2=0 $Y2=0
cc_45 N_A2_c_45_n A1 0.0229361f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_46 A2 A1 0.0176664f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_47 N_A2_c_47_n A1 2.80579e-19 $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_48 A2 A1 0.0261123f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_49 N_A2_c_47_n A1 0.0121593f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_50 N_A2_c_47_n N_A1_c_74_n 0.0214526f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A2_c_45_n N_A1_c_75_n 0.0373148f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A2_M1007_g N_A_56_297#_c_175_n 0.0176997f $X=0.62 $Y=1.985 $X2=0 $Y2=0
cc_53 A2 N_A_56_297#_c_174_n 0.0140264f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_54 N_A2_c_47_n N_A_56_297#_c_174_n 0.00398542f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A2_M1007_g N_VPWR_c_190_n 0.0121357f $X=0.62 $Y=1.985 $X2=0 $Y2=0
cc_56 N_A2_M1007_g N_VPWR_c_189_n 0.00938618f $X=0.62 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A2_M1007_g N_VPWR_c_193_n 0.00486043f $X=0.62 $Y=1.985 $X2=0 $Y2=0
cc_58 A2 N_VGND_M1002_s 0.00514774f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_59 N_A2_c_45_n N_VGND_c_257_n 0.0120356f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_60 A2 N_VGND_c_257_n 0.0283822f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A2_c_47_n N_VGND_c_257_n 9.79086e-19 $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A2_c_45_n N_VGND_c_259_n 0.00451512f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A2_c_45_n N_VGND_c_261_n 0.00868629f $X=0.62 $Y=0.995 $X2=0 $Y2=0
cc_64 A2 N_VGND_c_261_n 0.00171493f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A1_M1000_g N_B1_M1005_g 0.0246394f $X=1.05 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A1_M1000_g B1 0.00110332f $X=1.05 $Y=1.985 $X2=0 $Y2=0
cc_67 A1 N_B1_c_108_n 0.00211592f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A1_c_74_n N_B1_c_108_n 0.0202452f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_69 A1 N_B1_c_109_n 0.026361f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A1_c_74_n N_B1_c_109_n 3.35397e-19 $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A1_c_75_n N_B1_c_110_n 0.0223771f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A1_M1000_g N_A_56_297#_c_175_n 0.0145078f $X=1.05 $Y=1.985 $X2=0 $Y2=0
cc_73 A1 N_A_56_297#_c_175_n 0.0375417f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A1_c_74_n N_A_56_297#_c_175_n 0.00140323f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A1_M1000_g N_VPWR_c_190_n 0.0112076f $X=1.05 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A1_M1000_g N_VPWR_c_191_n 0.00486043f $X=1.05 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A1_M1000_g N_VPWR_c_189_n 0.0083285f $X=1.05 $Y=1.985 $X2=0 $Y2=0
cc_78 A1 N_Y_c_225_n 0.00523492f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_79 A1 N_VGND_c_257_n 0.0240748f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_80 N_A1_c_75_n N_VGND_c_258_n 0.00118446f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_81 A1 N_VGND_c_259_n 0.0143434f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_82 N_A1_c_75_n N_VGND_c_259_n 0.00585385f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_83 A1 N_VGND_c_261_n 0.00909608f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_84 N_A1_c_75_n N_VGND_c_261_n 0.010919f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_85 A1 A_139_47# 0.00780089f $X=0.605 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_86 N_B1_c_110_n N_C1_c_143_n 0.0235362f $X=1.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_87 N_B1_M1005_g N_C1_M1006_g 0.0467741f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_88 B1 N_C1_M1006_g 0.00647125f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_89 N_B1_M1005_g C1 2.46639e-19 $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_90 N_B1_c_108_n C1 3.06227e-19 $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B1_c_109_n C1 0.0458027f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B1_c_108_n N_C1_c_145_n 0.0208083f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B1_c_109_n N_C1_c_145_n 0.00647125f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_M1005_g N_VPWR_c_190_n 0.00131861f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_95 N_B1_M1005_g N_VPWR_c_191_n 0.00541763f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_96 B1 N_VPWR_c_191_n 0.0131481f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_97 N_B1_M1005_g N_VPWR_c_189_n 0.00992051f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_98 B1 N_VPWR_c_189_n 0.00860568f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_99 B1 A_311_297# 0.0111621f $X=1.525 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_100 N_B1_c_108_n N_Y_c_226_n 5.70186e-19 $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B1_c_109_n N_Y_c_226_n 0.0225453f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B1_c_110_n N_Y_c_226_n 0.011863f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B1_M1005_g N_Y_c_224_n 5.65891e-19 $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_104 B1 N_Y_c_224_n 0.0512973f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_105 N_B1_c_110_n N_VGND_c_258_n 0.00686288f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B1_c_110_n N_VGND_c_259_n 0.00394671f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_c_110_n N_VGND_c_261_n 0.00458871f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_108 N_C1_M1006_g N_VPWR_c_191_n 0.00465161f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_109 N_C1_M1006_g N_VPWR_c_189_n 0.00935851f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_110 C1 N_Y_M1006_d 0.00357431f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_111 N_C1_c_143_n N_Y_c_226_n 0.0146835f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_112 C1 N_Y_c_226_n 0.02019f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_113 N_C1_c_145_n N_Y_c_221_n 0.00332372f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_114 N_C1_c_143_n Y 0.00480251f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C1_M1006_g Y 0.00440033f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_116 C1 Y 0.0412166f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_117 N_C1_c_145_n Y 0.00807521f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C1_M1006_g N_Y_c_224_n 0.0115016f $X=1.94 $Y=1.985 $X2=0 $Y2=0
cc_119 C1 N_Y_c_224_n 0.0209818f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_120 N_C1_c_145_n N_Y_c_224_n 0.00247125f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C1_c_143_n N_VGND_c_258_n 0.00759606f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_122 N_C1_c_143_n N_VGND_c_260_n 0.00394671f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_123 N_C1_c_143_n N_VGND_c_261_n 0.00591208f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_56_297#_c_175_n N_VPWR_M1007_d 0.00369081f $X=1.17 $Y=1.625 $X2=-0.19
+ $Y2=1.305
cc_125 N_A_56_297#_c_175_n N_VPWR_c_190_n 0.0165341f $X=1.17 $Y=1.625 $X2=0
+ $Y2=0
cc_126 N_A_56_297#_c_183_p N_VPWR_c_191_n 0.0115386f $X=1.265 $Y=1.85 $X2=0
+ $Y2=0
cc_127 N_A_56_297#_M1007_s N_VPWR_c_189_n 0.00374186f $X=0.28 $Y=1.485 $X2=0
+ $Y2=0
cc_128 N_A_56_297#_M1000_d N_VPWR_c_189_n 0.00561807f $X=1.125 $Y=1.485 $X2=0
+ $Y2=0
cc_129 N_A_56_297#_c_173_n N_VPWR_c_189_n 0.00950576f $X=0.405 $Y=1.85 $X2=0
+ $Y2=0
cc_130 N_A_56_297#_c_183_p N_VPWR_c_189_n 0.00701433f $X=1.265 $Y=1.85 $X2=0
+ $Y2=0
cc_131 N_A_56_297#_c_173_n N_VPWR_c_193_n 0.0160687f $X=0.405 $Y=1.85 $X2=0
+ $Y2=0
cc_132 N_VPWR_c_189_n A_311_297# 0.00634519f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_133 N_VPWR_c_189_n N_Y_M1006_d 0.00214593f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_134 N_VPWR_c_191_n N_Y_c_224_n 0.0459704f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_c_189_n N_Y_c_224_n 0.0273732f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_136 N_Y_c_226_n N_VGND_M1004_d 0.00554698f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_137 N_Y_c_226_n N_VGND_c_258_n 0.0162239f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_138 N_Y_c_247_p N_VGND_c_259_n 0.0113711f $X=1.265 $Y=0.53 $X2=0 $Y2=0
cc_139 N_Y_c_226_n N_VGND_c_259_n 0.00274625f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_140 N_Y_c_226_n N_VGND_c_260_n 0.00992518f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_141 N_Y_c_250_p N_VGND_c_260_n 0.0136074f $X=2.155 $Y=0.53 $X2=0 $Y2=0
cc_142 N_Y_M1003_d N_VGND_c_261_n 0.00432688f $X=1.125 $Y=0.235 $X2=0 $Y2=0
cc_143 N_Y_M1001_d N_VGND_c_261_n 0.00228064f $X=2.015 $Y=0.235 $X2=0 $Y2=0
cc_144 N_Y_c_247_p N_VGND_c_261_n 0.00696927f $X=1.265 $Y=0.53 $X2=0 $Y2=0
cc_145 N_Y_c_226_n N_VGND_c_261_n 0.0214052f $X=2.055 $Y=0.72 $X2=0 $Y2=0
cc_146 N_Y_c_250_p N_VGND_c_261_n 0.00840761f $X=2.155 $Y=0.53 $X2=0 $Y2=0
cc_147 N_VGND_c_261_n A_139_47# 0.00645095f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

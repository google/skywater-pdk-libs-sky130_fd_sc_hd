* File: sky130_fd_sc_hd__or2_1.spice
* Created: Thu Aug 27 14:42:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or2_1.pex.spice"
.subckt sky130_fd_sc_hd__or2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_A_68_297#_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_68_297#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.0567 PD=0.773271 PS=0.69 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_68_297#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.121799 PD=1.82 PS=1.19673 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 A_150_297# N_B_M1004_g N_A_68_297#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_150_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.0441 PD=0.789718 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8
+ SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_68_297#_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.34 AS=0.205282 PD=2.68 PS=1.88028 NRD=14.7553 NRS=0 M=1 R=6.66667
+ SA=75000.5 SB=75000.3 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_160 A_150_297# 0 1.0136e-19 $X=0.75 $Y=1.485
*
.include "sky130_fd_sc_hd__or2_1.pxi.spice"
*
.ends
*
*

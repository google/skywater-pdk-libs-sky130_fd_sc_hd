* File: sky130_fd_sc_hd__nand4b_4.pex.spice
* Created: Tue Sep  1 19:17:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4B_4%A_N 1 3 6 8 13
c30 8 0 1.2849e-19 $X=0.235 $Y=1.19
r31 11 13 30.8164 $w=3.05e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r33 4 13 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r34 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r35 1 13 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 41 43
+ 45 47 48 49 52 54 60 65 66 73
c129 66 0 1.2849e-19 $X=1.335 $Y=1.16
r130 72 73 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.67 $Y2=1.16
r131 69 70 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.41 $Y=1.16
+ $X2=1.83 $Y2=1.16
r132 66 69 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.41 $Y2=1.16
r133 61 72 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.04 $Y=1.16
+ $X2=2.25 $Y2=1.16
r134 61 70 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.04 $Y=1.16
+ $X2=1.83 $Y2=1.16
r135 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.16 $X2=2.04 $Y2=1.16
r136 58 66 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.335 $Y2=1.16
r137 57 60 48.2455 $w=1.98e-07 $l=8.7e-07 $layer=LI1_cond $X=1.17 $Y=1.175
+ $X2=2.04 $Y2=1.175
r138 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r139 55 65 1.25155 $w=2e-07 $l=9.8e-08 $layer=LI1_cond $X=0.805 $Y=1.175
+ $X2=0.707 $Y2=1.175
r140 55 57 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=0.805 $Y=1.175
+ $X2=1.17 $Y2=1.175
r141 53 65 5.27577 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=0.707 $Y=1.275
+ $X2=0.707 $Y2=1.175
r142 53 54 12.5128 $w=1.93e-07 $l=2.2e-07 $layer=LI1_cond $X=0.707 $Y=1.275
+ $X2=0.707 $Y2=1.495
r143 52 65 5.27577 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=0.707 $Y=1.075
+ $X2=0.707 $Y2=1.175
r144 51 52 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.707 $Y=0.905
+ $X2=0.707 $Y2=1.075
r145 50 64 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=1.58
+ $X2=0.257 $Y2=1.58
r146 49 54 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.61 $Y=1.58
+ $X2=0.707 $Y2=1.495
r147 49 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.61 $Y=1.58
+ $X2=0.425 $Y2=1.58
r148 47 51 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.61 $Y=0.82
+ $X2=0.707 $Y2=0.905
r149 47 48 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.61 $Y=0.82
+ $X2=0.425 $Y2=0.82
r150 43 64 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=1.58
r151 43 45 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.34
r152 39 48 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r153 39 41 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.38
r154 35 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.16
r155 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r156 31 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=1.16
r157 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=0.56
r158 27 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.16
r159 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.985
r160 23 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=1.16
r161 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r162 19 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.16
r163 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.985
r164 15 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=1.16
r165 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=0.56
r166 11 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.16
r167 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.985
r168 7 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.16
r169 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r170 2 64 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r171 2 45 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r172 1 41 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%B 3 7 11 15 19 23 27 31 33 34 35 36 47
r86 47 49 13.2418 $w=2.73e-07 $l=7.5e-08 $layer=POLY_cond $X=4.35 $Y=1.16
+ $X2=4.425 $Y2=1.16
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.12
+ $Y=1.16 $X2=3.12 $Y2=1.16
r88 36 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.425
+ $Y=1.16 $X2=4.425 $Y2=1.16
r89 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=4.395 $Y2=1.175
r90 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.935 $Y2=1.175
r91 34 44 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.12 $Y2=1.175
r92 33 44 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.12 $Y2=1.175
r93 29 47 16.7618 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.35 $Y=1.305
+ $X2=4.35 $Y2=1.16
r94 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.35 $Y=1.305
+ $X2=4.35 $Y2=1.985
r95 25 47 16.7618 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.35 $Y=1.015
+ $X2=4.35 $Y2=1.16
r96 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.35 $Y=1.015
+ $X2=4.35 $Y2=0.56
r97 17 47 74.1538 $w=2.73e-07 $l=4.2e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.35 $Y2=1.16
r98 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.985
r99 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=0.56
r100 9 17 74.1538 $w=2.73e-07 $l=4.2e-07 $layer=POLY_cond $X=3.51 $Y=1.16
+ $X2=3.93 $Y2=1.16
r101 9 43 68.8571 $w=2.73e-07 $l=3.9e-07 $layer=POLY_cond $X=3.51 $Y=1.16
+ $X2=3.12 $Y2=1.16
r102 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.985
r103 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=0.56
r104 1 43 5.2967 $w=2.73e-07 $l=3e-08 $layer=POLY_cond $X=3.09 $Y=1.16 $X2=3.12
+ $Y2=1.16
r105 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r106 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%C 3 7 11 15 19 23 27 31 33 34 35 36 41 51
+ 52
c82 51 0 1.21049e-19 $X=6.345 $Y=1.16
c83 27 0 1.79953e-19 $X=6.55 $Y=0.56
r84 50 52 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=6.345 $Y=1.16
+ $X2=6.55 $Y2=1.16
r85 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.345
+ $Y=1.16 $X2=6.345 $Y2=1.16
r86 48 50 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=6.13 $Y=1.16
+ $X2=6.345 $Y2=1.16
r87 47 48 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.71 $Y=1.16 $X2=6.13
+ $Y2=1.16
r88 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.29 $Y=1.16 $X2=5.71
+ $Y2=1.16
r89 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.985
+ $Y=1.16 $X2=4.985 $Y2=1.16
r90 41 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.215 $Y=1.16
+ $X2=5.29 $Y2=1.16
r91 41 43 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=5.215 $Y=1.16 $X2=4.985
+ $Y2=1.16
r92 36 51 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=6.255 $Y=1.175
+ $X2=6.345 $Y2=1.175
r93 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=5.795 $Y=1.175
+ $X2=6.255 $Y2=1.175
r94 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=5.335 $Y=1.175
+ $X2=5.795 $Y2=1.175
r95 34 44 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=5.335 $Y=1.175
+ $X2=4.985 $Y2=1.175
r96 33 44 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=4.875 $Y=1.175 $X2=4.985
+ $Y2=1.175
r97 29 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.16
r98 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.985
r99 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.025
+ $X2=6.55 $Y2=1.16
r100 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.55 $Y=1.025
+ $X2=6.55 $Y2=0.56
r101 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.13 $Y=1.295
+ $X2=6.13 $Y2=1.16
r102 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.13 $Y=1.295
+ $X2=6.13 $Y2=1.985
r103 17 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.13 $Y=1.025
+ $X2=6.13 $Y2=1.16
r104 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.13 $Y=1.025
+ $X2=6.13 $Y2=0.56
r105 13 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.71 $Y=1.295
+ $X2=5.71 $Y2=1.16
r106 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.71 $Y=1.295
+ $X2=5.71 $Y2=1.985
r107 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.71 $Y=1.025
+ $X2=5.71 $Y2=1.16
r108 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.71 $Y=1.025
+ $X2=5.71 $Y2=0.56
r109 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.29 $Y=1.295
+ $X2=5.29 $Y2=1.16
r110 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.29 $Y=1.295
+ $X2=5.29 $Y2=1.985
r111 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.29 $Y=1.025
+ $X2=5.29 $Y2=1.16
r112 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.29 $Y=1.025
+ $X2=5.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%D 3 7 11 15 19 23 27 31 33 34 35 36 41 43
c90 3 0 8.56806e-20 $X=6.97 $Y=0.56
r91 41 52 12.7139 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=8.305 $Y=1.16
+ $X2=8.23 $Y2=1.16
r92 41 43 34.1305 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.305 $Y=1.16
+ $X2=8.47 $Y2=1.16
r93 36 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.47
+ $Y=1.16 $X2=8.47 $Y2=1.16
r94 35 36 20.7955 $w=1.98e-07 $l=3.75e-07 $layer=LI1_cond $X=8.095 $Y=1.175
+ $X2=8.47 $Y2=1.175
r95 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=7.635 $Y=1.175
+ $X2=8.095 $Y2=1.175
r96 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=7.175 $Y=1.175
+ $X2=7.635 $Y2=1.175
r97 33 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.18
+ $Y=1.16 $X2=7.18 $Y2=1.16
r98 29 52 16.6763 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.23 $Y=1.305
+ $X2=8.23 $Y2=1.16
r99 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.23 $Y=1.305
+ $X2=8.23 $Y2=1.985
r100 25 52 16.6763 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.23 $Y=1.015
+ $X2=8.23 $Y2=1.16
r101 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.23 $Y=1.015
+ $X2=8.23 $Y2=0.56
r102 17 52 74.4265 $w=2.72e-07 $l=4.2e-07 $layer=POLY_cond $X=7.81 $Y=1.16
+ $X2=8.23 $Y2=1.16
r103 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.81 $Y=1.295
+ $X2=7.81 $Y2=1.985
r104 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.81 $Y=1.025
+ $X2=7.81 $Y2=0.56
r105 9 17 74.4265 $w=2.72e-07 $l=4.2e-07 $layer=POLY_cond $X=7.39 $Y=1.16
+ $X2=7.81 $Y2=1.16
r106 9 48 37.2132 $w=2.72e-07 $l=2.1e-07 $layer=POLY_cond $X=7.39 $Y=1.16
+ $X2=7.18 $Y2=1.16
r107 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.39 $Y=1.295
+ $X2=7.39 $Y2=1.985
r108 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.39 $Y=1.025
+ $X2=7.39 $Y2=0.56
r109 1 48 37.2132 $w=2.72e-07 $l=2.1e-07 $layer=POLY_cond $X=6.97 $Y=1.16
+ $X2=7.18 $Y2=1.16
r110 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.985
r111 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.97 $Y=1.025
+ $X2=6.97 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%VPWR 1 2 3 4 5 6 7 8 9 10 34 37 41 45 49 53
+ 57 61 63 67 69 71 76 79 80 82 83 85 86 88 89 90 91 92 94 109 120 126 129 132
+ 136
r135 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r136 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r137 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 124 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r140 124 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r141 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r142 121 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=2.72
+ $X2=7.6 $Y2=2.72
r143 121 123 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.685 $Y=2.72
+ $X2=8.05 $Y2=2.72
r144 120 135 4.02932 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=8.355 $Y=2.72
+ $X2=8.547 $Y2=2.72
r145 120 123 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.355 $Y=2.72
+ $X2=8.05 $Y2=2.72
r146 119 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r147 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r148 116 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r149 116 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r150 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r151 113 129 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=5.165 $Y=2.72
+ $X2=4.82 $Y2=2.72
r152 113 115 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.165 $Y=2.72
+ $X2=5.75 $Y2=2.72
r153 112 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r154 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 109 129 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.475 $Y=2.72
+ $X2=4.82 $Y2=2.72
r156 109 111 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=2.72
+ $X2=4.37 $Y2=2.72
r157 108 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r158 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r159 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r161 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r162 102 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r163 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r164 99 126 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=0.94 $Y2=2.72
r165 99 101 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.61 $Y2=2.72
r166 94 126 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.94 $Y2=2.72
r167 94 96 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r168 92 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r169 92 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r170 90 118 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.67 $Y2=2.72
r171 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.76 $Y2=2.72
r172 88 115 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=2.72
+ $X2=5.75 $Y2=2.72
r173 88 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=2.72
+ $X2=5.92 $Y2=2.72
r174 87 118 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.005 $Y=2.72
+ $X2=6.67 $Y2=2.72
r175 87 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.72
+ $X2=5.92 $Y2=2.72
r176 85 107 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.45 $Y2=2.72
r177 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.72 $Y2=2.72
r178 84 111 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=4.37 $Y2=2.72
r179 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.72 $Y2=2.72
r180 82 104 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r181 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.88 $Y2=2.72
r182 81 107 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=3.45 $Y2=2.72
r183 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.88 $Y2=2.72
r184 79 101 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r185 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.04 $Y2=2.72
r186 78 104 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.53 $Y2=2.72
r187 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.04 $Y2=2.72
r188 76 77 6.97577 $w=6.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=2 $X2=0.94
+ $Y2=1.835
r189 71 74 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=8.482 $Y=1.66
+ $X2=8.482 $Y2=2.34
r190 69 135 3.14791 $w=2.55e-07 $l=1.12916e-07 $layer=LI1_cond $X=8.482 $Y=2.635
+ $X2=8.547 $Y2=2.72
r191 69 74 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=8.482 $Y=2.635
+ $X2=8.482 $Y2=2.34
r192 65 132 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=2.635
+ $X2=7.6 $Y2=2.72
r193 65 67 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.6 $Y=2.635
+ $X2=7.6 $Y2=2
r194 64 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=2.72
+ $X2=6.76 $Y2=2.72
r195 63 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=2.72
+ $X2=7.6 $Y2=2.72
r196 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.515 $Y=2.72
+ $X2=6.845 $Y2=2.72
r197 59 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=2.635
+ $X2=6.76 $Y2=2.72
r198 59 61 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.76 $Y=2.635
+ $X2=6.76 $Y2=2
r199 55 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.635
+ $X2=5.92 $Y2=2.72
r200 55 57 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.92 $Y=2.635
+ $X2=5.92 $Y2=2
r201 51 129 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.82 $Y=2.635
+ $X2=4.82 $Y2=2.72
r202 51 53 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=4.82 $Y=2.635
+ $X2=4.82 $Y2=2
r203 47 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2.72
r204 47 49 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2
r205 43 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2.72
r206 43 45 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2
r207 39 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r208 39 41 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2
r209 37 77 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=1.14 $Y=1.66
+ $X2=1.14 $Y2=1.835
r210 32 126 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.72
r211 32 34 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.34
r212 31 76 3.1202 $w=6.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.94 $Y=2.18
+ $X2=0.94 $Y2=2
r213 31 34 2.77352 $w=6.88e-07 $l=1.6e-07 $layer=LI1_cond $X=0.94 $Y=2.18
+ $X2=0.94 $Y2=2.34
r214 10 74 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=2.34
r215 10 71 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=1.66
r216 9 67 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.465
+ $Y=1.485 $X2=7.6 $Y2=2
r217 8 61 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.625
+ $Y=1.485 $X2=6.76 $Y2=2
r218 7 57 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.785
+ $Y=1.485 $X2=5.92 $Y2=2
r219 6 53 150 $w=1.7e-07 $l=7.91675e-07 $layer=licon1_PDIFF $count=4 $X=4.425
+ $Y=1.485 $X2=5 $Y2=2
r220 5 49 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2
r221 4 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2
r222 3 41 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2
r223 2 37 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.66
r224 2 34 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.34
r225 1 76 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%Y 1 2 3 4 5 6 7 8 9 10 31 35 37 39 43 47 49
+ 53 55 59 61 65 67 71 73 75 77 81 83 85 87 89 91 94 95 96 103
r174 95 96 8.50329 $w=4.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.507 $Y=1.19
+ $X2=2.507 $Y2=1.445
r175 94 103 3.44693 $w=2.65e-07 $l=1.35e-07 $layer=LI1_cond $X=2.507 $Y=0.77
+ $X2=2.507 $Y2=0.905
r176 94 95 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=2.507 $Y=0.92
+ $X2=2.507 $Y2=1.19
r177 94 103 0.652326 $w=2.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.507 $Y=0.92
+ $X2=2.507 $Y2=0.905
r178 81 96 15.9003 $w=3.88e-07 $l=4.95e-07 $layer=LI1_cond $X=3.135 $Y=1.555
+ $X2=2.64 $Y2=1.555
r179 81 83 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=1.555
+ $X2=3.3 $Y2=1.555
r180 75 93 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=8.02 $Y=1.665
+ $X2=8.02 $Y2=1.555
r181 75 77 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.02 $Y=1.665
+ $X2=8.02 $Y2=2.34
r182 74 91 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.345 $Y=1.555
+ $X2=7.18 $Y2=1.555
r183 73 93 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.855 $Y=1.555
+ $X2=8.02 $Y2=1.555
r184 73 74 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=7.855 $Y=1.555
+ $X2=7.345 $Y2=1.555
r185 69 91 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=7.18 $Y=1.665
+ $X2=7.18 $Y2=1.555
r186 69 71 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.18 $Y=1.665
+ $X2=7.18 $Y2=2.34
r187 68 89 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=1.555
+ $X2=6.34 $Y2=1.555
r188 67 91 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=1.555
+ $X2=7.18 $Y2=1.555
r189 67 68 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=7.015 $Y=1.555
+ $X2=6.505 $Y2=1.555
r190 63 89 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.34 $Y=1.665
+ $X2=6.34 $Y2=1.555
r191 63 65 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.34 $Y=1.665
+ $X2=6.34 $Y2=2.34
r192 62 87 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=1.555
+ $X2=5.5 $Y2=1.555
r193 61 89 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=1.555
+ $X2=6.34 $Y2=1.555
r194 61 62 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=6.175 $Y=1.555
+ $X2=5.665 $Y2=1.555
r195 57 87 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.5 $Y=1.665
+ $X2=5.5 $Y2=1.555
r196 57 59 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.5 $Y=1.665
+ $X2=5.5 $Y2=2.34
r197 56 85 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=1.555
+ $X2=4.14 $Y2=1.555
r198 55 87 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=1.555
+ $X2=5.5 $Y2=1.555
r199 55 56 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=5.335 $Y=1.555
+ $X2=4.305 $Y2=1.555
r200 51 85 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.14 $Y=1.665
+ $X2=4.14 $Y2=1.555
r201 51 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.14 $Y=1.665
+ $X2=4.14 $Y2=2.34
r202 50 83 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=1.555
+ $X2=3.3 $Y2=1.555
r203 49 85 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=1.555
+ $X2=4.14 $Y2=1.555
r204 49 50 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=3.975 $Y=1.555
+ $X2=3.465 $Y2=1.555
r205 45 83 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.3 $Y=1.665
+ $X2=3.3 $Y2=1.555
r206 45 47 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.3 $Y=1.665
+ $X2=3.3 $Y2=2.34
r207 41 96 2.18349 $w=3.3e-07 $l=1.13446e-07 $layer=LI1_cond $X=2.46 $Y=1.665
+ $X2=2.467 $Y2=1.555
r208 41 43 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.46 $Y=1.665
+ $X2=2.46 $Y2=2.34
r209 40 80 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=1.555
+ $X2=1.62 $Y2=1.555
r210 39 96 4.01688 $w=2.2e-07 $l=1.72e-07 $layer=LI1_cond $X=2.295 $Y=1.555
+ $X2=2.467 $Y2=1.555
r211 39 40 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.295 $Y=1.555
+ $X2=1.785 $Y2=1.555
r212 35 80 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.555
r213 35 37 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=2.34
r214 31 94 3.37033 $w=2.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.375 $Y=0.77
+ $X2=2.507 $Y2=0.77
r215 31 33 32.2257 $w=2.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.375 $Y=0.77
+ $X2=1.62 $Y2=0.77
r216 10 93 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=1.66
r217 10 77 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.34
r218 9 91 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.485 $X2=7.18 $Y2=1.66
r219 9 71 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.485 $X2=7.18 $Y2=2.34
r220 8 89 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=1.66
r221 8 65 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=2.34
r222 7 87 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.5 $Y2=1.66
r223 7 59 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.5 $Y2=2.34
r224 6 85 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=1.66
r225 6 53 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.34
r226 5 83 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.66
r227 5 47 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2.34
r228 4 96 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.66
r229 4 43 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.34
r230 3 80 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.66
r231 3 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2.34
r232 2 94 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.72
r233 1 33 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%VGND 1 2 3 12 16 20 23 24 25 27 32 42 43 46
+ 49
r101 49 50 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r102 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r103 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r104 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r105 40 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r106 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r107 37 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.265 $Y=0 $X2=7.18
+ $Y2=0
r108 37 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=7.59 $Y2=0
r109 36 50 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=7.13
+ $Y2=0
r110 36 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r111 35 36 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r112 33 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.72
+ $Y2=0
r113 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r114 32 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=0 $X2=7.18
+ $Y2=0
r115 32 35 387.856 $w=1.68e-07 $l=5.945e-06 $layer=LI1_cond $X=7.095 $Y=0
+ $X2=1.15 $Y2=0
r116 27 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.72
+ $Y2=0
r117 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r118 25 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 23 39 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.59
+ $Y2=0
r121 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=0 $X2=8.02
+ $Y2=0
r122 22 42 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=8.51 $Y2=0
r123 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.02
+ $Y2=0
r124 18 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0
r125 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0.38
r126 14 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=0.085
+ $X2=7.18 $Y2=0
r127 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.18 $Y=0.085
+ $X2=7.18 $Y2=0.38
r128 10 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r129 10 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.38
r130 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.38
r131 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.045
+ $Y=0.235 $X2=7.18 $Y2=0.38
r132 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%A_215_47# 1 2 3 4 5 16 18 28
r44 26 28 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=3.72 $Y=0.36
+ $X2=4.56 $Y2=0.36
r45 24 26 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=2.88 $Y=0.36
+ $X2=3.72 $Y2=0.36
r46 22 24 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=2.04 $Y=0.36
+ $X2=2.88 $Y2=0.36
r47 20 31 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=1.16 $Y2=0.36
r48 20 22 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=2.04 $Y2=0.36
r49 16 31 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.36
r50 16 18 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.72
r51 5 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.38
r52 4 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.38
r53 3 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.38
r54 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r55 1 31 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
r56 1 18 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%A_633_47# 1 2 3 4 21
c34 21 0 8.56806e-20 $X=6.34 $Y=0.72
r35 19 21 35.8538 $w=2.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.5 $Y=0.77 $X2=6.34
+ $Y2=0.77
r36 17 19 58.049 $w=2.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.14 $Y=0.77 $X2=5.5
+ $Y2=0.77
r37 14 17 35.8538 $w=2.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.3 $Y=0.77 $X2=4.14
+ $Y2=0.77
r38 4 21 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.205
+ $Y=0.235 $X2=6.34 $Y2=0.72
r39 3 19 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.235 $X2=5.5 $Y2=0.72
r40 2 17 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.72
r41 1 14 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_4%A_991_47# 1 2 3 4 5 16 22 25 26 27 30 32 36
+ 40
c65 27 0 1.79953e-19 $X=6.925 $Y=0.82
c66 16 0 1.21049e-19 $X=6.675 $Y=0.36
r67 34 36 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=8.442 $Y=0.735
+ $X2=8.442 $Y2=0.38
r68 33 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0.82
+ $X2=7.6 $Y2=0.82
r69 32 34 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=8.275 $Y=0.82
+ $X2=8.442 $Y2=0.735
r70 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.275 $Y=0.82
+ $X2=7.765 $Y2=0.82
r71 28 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=0.735 $X2=7.6
+ $Y2=0.82
r72 28 30 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.6 $Y=0.735
+ $X2=7.6 $Y2=0.38
r73 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=0.82
+ $X2=7.6 $Y2=0.82
r74 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.435 $Y=0.82
+ $X2=6.925 $Y2=0.82
r75 23 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.8 $Y=0.735
+ $X2=6.925 $Y2=0.82
r76 23 25 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=6.8 $Y=0.735
+ $X2=6.8 $Y2=0.72
r77 22 39 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=6.8 $Y=0.465 $X2=6.8
+ $Y2=0.36
r78 22 25 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.8 $Y=0.465
+ $X2=6.8 $Y2=0.72
r79 18 21 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=5.08 $Y=0.36
+ $X2=5.92 $Y2=0.36
r80 16 39 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.675 $Y=0.36
+ $X2=6.8 $Y2=0.36
r81 16 21 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=6.675 $Y=0.36
+ $X2=5.92 $Y2=0.36
r82 5 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.38
r83 4 30 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.465
+ $Y=0.235 $X2=7.6 $Y2=0.38
r84 3 39 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.235 $X2=6.76 $Y2=0.38
r85 3 25 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.235 $X2=6.76 $Y2=0.72
r86 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.235 $X2=5.92 $Y2=0.38
r87 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.08 $Y2=0.38
.ends


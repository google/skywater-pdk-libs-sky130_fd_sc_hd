* File: sky130_fd_sc_hd__o2bb2ai_1.pxi.spice
* Created: Thu Aug 27 14:38:34 2020
* 
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%A1_N N_A1_N_c_59_n N_A1_N_M1008_g N_A1_N_M1004_g
+ A1_N N_A1_N_c_61_n PM_SKY130_FD_SC_HD__O2BB2AI_1%A1_N
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%A2_N N_A2_N_M1006_g N_A2_N_M1009_g A2_N
+ N_A2_N_c_82_n N_A2_N_c_83_n N_A2_N_c_84_n N_A2_N_c_85_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_1%A2_N
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%A_112_297# N_A_112_297#_M1006_d
+ N_A_112_297#_M1004_d N_A_112_297#_c_122_n N_A_112_297#_M1000_g
+ N_A_112_297#_M1007_g N_A_112_297#_c_123_n N_A_112_297#_c_124_n
+ N_A_112_297#_c_159_p N_A_112_297#_c_136_n N_A_112_297#_c_139_n
+ N_A_112_297#_c_125_n N_A_112_297#_c_132_n N_A_112_297#_c_126_n
+ N_A_112_297#_c_127_n N_A_112_297#_c_128_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_1%A_112_297#
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%B2 N_B2_c_182_n N_B2_M1003_g N_B2_M1005_g
+ N_B2_c_183_n N_B2_c_184_n B2 PM_SKY130_FD_SC_HD__O2BB2AI_1%B2
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%B1 N_B1_c_223_n N_B1_M1001_g N_B1_M1002_g B1
+ N_B1_c_225_n PM_SKY130_FD_SC_HD__O2BB2AI_1%B1
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%VPWR N_VPWR_M1004_s N_VPWR_M1009_d
+ N_VPWR_M1002_d N_VPWR_c_249_n N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n
+ N_VPWR_c_253_n VPWR N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n
+ N_VPWR_c_248_n PM_SKY130_FD_SC_HD__O2BB2AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%Y N_Y_M1000_s N_Y_M1007_d N_Y_c_294_n
+ N_Y_c_303_n N_Y_c_296_n Y PM_SKY130_FD_SC_HD__O2BB2AI_1%Y
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%VGND N_VGND_M1008_s N_VGND_M1003_d
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n N_VGND_c_334_n
+ VGND N_VGND_c_335_n N_VGND_c_336_n PM_SKY130_FD_SC_HD__O2BB2AI_1%VGND
x_PM_SKY130_FD_SC_HD__O2BB2AI_1%A_394_47# N_A_394_47#_M1000_d
+ N_A_394_47#_M1001_d N_A_394_47#_c_379_n N_A_394_47#_c_375_n
+ N_A_394_47#_c_376_n N_A_394_47#_c_377_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_1%A_394_47#
cc_1 VNB N_A1_N_c_59_n 0.0206444f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB A1_N 0.0151055f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A1_N_c_61_n 0.0382042f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_4 VNB N_A2_N_c_82_n 0.022462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A2_N_c_83_n 0.00236211f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_6 VNB N_A2_N_c_84_n 0.0183631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A2_N_c_85_n 0.00145567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_112_297#_c_122_n 0.0193916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_112_297#_c_123_n 0.0400467f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_10 VNB N_A_112_297#_c_124_n 0.0101887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_112_297#_c_125_n 0.00484836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_112_297#_c_126_n 0.0016501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_112_297#_c_127_n 0.00665212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_112_297#_c_128_n 0.00231983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B2_c_182_n 0.0162183f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_16 VNB N_B2_c_183_n 0.00584658f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_17 VNB N_B2_c_184_n 0.0190143f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_18 VNB N_B1_c_223_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_19 VNB B1 0.0092237f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_20 VNB N_B1_c_225_n 0.0387151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_248_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_294_n 0.0021772f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_23 VNB N_VGND_c_330_n 0.0103615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_331_n 0.0257225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_332_n 0.00467422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_333_n 0.0537918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_334_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_335_n 0.0179469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_336_n 0.190848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_394_47#_c_375_n 0.0128186f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_31 VNB N_A_394_47#_c_376_n 0.00268834f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_32 VNB N_A_394_47#_c_377_n 0.0176751f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A1_N_M1004_g 0.0255341f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_34 VPB N_A1_N_c_61_n 0.0111135f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_35 VPB N_A2_N_M1009_g 0.0224136f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_36 VPB N_A2_N_c_82_n 0.00411535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A2_N_c_83_n 0.00172123f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_38 VPB N_A_112_297#_M1007_g 0.0221836f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_39 VPB N_A_112_297#_c_123_n 0.0179747f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_40 VPB N_A_112_297#_c_124_n 6.39329e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_112_297#_c_132_n 0.00291982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_112_297#_c_127_n 0.00202528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B2_M1005_g 0.0191064f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_44 VPB N_B2_c_183_n 0.00170932f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_45 VPB N_B2_c_184_n 0.00537013f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_46 VPB B2 0.00281798f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_47 VPB N_B1_M1002_g 0.0254848f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_48 VPB N_B1_c_225_n 0.0111302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_249_n 0.0117686f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_50 VPB N_VPWR_c_250_n 0.00760593f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_51 VPB N_VPWR_c_251_n 0.00744134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_252_n 0.0117686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_253_n 0.00812731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_254_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_255_n 0.0285636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_256_n 0.0149739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_248_n 0.0462699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_Y_c_294_n 0.0029742f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_59 N_A1_N_M1004_g N_A2_N_M1009_g 0.0257189f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_60 A1_N N_A2_N_c_82_n 2.19072e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_61 N_A1_N_c_61_n N_A2_N_c_82_n 0.0370785f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_62 A1_N N_A2_N_c_83_n 0.0234435f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A1_N_c_61_n N_A2_N_c_83_n 0.00335835f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A1_N_c_59_n N_A2_N_c_84_n 0.0370785f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A1_N_c_59_n N_A2_N_c_85_n 0.00450768f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_66 A1_N N_A2_N_c_85_n 6.58212e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A1_N_M1004_g N_VPWR_c_250_n 0.00463996f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_68 A1_N N_VPWR_c_250_n 0.020778f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A1_N_c_61_n N_VPWR_c_250_n 0.00606334f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A1_N_M1004_g N_VPWR_c_254_n 0.00585385f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A1_N_M1004_g N_VPWR_c_248_n 0.0114323f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A1_N_c_59_n N_VGND_c_331_n 0.0116313f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_73 A1_N N_VGND_c_331_n 0.0260499f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A1_N_c_61_n N_VGND_c_331_n 0.00218111f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A1_N_c_59_n N_VGND_c_333_n 0.00525069f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A1_N_c_59_n N_VGND_c_336_n 0.00875452f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A2_N_c_82_n N_A_112_297#_c_123_n 0.0203089f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A2_N_c_83_n N_A_112_297#_c_123_n 3.23394e-19 $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_79 N_A2_N_M1009_g N_A_112_297#_c_136_n 0.0161808f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_80 N_A2_N_c_82_n N_A_112_297#_c_136_n 0.00123493f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_81 N_A2_N_c_83_n N_A_112_297#_c_136_n 0.0118376f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A2_N_c_82_n N_A_112_297#_c_139_n 0.00121878f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_83 N_A2_N_c_83_n N_A_112_297#_c_139_n 0.0157851f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A2_N_c_84_n N_A_112_297#_c_125_n 0.011884f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A2_N_c_85_n N_A_112_297#_c_125_n 0.0402206f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A2_N_M1009_g N_A_112_297#_c_132_n 0.00564554f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_87 N_A2_N_c_82_n N_A_112_297#_c_126_n 0.00115304f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_88 N_A2_N_c_82_n N_A_112_297#_c_127_n 0.00197689f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A2_N_c_83_n N_A_112_297#_c_127_n 0.0262303f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A2_N_c_84_n N_A_112_297#_c_128_n 0.00321851f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_91 N_A2_N_c_85_n N_A_112_297#_c_128_n 0.00716273f $X=0.715 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A2_N_M1009_g N_VPWR_c_251_n 0.00352998f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A2_N_M1009_g N_VPWR_c_254_n 0.00585385f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A2_N_M1009_g N_VPWR_c_248_n 0.01179f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A2_N_M1009_g N_Y_c_296_n 6.51986e-19 $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A2_N_c_84_n N_VGND_c_331_n 0.00172438f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A2_N_c_84_n N_VGND_c_333_n 0.00505274f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A2_N_c_85_n N_VGND_c_333_n 0.0111129f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A2_N_c_84_n N_VGND_c_336_n 0.0100595f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A2_N_c_85_n N_VGND_c_336_n 0.0080551f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A2_N_c_85_n A_112_47# 9.93238e-19 $X=0.715 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_102 N_A_112_297#_c_122_n N_B2_c_182_n 0.0238836f $X=1.895 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_112_297#_M1007_g N_B2_M1005_g 0.013692f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_112_297#_c_124_n N_B2_c_183_n 0.00228667f $X=1.895 $Y=1.16 $X2=0
+ $Y2=0
cc_105 N_A_112_297#_c_124_n N_B2_c_184_n 0.022209f $X=1.895 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_112_297#_c_136_n N_VPWR_M1009_d 0.00952422f $X=1.17 $Y=1.58 $X2=0
+ $Y2=0
cc_107 N_A_112_297#_c_132_n N_VPWR_M1009_d 2.13521e-19 $X=1.255 $Y=1.495 $X2=0
+ $Y2=0
cc_108 N_A_112_297#_M1007_g N_VPWR_c_251_n 0.0173285f $X=1.895 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_112_297#_c_123_n N_VPWR_c_251_n 0.00654341f $X=1.82 $Y=1.16 $X2=0
+ $Y2=0
cc_110 N_A_112_297#_c_136_n N_VPWR_c_251_n 0.0260215f $X=1.17 $Y=1.58 $X2=0
+ $Y2=0
cc_111 N_A_112_297#_c_127_n N_VPWR_c_251_n 0.00454295f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_112 N_A_112_297#_c_159_p N_VPWR_c_254_n 0.0142343f $X=0.695 $Y=1.96 $X2=0
+ $Y2=0
cc_113 N_A_112_297#_M1007_g N_VPWR_c_255_n 0.00541359f $X=1.895 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_112_297#_M1004_d N_VPWR_c_248_n 0.00284632f $X=0.56 $Y=1.485 $X2=0
+ $Y2=0
cc_115 N_A_112_297#_M1007_g N_VPWR_c_248_n 0.0109815f $X=1.895 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_112_297#_c_159_p N_VPWR_c_248_n 0.00955092f $X=0.695 $Y=1.96 $X2=0
+ $Y2=0
cc_117 N_A_112_297#_c_122_n N_Y_c_294_n 0.00582248f $X=1.895 $Y=0.995 $X2=0
+ $Y2=0
cc_118 N_A_112_297#_M1007_g N_Y_c_294_n 0.00487298f $X=1.895 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_112_297#_c_123_n N_Y_c_294_n 0.0200293f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_112_297#_c_132_n N_Y_c_294_n 0.00855475f $X=1.255 $Y=1.495 $X2=0
+ $Y2=0
cc_121 N_A_112_297#_c_126_n N_Y_c_294_n 0.0102948f $X=1.17 $Y=0.825 $X2=0 $Y2=0
cc_122 N_A_112_297#_c_127_n N_Y_c_294_n 0.0233867f $X=1.385 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_112_297#_c_123_n N_Y_c_303_n 0.00311175f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_112_297#_c_125_n N_Y_c_303_n 0.0239842f $X=1.165 $Y=0.39 $X2=0 $Y2=0
cc_125 N_A_112_297#_M1007_g N_Y_c_296_n 0.0174092f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_112_297#_c_123_n N_Y_c_296_n 8.19407e-19 $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_112_297#_c_136_n N_Y_c_296_n 0.0098813f $X=1.17 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_112_297#_M1007_g Y 0.0146918f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_112_297#_c_122_n N_VGND_c_333_n 0.00585385f $X=1.895 $Y=0.995 $X2=0
+ $Y2=0
cc_130 N_A_112_297#_c_125_n N_VGND_c_333_n 0.0203781f $X=1.165 $Y=0.39 $X2=0
+ $Y2=0
cc_131 N_A_112_297#_M1006_d N_VGND_c_336_n 0.00582732f $X=0.92 $Y=0.235 $X2=0
+ $Y2=0
cc_132 N_A_112_297#_c_122_n N_VGND_c_336_n 0.0122169f $X=1.895 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_112_297#_c_125_n N_VGND_c_336_n 0.0128195f $X=1.165 $Y=0.39 $X2=0
+ $Y2=0
cc_134 N_A_112_297#_c_122_n N_A_394_47#_c_376_n 5.52151e-19 $X=1.895 $Y=0.995
+ $X2=0 $Y2=0
cc_135 N_B2_c_182_n N_B1_c_223_n 0.0258694f $X=2.315 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_136 N_B2_M1005_g N_B1_M1002_g 0.0499138f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_137 B2 N_B1_M1002_g 0.00723463f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_138 N_B2_c_183_n B1 0.0174773f $X=2.445 $Y=1.2 $X2=0 $Y2=0
cc_139 N_B2_c_183_n N_B1_c_225_n 0.00296314f $X=2.445 $Y=1.2 $X2=0 $Y2=0
cc_140 N_B2_c_184_n N_B1_c_225_n 0.0217754f $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_141 B2 N_VPWR_c_253_n 0.00197059f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_142 N_B2_M1005_g N_VPWR_c_255_n 0.00541359f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_143 B2 N_VPWR_c_255_n 0.00906544f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_144 N_B2_M1005_g N_VPWR_c_248_n 0.00975563f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_145 B2 N_VPWR_c_248_n 0.00633628f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_146 N_B2_c_183_n N_Y_c_294_n 0.0162871f $X=2.445 $Y=1.2 $X2=0 $Y2=0
cc_147 N_B2_c_184_n N_Y_c_294_n 5.96318e-19 $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_148 B2 N_Y_c_294_n 0.0046733f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_149 N_B2_M1005_g N_Y_c_296_n 0.00226417f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B2_c_183_n N_Y_c_296_n 0.0157638f $X=2.445 $Y=1.2 $X2=0 $Y2=0
cc_151 N_B2_c_184_n N_Y_c_296_n 0.00122018f $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_152 N_B2_M1005_g Y 0.00906361f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_153 B2 A_478_297# 0.00948631f $X=2.445 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_154 N_B2_c_182_n N_VGND_c_332_n 0.00268723f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_182_n N_VGND_c_333_n 0.00429718f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B2_c_182_n N_VGND_c_336_n 0.00584248f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B2_c_182_n N_A_394_47#_c_379_n 0.00473705f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_158 N_B2_c_182_n N_A_394_47#_c_375_n 0.00865686f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_B2_c_183_n N_A_394_47#_c_375_n 0.0268047f $X=2.445 $Y=1.2 $X2=0 $Y2=0
cc_160 N_B2_c_184_n N_A_394_47#_c_375_n 0.00148082f $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B2_c_182_n N_A_394_47#_c_376_n 0.00191187f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_B2_c_183_n N_A_394_47#_c_376_n 0.0197611f $X=2.445 $Y=1.2 $X2=0 $Y2=0
cc_163 N_B2_c_184_n N_A_394_47#_c_376_n 0.00152154f $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B2_c_182_n N_A_394_47#_c_377_n 5.16334e-19 $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_B1_M1002_g N_VPWR_c_253_n 0.00554249f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_166 B1 N_VPWR_c_253_n 0.0202873f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_167 N_B1_c_225_n N_VPWR_c_253_n 0.00606334f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_M1002_g N_VPWR_c_255_n 0.00585385f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_169 N_B1_M1002_g N_VPWR_c_248_n 0.0115092f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_170 N_B1_M1002_g Y 3.49602e-19 $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B1_c_223_n N_VGND_c_332_n 0.00268723f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_223_n N_VGND_c_335_n 0.00424138f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B1_c_223_n N_VGND_c_336_n 0.0067128f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B1_c_223_n N_A_394_47#_c_379_n 4.72684e-19 $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_B1_c_223_n N_A_394_47#_c_375_n 0.0135592f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_176 B1 N_A_394_47#_c_375_n 0.026301f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_177 N_B1_c_225_n N_A_394_47#_c_375_n 0.0076706f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B1_c_223_n N_A_394_47#_c_377_n 0.00612654f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_248_n N_Y_M1007_d 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_180 N_VPWR_M1009_d N_Y_c_294_n 4.87112e-19 $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_181 N_VPWR_M1009_d N_Y_c_296_n 0.00379869f $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_182 N_VPWR_c_251_n N_Y_c_296_n 0.00997062f $X=1.605 $Y=1.96 $X2=0 $Y2=0
cc_183 N_VPWR_c_255_n Y 0.0189039f $X=2.82 $Y=2.72 $X2=0 $Y2=0
cc_184 N_VPWR_c_248_n Y 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_185 N_VPWR_c_248_n A_478_297# 0.00572363f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_186 N_Y_c_303_n N_VGND_c_333_n 0.00729741f $X=1.685 $Y=0.605 $X2=0 $Y2=0
cc_187 N_Y_M1000_s N_VGND_c_336_n 0.00272996f $X=1.56 $Y=0.235 $X2=0 $Y2=0
cc_188 N_Y_c_303_n N_VGND_c_336_n 0.00856237f $X=1.685 $Y=0.605 $X2=0 $Y2=0
cc_189 N_Y_c_294_n N_A_394_47#_c_376_n 0.00160357f $X=1.725 $Y=1.495 $X2=0 $Y2=0
cc_190 N_Y_c_296_n N_A_394_47#_c_376_n 9.73798e-19 $X=2.105 $Y=1.62 $X2=0 $Y2=0
cc_191 N_VGND_c_336_n A_112_47# 0.00329021f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_192 N_VGND_c_336_n N_A_394_47#_M1000_d 0.00280325f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_193 N_VGND_c_336_n N_A_394_47#_M1001_d 0.00210124f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_333_n N_A_394_47#_c_379_n 0.00776949f $X=2.44 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_336_n N_A_394_47#_c_379_n 0.0097648f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_M1003_d N_A_394_47#_c_375_n 0.00162089f $X=2.39 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_VGND_c_332_n N_A_394_47#_c_375_n 0.0122559f $X=2.525 $Y=0.39 $X2=0
+ $Y2=0
cc_198 N_VGND_c_333_n N_A_394_47#_c_375_n 0.00198695f $X=2.44 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_335_n N_A_394_47#_c_375_n 0.00198695f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_336_n N_A_394_47#_c_375_n 0.00835832f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_201 N_VGND_c_335_n N_A_394_47#_c_377_n 0.018566f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_336_n N_A_394_47#_c_377_n 0.0122779f $X=2.99 $Y=0 $X2=0 $Y2=0

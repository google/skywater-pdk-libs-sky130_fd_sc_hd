* NGSPICE file created from sky130_fd_sc_hd__a41o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_381_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=9.6e+11p pd=7.92e+06u as=1.06e+12p ps=1.012e+07u
M1001 VPWR A2 a_381_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=3.38e+11p ps=3.64e+06u
M1003 a_665_47# A2 a_549_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.795e+11p ps=2.16e+06u
M1004 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 a_465_47# A4 VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1006 a_79_21# A1 a_665_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1008 a_549_47# A3 a_465_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_381_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A4 a_381_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_381_297# B1 a_79_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1013 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a2111oi_4.spice.SKY130_FD_SC_HD__A2111OI_4.pxi
* Created: Thu Aug 27 13:59:11 2020
* 
x_PM_SKY130_FD_SC_HD__A2111OI_4%D1 N_D1_M1003_g N_D1_c_132_n N_D1_M1007_g
+ N_D1_c_133_n N_D1_M1009_g N_D1_M1014_g N_D1_c_134_n N_D1_M1016_g N_D1_M1015_g
+ N_D1_c_135_n N_D1_M1027_g N_D1_M1032_g D1 N_D1_c_136_n N_D1_c_137_n
+ PM_SKY130_FD_SC_HD__A2111OI_4%D1
x_PM_SKY130_FD_SC_HD__A2111OI_4%C1 N_C1_M1005_g N_C1_c_208_n N_C1_M1008_g
+ N_C1_M1011_g N_C1_c_209_n N_C1_M1010_g N_C1_M1023_g N_C1_c_210_n N_C1_M1021_g
+ N_C1_M1028_g N_C1_c_211_n N_C1_M1036_g C1 N_C1_c_212_n N_C1_c_213_n
+ PM_SKY130_FD_SC_HD__A2111OI_4%C1
x_PM_SKY130_FD_SC_HD__A2111OI_4%B1 N_B1_c_293_n N_B1_M1001_g N_B1_M1012_g
+ N_B1_c_294_n N_B1_M1002_g N_B1_M1013_g N_B1_c_295_n N_B1_M1029_g N_B1_M1025_g
+ N_B1_c_296_n N_B1_M1037_g N_B1_M1031_g B1 N_B1_c_297_n N_B1_c_298_n
+ PM_SKY130_FD_SC_HD__A2111OI_4%B1
x_PM_SKY130_FD_SC_HD__A2111OI_4%A1 N_A1_M1018_g N_A1_c_376_n N_A1_M1017_g
+ N_A1_M1026_g N_A1_c_377_n N_A1_M1020_g N_A1_M1033_g N_A1_c_378_n N_A1_M1034_g
+ N_A1_M1035_g N_A1_c_379_n N_A1_M1038_g A1 N_A1_c_380_n N_A1_c_381_n
+ PM_SKY130_FD_SC_HD__A2111OI_4%A1
x_PM_SKY130_FD_SC_HD__A2111OI_4%A2 N_A2_M1000_g N_A2_c_448_n N_A2_M1006_g
+ N_A2_M1004_g N_A2_c_449_n N_A2_M1022_g N_A2_M1019_g N_A2_c_450_n N_A2_M1024_g
+ N_A2_M1030_g N_A2_c_451_n N_A2_M1039_g A2 N_A2_c_452_n N_A2_c_453_n
+ N_A2_c_464_n PM_SKY130_FD_SC_HD__A2111OI_4%A2
x_PM_SKY130_FD_SC_HD__A2111OI_4%A_28_297# N_A_28_297#_M1003_d
+ N_A_28_297#_M1014_d N_A_28_297#_M1032_d N_A_28_297#_M1011_d
+ N_A_28_297#_M1028_d N_A_28_297#_c_518_n N_A_28_297#_c_519_n
+ N_A_28_297#_c_522_n N_A_28_297#_c_541_p N_A_28_297#_c_524_n
+ N_A_28_297#_c_526_n N_A_28_297#_c_528_n N_A_28_297#_c_549_p
+ N_A_28_297#_c_530_n N_A_28_297#_c_520_n N_A_28_297#_c_521_n
+ N_A_28_297#_c_564_p N_A_28_297#_c_565_p N_A_28_297#_c_566_p
+ PM_SKY130_FD_SC_HD__A2111OI_4%A_28_297#
x_PM_SKY130_FD_SC_HD__A2111OI_4%Y N_Y_M1007_s N_Y_M1016_s N_Y_M1008_d
+ N_Y_M1021_d N_Y_M1001_d N_Y_M1029_d N_Y_M1017_s N_Y_M1034_s N_Y_M1003_s
+ N_Y_M1015_s N_Y_c_583_n N_Y_c_584_n N_Y_c_591_n N_Y_c_585_n N_Y_c_599_n
+ N_Y_c_622_n N_Y_c_626_n N_Y_c_639_n N_Y_c_581_n N_Y_c_586_n N_Y_c_606_n
+ N_Y_c_587_n N_Y_c_614_n N_Y_c_630_n N_Y_c_632_n N_Y_c_635_n N_Y_c_650_n Y
+ N_Y_c_677_p Y PM_SKY130_FD_SC_HD__A2111OI_4%Y
x_PM_SKY130_FD_SC_HD__A2111OI_4%A_455_297# N_A_455_297#_M1005_s
+ N_A_455_297#_M1023_s N_A_455_297#_M1012_s N_A_455_297#_M1025_s
+ N_A_455_297#_c_738_n N_A_455_297#_c_739_n N_A_455_297#_c_740_n
+ N_A_455_297#_c_741_n N_A_455_297#_c_742_n N_A_455_297#_c_743_n
+ N_A_455_297#_c_744_n PM_SKY130_FD_SC_HD__A2111OI_4%A_455_297#
x_PM_SKY130_FD_SC_HD__A2111OI_4%A_821_297# N_A_821_297#_M1012_d
+ N_A_821_297#_M1013_d N_A_821_297#_M1031_d N_A_821_297#_M1026_d
+ N_A_821_297#_M1035_d N_A_821_297#_M1004_s N_A_821_297#_M1030_s
+ N_A_821_297#_c_808_n N_A_821_297#_c_809_n N_A_821_297#_c_819_n
+ N_A_821_297#_c_857_n N_A_821_297#_c_821_n N_A_821_297#_c_810_n
+ N_A_821_297#_c_811_n N_A_821_297#_c_867_p N_A_821_297#_c_812_n
+ N_A_821_297#_c_813_n N_A_821_297#_c_870_p N_A_821_297#_c_814_n
+ N_A_821_297#_c_815_n N_A_821_297#_c_875_p N_A_821_297#_c_816_n
+ N_A_821_297#_c_817_n N_A_821_297#_c_818_n
+ PM_SKY130_FD_SC_HD__A2111OI_4%A_821_297#
x_PM_SKY130_FD_SC_HD__A2111OI_4%VPWR N_VPWR_M1018_s N_VPWR_M1033_s
+ N_VPWR_M1000_d N_VPWR_M1019_d N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n
+ N_VPWR_c_900_n N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n
+ N_VPWR_c_905_n N_VPWR_c_906_n N_VPWR_c_907_n VPWR N_VPWR_c_908_n
+ N_VPWR_c_896_n N_VPWR_c_910_n PM_SKY130_FD_SC_HD__A2111OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A2111OI_4%VGND N_VGND_M1007_d N_VGND_M1009_d
+ N_VGND_M1027_d N_VGND_M1010_s N_VGND_M1036_s N_VGND_M1002_s N_VGND_M1037_s
+ N_VGND_M1006_d N_VGND_M1024_d N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n
+ N_VGND_c_1030_n N_VGND_c_1031_n N_VGND_c_1032_n N_VGND_c_1033_n
+ N_VGND_c_1034_n N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n
+ N_VGND_c_1038_n N_VGND_c_1039_n VGND N_VGND_c_1040_n N_VGND_c_1041_n
+ N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n VGND
+ PM_SKY130_FD_SC_HD__A2111OI_4%VGND
x_PM_SKY130_FD_SC_HD__A2111OI_4%A_1205_47# N_A_1205_47#_M1017_d
+ N_A_1205_47#_M1020_d N_A_1205_47#_M1038_d N_A_1205_47#_M1022_s
+ N_A_1205_47#_M1039_s N_A_1205_47#_c_1202_n N_A_1205_47#_c_1210_n
+ N_A_1205_47#_c_1212_n N_A_1205_47#_c_1211_n N_A_1205_47#_c_1246_n
+ N_A_1205_47#_c_1203_n N_A_1205_47#_c_1204_n N_A_1205_47#_c_1223_n
+ PM_SKY130_FD_SC_HD__A2111OI_4%A_1205_47#
cc_1 VNB N_D1_c_132_n 0.0183006f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_D1_c_133_n 0.0159028f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_D1_c_134_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.995
cc_4 VNB N_D1_c_135_n 0.0169004f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=0.995
cc_5 VNB N_D1_c_136_n 0.00168995f $X=-0.19 $Y=-0.24 $X2=1.68 $Y2=1.16
cc_6 VNB N_D1_c_137_n 0.0661711f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_7 VNB N_C1_c_208_n 0.0169004f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_C1_c_209_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_9 VNB N_C1_c_210_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=1.985
cc_10 VNB N_C1_c_211_n 0.0173848f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.985
cc_11 VNB N_C1_c_212_n 0.0769621f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.147
cc_12 VNB N_C1_c_213_n 0.0033799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B1_c_293_n 0.0173848f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_14 VNB N_B1_c_294_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_15 VNB N_B1_c_295_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.995
cc_16 VNB N_B1_c_296_n 0.0211871f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=0.995
cc_17 VNB N_B1_c_297_n 0.00168995f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.147
cc_18 VNB N_B1_c_298_n 0.0892075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A1_c_376_n 0.0220814f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_20 VNB N_A1_c_377_n 0.0162054f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_21 VNB N_A1_c_378_n 0.0162054f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=1.985
cc_22 VNB N_A1_c_379_n 0.0172663f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.985
cc_23 VNB N_A1_c_380_n 0.00405118f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.147
cc_24 VNB N_A1_c_381_n 0.0761397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A2_c_448_n 0.0170672f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_26 VNB N_A2_c_449_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_27 VNB N_A2_c_450_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=1.985
cc_28 VNB N_A2_c_451_n 0.0218823f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.985
cc_29 VNB N_A2_c_452_n 0.0704371f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_30 VNB N_A2_c_453_n 0.0451522f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_31 VNB N_Y_c_581_n 0.00988648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB Y 0.0198674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_896_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_1027_n 0.0109397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_1028_n 0.0113283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_1029_n 3.06362e-19 $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_37 VNB N_VGND_c_1030_n 3.19317e-19 $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=1.16
cc_38 VNB N_VGND_c_1031_n 0.00435991f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_39 VNB N_VGND_c_1032_n 3.16793e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_1033_n 0.00499481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_1034_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_1035_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_1036_n 0.0567094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_1037_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_1038_n 0.0115005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_1039_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_1040_n 0.0115433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_1041_n 0.0119466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1042_n 0.0119466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1043_n 0.0145001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1044_n 0.0142196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1045_n 0.011798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1046_n 0.0198338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1047_n 0.476259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1048_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1049_n 0.00574824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1050_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1051_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1052_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1053_n 0.00516648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1205_47#_c_1202_n 0.00232422f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.56
cc_62 VNB N_A_1205_47#_c_1203_n 0.00744431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1205_47#_c_1204_n 0.012495f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_64 VPB N_D1_M1003_g 0.0219723f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_65 VPB N_D1_M1014_g 0.0186211f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_66 VPB N_D1_M1015_g 0.0186263f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_67 VPB N_D1_M1032_g 0.019013f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_68 VPB N_D1_c_137_n 0.0110908f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_69 VPB N_C1_M1005_g 0.019013f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_70 VPB N_C1_M1011_g 0.0186263f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_71 VPB N_C1_M1023_g 0.0186263f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.56
cc_72 VPB N_C1_M1028_g 0.0258394f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_73 VPB N_C1_c_212_n 0.0194745f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.147
cc_74 VPB N_B1_M1012_g 0.0258394f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_75 VPB N_B1_M1013_g 0.0186263f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_76 VPB N_B1_M1025_g 0.018625f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_77 VPB N_B1_M1031_g 0.0191108f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_78 VPB N_B1_c_298_n 0.0225399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A1_M1018_g 0.0185528f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_80 VPB N_A1_M1026_g 0.0181805f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_81 VPB N_A1_M1033_g 0.0184149f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.56
cc_82 VPB N_A1_M1035_g 0.019898f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_83 VPB N_A1_c_381_n 0.0172641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A2_M1000_g 0.0196662f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_85 VPB N_A2_M1004_g 0.0191741f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_86 VPB N_A2_M1019_g 0.0191741f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.56
cc_87 VPB N_A2_M1030_g 0.0249657f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_88 VPB N_A2_c_452_n 0.015514f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_89 VPB N_A2_c_453_n 0.0181664f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_90 VPB N_A_28_297#_c_518_n 0.00831299f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.56
cc_91 VPB N_A_28_297#_c_519_n 0.0173377f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.325
cc_92 VPB N_A_28_297#_c_520_n 0.00206763f $X=-0.19 $Y=1.305 $X2=1.68 $Y2=1.16
cc_93 VPB N_A_28_297#_c_521_n 0.00422673f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_94 VPB N_Y_c_583_n 0.00290608f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_95 VPB N_Y_c_584_n 4.36864e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_Y_c_585_n 0.00238451f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_97 VPB N_Y_c_586_n 0.00242529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_587_n 0.00242529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB Y 0.00787544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_455_297#_c_738_n 0.00238451f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.995
cc_101 VPB N_A_455_297#_c_739_n 0.0203254f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_102 VPB N_A_455_297#_c_740_n 0.00238451f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_103 VPB N_A_455_297#_c_741_n 0.00242529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_455_297#_c_742_n 0.00242529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_455_297#_c_743_n 0.00242529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_455_297#_c_744_n 0.00257664f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_107 VPB N_A_821_297#_c_808_n 0.00206763f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.995
cc_108 VPB N_A_821_297#_c_809_n 0.00413519f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_109 VPB N_A_821_297#_c_810_n 0.00338003f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.16
cc_110 VPB N_A_821_297#_c_811_n 0.00372869f $X=-0.19 $Y=1.305 $X2=1.68 $Y2=1.16
cc_111 VPB N_A_821_297#_c_812_n 0.00290574f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.147
cc_112 VPB N_A_821_297#_c_813_n 0.00339073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_821_297#_c_814_n 0.0139575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_821_297#_c_815_n 0.0217206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_821_297#_c_816_n 0.001447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_821_297#_c_817_n 0.00717074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_821_297#_c_818_n 0.00180864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_897_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.995
cc_119 VPB N_VPWR_c_898_n 0.01339f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.56
cc_120 VPB N_VPWR_c_899_n 3.31161e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_900_n 3.46032e-19 $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.325
cc_122 VPB N_VPWR_c_901_n 4.14e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_123 VPB N_VPWR_c_902_n 0.146989f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_124 VPB N_VPWR_c_903_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_904_n 0.0168633f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_126 VPB N_VPWR_c_905_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_127 VPB N_VPWR_c_906_n 0.0158499f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_128 VPB N_VPWR_c_907_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.16
cc_129 VPB N_VPWR_c_908_n 0.0237833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_896_n 0.0647233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_910_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 N_D1_M1032_g N_C1_M1005_g 0.0282574f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_133 N_D1_c_135_n N_C1_c_208_n 0.0251544f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_134 N_D1_c_136_n N_C1_c_212_n 3.13866e-19 $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_135 N_D1_c_137_n N_C1_c_212_n 0.0229865f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_136 N_D1_c_136_n N_C1_c_213_n 0.0180521f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_137 N_D1_c_137_n N_C1_c_213_n 3.13866e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_138 N_D1_M1003_g N_A_28_297#_c_522_n 0.0100325f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_139 N_D1_M1014_g N_A_28_297#_c_522_n 0.00994206f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_140 N_D1_M1015_g N_A_28_297#_c_524_n 0.00994206f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_141 N_D1_M1032_g N_A_28_297#_c_524_n 0.012231f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_142 N_D1_M1003_g N_Y_c_583_n 0.0134271f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_143 N_D1_c_136_n N_Y_c_583_n 0.00212907f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_144 N_D1_c_133_n N_Y_c_591_n 0.0098261f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_145 N_D1_c_134_n N_Y_c_591_n 0.0098261f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_146 N_D1_c_136_n N_Y_c_591_n 0.0312007f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_147 N_D1_c_137_n N_Y_c_591_n 0.00221013f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_148 N_D1_M1014_g N_Y_c_585_n 0.0101046f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_149 N_D1_M1015_g N_Y_c_585_n 0.0101046f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_150 N_D1_c_136_n N_Y_c_585_n 0.034118f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_151 N_D1_c_137_n N_Y_c_585_n 0.00234522f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_152 N_D1_c_135_n N_Y_c_599_n 0.010254f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_153 N_D1_c_136_n N_Y_c_599_n 0.00932844f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_154 N_D1_M1003_g N_Y_c_586_n 0.0117535f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_155 N_D1_M1014_g N_Y_c_586_n 0.00655853f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_156 N_D1_M1015_g N_Y_c_586_n 4.99919e-19 $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_157 N_D1_c_136_n N_Y_c_586_n 0.0237666f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_158 N_D1_c_137_n N_Y_c_586_n 0.00246427f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_159 N_D1_c_132_n N_Y_c_606_n 0.0133602f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_160 N_D1_c_136_n N_Y_c_606_n 0.0149269f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_161 N_D1_c_137_n N_Y_c_606_n 0.00203131f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_162 N_D1_M1014_g N_Y_c_587_n 4.99919e-19 $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_163 N_D1_M1015_g N_Y_c_587_n 0.00656102f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_164 N_D1_M1032_g N_Y_c_587_n 0.00975779f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_165 N_D1_c_136_n N_Y_c_587_n 0.0237666f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_166 N_D1_c_137_n N_Y_c_587_n 0.00242396f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_167 N_D1_c_136_n N_Y_c_614_n 0.0105162f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_168 N_D1_c_137_n N_Y_c_614_n 0.00225701f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_169 N_D1_c_132_n Y 0.00778975f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_170 N_D1_c_136_n Y 0.0198164f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_171 N_D1_c_137_n Y 0.0165154f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_172 N_D1_M1032_g N_A_455_297#_c_741_n 0.00111563f $X=1.77 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_D1_M1003_g N_VPWR_c_902_n 0.00362032f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_174 N_D1_M1014_g N_VPWR_c_902_n 0.00362032f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_175 N_D1_M1015_g N_VPWR_c_902_n 0.00362032f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_176 N_D1_M1032_g N_VPWR_c_902_n 0.00362032f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_177 N_D1_M1003_g N_VPWR_c_896_n 0.00622166f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_178 N_D1_M1014_g N_VPWR_c_896_n 0.00528435f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_179 N_D1_M1015_g N_VPWR_c_896_n 0.00528435f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_180 N_D1_M1032_g N_VPWR_c_896_n 0.00530968f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_181 N_D1_c_132_n N_VGND_c_1028_n 0.00888944f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_182 N_D1_c_133_n N_VGND_c_1028_n 0.00100453f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_183 N_D1_c_132_n N_VGND_c_1029_n 9.93364e-19 $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_184 N_D1_c_133_n N_VGND_c_1029_n 0.00755691f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_185 N_D1_c_134_n N_VGND_c_1029_n 0.00765006f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_186 N_D1_c_135_n N_VGND_c_1029_n 0.00100064f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_187 N_D1_c_132_n N_VGND_c_1040_n 0.00337001f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_188 N_D1_c_133_n N_VGND_c_1040_n 0.00351072f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_189 N_D1_c_134_n N_VGND_c_1041_n 0.00351072f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_190 N_D1_c_135_n N_VGND_c_1041_n 0.0035176f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_191 N_D1_c_132_n N_VGND_c_1047_n 0.00394833f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_192 N_D1_c_133_n N_VGND_c_1047_n 0.00408938f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_193 N_D1_c_134_n N_VGND_c_1047_n 0.00411677f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_194 N_D1_c_135_n N_VGND_c_1047_n 0.00411682f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_195 N_D1_c_134_n N_VGND_c_1049_n 0.00100466f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_196 N_D1_c_135_n N_VGND_c_1049_n 0.010976f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_197 N_C1_c_211_n N_B1_c_293_n 0.0227346f $X=3.57 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_198 N_C1_c_212_n N_B1_c_297_n 3.13866e-19 $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_199 N_C1_c_213_n N_B1_c_297_n 0.0180521f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_200 N_C1_c_212_n N_B1_c_298_n 0.0229865f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_201 N_C1_c_213_n N_B1_c_298_n 3.13866e-19 $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_202 N_C1_c_212_n N_A_28_297#_c_526_n 3.92719e-19 $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_203 N_C1_c_213_n N_A_28_297#_c_526_n 5.43064e-19 $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_204 N_C1_M1005_g N_A_28_297#_c_528_n 0.012231f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_205 N_C1_M1011_g N_A_28_297#_c_528_n 0.00994206f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_206 N_C1_M1023_g N_A_28_297#_c_530_n 0.00994206f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_207 N_C1_M1028_g N_A_28_297#_c_530_n 0.0100325f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_208 N_C1_c_208_n N_Y_c_599_n 0.010254f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_209 N_C1_c_212_n N_Y_c_599_n 0.00346164f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_210 N_C1_c_213_n N_Y_c_599_n 0.0161647f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_211 N_C1_c_209_n N_Y_c_622_n 0.0098261f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_212 N_C1_c_210_n N_Y_c_622_n 0.0098261f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_213 N_C1_c_212_n N_Y_c_622_n 0.00251203f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_214 N_C1_c_213_n N_Y_c_622_n 0.0312007f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_215 N_C1_c_211_n N_Y_c_626_n 0.0103625f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_216 N_C1_c_212_n N_Y_c_626_n 0.00205467f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_217 N_C1_c_213_n N_Y_c_626_n 0.0113056f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_218 N_C1_M1005_g N_Y_c_587_n 0.00111563f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_219 N_C1_c_212_n N_Y_c_630_n 0.00255924f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_220 N_C1_c_213_n N_Y_c_630_n 0.0105162f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_221 N_C1_c_211_n N_Y_c_632_n 0.00430183f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_222 N_C1_c_212_n N_Y_c_632_n 0.00255924f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_223 N_C1_c_213_n N_Y_c_632_n 0.0125709f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_224 N_C1_c_211_n N_Y_c_635_n 5.62912e-19 $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_225 N_C1_M1011_g N_A_455_297#_c_738_n 0.0101046f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_226 N_C1_M1023_g N_A_455_297#_c_738_n 0.0101046f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_227 N_C1_c_212_n N_A_455_297#_c_738_n 0.00266731f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_228 N_C1_c_213_n N_A_455_297#_c_738_n 0.034118f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_229 N_C1_M1028_g N_A_455_297#_c_739_n 0.0116119f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_230 N_C1_c_212_n N_A_455_297#_c_739_n 0.004526f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_231 N_C1_c_213_n N_A_455_297#_c_739_n 0.0194763f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_232 N_C1_M1005_g N_A_455_297#_c_741_n 0.00975779f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_233 N_C1_M1011_g N_A_455_297#_c_741_n 0.00656102f $X=2.63 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_C1_M1023_g N_A_455_297#_c_741_n 4.99919e-19 $X=3.06 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_C1_c_212_n N_A_455_297#_c_741_n 0.0027464f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_236 N_C1_c_213_n N_A_455_297#_c_741_n 0.0237666f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_237 N_C1_M1011_g N_A_455_297#_c_742_n 4.99919e-19 $X=2.63 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_C1_M1023_g N_A_455_297#_c_742_n 0.00656102f $X=3.06 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_C1_M1028_g N_A_455_297#_c_742_n 0.0117535f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_240 N_C1_c_212_n N_A_455_297#_c_742_n 0.0027464f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_241 N_C1_c_213_n N_A_455_297#_c_742_n 0.0237666f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_242 N_C1_M1005_g N_VPWR_c_902_n 0.00362032f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_243 N_C1_M1011_g N_VPWR_c_902_n 0.00362032f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_244 N_C1_M1023_g N_VPWR_c_902_n 0.00362032f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_245 N_C1_M1028_g N_VPWR_c_902_n 0.00362032f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_246 N_C1_M1005_g N_VPWR_c_896_n 0.00530968f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_247 N_C1_M1011_g N_VPWR_c_896_n 0.00528435f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_248 N_C1_M1023_g N_VPWR_c_896_n 0.00528435f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_249 N_C1_M1028_g N_VPWR_c_896_n 0.00658404f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_250 N_C1_c_208_n N_VGND_c_1030_n 0.00100064f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_251 N_C1_c_209_n N_VGND_c_1030_n 0.00765006f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_252 N_C1_c_210_n N_VGND_c_1030_n 0.00796708f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_253 N_C1_c_211_n N_VGND_c_1030_n 0.00103817f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_254 N_C1_c_211_n N_VGND_c_1031_n 0.00291058f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_255 N_C1_c_208_n N_VGND_c_1042_n 0.0035176f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_256 N_C1_c_209_n N_VGND_c_1042_n 0.00351072f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_257 N_C1_c_210_n N_VGND_c_1043_n 0.00351072f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_258 N_C1_c_211_n N_VGND_c_1043_n 0.00420764f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_259 N_C1_c_208_n N_VGND_c_1047_n 0.00411682f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_260 N_C1_c_209_n N_VGND_c_1047_n 0.00411677f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_261 N_C1_c_210_n N_VGND_c_1047_n 0.00411677f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_262 N_C1_c_211_n N_VGND_c_1047_n 0.00595561f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_263 N_C1_c_208_n N_VGND_c_1049_n 0.00794284f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_264 N_C1_c_209_n N_VGND_c_1049_n 0.00100466f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B1_M1031_g N_A1_M1018_g 0.0194752f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B1_c_297_n N_A1_c_380_n 0.00976766f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B1_c_298_n N_A1_c_380_n 0.00122736f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B1_c_297_n N_A1_c_381_n 2.53861e-19 $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B1_c_298_n N_A1_c_381_n 0.0194752f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B1_c_293_n N_Y_c_626_n 0.0109052f $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B1_c_297_n N_Y_c_626_n 0.0107168f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_298_n N_Y_c_626_n 0.00161264f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B1_c_294_n N_Y_c_639_n 0.0098261f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B1_c_295_n N_Y_c_639_n 0.0098261f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B1_c_297_n N_Y_c_639_n 0.0312007f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B1_c_298_n N_Y_c_639_n 0.00258751f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_277 N_B1_c_296_n N_Y_c_581_n 0.0118691f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B1_c_297_n N_Y_c_581_n 0.0177149f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_279 N_B1_c_298_n N_Y_c_581_n 0.0101953f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B1_c_293_n N_Y_c_632_n 3.36045e-19 $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B1_c_293_n N_Y_c_635_n 0.00359681f $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B1_c_297_n N_Y_c_635_n 0.0120005f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_283 N_B1_c_298_n N_Y_c_635_n 0.00229479f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_284 N_B1_c_297_n N_Y_c_650_n 0.0103765f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B1_c_298_n N_Y_c_650_n 0.00263479f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B1_M1012_g N_A_455_297#_c_739_n 0.0116119f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_287 N_B1_c_297_n N_A_455_297#_c_739_n 0.0345481f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_288 N_B1_c_298_n N_A_455_297#_c_739_n 0.0105418f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B1_M1013_g N_A_455_297#_c_740_n 0.0101046f $X=4.87 $Y=1.985 $X2=0 $Y2=0
cc_290 N_B1_M1025_g N_A_455_297#_c_740_n 0.0101656f $X=5.3 $Y=1.985 $X2=0 $Y2=0
cc_291 N_B1_c_297_n N_A_455_297#_c_740_n 0.034118f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_298_n N_A_455_297#_c_740_n 0.00274783f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_293 N_B1_M1012_g N_A_455_297#_c_743_n 0.0117535f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_294 N_B1_M1013_g N_A_455_297#_c_743_n 0.00656102f $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_B1_M1025_g N_A_455_297#_c_743_n 4.99919e-19 $X=5.3 $Y=1.985 $X2=0 $Y2=0
cc_296 N_B1_c_297_n N_A_455_297#_c_743_n 0.0237666f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_297 N_B1_c_298_n N_A_455_297#_c_743_n 0.00282701f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_298 N_B1_M1013_g N_A_455_297#_c_744_n 4.99919e-19 $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_B1_M1025_g N_A_455_297#_c_744_n 0.00658023f $X=5.3 $Y=1.985 $X2=0 $Y2=0
cc_300 N_B1_M1031_g N_A_455_297#_c_744_n 0.00791191f $X=5.73 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_B1_c_297_n N_A_455_297#_c_744_n 0.0216987f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_302 N_B1_c_298_n N_A_455_297#_c_744_n 0.00246427f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_303 N_B1_M1012_g N_A_821_297#_c_819_n 0.0100272f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_304 N_B1_M1013_g N_A_821_297#_c_819_n 0.00994206f $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_B1_M1025_g N_A_821_297#_c_821_n 0.00943721f $X=5.3 $Y=1.985 $X2=0 $Y2=0
cc_306 N_B1_M1031_g N_A_821_297#_c_821_n 0.0116577f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_307 N_B1_M1031_g N_A_821_297#_c_811_n 0.00103319f $X=5.73 $Y=1.985 $X2=0
+ $Y2=0
cc_308 N_B1_M1031_g N_VPWR_c_897_n 0.00113191f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_309 N_B1_M1012_g N_VPWR_c_902_n 0.00362032f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_310 N_B1_M1013_g N_VPWR_c_902_n 0.00362032f $X=4.87 $Y=1.985 $X2=0 $Y2=0
cc_311 N_B1_M1025_g N_VPWR_c_902_n 0.00362032f $X=5.3 $Y=1.985 $X2=0 $Y2=0
cc_312 N_B1_M1031_g N_VPWR_c_902_n 0.00362032f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_313 N_B1_M1012_g N_VPWR_c_896_n 0.00658404f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_314 N_B1_M1013_g N_VPWR_c_896_n 0.00528435f $X=4.87 $Y=1.985 $X2=0 $Y2=0
cc_315 N_B1_M1025_g N_VPWR_c_896_n 0.00528435f $X=5.3 $Y=1.985 $X2=0 $Y2=0
cc_316 N_B1_M1031_g N_VPWR_c_896_n 0.00537559f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_317 N_B1_c_293_n N_VGND_c_1031_n 0.00172216f $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_293_n N_VGND_c_1032_n 0.00103201f $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B1_c_294_n N_VGND_c_1032_n 0.00791591f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_320 N_B1_c_295_n N_VGND_c_1032_n 0.00762255f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B1_c_296_n N_VGND_c_1032_n 9.97443e-19 $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B1_c_295_n N_VGND_c_1033_n 0.00100884f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B1_c_296_n N_VGND_c_1033_n 0.0089652f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B1_c_293_n N_VGND_c_1044_n 0.00422505f $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_325 N_B1_c_294_n N_VGND_c_1044_n 0.00351072f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B1_c_295_n N_VGND_c_1045_n 0.00351072f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B1_c_296_n N_VGND_c_1045_n 0.00337001f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B1_c_293_n N_VGND_c_1047_n 0.00585788f $X=4.11 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B1_c_294_n N_VGND_c_1047_n 0.00411677f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B1_c_295_n N_VGND_c_1047_n 0.00411677f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B1_c_296_n N_VGND_c_1047_n 0.00397572f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A1_M1035_g N_A2_M1000_g 0.0245668f $X=7.48 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A1_c_379_n N_A2_c_448_n 0.0224354f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A1_c_380_n N_A2_c_452_n 0.00102338f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A1_c_381_n N_A2_c_452_n 0.0233834f $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A1_c_380_n N_A2_c_464_n 0.0176471f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A1_c_381_n N_A2_c_464_n 3.1084e-19 $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A1_c_376_n N_Y_c_581_n 0.0108392f $X=6.38 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A1_c_377_n N_Y_c_581_n 0.00879865f $X=6.81 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A1_c_378_n N_Y_c_581_n 0.00879865f $X=7.24 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A1_c_379_n N_Y_c_581_n 0.00281687f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A1_c_380_n N_Y_c_581_n 0.0734043f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A1_c_381_n N_Y_c_581_n 0.0130408f $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A1_M1018_g N_A_821_297#_c_810_n 0.0126379f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A1_M1026_g N_A_821_297#_c_810_n 0.0126841f $X=6.6 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A1_c_380_n N_A_821_297#_c_810_n 0.0449067f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A1_c_381_n N_A_821_297#_c_810_n 0.00279407f $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A1_M1033_g N_A_821_297#_c_812_n 0.0128702f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A1_M1035_g N_A_821_297#_c_812_n 0.0135353f $X=7.48 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A1_c_380_n N_A_821_297#_c_812_n 0.0481855f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A1_c_381_n N_A_821_297#_c_812_n 0.00404898f $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A1_c_380_n N_A_821_297#_c_816_n 0.015747f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A1_c_381_n N_A_821_297#_c_816_n 0.00289127f $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A1_c_380_n N_A_821_297#_c_817_n 0.013673f $X=7.55 $Y=1.16 $X2=0 $Y2=0
cc_355 N_A1_c_381_n N_A_821_297#_c_817_n 0.00477059f $X=7.67 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A1_M1018_g N_VPWR_c_897_n 0.0134872f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A1_M1026_g N_VPWR_c_897_n 0.0132743f $X=6.6 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A1_M1033_g N_VPWR_c_897_n 0.00107604f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A1_M1026_g N_VPWR_c_898_n 0.00486043f $X=6.6 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A1_M1033_g N_VPWR_c_898_n 0.00486043f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A1_M1026_g N_VPWR_c_899_n 0.00107038f $X=6.6 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A1_M1033_g N_VPWR_c_899_n 0.0132414f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A1_M1035_g N_VPWR_c_899_n 0.0121529f $X=7.48 $Y=1.985 $X2=0 $Y2=0
cc_364 N_A1_M1035_g N_VPWR_c_900_n 0.00101684f $X=7.48 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A1_M1018_g N_VPWR_c_902_n 0.00486043f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A1_M1035_g N_VPWR_c_904_n 0.00564095f $X=7.48 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A1_M1018_g N_VPWR_c_896_n 0.00835349f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A1_M1026_g N_VPWR_c_896_n 0.00830219f $X=6.6 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A1_M1033_g N_VPWR_c_896_n 0.00830219f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_370 N_A1_M1035_g N_VPWR_c_896_n 0.00982899f $X=7.48 $Y=1.985 $X2=0 $Y2=0
cc_371 N_A1_c_376_n N_VGND_c_1033_n 0.00251113f $X=6.38 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A1_c_379_n N_VGND_c_1034_n 0.00119703f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A1_c_376_n N_VGND_c_1036_n 0.00362032f $X=6.38 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A1_c_377_n N_VGND_c_1036_n 0.00362032f $X=6.81 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A1_c_378_n N_VGND_c_1036_n 0.00362032f $X=7.24 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A1_c_379_n N_VGND_c_1036_n 0.00362032f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A1_c_376_n N_VGND_c_1047_n 0.00658404f $X=6.38 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A1_c_377_n N_VGND_c_1047_n 0.00528435f $X=6.81 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A1_c_378_n N_VGND_c_1047_n 0.00528435f $X=7.24 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A1_c_379_n N_VGND_c_1047_n 0.00557067f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A1_c_376_n N_A_1205_47#_c_1202_n 0.00782153f $X=6.38 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A1_c_377_n N_A_1205_47#_c_1202_n 0.00782153f $X=6.81 $Y=0.995 $X2=0
+ $Y2=0
cc_383 N_A1_c_378_n N_A_1205_47#_c_1202_n 0.00782153f $X=7.24 $Y=0.995 $X2=0
+ $Y2=0
cc_384 N_A1_c_379_n N_A_1205_47#_c_1202_n 0.0116522f $X=7.67 $Y=0.995 $X2=0
+ $Y2=0
cc_385 N_A1_c_380_n N_A_1205_47#_c_1202_n 0.00320389f $X=7.55 $Y=1.16 $X2=0
+ $Y2=0
cc_386 N_A1_c_379_n N_A_1205_47#_c_1210_n 0.00386499f $X=7.67 $Y=0.995 $X2=0
+ $Y2=0
cc_387 N_A1_c_379_n N_A_1205_47#_c_1211_n 0.00164103f $X=7.67 $Y=0.995 $X2=0
+ $Y2=0
cc_388 N_A2_M1000_g N_A_821_297#_c_813_n 0.0172236f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_389 N_A2_M1004_g N_A_821_297#_c_813_n 0.0150755f $X=8.46 $Y=1.985 $X2=0 $Y2=0
cc_390 N_A2_c_452_n N_A_821_297#_c_813_n 0.00280754f $X=9.56 $Y=1.16 $X2=0 $Y2=0
cc_391 N_A2_c_464_n N_A_821_297#_c_813_n 0.0456123f $X=8.125 $Y=1.16 $X2=0 $Y2=0
cc_392 N_A2_M1019_g N_A_821_297#_c_814_n 0.0151745f $X=8.98 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A2_M1030_g N_A_821_297#_c_814_n 0.0156575f $X=9.41 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A2_c_452_n N_A_821_297#_c_814_n 0.0100051f $X=9.56 $Y=1.16 $X2=0 $Y2=0
cc_395 N_A2_c_464_n N_A_821_297#_c_814_n 0.070956f $X=8.125 $Y=1.16 $X2=0 $Y2=0
cc_396 N_A2_c_452_n N_A_821_297#_c_818_n 0.00538582f $X=9.56 $Y=1.16 $X2=0 $Y2=0
cc_397 N_A2_c_464_n N_A_821_297#_c_818_n 0.0216546f $X=8.125 $Y=1.16 $X2=0 $Y2=0
cc_398 N_A2_M1000_g N_VPWR_c_899_n 0.00100501f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_399 N_A2_M1000_g N_VPWR_c_900_n 0.0120718f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A2_M1004_g N_VPWR_c_900_n 0.0120394f $X=8.46 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A2_M1019_g N_VPWR_c_900_n 0.0010788f $X=8.98 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A2_M1004_g N_VPWR_c_901_n 0.00108355f $X=8.46 $Y=1.985 $X2=0 $Y2=0
cc_403 N_A2_M1019_g N_VPWR_c_901_n 0.0120258f $X=8.98 $Y=1.985 $X2=0 $Y2=0
cc_404 N_A2_M1030_g N_VPWR_c_901_n 0.0185012f $X=9.41 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A2_M1000_g N_VPWR_c_904_n 0.00486043f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_406 N_A2_M1004_g N_VPWR_c_906_n 0.00486043f $X=8.46 $Y=1.985 $X2=0 $Y2=0
cc_407 N_A2_M1019_g N_VPWR_c_906_n 0.00486043f $X=8.98 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A2_M1030_g N_VPWR_c_908_n 0.00486043f $X=9.41 $Y=1.985 $X2=0 $Y2=0
cc_409 N_A2_M1000_g N_VPWR_c_896_n 0.00860044f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_410 N_A2_M1004_g N_VPWR_c_896_n 0.00852643f $X=8.46 $Y=1.985 $X2=0 $Y2=0
cc_411 N_A2_M1019_g N_VPWR_c_896_n 0.00852643f $X=8.98 $Y=1.985 $X2=0 $Y2=0
cc_412 N_A2_M1030_g N_VPWR_c_896_n 0.00943606f $X=9.41 $Y=1.985 $X2=0 $Y2=0
cc_413 N_A2_c_448_n N_VGND_c_1034_n 0.00762713f $X=8.195 $Y=0.995 $X2=0 $Y2=0
cc_414 N_A2_c_449_n N_VGND_c_1034_n 0.00658529f $X=8.625 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A2_c_450_n N_VGND_c_1034_n 6.58014e-19 $X=9.055 $Y=0.995 $X2=0 $Y2=0
cc_416 N_A2_c_449_n N_VGND_c_1035_n 6.58014e-19 $X=8.625 $Y=0.995 $X2=0 $Y2=0
cc_417 N_A2_c_450_n N_VGND_c_1035_n 0.00658529f $X=9.055 $Y=0.995 $X2=0 $Y2=0
cc_418 N_A2_c_451_n N_VGND_c_1035_n 0.00903352f $X=9.485 $Y=0.995 $X2=0 $Y2=0
cc_419 N_A2_c_448_n N_VGND_c_1036_n 0.00351072f $X=8.195 $Y=0.995 $X2=0 $Y2=0
cc_420 N_A2_c_449_n N_VGND_c_1038_n 0.00351072f $X=8.625 $Y=0.995 $X2=0 $Y2=0
cc_421 N_A2_c_450_n N_VGND_c_1038_n 0.00351072f $X=9.055 $Y=0.995 $X2=0 $Y2=0
cc_422 N_A2_c_451_n N_VGND_c_1046_n 0.00351072f $X=9.485 $Y=0.995 $X2=0 $Y2=0
cc_423 N_A2_c_448_n N_VGND_c_1047_n 0.00436315f $X=8.195 $Y=0.995 $X2=0 $Y2=0
cc_424 N_A2_c_449_n N_VGND_c_1047_n 0.00411677f $X=8.625 $Y=0.995 $X2=0 $Y2=0
cc_425 N_A2_c_450_n N_VGND_c_1047_n 0.00411677f $X=9.055 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A2_c_451_n N_VGND_c_1047_n 0.00521005f $X=9.485 $Y=0.995 $X2=0 $Y2=0
cc_427 N_A2_c_448_n N_A_1205_47#_c_1212_n 0.0107826f $X=8.195 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A2_c_449_n N_A_1205_47#_c_1212_n 0.0107877f $X=8.625 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_A2_c_452_n N_A_1205_47#_c_1212_n 0.00258646f $X=9.56 $Y=1.16 $X2=0
+ $Y2=0
cc_430 N_A2_c_464_n N_A_1205_47#_c_1212_n 0.0313807f $X=8.125 $Y=1.16 $X2=0
+ $Y2=0
cc_431 N_A2_c_452_n N_A_1205_47#_c_1211_n 0.00318766f $X=9.56 $Y=1.16 $X2=0
+ $Y2=0
cc_432 N_A2_c_464_n N_A_1205_47#_c_1211_n 0.00666045f $X=8.125 $Y=1.16 $X2=0
+ $Y2=0
cc_433 N_A2_c_450_n N_A_1205_47#_c_1203_n 0.0108343f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_434 N_A2_c_451_n N_A_1205_47#_c_1203_n 0.0114867f $X=9.485 $Y=0.995 $X2=0
+ $Y2=0
cc_435 N_A2_c_452_n N_A_1205_47#_c_1203_n 0.00249211f $X=9.56 $Y=1.16 $X2=0
+ $Y2=0
cc_436 N_A2_c_453_n N_A_1205_47#_c_1203_n 0.00590339f $X=9.825 $Y=1.16 $X2=0
+ $Y2=0
cc_437 N_A2_c_464_n N_A_1205_47#_c_1203_n 0.0470987f $X=8.125 $Y=1.16 $X2=0
+ $Y2=0
cc_438 N_A2_c_452_n N_A_1205_47#_c_1223_n 0.00256816f $X=9.56 $Y=1.16 $X2=0
+ $Y2=0
cc_439 N_A2_c_464_n N_A_1205_47#_c_1223_n 0.0109235f $X=8.125 $Y=1.16 $X2=0
+ $Y2=0
cc_440 N_A_28_297#_c_522_n N_Y_M1003_s 0.00340502f $X=1.03 $Y=2.35 $X2=0 $Y2=0
cc_441 N_A_28_297#_c_524_n N_Y_M1015_s 0.00340502f $X=1.89 $Y=2.35 $X2=0 $Y2=0
cc_442 N_A_28_297#_M1003_d N_Y_c_583_n 2.94505e-19 $X=0.14 $Y=1.485 $X2=0 $Y2=0
cc_443 N_A_28_297#_c_519_n N_Y_c_583_n 0.00213663f $X=0.265 $Y=2 $X2=0 $Y2=0
cc_444 N_A_28_297#_c_522_n N_Y_c_583_n 0.0030004f $X=1.03 $Y=2.35 $X2=0 $Y2=0
cc_445 N_A_28_297#_M1003_d N_Y_c_584_n 0.0104056f $X=0.14 $Y=1.485 $X2=0 $Y2=0
cc_446 N_A_28_297#_c_519_n N_Y_c_584_n 0.0149932f $X=0.265 $Y=2 $X2=0 $Y2=0
cc_447 N_A_28_297#_M1014_d N_Y_c_585_n 0.00177615f $X=0.985 $Y=1.485 $X2=0 $Y2=0
cc_448 N_A_28_297#_c_522_n N_Y_c_585_n 0.00318184f $X=1.03 $Y=2.35 $X2=0 $Y2=0
cc_449 N_A_28_297#_c_541_p N_Y_c_585_n 0.0135452f $X=1.125 $Y=2.02 $X2=0 $Y2=0
cc_450 N_A_28_297#_c_524_n N_Y_c_585_n 0.00318184f $X=1.89 $Y=2.35 $X2=0 $Y2=0
cc_451 N_A_28_297#_c_522_n N_Y_c_586_n 0.0161241f $X=1.03 $Y=2.35 $X2=0 $Y2=0
cc_452 N_A_28_297#_c_524_n N_Y_c_587_n 0.0161241f $X=1.89 $Y=2.35 $X2=0 $Y2=0
cc_453 N_A_28_297#_c_528_n N_A_455_297#_M1005_s 0.00340502f $X=2.75 $Y=2.35
+ $X2=-0.19 $Y2=1.305
cc_454 N_A_28_297#_c_530_n N_A_455_297#_M1023_s 0.00340502f $X=3.61 $Y=2.35
+ $X2=0 $Y2=0
cc_455 N_A_28_297#_M1011_d N_A_455_297#_c_738_n 0.00177615f $X=2.705 $Y=1.485
+ $X2=0 $Y2=0
cc_456 N_A_28_297#_c_528_n N_A_455_297#_c_738_n 0.00318184f $X=2.75 $Y=2.35
+ $X2=0 $Y2=0
cc_457 N_A_28_297#_c_549_p N_A_455_297#_c_738_n 0.0135452f $X=2.845 $Y=2.02
+ $X2=0 $Y2=0
cc_458 N_A_28_297#_c_530_n N_A_455_297#_c_738_n 0.00318184f $X=3.61 $Y=2.35
+ $X2=0 $Y2=0
cc_459 N_A_28_297#_M1028_d N_A_455_297#_c_739_n 0.00296258f $X=3.565 $Y=1.485
+ $X2=0 $Y2=0
cc_460 N_A_28_297#_c_530_n N_A_455_297#_c_739_n 0.0030004f $X=3.61 $Y=2.35 $X2=0
+ $Y2=0
cc_461 N_A_28_297#_c_521_n N_A_455_297#_c_739_n 0.0192968f $X=3.7 $Y=2 $X2=0
+ $Y2=0
cc_462 N_A_28_297#_c_528_n N_A_455_297#_c_741_n 0.0161241f $X=2.75 $Y=2.35 $X2=0
+ $Y2=0
cc_463 N_A_28_297#_c_530_n N_A_455_297#_c_742_n 0.0161241f $X=3.61 $Y=2.35 $X2=0
+ $Y2=0
cc_464 N_A_28_297#_c_520_n N_A_821_297#_c_808_n 0.016447f $X=3.74 $Y=2.255 $X2=0
+ $Y2=0
cc_465 N_A_28_297#_c_521_n N_A_821_297#_c_809_n 0.0311202f $X=3.7 $Y=2 $X2=0
+ $Y2=0
cc_466 N_A_28_297#_c_518_n N_VPWR_c_902_n 0.0157654f $X=0.23 $Y=2.255 $X2=0
+ $Y2=0
cc_467 N_A_28_297#_c_522_n N_VPWR_c_902_n 0.032265f $X=1.03 $Y=2.35 $X2=0 $Y2=0
cc_468 N_A_28_297#_c_524_n N_VPWR_c_902_n 0.032265f $X=1.89 $Y=2.35 $X2=0 $Y2=0
cc_469 N_A_28_297#_c_528_n N_VPWR_c_902_n 0.032265f $X=2.75 $Y=2.35 $X2=0 $Y2=0
cc_470 N_A_28_297#_c_530_n N_VPWR_c_902_n 0.032265f $X=3.61 $Y=2.35 $X2=0 $Y2=0
cc_471 N_A_28_297#_c_520_n N_VPWR_c_902_n 0.0157719f $X=3.74 $Y=2.255 $X2=0
+ $Y2=0
cc_472 N_A_28_297#_c_564_p N_VPWR_c_902_n 0.0109994f $X=1.125 $Y=2.36 $X2=0
+ $Y2=0
cc_473 N_A_28_297#_c_565_p N_VPWR_c_902_n 0.0109994f $X=1.985 $Y=2.36 $X2=0
+ $Y2=0
cc_474 N_A_28_297#_c_566_p N_VPWR_c_902_n 0.0109994f $X=2.845 $Y=2.36 $X2=0
+ $Y2=0
cc_475 N_A_28_297#_M1003_d N_VPWR_c_896_n 0.00214249f $X=0.14 $Y=1.485 $X2=0
+ $Y2=0
cc_476 N_A_28_297#_M1014_d N_VPWR_c_896_n 0.00224115f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_477 N_A_28_297#_M1032_d N_VPWR_c_896_n 0.00224115f $X=1.845 $Y=1.485 $X2=0
+ $Y2=0
cc_478 N_A_28_297#_M1011_d N_VPWR_c_896_n 0.00224115f $X=2.705 $Y=1.485 $X2=0
+ $Y2=0
cc_479 N_A_28_297#_M1028_d N_VPWR_c_896_n 0.00210134f $X=3.565 $Y=1.485 $X2=0
+ $Y2=0
cc_480 N_A_28_297#_c_518_n N_VPWR_c_896_n 0.00988695f $X=0.23 $Y=2.255 $X2=0
+ $Y2=0
cc_481 N_A_28_297#_c_522_n N_VPWR_c_896_n 0.0231894f $X=1.03 $Y=2.35 $X2=0 $Y2=0
cc_482 N_A_28_297#_c_524_n N_VPWR_c_896_n 0.0231894f $X=1.89 $Y=2.35 $X2=0 $Y2=0
cc_483 N_A_28_297#_c_528_n N_VPWR_c_896_n 0.0231894f $X=2.75 $Y=2.35 $X2=0 $Y2=0
cc_484 N_A_28_297#_c_530_n N_VPWR_c_896_n 0.0231894f $X=3.61 $Y=2.35 $X2=0 $Y2=0
cc_485 N_A_28_297#_c_520_n N_VPWR_c_896_n 0.00988695f $X=3.74 $Y=2.255 $X2=0
+ $Y2=0
cc_486 N_A_28_297#_c_564_p N_VPWR_c_896_n 0.00721854f $X=1.125 $Y=2.36 $X2=0
+ $Y2=0
cc_487 N_A_28_297#_c_565_p N_VPWR_c_896_n 0.00721854f $X=1.985 $Y=2.36 $X2=0
+ $Y2=0
cc_488 N_A_28_297#_c_566_p N_VPWR_c_896_n 0.00721854f $X=2.845 $Y=2.36 $X2=0
+ $Y2=0
cc_489 N_Y_c_587_n N_A_455_297#_c_741_n 0.0119588f $X=1.555 $Y=1.655 $X2=0 $Y2=0
cc_490 N_Y_c_581_n N_A_821_297#_c_810_n 0.00123169f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_491 N_Y_c_581_n N_A_821_297#_c_811_n 0.00616906f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_492 N_Y_M1003_s N_VPWR_c_896_n 0.00225769f $X=0.555 $Y=1.485 $X2=0 $Y2=0
cc_493 N_Y_M1015_s N_VPWR_c_896_n 0.00225769f $X=1.415 $Y=1.485 $X2=0 $Y2=0
cc_494 N_Y_c_606_n N_VGND_M1007_d 0.00178868f $X=0.7 $Y=0.62 $X2=-0.19 $Y2=-0.24
cc_495 N_Y_c_677_p N_VGND_M1007_d 0.00995319f $X=0.232 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_496 Y N_VGND_M1007_d 0.00538444f $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_497 N_Y_c_591_n N_VGND_M1009_d 0.00346729f $X=1.46 $Y=0.7 $X2=0 $Y2=0
cc_498 N_Y_c_599_n N_VGND_M1027_d 0.00924122f $X=2.4 $Y=0.7 $X2=0 $Y2=0
cc_499 N_Y_c_622_n N_VGND_M1010_s 0.00346729f $X=3.26 $Y=0.7 $X2=0 $Y2=0
cc_500 N_Y_c_626_n N_VGND_M1036_s 0.0117401f $X=4.18 $Y=0.7 $X2=0 $Y2=0
cc_501 N_Y_c_639_n N_VGND_M1002_s 0.00346729f $X=5.09 $Y=0.7 $X2=0 $Y2=0
cc_502 N_Y_c_581_n N_VGND_M1037_s 0.00559329f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_503 N_Y_c_606_n N_VGND_c_1028_n 0.00486505f $X=0.7 $Y=0.62 $X2=0 $Y2=0
cc_504 N_Y_c_677_p N_VGND_c_1028_n 0.0146521f $X=0.232 $Y=0.785 $X2=0 $Y2=0
cc_505 N_Y_c_591_n N_VGND_c_1029_n 0.0159085f $X=1.46 $Y=0.7 $X2=0 $Y2=0
cc_506 N_Y_c_622_n N_VGND_c_1030_n 0.0159085f $X=3.26 $Y=0.7 $X2=0 $Y2=0
cc_507 N_Y_c_626_n N_VGND_c_1031_n 0.020923f $X=4.18 $Y=0.7 $X2=0 $Y2=0
cc_508 N_Y_c_639_n N_VGND_c_1032_n 0.0159085f $X=5.09 $Y=0.7 $X2=0 $Y2=0
cc_509 N_Y_c_581_n N_VGND_c_1033_n 0.0208104f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_510 N_Y_c_581_n N_VGND_c_1036_n 0.00380563f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_511 N_Y_c_591_n N_VGND_c_1040_n 0.0025909f $X=1.46 $Y=0.7 $X2=0 $Y2=0
cc_512 N_Y_c_606_n N_VGND_c_1040_n 0.0073321f $X=0.7 $Y=0.62 $X2=0 $Y2=0
cc_513 N_Y_c_591_n N_VGND_c_1041_n 0.0025909f $X=1.46 $Y=0.7 $X2=0 $Y2=0
cc_514 N_Y_c_599_n N_VGND_c_1041_n 0.00260121f $X=2.4 $Y=0.7 $X2=0 $Y2=0
cc_515 N_Y_c_614_n N_VGND_c_1041_n 0.00514479f $X=1.555 $Y=0.62 $X2=0 $Y2=0
cc_516 N_Y_c_599_n N_VGND_c_1042_n 0.00260121f $X=2.4 $Y=0.7 $X2=0 $Y2=0
cc_517 N_Y_c_622_n N_VGND_c_1042_n 0.0025909f $X=3.26 $Y=0.7 $X2=0 $Y2=0
cc_518 N_Y_c_630_n N_VGND_c_1042_n 0.00514479f $X=2.495 $Y=0.62 $X2=0 $Y2=0
cc_519 N_Y_c_622_n N_VGND_c_1043_n 0.0025909f $X=3.26 $Y=0.7 $X2=0 $Y2=0
cc_520 N_Y_c_626_n N_VGND_c_1043_n 0.00266609f $X=4.18 $Y=0.7 $X2=0 $Y2=0
cc_521 N_Y_c_632_n N_VGND_c_1043_n 0.00626203f $X=3.355 $Y=0.62 $X2=0 $Y2=0
cc_522 N_Y_c_626_n N_VGND_c_1044_n 0.00273445f $X=4.18 $Y=0.7 $X2=0 $Y2=0
cc_523 N_Y_c_639_n N_VGND_c_1044_n 0.0025909f $X=5.09 $Y=0.7 $X2=0 $Y2=0
cc_524 N_Y_c_635_n N_VGND_c_1044_n 0.0059878f $X=4.325 $Y=0.62 $X2=0 $Y2=0
cc_525 N_Y_c_639_n N_VGND_c_1045_n 0.0025909f $X=5.09 $Y=0.7 $X2=0 $Y2=0
cc_526 N_Y_c_581_n N_VGND_c_1045_n 0.00255672f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_527 N_Y_c_650_n N_VGND_c_1045_n 0.00506386f $X=5.185 $Y=0.62 $X2=0 $Y2=0
cc_528 N_Y_M1007_s N_VGND_c_1047_n 0.00269459f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_529 N_Y_M1016_s N_VGND_c_1047_n 0.00277743f $X=1.415 $Y=0.235 $X2=0 $Y2=0
cc_530 N_Y_M1008_d N_VGND_c_1047_n 0.00277743f $X=2.355 $Y=0.235 $X2=0 $Y2=0
cc_531 N_Y_M1021_d N_VGND_c_1047_n 0.00269352f $X=3.215 $Y=0.235 $X2=0 $Y2=0
cc_532 N_Y_M1001_d N_VGND_c_1047_n 0.00269352f $X=4.185 $Y=0.235 $X2=0 $Y2=0
cc_533 N_Y_M1029_d N_VGND_c_1047_n 0.00278779f $X=5.045 $Y=0.235 $X2=0 $Y2=0
cc_534 N_Y_M1017_s N_VGND_c_1047_n 0.00225769f $X=6.455 $Y=0.235 $X2=0 $Y2=0
cc_535 N_Y_M1034_s N_VGND_c_1047_n 0.00225769f $X=7.315 $Y=0.235 $X2=0 $Y2=0
cc_536 N_Y_c_591_n N_VGND_c_1047_n 0.010077f $X=1.46 $Y=0.7 $X2=0 $Y2=0
cc_537 N_Y_c_599_n N_VGND_c_1047_n 0.0104456f $X=2.4 $Y=0.7 $X2=0 $Y2=0
cc_538 N_Y_c_622_n N_VGND_c_1047_n 0.010077f $X=3.26 $Y=0.7 $X2=0 $Y2=0
cc_539 N_Y_c_626_n N_VGND_c_1047_n 0.00984546f $X=4.18 $Y=0.7 $X2=0 $Y2=0
cc_540 N_Y_c_639_n N_VGND_c_1047_n 0.010077f $X=5.09 $Y=0.7 $X2=0 $Y2=0
cc_541 N_Y_c_581_n N_VGND_c_1047_n 0.014747f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_542 N_Y_c_606_n N_VGND_c_1047_n 0.0106264f $X=0.7 $Y=0.62 $X2=0 $Y2=0
cc_543 N_Y_c_614_n N_VGND_c_1047_n 0.00625591f $X=1.555 $Y=0.62 $X2=0 $Y2=0
cc_544 N_Y_c_630_n N_VGND_c_1047_n 0.00625591f $X=2.495 $Y=0.62 $X2=0 $Y2=0
cc_545 N_Y_c_632_n N_VGND_c_1047_n 0.00817182f $X=3.355 $Y=0.62 $X2=0 $Y2=0
cc_546 N_Y_c_635_n N_VGND_c_1047_n 0.00788856f $X=4.325 $Y=0.62 $X2=0 $Y2=0
cc_547 N_Y_c_650_n N_VGND_c_1047_n 0.00608953f $X=5.185 $Y=0.62 $X2=0 $Y2=0
cc_548 N_Y_c_677_p N_VGND_c_1047_n 9.15151e-19 $X=0.232 $Y=0.785 $X2=0 $Y2=0
cc_549 N_Y_c_599_n N_VGND_c_1049_n 0.0220137f $X=2.4 $Y=0.7 $X2=0 $Y2=0
cc_550 N_Y_c_581_n N_A_1205_47#_M1017_d 0.00614851f $X=7.455 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_551 N_Y_c_581_n N_A_1205_47#_M1020_d 0.00347122f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_552 N_Y_M1017_s N_A_1205_47#_c_1202_n 0.00329338f $X=6.455 $Y=0.235 $X2=0
+ $Y2=0
cc_553 N_Y_M1034_s N_A_1205_47#_c_1202_n 0.00329338f $X=7.315 $Y=0.235 $X2=0
+ $Y2=0
cc_554 N_Y_c_581_n N_A_1205_47#_c_1202_n 0.0829405f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_555 N_Y_c_581_n N_A_1205_47#_c_1211_n 0.0104127f $X=7.455 $Y=0.7 $X2=0 $Y2=0
cc_556 N_A_455_297#_c_739_n N_A_821_297#_M1012_d 0.00296258f $X=4.49 $Y=1.565
+ $X2=-0.19 $Y2=1.305
cc_557 N_A_455_297#_c_740_n N_A_821_297#_M1013_d 0.00177615f $X=5.35 $Y=1.58
+ $X2=0 $Y2=0
cc_558 N_A_455_297#_c_739_n N_A_821_297#_c_809_n 0.0192967f $X=4.49 $Y=1.565
+ $X2=0 $Y2=0
cc_559 N_A_455_297#_M1012_s N_A_821_297#_c_819_n 0.00340502f $X=4.515 $Y=1.485
+ $X2=0 $Y2=0
cc_560 N_A_455_297#_c_739_n N_A_821_297#_c_819_n 0.0030004f $X=4.49 $Y=1.565
+ $X2=0 $Y2=0
cc_561 N_A_455_297#_c_740_n N_A_821_297#_c_819_n 0.00318184f $X=5.35 $Y=1.58
+ $X2=0 $Y2=0
cc_562 N_A_455_297#_c_743_n N_A_821_297#_c_819_n 0.0161241f $X=4.655 $Y=1.655
+ $X2=0 $Y2=0
cc_563 N_A_455_297#_c_740_n N_A_821_297#_c_857_n 0.0135452f $X=5.35 $Y=1.58
+ $X2=0 $Y2=0
cc_564 N_A_455_297#_M1025_s N_A_821_297#_c_821_n 0.00347863f $X=5.375 $Y=1.485
+ $X2=0 $Y2=0
cc_565 N_A_455_297#_c_740_n N_A_821_297#_c_821_n 0.00305748f $X=5.35 $Y=1.58
+ $X2=0 $Y2=0
cc_566 N_A_455_297#_c_744_n N_A_821_297#_c_821_n 0.0144667f $X=5.515 $Y=1.655
+ $X2=0 $Y2=0
cc_567 N_A_455_297#_c_744_n N_A_821_297#_c_811_n 0.00606143f $X=5.515 $Y=1.655
+ $X2=0 $Y2=0
cc_568 N_A_455_297#_M1005_s N_VPWR_c_896_n 0.00225769f $X=2.275 $Y=1.485 $X2=0
+ $Y2=0
cc_569 N_A_455_297#_M1023_s N_VPWR_c_896_n 0.00225769f $X=3.135 $Y=1.485 $X2=0
+ $Y2=0
cc_570 N_A_455_297#_M1012_s N_VPWR_c_896_n 0.00225769f $X=4.515 $Y=1.485 $X2=0
+ $Y2=0
cc_571 N_A_455_297#_M1025_s N_VPWR_c_896_n 0.00225769f $X=5.375 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_821_297#_c_810_n N_VPWR_M1018_s 0.00176461f $X=6.72 $Y=1.53 $X2=-0.19
+ $Y2=1.305
cc_573 N_A_821_297#_c_812_n N_VPWR_M1033_s 0.00207281f $X=7.58 $Y=1.53 $X2=0
+ $Y2=0
cc_574 N_A_821_297#_c_813_n N_VPWR_M1000_d 0.00203249f $X=8.58 $Y=1.555 $X2=0
+ $Y2=0
cc_575 N_A_821_297#_c_814_n N_VPWR_M1019_d 0.00209536f $X=9.53 $Y=1.557 $X2=0
+ $Y2=0
cc_576 N_A_821_297#_c_810_n N_VPWR_c_897_n 0.0170777f $X=6.72 $Y=1.53 $X2=0
+ $Y2=0
cc_577 N_A_821_297#_c_867_p N_VPWR_c_898_n 0.00630278f $X=6.815 $Y=1.63 $X2=0
+ $Y2=0
cc_578 N_A_821_297#_c_812_n N_VPWR_c_899_n 0.0157999f $X=7.58 $Y=1.53 $X2=0
+ $Y2=0
cc_579 N_A_821_297#_c_813_n N_VPWR_c_900_n 0.0138355f $X=8.58 $Y=1.555 $X2=0
+ $Y2=0
cc_580 N_A_821_297#_c_870_p N_VPWR_c_901_n 0.0262333f $X=8.71 $Y=1.725 $X2=0
+ $Y2=0
cc_581 N_A_821_297#_c_814_n N_VPWR_c_901_n 0.0132165f $X=9.53 $Y=1.557 $X2=0
+ $Y2=0
cc_582 N_A_821_297#_c_808_n N_VPWR_c_902_n 0.0157719f $X=4.19 $Y=2.255 $X2=0
+ $Y2=0
cc_583 N_A_821_297#_c_819_n N_VPWR_c_902_n 0.032265f $X=4.99 $Y=2.35 $X2=0 $Y2=0
cc_584 N_A_821_297#_c_821_n N_VPWR_c_902_n 0.0438049f $X=5.86 $Y=2.36 $X2=0
+ $Y2=0
cc_585 N_A_821_297#_c_875_p N_VPWR_c_902_n 0.0109994f $X=5.085 $Y=2.36 $X2=0
+ $Y2=0
cc_586 N_A_821_297#_c_817_n N_VPWR_c_904_n 0.0109365f $X=7.695 $Y=1.63 $X2=0
+ $Y2=0
cc_587 N_A_821_297#_c_870_p N_VPWR_c_906_n 0.00826453f $X=8.71 $Y=1.725 $X2=0
+ $Y2=0
cc_588 N_A_821_297#_c_815_n N_VPWR_c_908_n 0.0069691f $X=9.625 $Y=1.725 $X2=0
+ $Y2=0
cc_589 N_A_821_297#_M1012_d N_VPWR_c_896_n 0.00210134f $X=4.105 $Y=1.485 $X2=0
+ $Y2=0
cc_590 N_A_821_297#_M1013_d N_VPWR_c_896_n 0.00224115f $X=4.945 $Y=1.485 $X2=0
+ $Y2=0
cc_591 N_A_821_297#_M1031_d N_VPWR_c_896_n 0.00389862f $X=5.805 $Y=1.485 $X2=0
+ $Y2=0
cc_592 N_A_821_297#_M1026_d N_VPWR_c_896_n 0.0055905f $X=6.675 $Y=1.485 $X2=0
+ $Y2=0
cc_593 N_A_821_297#_M1035_d N_VPWR_c_896_n 0.0059702f $X=7.555 $Y=1.485 $X2=0
+ $Y2=0
cc_594 N_A_821_297#_M1004_s N_VPWR_c_896_n 0.00712439f $X=8.535 $Y=1.485 $X2=0
+ $Y2=0
cc_595 N_A_821_297#_M1030_s N_VPWR_c_896_n 0.00403373f $X=9.485 $Y=1.485 $X2=0
+ $Y2=0
cc_596 N_A_821_297#_c_808_n N_VPWR_c_896_n 0.00988695f $X=4.19 $Y=2.255 $X2=0
+ $Y2=0
cc_597 N_A_821_297#_c_819_n N_VPWR_c_896_n 0.0231894f $X=4.99 $Y=2.35 $X2=0
+ $Y2=0
cc_598 N_A_821_297#_c_821_n N_VPWR_c_896_n 0.0307932f $X=5.86 $Y=2.36 $X2=0
+ $Y2=0
cc_599 N_A_821_297#_c_867_p N_VPWR_c_896_n 0.00664749f $X=6.815 $Y=1.63 $X2=0
+ $Y2=0
cc_600 N_A_821_297#_c_870_p N_VPWR_c_896_n 0.00897434f $X=8.71 $Y=1.725 $X2=0
+ $Y2=0
cc_601 N_A_821_297#_c_815_n N_VPWR_c_896_n 0.00811321f $X=9.625 $Y=1.725 $X2=0
+ $Y2=0
cc_602 N_A_821_297#_c_875_p N_VPWR_c_896_n 0.00721854f $X=5.085 $Y=2.36 $X2=0
+ $Y2=0
cc_603 N_A_821_297#_c_817_n N_VPWR_c_896_n 0.0115978f $X=7.695 $Y=1.63 $X2=0
+ $Y2=0
cc_604 N_A_821_297#_c_813_n N_A_1205_47#_c_1211_n 0.00152474f $X=8.58 $Y=1.555
+ $X2=0 $Y2=0
cc_605 N_A_821_297#_c_817_n N_A_1205_47#_c_1211_n 8.38391e-19 $X=7.695 $Y=1.63
+ $X2=0 $Y2=0
cc_606 N_VGND_c_1047_n N_A_1205_47#_M1017_d 0.00226644f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_607 N_VGND_c_1047_n N_A_1205_47#_M1020_d 0.00224157f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1047_n N_A_1205_47#_M1038_d 0.00317306f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_c_1047_n N_A_1205_47#_M1022_s 0.00255449f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_610 N_VGND_c_1047_n N_A_1205_47#_M1039_s 0.00230091f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1033_n N_A_1205_47#_c_1202_n 0.0132643f $X=5.61 $Y=0.36 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1036_n N_A_1205_47#_c_1202_n 0.106051f $X=8.245 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1047_n N_A_1205_47#_c_1202_n 0.0743189f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_M1006_d N_A_1205_47#_c_1212_n 0.00346397f $X=8.27 $Y=0.235 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1034_n N_A_1205_47#_c_1212_n 0.0159085f $X=8.41 $Y=0.36 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1036_n N_A_1205_47#_c_1212_n 0.0025909f $X=8.245 $Y=0 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1038_n N_A_1205_47#_c_1212_n 0.0025909f $X=9.105 $Y=0 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1047_n N_A_1205_47#_c_1212_n 0.0100658f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1038_n N_A_1205_47#_c_1246_n 0.00945039f $X=9.105 $Y=0 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1047_n N_A_1205_47#_c_1246_n 0.0070077f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_M1024_d N_A_1205_47#_c_1203_n 0.00346397f $X=9.13 $Y=0.235 $X2=0
+ $Y2=0
cc_622 N_VGND_c_1035_n N_A_1205_47#_c_1203_n 0.0159085f $X=9.27 $Y=0.36 $X2=0
+ $Y2=0
cc_623 N_VGND_c_1038_n N_A_1205_47#_c_1203_n 0.0025909f $X=9.105 $Y=0 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1046_n N_A_1205_47#_c_1203_n 0.0025909f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_625 N_VGND_c_1047_n N_A_1205_47#_c_1203_n 0.0100658f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_626 N_VGND_c_1046_n N_A_1205_47#_c_1204_n 0.0142273f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_627 N_VGND_c_1047_n N_A_1205_47#_c_1204_n 0.00967631f $X=9.89 $Y=0 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__clkdlybuf4s25_2.spice
* Created: Thu Aug 27 14:11:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s25_2.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s25_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1113 PD=0.765421 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_225_47#_M1007_d N_A_27_47#_M1007_g N_VGND_M1003_d VNB NSHORT L=0.25
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=2.6 SA=125000
+ SB=125000 A=0.1625 P=1.8 MULT=1
MM1008 N_VGND_M1008_d N_A_225_47#_M1008_g N_A_331_47#_M1008_s VNB NSHORT L=0.25
+ W=0.65 AD=0.11785 AS=0.169 PD=1.18458 PS=1.82 NRD=0 NRS=0 M=1 R=2.6 SA=125000
+ SB=125001 A=0.1625 P=1.8 MULT=1
MM1000 N_X_M1000_d N_A_331_47#_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0761495 PD=0.77 PS=0.765421 NRD=21.42 NRS=14.28 M=1 R=2.8
+ SA=75000.8 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1000_d N_A_331_47#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1407 PD=0.77 PS=1.51 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.171154 AS=0.265 PD=1.45604 PS=2.53 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1006 N_A_225_47#_M1006_d N_A_27_47#_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.25
+ W=0.82 AD=0.2132 AS=0.140346 PD=2.16 PS=1.19396 NRD=0 NRS=0 M=1 R=3.28
+ SA=125001 SB=125000 A=0.205 P=2.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_225_47#_M1001_g N_A_331_47#_M1001_s VPB PHIGHVT L=0.25
+ W=0.82 AD=0.140346 AS=0.2132 PD=1.19396 PS=2.16 NRD=0 NRS=0 M=1 R=3.28
+ SA=125000 SB=125001 A=0.205 P=2.14 MULT=1
MM1002 N_X_M1002_d N_A_331_47#_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.171154 PD=1.35 PS=1.45604 NRD=14.7553 NRS=9.8303 M=1 R=6.66667
+ SA=75000.7 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1002_d N_A_331_47#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.335 PD=1.35 PS=2.67 NRD=0 NRS=13.7703 M=1 R=6.66667 SA=75001.2
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_65 VPB 0 2.38063e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__clkdlybuf4s25_2.pxi.spice"
*
.ends
*
*

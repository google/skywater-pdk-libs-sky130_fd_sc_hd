* File: sky130_fd_sc_hd__and4_2.spice.pex
* Created: Thu Aug 27 14:08:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4_2%A 3 7 9 10 11 12 21
r31 18 21 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r32 11 12 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.227 $Y=1.53
+ $X2=0.227 $Y2=1.87
r33 10 11 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.227 $Y=1.16
+ $X2=0.227 $Y2=1.53
r34 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r35 9 10 16.7716 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=0.227 $Y=0.85
+ $X2=0.227 $Y2=1.16
r36 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r37 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r38 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r39 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%B 3 7 9 10 14
c36 14 0 3.07319e-19 $X=0.975 $Y=1.16
r37 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=0.975 $Y2=0.995
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.16 $X2=0.975 $Y2=1.16
r39 10 15 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=1.067 $Y=0.85
+ $X2=1.067 $Y2=1.16
r40 9 10 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=1.067 $Y=0.51
+ $X2=1.067 $Y2=0.85
r41 5 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.16
r42 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=2.275
r43 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.915 $Y=0.445
+ $X2=0.915 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%C 3 7 9 10 11 17 30
c37 30 0 1.58629e-19 $X=1.615 $Y=1.19
c38 9 0 1.48689e-19 $X=1.615 $Y=0.51
r39 18 30 1.28873 $w=2.84e-07 $l=3e-08 $layer=LI1_cond $X=1.57 $Y=1.16 $X2=1.57
+ $Y2=1.19
r40 18 21 0.25114 $w=3e-07 $l=5e-09 $layer=LI1_cond $X=1.57 $Y=1.16 $X2=1.57
+ $Y2=1.155
r41 17 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.16
+ $X2=1.505 $Y2=1.325
r42 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.16
+ $X2=1.505 $Y2=0.995
r43 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.16 $X2=1.505 $Y2=1.16
r44 11 30 1.07394 $w=2.84e-07 $l=2.5e-08 $layer=LI1_cond $X=1.57 $Y=1.215
+ $X2=1.57 $Y2=1.19
r45 11 21 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=1.57 $Y=1.13
+ $X2=1.57 $Y2=1.155
r46 10 11 10.7561 $w=2.98e-07 $l=2.8e-07 $layer=LI1_cond $X=1.57 $Y=0.85
+ $X2=1.57 $Y2=1.13
r47 9 10 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.57 $Y=0.51 $X2=1.57
+ $Y2=0.85
r48 7 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.495 $Y=2.275
+ $X2=1.495 $Y2=1.325
r49 3 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.445 $Y=0.445
+ $X2=1.445 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%D 3 7 9 10 11 16
c38 16 0 6.10995e-20 $X=1.985 $Y=1.16
r39 16 19 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.16
+ $X2=2.01 $Y2=1.325
r40 16 18 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.16
+ $X2=2.01 $Y2=0.995
r41 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.985
+ $Y=1.16 $X2=1.985 $Y2=1.16
r42 11 17 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=2.03 $Y=1.19 $X2=2.03
+ $Y2=1.16
r43 10 17 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.03 $Y=0.85
+ $X2=2.03 $Y2=1.16
r44 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.03 $Y=0.51 $X2=2.03
+ $Y2=0.85
r45 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.925 $Y=2.275
+ $X2=1.925 $Y2=1.325
r46 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.925 $Y=0.445
+ $X2=1.925 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%A_27_47# 1 2 3 10 12 15 17 19 22 25 28 30 34
+ 36 39 43 45 46 50 56
c104 39 0 6.10995e-20 $X=2.442 $Y=1.495
r105 55 56 83.9334 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=3.17 $Y2=1.16
r106 51 55 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.56 $Y=1.16
+ $X2=2.69 $Y2=1.16
r107 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.16 $X2=2.56 $Y2=1.16
r108 47 50 5.66618 $w=2.38e-07 $l=1.18e-07 $layer=LI1_cond $X=2.442 $Y=1.195
+ $X2=2.56 $Y2=1.195
r109 41 43 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.26 $Y=0.42
+ $X2=0.585 $Y2=0.42
r110 38 47 1.13239 $w=2.25e-07 $l=1.2e-07 $layer=LI1_cond $X=2.442 $Y=1.315
+ $X2=2.442 $Y2=1.195
r111 38 39 9.21954 $w=2.23e-07 $l=1.8e-07 $layer=LI1_cond $X=2.442 $Y=1.315
+ $X2=2.442 $Y2=1.495
r112 37 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.71 $Y2=1.58
r113 36 39 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.33 $Y=1.58
+ $X2=2.442 $Y2=1.495
r114 36 37 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.33 $Y=1.58
+ $X2=1.835 $Y2=1.58
r115 32 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.58
r116 32 34 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=2.3
r117 31 45 2.11342 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.85 $Y=1.58
+ $X2=0.675 $Y2=1.58
r118 30 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.585 $Y=1.58
+ $X2=1.71 $Y2=1.58
r119 30 31 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.585 $Y=1.58
+ $X2=0.85 $Y2=1.58
r120 26 45 4.3182 $w=2.1e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.675 $Y2=1.58
r121 26 28 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=2.3
r122 25 45 4.3182 $w=2.1e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.585 $Y=1.495
+ $X2=0.675 $Y2=1.58
r123 24 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0.585
+ $X2=0.585 $Y2=0.42
r124 24 25 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.585 $Y=0.585
+ $X2=0.585 $Y2=1.495
r125 20 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.325
+ $X2=3.17 $Y2=1.16
r126 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.17 $Y=1.325
+ $X2=3.17 $Y2=1.985
r127 17 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=0.995
+ $X2=3.17 $Y2=1.16
r128 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.17 $Y=0.995
+ $X2=3.17 $Y2=0.56
r129 13 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.16
r130 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.985
r131 10 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=0.995
+ $X2=2.69 $Y2=1.16
r132 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.69 $Y=0.995
+ $X2=2.69 $Y2=0.56
r133 3 34 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=2.065 $X2=1.71 $Y2=2.3
r134 2 28 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.725 $Y2=2.3
r135 1 41 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%VPWR 1 2 3 4 13 15 17 21 25 27 29 32 33 34 40
+ 48 52
r53 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 40 51 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.462 $Y2=2.72
r58 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 39 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=2.72
+ $X2=1.235 $Y2=2.72
r63 36 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.4 $Y=2.72 $X2=2.07
+ $Y2=2.72
r64 34 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 34 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 32 38 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.4 $Y2=2.72
r68 31 42 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.4 $Y2=2.72
r70 27 51 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.41 $Y=2.635
+ $X2=3.462 $Y2=2.72
r71 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.41 $Y=2.635
+ $X2=3.41 $Y2=2
r72 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.635 $X2=2.4
+ $Y2=2.72
r73 23 25 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2
r74 19 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.635
+ $X2=1.235 $Y2=2.72
r75 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.235 $Y=2.635
+ $X2=1.235 $Y2=2.34
r76 18 45 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r77 17 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.72
+ $X2=1.235 $Y2=2.72
r78 17 18 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.07 $Y=2.72
+ $X2=0.425 $Y2=2.72
r79 13 45 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r80 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r81 4 29 300 $w=1.7e-07 $l=5.91777e-07 $layer=licon1_PDIFF $count=2 $X=3.245
+ $Y=1.485 $X2=3.41 $Y2=2
r82 3 25 300 $w=1.7e-07 $l=4.31277e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=2.065 $X2=2.4 $Y2=2
r83 2 21 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=2.065 $X2=1.235 $Y2=2.34
r84 1 15 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%X 1 2 7 8 9 10 11 12 21 24 44
r22 44 45 3.82115 $w=3.33e-07 $l=3.5e-08 $layer=LI1_cond $X=2.902 $Y=1.53
+ $X2=2.902 $Y2=1.495
r23 29 48 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=2.902 $Y=1.662
+ $X2=2.902 $Y2=1.66
r24 21 24 2.85195 $w=1.73e-07 $l=4.5e-08 $layer=LI1_cond $X=2.982 $Y=0.805
+ $X2=2.982 $Y2=0.85
r25 12 35 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=2.902 $Y=2.21
+ $X2=2.902 $Y2=2.34
r26 11 12 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.902 $Y=1.87
+ $X2=2.902 $Y2=2.21
r27 11 29 7.15547 $w=3.33e-07 $l=2.08e-07 $layer=LI1_cond $X=2.902 $Y=1.87
+ $X2=2.902 $Y2=1.662
r28 10 48 3.61213 $w=3.33e-07 $l=1.05e-07 $layer=LI1_cond $X=2.902 $Y=1.555
+ $X2=2.902 $Y2=1.66
r29 10 44 0.860032 $w=3.33e-07 $l=2.5e-08 $layer=LI1_cond $X=2.902 $Y=1.555
+ $X2=2.902 $Y2=1.53
r30 10 45 1.58442 $w=1.73e-07 $l=2.5e-08 $layer=LI1_cond $X=2.982 $Y=1.47
+ $X2=2.982 $Y2=1.495
r31 9 10 17.7455 $w=1.73e-07 $l=2.8e-07 $layer=LI1_cond $X=2.982 $Y=1.19
+ $X2=2.982 $Y2=1.47
r32 8 21 5.85659 $w=3.34e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.902 $Y=0.72
+ $X2=2.982 $Y2=0.805
r33 8 9 20.2805 $w=1.73e-07 $l=3.2e-07 $layer=LI1_cond $X=2.982 $Y=0.87
+ $X2=2.982 $Y2=1.19
r34 8 24 1.26753 $w=1.73e-07 $l=2e-08 $layer=LI1_cond $X=2.982 $Y=0.87 $X2=2.982
+ $Y2=0.85
r35 7 8 7.67066 $w=3.34e-07 $l=2.1e-07 $layer=LI1_cond $X=2.902 $Y=0.51
+ $X2=2.902 $Y2=0.72
r36 7 38 4.7485 $w=3.34e-07 $l=1.3e-07 $layer=LI1_cond $X=2.902 $Y=0.51
+ $X2=2.902 $Y2=0.38
r37 2 48 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=1.66
r38 2 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=2.34
r39 1 8 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.765
+ $Y=0.235 $X2=2.9 $Y2=0.72
r40 1 38 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.765
+ $Y=0.235 $X2=2.9 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_2%VGND 1 2 9 11 13 16 17 18 27 33
r44 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r45 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r47 27 32 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r48 27 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r49 26 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r50 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r51 21 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r52 18 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r53 18 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r54 16 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.07
+ $Y2=0
r55 16 17 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.447
+ $Y2=0
r56 15 29 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.99
+ $Y2=0
r57 15 17 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.447
+ $Y2=0
r58 11 32 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.467 $Y2=0
r59 11 13 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.42 $Y=0.085 $X2=3.42
+ $Y2=0.385
r60 7 17 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.447 $Y=0.085
+ $X2=2.447 $Y2=0
r61 7 9 14.712 $w=2.33e-07 $l=3e-07 $layer=LI1_cond $X=2.447 $Y=0.085 $X2=2.447
+ $Y2=0.385
r62 2 13 91 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_NDIFF $count=2 $X=3.245
+ $Y=0.235 $X2=3.42 $Y2=0.385
r63 1 9 91 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.235
+ $X2=2.47 $Y2=0.385
.ends


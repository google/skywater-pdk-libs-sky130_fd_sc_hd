* NGSPICE file created from sky130_fd_sc_hd__or3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
M1000 a_542_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=8.315e+11p ps=7.75e+06u
M1001 a_176_21# a_27_47# a_626_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=3.3e+11p ps=2.66e+06u
M1002 VGND a_176_21# X VNB nshort w=650000u l=150000u
+  ad=7.66e+11p pd=7.61e+06u as=3.51e+11p ps=3.68e+06u
M1003 X a_176_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_176_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1005 X a_176_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B a_176_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.445e+11p ps=3.66e+06u
M1007 X a_176_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_176_21# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_176_21# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_176_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_626_297# B a_542_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_176_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1014 VPWR C_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 X a_176_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_8.spice
* Created: Thu Aug 27 14:23:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_8.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_8  VNB VPB A KAPWR X VGND VPWR
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_A_110_47#_M1004_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75004.1
+ A=0.063 P=1.14 MULT=1
MM1012 N_A_110_47#_M1004_d N_A_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75003.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1012_s N_A_110_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75003.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_110_47#_M1006_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1006_d N_A_110_47#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_110_47#_M1010_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1010_d N_A_110_47#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_110_47#_M1016_g N_X_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1016_d N_A_110_47#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_110_47#_M1019_g N_X_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0588 PD=1.38 PS=0.7 NRD=1.428 NRS=0 M=1 R=2.8 SA=75004.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_110_47#_M1007_d N_A_M1007_g N_KAPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1018 N_A_110_47#_M1007_d N_A_M1018_g N_KAPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_110_47#_M1000_g N_KAPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75003.2
+ A=0.15 P=2.3 MULT=1
MM1002 N_X_M1000_d N_A_110_47#_M1002_g N_KAPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_110_47#_M1003_g N_KAPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1003_d N_A_110_47#_M1005_g N_KAPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1009_d N_A_110_47#_M1009_g N_KAPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1009_d N_A_110_47#_M1011_g N_KAPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1013 N_X_M1013_d N_A_110_47#_M1013_g N_KAPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_X_M1013_d N_A_110_47#_M1015_g N_KAPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_8.pxi.spice"
*
.ends
*
*

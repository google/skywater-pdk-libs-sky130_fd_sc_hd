* File: sky130_fd_sc_hd__nor4_4.spice
* Created: Thu Aug 27 14:32:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor4_4.spice.pex"
.subckt sky130_fd_sc_hd__nor4_4  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75007 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1006_d N_A_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75006.2 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1018_d N_A_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75005.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1019_s N_B_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_B_M1020_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1020_d N_B_M1023_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1027_d N_B_M1027_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1027_d N_C_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1007_d N_C_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_C_M1011_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_D_M1000_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.8
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1000_d N_D_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1009_d N_D_M1009_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1009_d N_D_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75007
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1003_d N_A_M1021_g N_A_27_297#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g N_A_27_297#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1029 N_VPWR_M1024_d N_A_M1029_g N_A_27_297#_M1029_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1002 N_A_27_297#_M1029_s N_B_M1002_g N_A_449_297#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1014 N_A_27_297#_M1014_d N_B_M1014_g N_A_449_297#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1015 N_A_27_297#_M1014_d N_B_M1015_g N_A_449_297#_M1015_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1025 N_A_27_297#_M1025_d N_B_M1025_g N_A_449_297#_M1015_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_449_297#_M1001_d N_C_M1001_g N_A_807_297#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1016 N_A_449_297#_M1001_d N_C_M1016_g N_A_807_297#_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1026 N_A_449_297#_M1026_d N_C_M1026_g N_A_807_297#_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1030 N_A_449_297#_M1026_d N_C_M1030_g N_A_807_297#_M1030_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1017 N_A_807_297#_M1030_s N_D_M1017_g N_Y_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1022 N_A_807_297#_M1022_d N_D_M1022_g N_Y_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1028 N_A_807_297#_M1022_d N_D_M1028_g N_Y_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1031 N_A_807_297#_M1031_d N_D_M1031_g N_Y_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__nor4_4.spice.SKY130_FD_SC_HD__NOR4_4.pxi"
*
.ends
*
*

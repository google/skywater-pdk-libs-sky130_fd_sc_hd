* File: sky130_fd_sc_hd__o21ai_4.spice.SKY130_FD_SC_HD__O21AI_4.pxi
* Created: Thu Aug 27 14:35:52 2020
* 
x_PM_SKY130_FD_SC_HD__O21AI_4%A1 N_A1_c_82_n N_A1_M1012_g N_A1_M1002_g
+ N_A1_c_83_n N_A1_M1017_g N_A1_M1004_g N_A1_c_84_n N_A1_M1021_g N_A1_M1007_g
+ N_A1_M1020_g N_A1_M1022_g N_A1_c_102_p N_A1_c_85_n N_A1_c_86_n A1 N_A1_c_87_n
+ N_A1_c_88_n N_A1_c_89_n N_A1_c_90_n PM_SKY130_FD_SC_HD__O21AI_4%A1
x_PM_SKY130_FD_SC_HD__O21AI_4%A2 N_A2_c_192_n N_A2_M1005_g N_A2_M1000_g
+ N_A2_c_193_n N_A2_M1009_g N_A2_M1008_g N_A2_c_194_n N_A2_M1018_g N_A2_M1013_g
+ N_A2_c_195_n N_A2_M1019_g N_A2_M1016_g A2 N_A2_c_196_n N_A2_c_197_n
+ PM_SKY130_FD_SC_HD__O21AI_4%A2
x_PM_SKY130_FD_SC_HD__O21AI_4%B1 N_B1_c_263_n N_B1_M1001_g N_B1_M1006_g
+ N_B1_c_264_n N_B1_M1003_g N_B1_M1011_g N_B1_c_265_n N_B1_M1010_g N_B1_M1014_g
+ N_B1_c_266_n N_B1_M1015_g N_B1_M1023_g B1 N_B1_c_267_n N_B1_c_268_n
+ PM_SKY130_FD_SC_HD__O21AI_4%B1
x_PM_SKY130_FD_SC_HD__O21AI_4%VPWR N_VPWR_M1002_s N_VPWR_M1004_s N_VPWR_M1020_s
+ N_VPWR_M1011_d N_VPWR_M1023_d N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n VPWR
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_332_n N_VPWR_c_348_n
+ PM_SKY130_FD_SC_HD__O21AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O21AI_4%A_115_297# N_A_115_297#_M1002_d
+ N_A_115_297#_M1007_d N_A_115_297#_M1008_s N_A_115_297#_M1016_s
+ N_A_115_297#_c_451_n N_A_115_297#_c_433_n N_A_115_297#_c_438_n
+ N_A_115_297#_c_458_n N_A_115_297#_c_441_n
+ PM_SKY130_FD_SC_HD__O21AI_4%A_115_297#
x_PM_SKY130_FD_SC_HD__O21AI_4%Y N_Y_M1001_d N_Y_M1010_d N_Y_M1000_d N_Y_M1013_d
+ N_Y_M1006_s N_Y_M1014_s N_Y_c_476_n N_Y_c_480_n N_Y_c_518_n N_Y_c_469_n
+ N_Y_c_470_n N_Y_c_527_n N_Y_c_471_n N_Y_c_472_n Y N_Y_c_467_n Y
+ PM_SKY130_FD_SC_HD__O21AI_4%Y
x_PM_SKY130_FD_SC_HD__O21AI_4%A_32_47# N_A_32_47#_M1012_s N_A_32_47#_M1017_s
+ N_A_32_47#_M1005_s N_A_32_47#_M1018_s N_A_32_47#_M1022_s N_A_32_47#_M1003_s
+ N_A_32_47#_M1015_s N_A_32_47#_c_548_n N_A_32_47#_c_590_p N_A_32_47#_c_549_n
+ PM_SKY130_FD_SC_HD__O21AI_4%A_32_47#
x_PM_SKY130_FD_SC_HD__O21AI_4%VGND N_VGND_M1012_d N_VGND_M1021_d N_VGND_M1009_d
+ N_VGND_M1019_d N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n N_VGND_c_605_n
+ N_VGND_c_606_n N_VGND_c_607_n VGND N_VGND_c_608_n N_VGND_c_609_n
+ N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n N_VGND_c_614_n
+ N_VGND_c_615_n PM_SKY130_FD_SC_HD__O21AI_4%VGND
cc_1 VNB N_A1_c_82_n 0.0218823f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_2 VNB N_A1_c_83_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.995
cc_3 VNB N_A1_c_84_n 0.016201f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=0.995
cc_4 VNB N_A1_c_85_n 0.00102663f $X=-0.19 $Y=-0.24 $X2=3.53 $Y2=1.16
cc_5 VNB N_A1_c_86_n 0.0259364f $X=-0.19 $Y=-0.24 $X2=3.53 $Y2=1.16
cc_6 VNB N_A1_c_87_n 0.0117702f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_7 VNB N_A1_c_88_n 0.070642f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=1.16
cc_8 VNB N_A1_c_89_n 0.016885f $X=-0.19 $Y=-0.24 $X2=3.53 $Y2=0.995
cc_9 VNB N_A1_c_90_n 0.00288578f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=1.35
cc_10 VNB N_A2_c_192_n 0.016201f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_11 VNB N_A2_c_193_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.995
cc_12 VNB N_A2_c_194_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=0.995
cc_13 VNB N_A2_c_195_n 0.0164823f $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.325
cc_14 VNB N_A2_c_196_n 0.0026767f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_15 VNB N_A2_c_197_n 0.063975f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_16 VNB N_B1_c_263_n 0.0163671f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_17 VNB N_B1_c_264_n 0.0161356f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.995
cc_18 VNB N_B1_c_265_n 0.0162015f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=0.995
cc_19 VNB N_B1_c_266_n 0.0192832f $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.325
cc_20 VNB N_B1_c_267_n 0.00172607f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_21 VNB N_B1_c_268_n 0.0658413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_332_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_467_n 0.0136716f $X=-0.19 $Y=-0.24 $X2=3.53 $Y2=0.995
cc_24 VNB Y 0.0266401f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.35
cc_25 VNB N_A_32_47#_c_548_n 0.00946883f $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.325
cc_26 VNB N_A_32_47#_c_549_n 0.00812227f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_27 VNB N_VGND_c_602_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=0.995
cc_28 VNB N_VGND_c_603_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=1.985
cc_29 VNB N_VGND_c_604_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.985
cc_30 VNB N_VGND_c_605_n 0.00274151f $X=-0.19 $Y=-0.24 $X2=3.55 $Y2=0.56
cc_31 VNB N_VGND_c_606_n 0.0122674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_607_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=3.445 $Y2=1.6
cc_33 VNB N_VGND_c_608_n 0.0166153f $X=-0.19 $Y=-0.24 $X2=3.57 $Y2=1.16
cc_34 VNB N_VGND_c_609_n 0.0122674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_610_n 0.0122674f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_36 VNB N_VGND_c_611_n 0.0611935f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.35
cc_37 VNB N_VGND_c_612_n 0.300469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_613_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.35
cc_39 VNB N_VGND_c_614_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_615_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VPB N_A1_M1002_g 0.025427f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_42 VPB N_A1_M1004_g 0.0171771f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.985
cc_43 VPB N_A1_M1007_g 0.0172416f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.985
cc_44 VPB N_A1_M1020_g 0.0188845f $X=-0.19 $Y=1.305 $X2=3.51 $Y2=1.985
cc_45 VPB N_A1_c_85_n 0.00151152f $X=-0.19 $Y=1.305 $X2=3.53 $Y2=1.16
cc_46 VPB N_A1_c_86_n 0.00619181f $X=-0.19 $Y=1.305 $X2=3.53 $Y2=1.16
cc_47 VPB N_A1_c_87_n 5.70185e-19 $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_48 VPB N_A1_c_88_n 0.0202636f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.16
cc_49 VPB N_A1_c_90_n 0.00204956f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=1.35
cc_50 VPB N_A2_M1000_g 0.0190346f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_51 VPB N_A2_M1008_g 0.0185962f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.985
cc_52 VPB N_A2_M1013_g 0.0185977f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.985
cc_53 VPB N_A2_M1016_g 0.0188697f $X=-0.19 $Y=1.305 $X2=3.55 $Y2=0.56
cc_54 VPB N_A2_c_196_n 0.00818697f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_55 VPB N_A2_c_197_n 0.0120771f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_56 VPB N_B1_M1006_g 0.0190237f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_57 VPB N_B1_M1011_g 0.0181789f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.985
cc_58 VPB N_B1_M1014_g 0.0181588f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.985
cc_59 VPB N_B1_M1023_g 0.0211964f $X=-0.19 $Y=1.305 $X2=3.55 $Y2=0.56
cc_60 VPB N_B1_c_268_n 0.0109651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_333_n 0.0114848f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=0.56
cc_62 VPB N_VPWR_c_334_n 0.0303061f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.325
cc_63 VPB N_VPWR_c_335_n 4.06898e-19 $X=-0.19 $Y=1.305 $X2=3.51 $Y2=1.325
cc_64 VPB N_VPWR_c_336_n 0.00252906f $X=-0.19 $Y=1.305 $X2=3.55 $Y2=0.995
cc_65 VPB N_VPWR_c_337_n 3.12649e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_338_n 0.0264268f $X=-0.19 $Y=1.305 $X2=3.57 $Y2=1.16
cc_67 VPB N_VPWR_c_339_n 0.0520859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_340_n 0.0042586f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.445
cc_69 VPB N_VPWR_c_341_n 0.0119442f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.16
cc_70 VPB N_VPWR_c_342_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_343_n 0.0121761f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_72 VPB N_VPWR_c_344_n 0.00510842f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_73 VPB N_VPWR_c_345_n 0.0142188f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_74 VPB N_VPWR_c_346_n 0.0126445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_332_n 0.0541738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_348_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_Y_c_469_n 0.00312134f $X=-0.19 $Y=1.305 $X2=3.53 $Y2=1.16
cc_78 VPB N_Y_c_470_n 0.00186893f $X=-0.19 $Y=1.305 $X2=3.53 $Y2=1.16
cc_79 VPB N_Y_c_471_n 0.0220671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_Y_c_472_n 0.001447f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_81 VPB Y 0.00832566f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.35
cc_82 N_A1_c_84_n N_A2_c_192_n 0.0269803f $X=1.36 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_83 N_A1_M1007_g N_A2_M1000_g 0.040849f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A1_c_102_p N_A2_M1000_g 0.016698f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_85 N_A1_c_90_n N_A2_M1000_g 0.00382797f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_86 N_A1_c_102_p N_A2_M1008_g 0.0104926f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_87 N_A1_c_102_p N_A2_M1013_g 0.0104926f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_88 N_A1_c_89_n N_A2_c_195_n 0.0232572f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A1_M1020_g N_A2_M1016_g 0.0459592f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A1_c_102_p N_A2_M1016_g 0.010446f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_91 N_A1_c_85_n N_A2_M1016_g 0.00104941f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A1_c_102_p N_A2_c_196_n 0.0837773f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_93 N_A1_c_85_n N_A2_c_196_n 0.0225557f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A1_c_86_n N_A2_c_196_n 0.00183217f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A1_c_88_n N_A2_c_196_n 2.1924e-19 $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A1_c_90_n N_A2_c_196_n 0.00953092f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_97 N_A1_c_102_p N_A2_c_197_n 0.00290276f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_98 N_A1_c_85_n N_A2_c_197_n 7.26125e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A1_c_86_n N_A2_c_197_n 0.0212933f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A1_c_88_n N_A2_c_197_n 0.0191171f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_c_90_n N_A2_c_197_n 0.00164529f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A1_c_89_n N_B1_c_263_n 0.0231424f $X=3.53 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_103 N_A1_M1020_g N_B1_M1006_g 0.0362349f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A1_c_102_p N_B1_M1006_g 0.00124789f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_105 N_A1_c_85_n N_B1_M1006_g 0.00304502f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A1_c_85_n N_B1_c_267_n 0.0170338f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_c_86_n N_B1_c_267_n 8.96733e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A1_c_85_n N_B1_c_268_n 8.79736e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A1_c_86_n N_B1_c_268_n 0.02144f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A1_c_90_n N_VPWR_M1004_s 0.0021089f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_111 N_A1_c_102_p N_VPWR_M1020_s 0.00229926f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_112 N_A1_c_85_n N_VPWR_M1020_s 2.85254e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A1_M1002_g N_VPWR_c_334_n 0.00331f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A1_c_87_n N_VPWR_c_334_n 0.00925631f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A1_c_88_n N_VPWR_c_334_n 0.00509813f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_M1002_g N_VPWR_c_335_n 5.22097e-19 $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A1_M1004_g N_VPWR_c_335_n 0.00656071f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A1_M1007_g N_VPWR_c_335_n 0.00759172f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A1_M1020_g N_VPWR_c_336_n 0.00293166f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A1_M1007_g N_VPWR_c_339_n 0.00353537f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A1_M1020_g N_VPWR_c_339_n 0.00421077f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A1_M1002_g N_VPWR_c_345_n 0.00585385f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A1_M1004_g N_VPWR_c_345_n 0.00353537f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A1_M1002_g N_VPWR_c_332_n 0.01147f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A1_M1004_g N_VPWR_c_332_n 0.00411309f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A1_M1007_g N_VPWR_c_332_n 0.00413843f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A1_M1020_g N_VPWR_c_332_n 0.00587621f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A1_c_90_n N_A_115_297#_M1002_d 0.00253064f $X=1.475 $Y=1.35 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A1_c_102_p N_A_115_297#_M1007_d 0.00834989f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_130 N_A1_c_102_p N_A_115_297#_M1008_s 0.00331496f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_131 N_A1_c_102_p N_A_115_297#_M1016_s 0.00602712f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_132 N_A1_M1004_g N_A_115_297#_c_433_n 0.0118869f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A1_M1007_g N_A_115_297#_c_433_n 0.0114839f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A1_c_102_p N_A_115_297#_c_433_n 0.0106067f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_135 N_A1_c_88_n N_A_115_297#_c_433_n 3.31919e-19 $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A1_c_90_n N_A_115_297#_c_433_n 0.0285775f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_137 N_A1_M1002_g N_A_115_297#_c_438_n 0.00154364f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_c_88_n N_A_115_297#_c_438_n 3.74059e-19 $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A1_c_90_n N_A_115_297#_c_438_n 0.0117058f $X=1.475 $Y=1.35 $X2=0 $Y2=0
cc_140 N_A1_M1020_g N_A_115_297#_c_441_n 0.00251621f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A1_c_102_p N_A_115_297#_c_441_n 0.00304589f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_142 N_A1_c_102_p N_Y_M1000_d 0.00432239f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_143 N_A1_c_102_p N_Y_M1013_d 0.00331496f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_144 N_A1_M1007_g N_Y_c_476_n 3.6643e-19 $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1020_g N_Y_c_476_n 0.012038f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_c_102_p N_Y_c_476_n 0.0958491f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_147 N_A1_c_86_n N_Y_c_476_n 2.92808e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A1_c_89_n N_Y_c_480_n 2.12504e-19 $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A1_M1020_g N_Y_c_470_n 0.00121728f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A1_c_102_p N_Y_c_470_n 0.0113729f $X=3.445 $Y=1.6 $X2=0 $Y2=0
cc_151 N_A1_c_85_n N_Y_c_470_n 0.00436123f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A1_c_82_n N_A_32_47#_c_548_n 0.0105709f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_83_n N_A_32_47#_c_548_n 0.0105709f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_84_n N_A_32_47#_c_548_n 0.0105146f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A1_c_85_n N_A_32_47#_c_548_n 0.0167224f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A1_c_86_n N_A_32_47#_c_548_n 0.0029684f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_87_n N_A_32_47#_c_548_n 0.0820457f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A1_c_88_n N_A_32_47#_c_548_n 0.0111987f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_c_89_n N_A_32_47#_c_548_n 0.0116597f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A1_c_82_n N_VGND_c_602_n 0.0141001f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_c_83_n N_VGND_c_602_n 0.00765006f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A1_c_84_n N_VGND_c_602_n 0.00104385f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_83_n N_VGND_c_603_n 0.00104385f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_84_n N_VGND_c_603_n 0.0076143f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_89_n N_VGND_c_605_n 0.00315951f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_82_n N_VGND_c_608_n 0.00351072f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_c_83_n N_VGND_c_609_n 0.00351072f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_84_n N_VGND_c_609_n 0.00351072f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_89_n N_VGND_c_611_n 0.00422112f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_82_n N_VGND_c_612_n 0.00510895f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_83_n N_VGND_c_612_n 0.00411677f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A1_c_84_n N_VGND_c_612_n 0.00411677f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_89_n N_VGND_c_612_n 0.00577486f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_M1000_g N_VPWR_c_335_n 0.00107483f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A2_M1000_g N_VPWR_c_339_n 0.00357877f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A2_M1008_g N_VPWR_c_339_n 0.00357877f $X=2.22 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1013_g N_VPWR_c_339_n 0.00357877f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_M1016_g N_VPWR_c_339_n 0.00357877f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_M1000_g N_VPWR_c_332_n 0.00530427f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A2_M1008_g N_VPWR_c_332_n 0.00527894f $X=2.22 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A2_M1013_g N_VPWR_c_332_n 0.00527894f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A2_M1016_g N_VPWR_c_332_n 0.00530427f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A2_M1000_g N_A_115_297#_c_441_n 0.00996109f $X=1.79 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A2_M1008_g N_A_115_297#_c_441_n 0.00863252f $X=2.22 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A2_M1013_g N_A_115_297#_c_441_n 0.00868463f $X=2.65 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A2_M1016_g N_A_115_297#_c_441_n 0.00868463f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A2_M1000_g N_Y_c_476_n 0.00299008f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_M1008_g N_Y_c_476_n 0.00888044f $X=2.22 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A2_M1013_g N_Y_c_476_n 0.00888044f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A2_M1016_g N_Y_c_476_n 0.00883388f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A2_c_192_n N_A_32_47#_c_548_n 0.0150408f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_193_n N_A_32_47#_c_548_n 0.0108891f $X=2.22 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_194_n N_A_32_47#_c_548_n 0.0108891f $X=2.65 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_195_n N_A_32_47#_c_548_n 0.0111048f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_196_n N_A_32_47#_c_548_n 0.0605407f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A2_c_197_n N_A_32_47#_c_548_n 0.0074458f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A2_c_192_n N_VGND_c_603_n 0.0076143f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_193_n N_VGND_c_603_n 0.00104385f $X=2.22 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_192_n N_VGND_c_604_n 0.00104385f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_193_n N_VGND_c_604_n 0.00765006f $X=2.22 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_c_194_n N_VGND_c_604_n 0.00765006f $X=2.65 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A2_c_195_n N_VGND_c_604_n 0.00104385f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_c_194_n N_VGND_c_605_n 0.00104385f $X=2.65 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_c_195_n N_VGND_c_605_n 0.00757635f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_c_192_n N_VGND_c_606_n 0.00351072f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A2_c_193_n N_VGND_c_606_n 0.00351072f $X=2.22 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A2_c_194_n N_VGND_c_610_n 0.00351072f $X=2.65 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A2_c_195_n N_VGND_c_610_n 0.00351072f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A2_c_192_n N_VGND_c_612_n 0.00411677f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A2_c_193_n N_VGND_c_612_n 0.00411677f $X=2.22 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A2_c_194_n N_VGND_c_612_n 0.00411677f $X=2.65 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A2_c_195_n N_VGND_c_612_n 0.00411677f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_M1006_g N_VPWR_c_336_n 0.00562133f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1011_g N_VPWR_c_336_n 5.00193e-19 $X=4.41 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1006_g N_VPWR_c_337_n 5.12235e-19 $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_M1011_g N_VPWR_c_337_n 0.00650396f $X=4.41 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B1_M1014_g N_VPWR_c_337_n 0.00645747f $X=4.84 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_M1023_g N_VPWR_c_337_n 5.0423e-19 $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B1_M1014_g N_VPWR_c_338_n 6.41224e-19 $X=4.84 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B1_M1023_g N_VPWR_c_338_n 0.0113107f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B1_M1006_g N_VPWR_c_341_n 0.00418382f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_222 N_B1_M1011_g N_VPWR_c_341_n 0.00353537f $X=4.41 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B1_M1014_g N_VPWR_c_343_n 0.00353537f $X=4.84 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B1_M1023_g N_VPWR_c_343_n 0.00486043f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B1_M1006_g N_VPWR_c_332_n 0.00482373f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B1_M1011_g N_VPWR_c_332_n 0.00411309f $X=4.41 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B1_M1014_g N_VPWR_c_332_n 0.00411309f $X=4.84 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B1_M1023_g N_VPWR_c_332_n 0.00822531f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B1_M1006_g N_Y_c_476_n 0.00401099f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_230 N_B1_c_267_n N_Y_c_476_n 7.51756e-19 $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B1_c_263_n N_Y_c_480_n 0.00319406f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B1_c_264_n N_Y_c_480_n 0.0100285f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_265_n N_Y_c_480_n 0.0100285f $X=4.84 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B1_c_266_n N_Y_c_480_n 0.0135749f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B1_c_267_n N_Y_c_480_n 0.0767656f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B1_c_268_n N_Y_c_480_n 0.00693528f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B1_M1011_g N_Y_c_469_n 0.0246931f $X=4.41 $Y=1.985 $X2=0 $Y2=0
cc_238 N_B1_M1014_g N_Y_c_469_n 0.0247479f $X=4.84 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B1_c_267_n N_Y_c_469_n 0.0536254f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B1_c_268_n N_Y_c_469_n 0.00246447f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B1_M1006_g N_Y_c_470_n 0.0178506f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_242 N_B1_c_267_n N_Y_c_470_n 0.0287708f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B1_c_268_n N_Y_c_470_n 0.00247486f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_244 N_B1_M1023_g N_Y_c_471_n 0.0208171f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_245 N_B1_c_267_n N_Y_c_471_n 0.00772446f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_246 N_B1_c_267_n N_Y_c_472_n 0.0157676f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B1_c_268_n N_Y_c_472_n 0.00247486f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B1_c_266_n Y 0.0225795f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B1_c_267_n Y 0.0220074f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B1_c_263_n N_A_32_47#_c_549_n 0.0107278f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B1_c_264_n N_A_32_47#_c_549_n 0.00816381f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_c_265_n N_A_32_47#_c_549_n 0.00821592f $X=4.84 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B1_c_266_n N_A_32_47#_c_549_n 0.00821592f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B1_c_267_n N_A_32_47#_c_549_n 0.00324863f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B1_c_263_n N_VGND_c_611_n 0.00357877f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_256 N_B1_c_264_n N_VGND_c_611_n 0.00357877f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B1_c_265_n N_VGND_c_611_n 0.00357877f $X=4.84 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B1_c_266_n N_VGND_c_611_n 0.00357877f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_259 N_B1_c_263_n N_VGND_c_612_n 0.00534514f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B1_c_264_n N_VGND_c_612_n 0.00527894f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B1_c_265_n N_VGND_c_612_n 0.00527894f $X=4.84 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B1_c_266_n N_VGND_c_612_n 0.00637081f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_263 N_VPWR_c_332_n N_A_115_297#_M1002_d 0.0023848f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_264 N_VPWR_c_332_n N_A_115_297#_M1007_d 0.00239287f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_332_n N_A_115_297#_M1008_s 0.00223258f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_332_n N_A_115_297#_M1016_s 0.00223258f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_345_n N_A_115_297#_c_451_n 0.0138713f $X=0.98 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_332_n N_A_115_297#_c_451_n 0.00892401f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_M1004_s N_A_115_297#_c_433_n 0.003602f $X=1.005 $Y=1.485 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_335_n N_A_115_297#_c_433_n 0.0160114f $X=1.145 $Y=2.34 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_339_n N_A_115_297#_c_433_n 0.00247598f $X=3.63 $Y=2.72 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_345_n N_A_115_297#_c_433_n 0.00247598f $X=0.98 $Y=2.72 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_332_n N_A_115_297#_c_433_n 0.00979637f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_339_n N_A_115_297#_c_458_n 0.0123456f $X=3.63 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_332_n N_A_115_297#_c_458_n 0.00727709f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_339_n N_A_115_297#_c_441_n 0.0986739f $X=3.63 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_332_n N_A_115_297#_c_441_n 0.0636286f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_332_n N_Y_M1000_d 0.00224864f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_332_n N_Y_M1013_d 0.00224864f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_332_n N_Y_M1006_s 0.00248504f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_332_n N_Y_M1014_s 0.00394701f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_M1020_s N_Y_c_476_n 0.00846156f $X=3.585 $Y=1.485 $X2=0 $Y2=0
cc_283 N_VPWR_c_336_n N_Y_c_476_n 0.0162461f $X=3.745 $Y=2.36 $X2=0 $Y2=0
cc_284 N_VPWR_c_339_n N_Y_c_476_n 0.00215462f $X=3.63 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_341_n N_Y_c_476_n 3.42949e-19 $X=4.46 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_332_n N_Y_c_476_n 0.00943415f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_287 N_VPWR_c_341_n N_Y_c_518_n 0.0131634f $X=4.46 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_332_n N_Y_c_518_n 0.00801045f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_M1011_d N_Y_c_469_n 0.0017682f $X=4.485 $Y=1.485 $X2=0 $Y2=0
cc_290 N_VPWR_c_337_n N_Y_c_469_n 0.0175341f $X=4.625 $Y=2.34 $X2=0 $Y2=0
cc_291 N_VPWR_c_341_n N_Y_c_469_n 0.00266112f $X=4.46 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_343_n N_Y_c_469_n 0.00266112f $X=5.32 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_332_n N_Y_c_469_n 0.0105156f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_341_n N_Y_c_470_n 0.00207595f $X=4.46 $Y=2.72 $X2=0 $Y2=0
cc_295 N_VPWR_c_332_n N_Y_c_470_n 0.00348792f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_343_n N_Y_c_527_n 0.0124538f $X=5.32 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_332_n N_Y_c_527_n 0.00724021f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_M1023_d N_Y_c_471_n 0.00335153f $X=5.345 $Y=1.485 $X2=0 $Y2=0
cc_299 N_VPWR_c_338_n N_Y_c_471_n 0.0230476f $X=5.485 $Y=1.965 $X2=0 $Y2=0
cc_300 N_A_115_297#_c_441_n N_Y_M1000_d 0.00367283f $X=3.295 $Y=2.36 $X2=0.5
+ $Y2=0.56
cc_301 N_A_115_297#_c_441_n N_Y_M1013_d 0.00367283f $X=3.295 $Y=2.36 $X2=0.5
+ $Y2=1.325
cc_302 N_A_115_297#_M1008_s N_Y_c_476_n 0.00368596f $X=2.295 $Y=1.485 $X2=1.36
+ $Y2=1.985
cc_303 N_A_115_297#_M1016_s N_Y_c_476_n 0.0037815f $X=3.155 $Y=1.485 $X2=1.36
+ $Y2=1.985
cc_304 N_A_115_297#_c_441_n N_Y_c_476_n 0.055936f $X=3.295 $Y=2.36 $X2=1.36
+ $Y2=1.985
cc_305 N_Y_c_480_n N_A_32_47#_M1003_s 0.00326005f $X=5.425 $Y=0.73 $X2=0 $Y2=0
cc_306 N_Y_c_480_n N_A_32_47#_M1015_s 6.38324e-19 $X=5.425 $Y=0.73 $X2=0 $Y2=0
cc_307 N_Y_c_467_n N_A_32_47#_M1015_s 0.00351563f $X=5.63 $Y=0.845 $X2=0 $Y2=0
cc_308 Y N_A_32_47#_M1015_s 7.06752e-19 $X=5.75 $Y=0.85 $X2=0 $Y2=0
cc_309 N_Y_M1001_d N_A_32_47#_c_549_n 0.00323484f $X=4.055 $Y=0.235 $X2=0 $Y2=0
cc_310 N_Y_M1010_d N_A_32_47#_c_549_n 0.00323484f $X=4.915 $Y=0.235 $X2=0 $Y2=0
cc_311 N_Y_c_480_n N_A_32_47#_c_549_n 0.0680193f $X=5.425 $Y=0.73 $X2=0 $Y2=0
cc_312 N_Y_c_467_n N_A_32_47#_c_549_n 0.0174133f $X=5.63 $Y=0.845 $X2=0 $Y2=0
cc_313 N_Y_c_467_n N_VGND_c_611_n 0.00391741f $X=5.63 $Y=0.845 $X2=0 $Y2=0
cc_314 N_Y_M1001_d N_VGND_c_612_n 0.00224864f $X=4.055 $Y=0.235 $X2=0 $Y2=0
cc_315 N_Y_M1010_d N_VGND_c_612_n 0.00224864f $X=4.915 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_c_467_n N_VGND_c_612_n 0.00624163f $X=5.63 $Y=0.845 $X2=0 $Y2=0
cc_317 N_A_32_47#_c_548_n N_VGND_M1012_d 0.00333948f $X=3.63 $Y=0.717 $X2=-0.19
+ $Y2=-0.24
cc_318 N_A_32_47#_c_548_n N_VGND_M1021_d 0.00817986f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_319 N_A_32_47#_c_548_n N_VGND_M1009_d 0.00352426f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_320 N_A_32_47#_c_548_n N_VGND_M1019_d 0.00705641f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_321 N_A_32_47#_c_548_n N_VGND_c_602_n 0.0161049f $X=3.63 $Y=0.717 $X2=0 $Y2=0
cc_322 N_A_32_47#_c_548_n N_VGND_c_603_n 0.0161049f $X=3.63 $Y=0.717 $X2=0 $Y2=0
cc_323 N_A_32_47#_c_548_n N_VGND_c_604_n 0.0161049f $X=3.63 $Y=0.717 $X2=0 $Y2=0
cc_324 N_A_32_47#_c_548_n N_VGND_c_605_n 0.0174908f $X=3.63 $Y=0.717 $X2=0 $Y2=0
cc_325 N_A_32_47#_c_548_n N_VGND_c_606_n 0.00855504f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_326 N_A_32_47#_c_548_n N_VGND_c_608_n 0.00736721f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_327 N_A_32_47#_c_548_n N_VGND_c_609_n 0.00855504f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_328 N_A_32_47#_c_548_n N_VGND_c_610_n 0.00855504f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_329 N_A_32_47#_c_548_n N_VGND_c_611_n 0.00279155f $X=3.63 $Y=0.717 $X2=0
+ $Y2=0
cc_330 N_A_32_47#_c_590_p N_VGND_c_611_n 0.0137873f $X=3.86 $Y=0.35 $X2=0 $Y2=0
cc_331 N_A_32_47#_c_549_n N_VGND_c_611_n 0.100426f $X=5.485 $Y=0.36 $X2=0 $Y2=0
cc_332 N_A_32_47#_M1012_s N_VGND_c_612_n 0.0030331f $X=0.16 $Y=0.235 $X2=0 $Y2=0
cc_333 N_A_32_47#_M1017_s N_VGND_c_612_n 0.00318969f $X=1.005 $Y=0.235 $X2=0
+ $Y2=0
cc_334 N_A_32_47#_M1005_s N_VGND_c_612_n 0.00318969f $X=1.865 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_A_32_47#_M1018_s N_VGND_c_612_n 0.00318969f $X=2.725 $Y=0.235 $X2=0
+ $Y2=0
cc_336 N_A_32_47#_M1022_s N_VGND_c_612_n 0.00226522f $X=3.625 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_A_32_47#_M1003_s N_VGND_c_612_n 0.00223258f $X=4.485 $Y=0.235 $X2=0
+ $Y2=0
cc_338 N_A_32_47#_M1015_s N_VGND_c_612_n 0.00229841f $X=5.345 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_32_47#_c_548_n N_VGND_c_612_n 0.0645215f $X=3.63 $Y=0.717 $X2=0 $Y2=0
cc_340 N_A_32_47#_c_590_p N_VGND_c_612_n 0.00881516f $X=3.86 $Y=0.35 $X2=0 $Y2=0
cc_341 N_A_32_47#_c_549_n N_VGND_c_612_n 0.0638826f $X=5.485 $Y=0.36 $X2=0 $Y2=0

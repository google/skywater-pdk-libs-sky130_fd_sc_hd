* File: sky130_fd_sc_hd__edfxbp_1.spice.pex
* Created: Thu Aug 27 14:19:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%CLK 1 2 3 5 6 8 11 13
c40 1 0 2.71124e-20 $X=0.31 $Y=1.325
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r42 9 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.47 $Y2=1.665
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r44 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r45 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r46 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r47 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r48 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r49 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_27_47# 1 2 9 13 17 21 25 27 31 35 39 40
+ 41 44 46 48 51 54 56 57 58 59 60 67 69 74 82 85 89
c250 89 0 1.92554e-19 $X=7.875 $Y=1.41
c251 51 0 1.74912e-19 $X=4.98 $Y=0.87
c252 48 0 1.43548e-19 $X=5.15 $Y=0.845
c253 44 0 1.8506e-19 $X=0.73 $Y=1.795
c254 41 0 5.65522e-20 $X=0.615 $Y=1.88
r255 88 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.875 $Y=1.41
+ $X2=7.875 $Y2=1.575
r256 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.875
+ $Y=1.41 $X2=7.875 $Y2=1.41
r257 85 88 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.875 $Y=1.32
+ $X2=7.875 $Y2=1.41
r258 79 82 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.31 $Y=1.74
+ $X2=5.405 $Y2=1.74
r259 70 89 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=7.885 $Y=1.87
+ $X2=7.885 $Y2=1.41
r260 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.885 $Y=1.87
+ $X2=7.885 $Y2=1.87
r261 67 96 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=5.295 $Y=1.83
+ $X2=5.235 $Y2=1.83
r262 67 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.74 $X2=5.405 $Y2=1.74
r263 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.295 $Y=1.87
+ $X2=5.295 $Y2=1.87
r264 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=1.87
r265 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.44 $Y=1.87
+ $X2=5.295 $Y2=1.87
r266 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.74 $Y=1.87
+ $X2=7.885 $Y2=1.87
r267 59 60 2.84653 $w=1.4e-07 $l=2.3e-06 $layer=MET1_cond $X=7.74 $Y=1.87
+ $X2=5.44 $Y2=1.87
r268 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=1.87
+ $X2=0.72 $Y2=1.87
r269 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.15 $Y=1.87
+ $X2=5.295 $Y2=1.87
r270 57 58 5.30321 $w=1.4e-07 $l=4.285e-06 $layer=MET1_cond $X=5.15 $Y=1.87
+ $X2=0.865 $Y2=1.87
r271 54 96 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.235 $Y=1.655
+ $X2=5.235 $Y2=1.83
r272 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.235 $Y=0.955
+ $X2=5.235 $Y2=1.655
r273 51 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.98 $Y=0.87
+ $X2=4.98 $Y2=0.735
r274 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=0.87 $X2=4.98 $Y2=0.87
r275 48 53 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.15 $Y=0.845
+ $X2=5.235 $Y2=0.955
r276 48 50 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=5.15 $Y=0.845
+ $X2=4.98 $Y2=0.845
r277 47 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r278 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r279 44 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r280 44 46 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r281 43 46 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.73 $Y=0.805
+ $X2=0.73 $Y2=1.235
r282 42 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r283 41 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r284 41 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.345 $Y2=1.88
r285 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.73 $Y2=0.805
r286 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r287 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r288 33 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r289 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=8.51 $Y=1.245
+ $X2=8.51 $Y2=0.415
r290 28 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.01 $Y=1.32
+ $X2=7.875 $Y2=1.32
r291 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.435 $Y=1.32
+ $X2=8.51 $Y2=1.245
r292 27 28 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=8.435 $Y=1.32
+ $X2=8.01 $Y2=1.32
r293 25 90 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=7.88 $Y=2.275
+ $X2=7.88 $Y2=1.575
r294 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.905
+ $X2=5.31 $Y2=1.74
r295 19 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.31 $Y=1.905
+ $X2=5.31 $Y2=2.275
r296 17 77 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.99 $Y=0.415
+ $X2=4.99 $Y2=0.735
r297 11 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r298 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r299 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r300 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r301 2 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r302 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%D 3 7 9 12 13 16
c51 7 0 5.26342e-20 $X=1.83 $Y=2.165
r52 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.78
+ $Y=1.145 $X2=1.78 $Y2=1.145
r53 11 16 70.9845 $w=3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.765 $Y=1.5
+ $X2=1.765 $Y2=1.145
r54 11 12 43.217 $w=3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.765 $Y=1.5 $X2=1.765
+ $Y2=1.65
r55 9 16 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.765 $Y=1.13 $X2=1.765
+ $Y2=1.145
r56 9 10 43.217 $w=3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.765 $Y=1.13 $X2=1.765
+ $Y2=0.98
r57 7 12 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.83 $Y=2.165
+ $X2=1.83 $Y2=1.65
r58 3 10 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_423_343# 1 2 7 9 12 16 20 23 26 27 36
c88 27 0 1.67735e-19 $X=3.55 $Y=1.01
c89 23 0 5.26342e-20 $X=2.932 $Y=1.355
c90 20 0 1.1082e-19 $X=2.92 $Y=0.51
r91 30 33 10.7351 $w=3.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.58 $Y=1.537
+ $X2=2.92 $Y2=1.537
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.52 $X2=2.58 $Y2=1.52
r93 27 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.01
+ $X2=3.55 $Y2=0.845
r94 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.01 $X2=3.55 $Y2=1.01
r95 24 36 0.565906 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=3.085 $Y=1.01
+ $X2=2.932 $Y2=1.01
r96 24 26 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.085 $Y=1.01
+ $X2=3.55 $Y2=1.01
r97 23 33 0.378885 $w=3.63e-07 $l=1.2e-08 $layer=LI1_cond $X=2.932 $Y=1.537
+ $X2=2.92 $Y2=1.537
r98 22 36 6.17543 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=2.932 $Y=1.175
+ $X2=2.932 $Y2=1.01
r99 22 23 6.8013 $w=3.03e-07 $l=1.8e-07 $layer=LI1_cond $X=2.932 $Y=1.175
+ $X2=2.932 $Y2=1.355
r100 18 36 6.17543 $w=2.65e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.892 $Y=0.845
+ $X2=2.932 $Y2=1.01
r101 18 20 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=2.892 $Y=0.845
+ $X2=2.892 $Y2=0.51
r102 14 33 1.32393 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=2.92 $Y=1.72
+ $X2=2.92 $Y2=1.537
r103 14 16 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.92 $Y=1.72
+ $X2=2.92 $Y2=1.99
r104 12 40 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.57 $Y=0.445
+ $X2=3.57 $Y2=0.845
r105 7 31 69.3653 $w=2.71e-07 $l=4.76833e-07 $layer=POLY_cond $X=2.19 $Y=1.77
+ $X2=2.58 $Y2=1.577
r106 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.19 $Y=1.77
+ $X2=2.19 $Y2=2.165
r107 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=1.845 $X2=2.92 $Y2=1.99
r108 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.92 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%DE 3 5 6 9 12 15 17 21 23 24 25
c85 6 0 1.1082e-19 $X=2.455 $Y=0.925
r86 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.01 $X2=2.29 $Y2=1.01
r87 27 29 13.5393 $w=3.56e-07 $l=1e-07 $layer=POLY_cond $X=2.19 $Y=0.992
+ $X2=2.29 $Y2=0.992
r88 25 30 5.12336 $w=3.81e-07 $l=1.6e-07 $layer=LI1_cond $X=2.337 $Y=0.85
+ $X2=2.337 $Y2=1.01
r89 19 21 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.57 $Y=1.61
+ $X2=3.57 $Y2=2.165
r90 18 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.205 $Y=1.535
+ $X2=3.13 $Y2=1.535
r91 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.495 $Y=1.535
+ $X2=3.57 $Y2=1.61
r92 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.495 $Y=1.535
+ $X2=3.205 $Y2=1.535
r93 13 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.61
+ $X2=3.13 $Y2=1.535
r94 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.13 $Y=1.61
+ $X2=3.13 $Y2=2.165
r95 12 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.46
+ $X2=3.13 $Y2=1.535
r96 11 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1 $X2=3.13
+ $Y2=0.925
r97 11 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.13 $Y=1 $X2=3.13
+ $Y2=1.46
r98 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=0.85 $X2=3.13
+ $Y2=0.925
r99 7 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.13 $Y=0.85 $X2=3.13
+ $Y2=0.445
r100 6 29 38.8573 $w=3.56e-07 $l=1.95653e-07 $layer=POLY_cond $X=2.455 $Y=0.925
+ $X2=2.29 $Y2=0.992
r101 5 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=0.925
+ $X2=3.13 $Y2=0.925
r102 5 6 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.055 $Y=0.925 $X2=2.455
+ $Y2=0.925
r103 1 27 23.0368 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.19 $Y=0.81
+ $X2=2.19 $Y2=0.992
r104 1 3 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.19 $Y=0.81 $X2=2.19
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_791_264# 1 2 9 13 17 21 23 24 27 31 33 34
+ 42 48 49 53 55 58 59 62 65 78
c195 53 0 1.11291e-19 $X=10.1 $Y=1.055
r196 66 78 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=10.47 $Y=0.85
+ $X2=10.47 $Y2=0.385
r197 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.475 $Y=0.85
+ $X2=10.475 $Y2=0.85
r198 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.89 $Y=0.85
+ $X2=3.89 $Y2=0.85
r199 59 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.035 $Y=0.85
+ $X2=3.89 $Y2=0.85
r200 58 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.33 $Y=0.85
+ $X2=10.475 $Y2=0.85
r201 58 59 7.79083 $w=1.4e-07 $l=6.295e-06 $layer=MET1_cond $X=10.33 $Y=0.85
+ $X2=4.035 $Y2=0.85
r202 56 66 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=10.47 $Y=0.89
+ $X2=10.47 $Y2=0.85
r203 55 56 0.533618 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=10.47 $Y=1.055
+ $X2=10.47 $Y2=0.89
r204 53 73 15.9965 $w=2.7e-07 $l=7.2e-08 $layer=POLY_cond $X=10.1 $Y=1.055
+ $X2=10.1 $Y2=1.127
r205 52 55 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.1 $Y=1.055
+ $X2=10.47 $Y2=1.055
r206 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.1
+ $Y=1.055 $X2=10.1 $Y2=1.055
r207 49 70 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.485
+ $X2=4.09 $Y2=1.65
r208 49 69 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.485
+ $X2=4.09 $Y2=1.32
r209 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.485 $X2=4.09 $Y2=1.485
r210 45 62 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.89 $Y=1.32
+ $X2=3.89 $Y2=0.85
r211 44 48 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.89 $Y=1.485 $X2=4.09
+ $Y2=1.485
r212 44 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=1.485
+ $X2=3.89 $Y2=1.32
r213 40 55 0.533618 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=10.47 $Y=1.22
+ $X2=10.47 $Y2=1.055
r214 40 42 26.0994 $w=3.38e-07 $l=7.7e-07 $layer=LI1_cond $X=10.47 $Y=1.22
+ $X2=10.47 $Y2=1.99
r215 33 73 11.7477 $w=1.85e-07 $l=1.35e-07 $layer=POLY_cond $X=9.965 $Y=1.127
+ $X2=10.1 $Y2=1.127
r216 33 34 155.158 $w=1.85e-07 $l=4.2e-07 $layer=POLY_cond $X=9.965 $Y=1.127
+ $X2=9.545 $Y2=1.127
r217 29 34 27.7067 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=9.47 $Y=1.127
+ $X2=9.545 $Y2=1.127
r218 29 38 42.4837 $w=1.85e-07 $l=1.15e-07 $layer=POLY_cond $X=9.47 $Y=1.127
+ $X2=9.355 $Y2=1.127
r219 29 31 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=9.47 $Y=1.035
+ $X2=9.47 $Y2=0.56
r220 25 38 7.77431 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=9.355 $Y=1.22
+ $X2=9.355 $Y2=1.127
r221 25 27 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=9.355 $Y=1.22
+ $X2=9.355 $Y2=1.985
r222 23 38 27.7067 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=9.28 $Y=1.127
+ $X2=9.355 $Y2=1.127
r223 23 24 81.2731 $w=1.85e-07 $l=2.2e-07 $layer=POLY_cond $X=9.28 $Y=1.127
+ $X2=9.06 $Y2=1.127
r224 19 24 27.7067 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=8.985 $Y=1.127
+ $X2=9.06 $Y2=1.127
r225 19 35 42.4837 $w=1.85e-07 $l=1.15e-07 $layer=POLY_cond $X=8.985 $Y=1.127
+ $X2=8.87 $Y2=1.127
r226 19 21 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.985 $Y=1.035
+ $X2=8.985 $Y2=0.445
r227 15 35 7.77431 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=8.87 $Y=1.22
+ $X2=8.87 $Y2=1.127
r228 15 17 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=8.87 $Y=1.22
+ $X2=8.87 $Y2=2.275
r229 13 70 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.08 $Y=2.165
+ $X2=4.08 $Y2=1.65
r230 9 69 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.08 $Y=0.445
+ $X2=4.08 $Y2=1.32
r231 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.34
+ $Y=1.845 $X2=10.465 $Y2=1.99
r232 1 78 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=10.35
+ $Y=0.235 $X2=10.475 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_193_47# 1 2 9 11 15 17 19 22 26 27 30 31
+ 32 33 42 43 45 49 58 62
c196 33 0 1.37287e-19 $X=5.03 $Y=1.53
c197 32 0 3.76247e-20 $X=8.16 $Y=1.53
c198 22 0 1.92554e-19 $X=8.3 $Y=2.275
c199 11 0 1.43548e-19 $X=5.355 $Y=1.29
r200 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.385
+ $Y=1.74 $X2=8.385 $Y2=1.74
r201 55 58 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=8.3 $Y=1.74
+ $X2=8.385 $Y2=1.74
r202 48 50 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.88 $Y=1.35
+ $X2=4.88 $Y2=1.485
r203 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.88
+ $Y=1.35 $X2=4.88 $Y2=1.35
r204 45 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.88 $Y=1.29 $X2=4.88
+ $Y2=1.35
r205 43 59 7.56291 $w=3.18e-07 $l=2.1e-07 $layer=LI1_cond $X=8.31 $Y=1.53
+ $X2=8.31 $Y2=1.74
r206 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.305 $Y=1.53
+ $X2=8.305 $Y2=1.53
r207 40 49 10.7912 $w=1.83e-07 $l=1.8e-07 $layer=LI1_cond $X=4.887 $Y=1.53
+ $X2=4.887 $Y2=1.35
r208 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.885 $Y=1.53
+ $X2=4.885 $Y2=1.53
r209 36 66 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.1 $Y=1.53 $X2=1.1
+ $Y2=1.96
r210 36 62 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.1 $Y=1.53
+ $X2=1.1 $Y2=0.51
r211 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.53 $X2=1.1
+ $Y2=1.53
r212 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.53
+ $X2=4.885 $Y2=1.53
r213 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.16 $Y=1.53
+ $X2=8.305 $Y2=1.53
r214 32 33 3.87375 $w=1.4e-07 $l=3.13e-06 $layer=MET1_cond $X=8.16 $Y=1.53
+ $X2=5.03 $Y2=1.53
r215 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.53
+ $X2=1.1 $Y2=1.53
r216 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.74 $Y=1.53
+ $X2=4.885 $Y2=1.53
r217 30 31 4.32549 $w=1.4e-07 $l=3.495e-06 $layer=MET1_cond $X=4.74 $Y=1.53
+ $X2=1.245 $Y2=1.53
r218 29 43 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=8.31 $Y=1.035
+ $X2=8.31 $Y2=1.53
r219 27 51 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.09 $Y=0.87
+ $X2=7.98 $Y2=0.87
r220 26 29 5.41706 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.237 $Y=0.87
+ $X2=8.237 $Y2=1.035
r221 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=0.87 $X2=8.09 $Y2=0.87
r222 20 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.3 $Y=1.875
+ $X2=8.3 $Y2=1.74
r223 20 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.3 $Y=1.875 $X2=8.3
+ $Y2=2.275
r224 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.98 $Y=0.705
+ $X2=7.98 $Y2=0.87
r225 17 19 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.98 $Y=0.705
+ $X2=7.98 $Y2=0.415
r226 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.43 $Y=1.215
+ $X2=5.43 $Y2=0.415
r227 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.045 $Y=1.29
+ $X2=4.88 $Y2=1.29
r228 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.355 $Y=1.29
+ $X2=5.43 $Y2=1.215
r229 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=5.355 $Y=1.29
+ $X2=5.045 $Y2=1.29
r230 9 50 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.855 $Y=2.275
+ $X2=4.855 $Y2=1.485
r231 2 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r232 1 62 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_1150_159# 1 2 9 13 17 21 25 27 28 32 36
+ 40 41 47 55
c118 40 0 6.28645e-20 $X=7.36 $Y=1.21
r119 49 50 5.12431 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=6.732 $Y=1.21
+ $X2=6.732 $Y2=1.375
r120 45 55 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=5.955 $Y=0.93
+ $X2=5.96 $Y2=0.93
r121 45 52 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=5.955 $Y=0.93
+ $X2=5.825 $Y2=0.93
r122 44 47 4.13427 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.955 $Y=0.93
+ $X2=6.07 $Y2=0.93
r123 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.955
+ $Y=0.93 $X2=5.955 $Y2=0.93
r124 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.36
+ $Y=1.21 $X2=7.36 $Y2=1.21
r125 38 49 1.93884 $w=3.3e-07 $l=2.03e-07 $layer=LI1_cond $X=6.935 $Y=1.21
+ $X2=6.732 $Y2=1.21
r126 38 40 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=6.935 $Y=1.21
+ $X2=7.36 $Y2=1.21
r127 36 50 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.695 $Y=1.88
+ $X2=6.695 $Y2=1.375
r128 30 32 10.6708 $w=4.03e-07 $l=3.75e-07 $layer=LI1_cond $X=6.732 $Y=0.765
+ $X2=6.732 $Y2=0.39
r129 28 49 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=6.732 $Y=0.915
+ $X2=6.732 $Y2=1.21
r130 28 30 4.26831 $w=4.03e-07 $l=1.5e-07 $layer=LI1_cond $X=6.732 $Y=0.915
+ $X2=6.732 $Y2=0.765
r131 28 47 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.53 $Y=0.915
+ $X2=6.07 $Y2=0.915
r132 26 41 6.10776 $w=2.75e-07 $l=2.8e-08 $layer=POLY_cond $X=7.362 $Y=1.238
+ $X2=7.362 $Y2=1.21
r133 26 27 42.1909 $w=2.75e-07 $l=1.37e-07 $layer=POLY_cond $X=7.362 $Y=1.238
+ $X2=7.362 $Y2=1.375
r134 25 41 35.9921 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.362 $Y=1.045
+ $X2=7.362 $Y2=1.21
r135 24 25 45.0266 $w=2.75e-07 $l=1.5e-07 $layer=POLY_cond $X=7.397 $Y=0.895
+ $X2=7.397 $Y2=1.045
r136 21 24 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.495 $Y=0.445
+ $X2=7.495 $Y2=0.895
r137 17 27 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=7.425 $Y=2.275
+ $X2=7.425 $Y2=1.375
r138 11 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.96 $Y=0.795
+ $X2=5.96 $Y2=0.93
r139 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.96 $Y=0.795
+ $X2=5.96 $Y2=0.445
r140 7 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.825 $Y=1.065
+ $X2=5.825 $Y2=0.93
r141 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.825 $Y=1.065
+ $X2=5.825 $Y2=2.275
r142 2 36 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.56
+ $Y=1.735 $X2=6.695 $Y2=1.88
r143 1 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.63
+ $Y=0.235 $X2=6.765 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_986_413# 1 2 8 11 15 16 17 18 19 20 24 29
+ 31 33
c106 29 0 1.40584e-19 $X=5.595 $Y=1.315
c107 17 0 6.28645e-20 $X=6.52 $Y=1.1
r108 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.275
+ $Y=1.41 $X2=6.275 $Y2=1.41
r109 33 35 20.25 $w=2.44e-07 $l=4.05e-07 $layer=LI1_cond $X=5.87 $Y=1.41
+ $X2=6.275 $Y2=1.41
r110 30 33 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.87 $Y=1.575
+ $X2=5.87 $Y2=1.41
r111 30 31 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.87 $Y=1.575
+ $X2=5.87 $Y2=2.175
r112 29 33 13.75 $w=2.44e-07 $l=2.75e-07 $layer=LI1_cond $X=5.595 $Y=1.41
+ $X2=5.87 $Y2=1.41
r113 28 29 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.595 $Y=0.565
+ $X2=5.595 $Y2=1.315
r114 24 28 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.51 $Y=0.41
+ $X2=5.595 $Y2=0.565
r115 24 26 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=5.51 $Y=0.41
+ $X2=5.2 $Y2=0.41
r116 20 31 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.785 $Y=2.275
+ $X2=5.87 $Y2=2.175
r117 20 22 39.0955 $w=1.98e-07 $l=7.05e-07 $layer=LI1_cond $X=5.785 $Y=2.275
+ $X2=5.08 $Y2=2.275
r118 18 36 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.41 $Y=1.41
+ $X2=6.275 $Y2=1.41
r119 18 19 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.41 $Y=1.41
+ $X2=6.485 $Y2=1.41
r120 16 17 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.52 $Y=0.95
+ $X2=6.52 $Y2=1.1
r121 15 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.555 $Y=0.555
+ $X2=6.555 $Y2=0.95
r122 9 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.485 $Y=1.545
+ $X2=6.485 $Y2=1.41
r123 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.485 $Y=1.545
+ $X2=6.485 $Y2=2.11
r124 8 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.485 $Y=1.275
+ $X2=6.485 $Y2=1.41
r125 8 17 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.485 $Y=1.275
+ $X2=6.485 $Y2=1.1
r126 2 22 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=2.065 $X2=5.08 $Y2=2.275
r127 1 26 182 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_NDIFF $count=1 $X=5.065
+ $Y=0.235 $X2=5.2 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_1591_413# 1 2 7 11 15 17 18 19 21 24 28
+ 29 33 39 40 43 46 49 53
c123 46 0 1.11291e-19 $X=10.015 $Y=1.87
r124 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.015
+ $Y=1.74 $X2=10.015 $Y2=1.74
r125 49 52 43.9904 $w=2.7e-07 $l=1.98e-07 $layer=POLY_cond $X=10.015 $Y=1.542
+ $X2=10.015 $Y2=1.74
r126 46 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.015 $Y=1.87
+ $X2=10.015 $Y2=1.87
r127 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.765 $Y=1.87
+ $X2=8.765 $Y2=1.87
r128 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.91 $Y=1.87
+ $X2=8.765 $Y2=1.87
r129 39 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.87 $Y=1.87
+ $X2=10.015 $Y2=1.87
r130 39 40 1.18812 $w=1.4e-07 $l=9.6e-07 $layer=MET1_cond $X=9.87 $Y=1.87
+ $X2=8.91 $Y2=1.87
r131 38 43 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.765 $Y=2.165
+ $X2=8.765 $Y2=1.87
r132 37 43 61.5405 $w=2.48e-07 $l=1.335e-06 $layer=LI1_cond $X=8.765 $Y=0.535
+ $X2=8.765 $Y2=1.87
r133 33 37 6.90357 $w=2.05e-07 $l=1.68819e-07 $layer=LI1_cond $X=8.64 $Y=0.432
+ $X2=8.765 $Y2=0.535
r134 33 35 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=8.64 $Y=0.432
+ $X2=8.205 $Y2=0.432
r135 29 38 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=8.64 $Y=2.26
+ $X2=8.765 $Y2=2.165
r136 29 31 32.1053 $w=1.88e-07 $l=5.5e-07 $layer=LI1_cond $X=8.64 $Y=2.26
+ $X2=8.09 $Y2=2.26
r137 22 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.17 $Y=1.325
+ $X2=11.17 $Y2=1.16
r138 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.17 $Y=1.325
+ $X2=11.17 $Y2=1.985
r139 19 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.17 $Y=0.995
+ $X2=11.17 $Y2=1.16
r140 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.17 $Y=0.995
+ $X2=11.17 $Y2=0.56
r141 17 28 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.095 $Y=1.16
+ $X2=11.17 $Y2=1.16
r142 17 18 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=11.095 $Y=1.16
+ $X2=10.76 $Y2=1.16
r143 13 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=10.685 $Y=1.655
+ $X2=10.685 $Y2=2.165
r144 9 18 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.685 $Y=0.995
+ $X2=10.685 $Y2=1.16
r145 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.685 $Y=0.995
+ $X2=10.685 $Y2=0.445
r146 8 49 7.22716 $w=2.25e-07 $l=1.35e-07 $layer=POLY_cond $X=10.15 $Y=1.542
+ $X2=10.015 $Y2=1.542
r147 7 13 57.9426 $w=1.5e-07 $l=1.13e-07 $layer=POLY_cond $X=10.685 $Y=1.542
+ $X2=10.685 $Y2=1.655
r148 7 18 195.877 $w=1.5e-07 $l=3.82e-07 $layer=POLY_cond $X=10.685 $Y=1.542
+ $X2=10.685 $Y2=1.16
r149 7 8 131.195 $w=2.25e-07 $l=4.6e-07 $layer=POLY_cond $X=10.61 $Y=1.542
+ $X2=10.15 $Y2=1.542
r150 2 31 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=7.955
+ $Y=2.065 $X2=8.09 $Y2=2.26
r151 1 35 182 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_NDIFF $count=1 $X=8.055
+ $Y=0.235 $X2=8.205 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 38 42 46 52
+ 57 58 60 61 62 64 76 80 92 98 99 102 105 108 111 114
c170 99 0 1.8506e-19 $X=11.73 $Y=2.72
c171 32 0 1.67735e-19 $X=3.35 $Y=1.99
c172 1 0 5.65522e-20 $X=0.545 $Y=1.815
r173 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r174 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r175 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r176 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r177 105 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r178 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r179 99 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=10.81 $Y2=2.72
r180 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r181 96 114 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=11.055 $Y=2.72
+ $X2=10.932 $Y2=2.72
r182 96 98 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=11.055 $Y=2.72
+ $X2=11.73 $Y2=2.72
r183 95 115 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.81 $Y2=2.72
r184 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r185 92 114 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=10.932 $Y2=2.72
r186 92 94 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=9.43 $Y2=2.72
r187 91 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r188 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r189 88 91 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.97 $Y2=2.72
r190 88 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r191 87 90 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=8.97 $Y2=2.72
r192 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r193 85 111 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.36 $Y=2.72
+ $X2=7.215 $Y2=2.72
r194 85 87 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.36 $Y=2.72
+ $X2=7.59 $Y2=2.72
r195 84 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r196 84 106 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.45 $Y2=2.72
r197 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r198 81 105 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.46 $Y=2.72
+ $X2=3.362 $Y2=2.72
r199 81 83 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=3.46 $Y=2.72
+ $X2=5.75 $Y2=2.72
r200 80 108 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.125 $Y=2.72
+ $X2=6.242 $Y2=2.72
r201 80 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.125 $Y=2.72
+ $X2=5.75 $Y2=2.72
r202 79 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r203 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r204 76 105 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.362 $Y2=2.72
r205 76 78 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=2.99 $Y2=2.72
r206 75 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r207 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r208 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r209 72 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r210 71 74 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r211 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r212 69 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r213 69 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r214 64 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r215 64 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r216 62 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r217 62 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r218 60 90 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=9.06 $Y=2.72 $X2=8.97
+ $Y2=2.72
r219 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.06 $Y=2.72
+ $X2=9.145 $Y2=2.72
r220 59 94 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.23 $Y=2.72 $X2=9.43
+ $Y2=2.72
r221 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.23 $Y=2.72
+ $X2=9.145 $Y2=2.72
r222 57 74 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r223 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.4 $Y2=2.72
r224 56 78 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.99 $Y2=2.72
r225 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.4 $Y2=2.72
r226 52 55 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=10.932 $Y=1.63
+ $X2=10.932 $Y2=1.97
r227 50 114 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.932 $Y=2.635
+ $X2=10.932 $Y2=2.72
r228 50 55 31.2806 $w=2.43e-07 $l=6.65e-07 $layer=LI1_cond $X=10.932 $Y=2.635
+ $X2=10.932 $Y2=1.97
r229 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.145 $Y=1.66
+ $X2=9.145 $Y2=2.34
r230 44 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=2.635
+ $X2=9.145 $Y2=2.72
r231 44 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.145 $Y=2.635
+ $X2=9.145 $Y2=2.34
r232 40 111 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=2.635
+ $X2=7.215 $Y2=2.72
r233 40 42 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.215 $Y=2.635
+ $X2=7.215 $Y2=2.275
r234 39 108 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.242 $Y2=2.72
r235 38 111 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.07 $Y=2.72
+ $X2=7.215 $Y2=2.72
r236 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.07 $Y=2.72
+ $X2=6.36 $Y2=2.72
r237 34 108 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.242 $Y=2.635
+ $X2=6.242 $Y2=2.72
r238 34 36 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=6.242 $Y=2.635
+ $X2=6.242 $Y2=2
r239 30 105 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.362 $Y=2.635
+ $X2=3.362 $Y2=2.72
r240 30 32 36.6853 $w=1.93e-07 $l=6.45e-07 $layer=LI1_cond $X=3.362 $Y=2.635
+ $X2=3.362 $Y2=1.99
r241 26 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.635 $X2=2.4
+ $Y2=2.72
r242 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2
r243 22 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r244 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r245 7 55 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=10.76
+ $Y=1.845 $X2=10.96 $Y2=1.97
r246 7 52 600 $w=1.7e-07 $l=2.98706e-07 $layer=licon1_PDIFF $count=1 $X=10.76
+ $Y=1.845 $X2=10.96 $Y2=1.63
r247 6 49 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=2.065 $X2=9.145 $Y2=2.34
r248 6 46 400 $w=1.7e-07 $l=4.95e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=2.065 $X2=9.145 $Y2=1.66
r249 5 42 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=7.09
+ $Y=2.065 $X2=7.215 $Y2=2.275
r250 4 36 300 $w=1.7e-07 $l=3.76098e-07 $layer=licon1_PDIFF $count=2 $X=5.9
+ $Y=2.065 $X2=6.245 $Y2=2
r251 3 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=1.845 $X2=3.35 $Y2=1.99
r252 2 28 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.845 $X2=2.4 $Y2=2
r253 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%A_299_47# 1 2 3 4 20 21 24 25 29 36 38 40
+ 43 48
c120 38 0 1.82232e-19 $X=4.27 $Y=0.51
r121 38 40 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.27 $Y=0.51
+ $X2=4.125 $Y2=0.51
r122 38 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.27 $Y=0.51
+ $X2=4.27 $Y2=0.51
r123 36 40 2.17465 $w=1.85e-07 $l=2.54e-06 $layer=MET1_cond $X=1.585 $Y=0.487
+ $X2=4.125 $Y2=0.487
r124 34 48 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.44 $Y=0.385
+ $X2=1.62 $Y2=0.385
r125 33 36 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.44 $Y=0.51
+ $X2=1.585 $Y2=0.51
r126 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.44 $Y=0.51
+ $X2=1.44 $Y2=0.51
r127 28 43 22.8354 $w=2.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.28 $Y=0.98
+ $X2=4.28 $Y2=0.445
r128 28 29 8.82932 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.33 $Y=0.98
+ $X2=4.33 $Y2=1.15
r129 25 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.43 $Y=1.82
+ $X2=4.43 $Y2=1.15
r130 24 25 9.05087 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=4.32 $Y=2 $X2=4.32
+ $Y2=1.82
r131 20 21 7.04283 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=1.57 $Y=1.99 $X2=1.57
+ $Y2=1.89
r132 13 34 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.44 $Y=0.515
+ $X2=1.44 $Y2=0.385
r133 13 21 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=1.44 $Y=0.515
+ $X2=1.44 $Y2=1.89
r134 4 24 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=4.155
+ $Y=1.845 $X2=4.29 $Y2=2
r135 3 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r136 2 43 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.235 $X2=4.29 $Y2=0.445
r137 1 48 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%Q_N 1 2 9 15 17
r36 17 22 6.49113 $w=4.43e-07 $l=2.2e-07 $layer=LI1_cond $X=9.622 $Y=1.19
+ $X2=9.622 $Y2=1.41
r37 17 20 4.03086 $w=4.43e-07 $l=1.25e-07 $layer=LI1_cond $X=9.622 $Y=1.19
+ $X2=9.622 $Y2=1.065
r38 15 20 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=9.68 $Y=0.395
+ $X2=9.68 $Y2=1.065
r39 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.565 $Y=1.63
+ $X2=9.565 $Y2=2.31
r40 9 22 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=9.565 $Y=1.63
+ $X2=9.565 $Y2=1.41
r41 2 11 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.43
+ $Y=1.485 $X2=9.565 $Y2=2.31
r42 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.43
+ $Y=1.485 $X2=9.565 $Y2=1.63
r43 1 15 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=9.545
+ $Y=0.235 $X2=9.68 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%Q 1 2 7 10
r18 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.39 $Y=1.63
+ $X2=11.39 $Y2=2.31
r19 7 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=11.39 $Y=1.19
+ $X2=11.39 $Y2=1.63
r20 7 10 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=11.39 $Y=1.19
+ $X2=11.39 $Y2=0.395
r21 2 17 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=1.485 $X2=11.39 $Y2=2.31
r22 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=1.485 $X2=11.39 $Y2=1.63
r23 1 10 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=11.245
+ $Y=0.235 $X2=11.39 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 50 55
+ 56 58 59 61 62 63 65 77 81 96 102 103 106 109 112 115
c175 103 0 2.71124e-20 $X=11.73 $Y=0
c176 81 0 1.82232e-19 $X=5.945 $Y=0
r177 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r178 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r179 109 110 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r180 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r181 103 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=10.81 $Y2=0
r182 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r183 100 115 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.932 $Y2=0
r184 100 102 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.73 $Y2=0
r185 99 116 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r186 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r187 96 115 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=10.81 $Y=0
+ $X2=10.932 $Y2=0
r188 96 98 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.81 $Y=0
+ $X2=9.43 $Y2=0
r189 95 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.43
+ $Y2=0
r190 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r191 92 95 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.97 $Y2=0
r192 91 94 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.59 $Y=0 $X2=8.97
+ $Y2=0
r193 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r194 89 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r195 89 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.21 $Y2=0
r196 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r197 86 112 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.142 $Y2=0
r198 86 88 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=7.13
+ $Y2=0
r199 85 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r200 85 110 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=3.45 $Y2=0
r201 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r202 82 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=3.35 $Y2=0
r203 82 84 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=5.75 $Y2=0
r204 81 112 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=6.142 $Y2=0
r205 81 84 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=5.75 $Y2=0
r206 80 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.45 $Y2=0
r207 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r208 77 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.35 $Y2=0
r209 77 79 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=2.99 $Y2=0
r210 76 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r211 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r212 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r213 73 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r214 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r215 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r216 70 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r217 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r218 65 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r219 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r220 63 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r221 63 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r222 61 94 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=8.97 $Y2=0
r223 61 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.095 $Y=0 $X2=9.22
+ $Y2=0
r224 60 98 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=0 $X2=9.43
+ $Y2=0
r225 60 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.345 $Y=0 $X2=9.22
+ $Y2=0
r226 58 88 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.165 $Y=0 $X2=7.13
+ $Y2=0
r227 58 59 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=7.302 $Y2=0
r228 57 91 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.59
+ $Y2=0
r229 57 59 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.302
+ $Y2=0
r230 55 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0
+ $X2=2.07 $Y2=0
r231 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.4
+ $Y2=0
r232 54 79 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=0
+ $X2=2.99 $Y2=0
r233 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.4
+ $Y2=0
r234 50 52 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=10.932 $Y=0.395
+ $X2=10.932 $Y2=0.735
r235 48 115 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.932 $Y=0.085
+ $X2=10.932 $Y2=0
r236 48 50 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=10.932 $Y=0.085
+ $X2=10.932 $Y2=0.395
r237 44 46 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=9.22 $Y=0.395
+ $X2=9.22 $Y2=0.735
r238 42 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0
r239 42 44 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0.395
r240 38 59 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.302 $Y=0.085
+ $X2=7.302 $Y2=0
r241 38 40 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=7.302 $Y=0.085
+ $X2=7.302 $Y2=0.45
r242 34 112 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.142 $Y=0.085
+ $X2=6.142 $Y2=0
r243 34 36 9.77388 $w=3.93e-07 $l=3.35e-07 $layer=LI1_cond $X=6.142 $Y=0.085
+ $X2=6.142 $Y2=0.42
r244 30 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r245 30 32 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.445
r246 26 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=0.085 $X2=2.4
+ $Y2=0
r247 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.4 $Y=0.085
+ $X2=2.4 $Y2=0.38
r248 22 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r249 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r250 7 52 182 $w=1.7e-07 $l=5.91608e-07 $layer=licon1_NDIFF $count=1 $X=10.76
+ $Y=0.235 $X2=10.96 $Y2=0.735
r251 7 50 182 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_NDIFF $count=1 $X=10.76
+ $Y=0.235 $X2=10.96 $Y2=0.395
r252 6 46 182 $w=1.7e-07 $l=5.91608e-07 $layer=licon1_NDIFF $count=1 $X=9.06
+ $Y=0.235 $X2=9.26 $Y2=0.735
r253 6 44 182 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_NDIFF $count=1 $X=9.06
+ $Y=0.235 $X2=9.26 $Y2=0.395
r254 5 40 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.235 $X2=7.285 $Y2=0.45
r255 4 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.035
+ $Y=0.235 $X2=6.175 $Y2=0.42
r256 3 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.35 $Y2=0.445
r257 2 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.38
r258 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__dlygate4sd1_1.pxi.spice
* Created: Thu Aug 27 14:18:38 2020
* 
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A N_A_M1006_g N_A_M1002_g A A N_A_c_68_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_27_47# N_A_27_47#_M1006_s
+ N_A_27_47#_M1002_s N_A_27_47#_M1004_g N_A_27_47#_M1007_g N_A_27_47#_c_106_n
+ N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_102_n N_A_27_47#_c_107_n
+ N_A_27_47#_c_108_n N_A_27_47#_c_103_n N_A_27_47#_c_110_n N_A_27_47#_c_104_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_193_47# N_A_193_47#_M1004_d
+ N_A_193_47#_M1007_d N_A_193_47#_c_170_n N_A_193_47#_M1000_g
+ N_A_193_47#_c_177_n N_A_193_47#_M1005_g N_A_193_47#_c_171_n
+ N_A_193_47#_c_172_n N_A_193_47#_c_173_n N_A_193_47#_c_174_n
+ N_A_193_47#_c_179_n N_A_193_47#_c_175_n N_A_193_47#_c_176_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_299_93# N_A_299_93#_M1000_s
+ N_A_299_93#_M1005_s N_A_299_93#_M1001_g N_A_299_93#_M1003_g
+ N_A_299_93#_c_240_n N_A_299_93#_c_234_n N_A_299_93#_c_241_n
+ N_A_299_93#_c_242_n N_A_299_93#_c_235_n N_A_299_93#_c_244_n
+ N_A_299_93#_c_236_n N_A_299_93#_c_237_n N_A_299_93#_c_238_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_299_93#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%VPWR N_VPWR_M1002_d N_VPWR_M1005_d
+ N_VPWR_c_302_n N_VPWR_c_303_n VPWR N_VPWR_c_304_n N_VPWR_c_305_n
+ N_VPWR_c_306_n N_VPWR_c_301_n N_VPWR_c_308_n N_VPWR_c_309_n VPWR
+ PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%VPWR
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%X N_X_M1001_d N_X_M1003_d N_X_c_344_n
+ N_X_c_347_n N_X_c_345_n X X X PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%X
x_PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%VGND N_VGND_M1006_d N_VGND_M1000_d
+ N_VGND_c_361_n N_VGND_c_362_n VGND N_VGND_c_363_n N_VGND_c_364_n
+ N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n VGND
+ PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%VGND
cc_1 VNB N_A_M1006_g 0.0353079f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.0124662f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_A_c_68_n 0.0311173f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_4 VNB N_A_27_47#_M1004_g 0.0310668f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_5 VNB N_A_27_47#_c_100_n 0.0184796f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.53
cc_6 VNB N_A_27_47#_c_101_n 0.00773781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_102_n 0.00959318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_103_n 0.00446609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_104_n 0.023062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_193_47#_c_170_n 0.0341166f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_11 VNB N_A_193_47#_c_171_n 0.0103069f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_12 VNB N_A_193_47#_c_172_n 5.78778e-19 $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=0.995
cc_13 VNB N_A_193_47#_c_173_n 0.0100937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_193_47#_c_174_n 0.00407265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_193_47#_c_175_n 0.00212837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_193_47#_c_176_n 0.0355467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_299_93#_c_234_n 0.00241192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_299_93#_c_235_n 0.00316925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_299_93#_c_236_n 0.00767985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_299_93#_c_237_n 0.0247766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_93#_c_238_n 0.0194144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_301_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_344_n 0.00558185f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.445
cc_24 VNB N_X_c_345_n 0.0216156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.0166789f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_26 VNB N_VGND_c_361_n 0.00491953f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_27 VNB N_VGND_c_362_n 0.00763671f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_28 VNB N_VGND_c_363_n 0.016294f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.325
cc_29 VNB N_VGND_c_364_n 0.0293903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_365_n 0.0306194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_366_n 0.20966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_367_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_368_n 0.00632006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_M1002_g 0.0597758f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_35 VPB A 0.0175395f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_36 VPB N_A_c_68_n 0.00784995f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_37 VPB N_A_27_47#_M1007_g 0.0515962f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_38 VPB N_A_27_47#_c_106_n 0.0187961f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.325
cc_39 VPB N_A_27_47#_c_107_n 0.00899275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_108_n 0.0123133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_103_n 6.80746e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_110_n 0.00337745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_104_n 0.00570466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_193_47#_c_177_n 0.0562899f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.445
cc_45 VPB N_A_193_47#_c_172_n 0.0180524f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=0.995
cc_46 VPB N_A_193_47#_c_179_n 0.0042109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_193_47#_c_176_n 0.0111291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_299_93#_M1003_g 0.0225543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_299_93#_c_240_n 0.00825106f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=0.995
cc_50 VPB N_A_299_93#_c_241_n 0.00123449f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.53
cc_51 VPB N_A_299_93#_c_242_n 0.00310093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_299_93#_c_235_n 2.01181e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_299_93#_c_244_n 0.00259665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_299_93#_c_237_n 0.00668369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_302_n 0.00491953f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_56 VPB N_VPWR_c_303_n 4.89488e-19 $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_57 VPB N_VPWR_c_304_n 0.0161999f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.325
cc_58 VPB N_VPWR_c_305_n 0.0291468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_306_n 0.0289002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_301_n 0.0732586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_308_n 0.00406576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_309_n 0.00476819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_X_c_347_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_345_n 0.00881722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB X 0.0322452f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_66 N_A_M1006_g N_A_27_47#_M1004_g 0.0256873f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_A_27_47#_M1007_g 0.0442697f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_68 A N_A_27_47#_M1007_g 8.69858e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_M1002_g N_A_27_47#_c_106_n 0.00375513f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_70 N_A_M1006_g N_A_27_47#_c_100_n 0.00374445f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1006_g N_A_27_47#_c_101_n 0.0134647f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_101_n 0.0131329f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A_c_68_n N_A_27_47#_c_101_n 3.58319e-19 $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_102_n 0.0252593f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_68_n N_A_27_47#_c_102_n 0.00511105f $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1002_g N_A_27_47#_c_107_n 0.0157992f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_77 A N_A_27_47#_c_107_n 0.0134407f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_108_n 0.0271506f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_c_68_n N_A_27_47#_c_108_n 8.59854e-19 $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_M1006_g N_A_27_47#_c_103_n 0.00355976f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_81 A N_A_27_47#_c_103_n 0.0227687f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_c_68_n N_A_27_47#_c_103_n 8.28474e-19 $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_A_27_47#_c_110_n 0.00432253f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_84 A N_A_27_47#_c_110_n 0.0236108f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_85 A N_A_27_47#_c_104_n 8.79072e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_68_n N_A_27_47#_c_104_n 0.0212951f $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VPWR_c_302_n 0.00300333f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_88 N_A_M1002_g N_VPWR_c_304_n 0.00436487f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_89 N_A_M1002_g N_VPWR_c_301_n 0.00681164f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_90 N_A_M1006_g N_VGND_c_361_n 0.00300333f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1006_g N_VGND_c_363_n 0.00436487f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_VGND_c_366_n 0.00681164f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1004_g N_A_193_47#_c_171_n 0.0107264f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_103_n N_A_193_47#_c_171_n 0.0217066f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_104_n N_A_193_47#_c_171_n 6.81659e-19 $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_M1007_g N_A_193_47#_c_172_n 0.01861f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_107_n N_A_193_47#_c_172_n 0.0129484f $X=0.725 $Y=1.895 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_103_n N_A_193_47#_c_172_n 0.00366575f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_110_n N_A_193_47#_c_172_n 0.0242721f $X=0.81 $Y=1.785 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_104_n N_A_193_47#_c_172_n 4.25141e-19 $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_M1004_g N_A_193_47#_c_174_n 0.00396006f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_103_n N_A_193_47#_c_174_n 0.00125522f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_104_n N_A_193_47#_c_174_n 7.21452e-19 $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_M1007_g N_A_193_47#_c_179_n 0.00463087f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_103_n N_A_193_47#_c_175_n 0.0166561f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_104_n N_A_193_47#_c_175_n 0.00189838f $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_104_n N_A_193_47#_c_176_n 0.00707105f $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_M1007_g N_VPWR_c_302_n 0.0027531f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_107_n N_VPWR_c_302_n 0.0149018f $X=0.725 $Y=1.895 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_c_106_n N_VPWR_c_304_n 0.0192429f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_107_n N_VPWR_c_304_n 0.00238773f $X=0.725 $Y=1.895 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_M1007_g N_VPWR_c_305_n 0.00460398f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_107_n N_VPWR_c_305_n 0.00206479f $X=0.725 $Y=1.895 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_M1002_s N_VPWR_c_301_n 0.00216553f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1007_g N_VPWR_c_301_n 0.00832113f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_106_n N_VPWR_c_301_n 0.0112839f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_107_n N_VPWR_c_301_n 0.00787286f $X=0.725 $Y=1.895 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_M1004_g N_VGND_c_361_n 0.0027531f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_101_n N_VGND_c_361_n 0.0115001f $X=0.725 $Y=0.8 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_103_n N_VGND_c_361_n 0.00316025f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_100_n N_VGND_c_363_n 0.0184302f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_101_n N_VGND_c_363_n 0.00234724f $X=0.725 $Y=0.8 $X2=0 $Y2=0
cc_123 N_A_27_47#_M1004_g N_VGND_c_364_n 0.00460398f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_103_n N_VGND_c_364_n 0.00206479f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1006_s N_VGND_c_366_n 0.00216553f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1004_g N_VGND_c_366_n 0.00832113f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_100_n N_VGND_c_366_n 0.010877f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_101_n N_VGND_c_366_n 0.00440284f $X=0.725 $Y=0.8 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_103_n N_VGND_c_366_n 0.00341021f $X=0.81 $Y=1.325 $X2=0
+ $Y2=0
cc_130 N_A_193_47#_c_177_n N_A_299_93#_M1003_g 0.032378f $X=1.84 $Y=1.325 $X2=0
+ $Y2=0
cc_131 N_A_193_47#_c_177_n N_A_299_93#_c_240_n 0.00858357f $X=1.84 $Y=1.325
+ $X2=0 $Y2=0
cc_132 N_A_193_47#_c_172_n N_A_299_93#_c_240_n 0.0294508f $X=1.235 $Y=2.175
+ $X2=0 $Y2=0
cc_133 N_A_193_47#_c_179_n N_A_299_93#_c_240_n 0.0189672f $X=1.235 $Y=2.32 $X2=0
+ $Y2=0
cc_134 N_A_193_47#_c_170_n N_A_299_93#_c_234_n 0.0109081f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_135 N_A_193_47#_c_173_n N_A_299_93#_c_234_n 0.0110006f $X=1.63 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_193_47#_c_176_n N_A_299_93#_c_234_n 0.0011681f $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_193_47#_c_177_n N_A_299_93#_c_241_n 0.016386f $X=1.84 $Y=1.325 $X2=0
+ $Y2=0
cc_138 N_A_193_47#_c_173_n N_A_299_93#_c_241_n 0.00704394f $X=1.63 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_193_47#_c_176_n N_A_299_93#_c_241_n 9.46666e-19 $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_193_47#_c_172_n N_A_299_93#_c_242_n 0.0129579f $X=1.235 $Y=2.175
+ $X2=0 $Y2=0
cc_141 N_A_193_47#_c_173_n N_A_299_93#_c_242_n 0.0120363f $X=1.63 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_193_47#_c_176_n N_A_299_93#_c_242_n 0.00516661f $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_193_47#_c_170_n N_A_299_93#_c_235_n 0.00192736f $X=1.83 $Y=0.995
+ $X2=0 $Y2=0
cc_144 N_A_193_47#_c_173_n N_A_299_93#_c_235_n 0.0165368f $X=1.63 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_193_47#_c_176_n N_A_299_93#_c_235_n 0.00436781f $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_193_47#_c_177_n N_A_299_93#_c_244_n 0.00534765f $X=1.84 $Y=1.325
+ $X2=0 $Y2=0
cc_147 N_A_193_47#_c_170_n N_A_299_93#_c_236_n 0.0064807f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_193_47#_c_171_n N_A_299_93#_c_236_n 0.0257188f $X=1.235 $Y=1.075
+ $X2=0 $Y2=0
cc_149 N_A_193_47#_c_173_n N_A_299_93#_c_236_n 0.0182754f $X=1.63 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_193_47#_c_174_n N_A_299_93#_c_236_n 0.0213903f $X=1.235 $Y=0.4 $X2=0
+ $Y2=0
cc_151 N_A_193_47#_c_176_n N_A_299_93#_c_236_n 0.00575864f $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_193_47#_c_173_n N_A_299_93#_c_237_n 2.02753e-19 $X=1.63 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A_193_47#_c_176_n N_A_299_93#_c_237_n 0.0210524f $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_193_47#_c_170_n N_A_299_93#_c_238_n 0.0242005f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_A_193_47#_c_177_n N_VPWR_c_303_n 0.015266f $X=1.84 $Y=1.325 $X2=0 $Y2=0
cc_156 N_A_193_47#_c_179_n N_VPWR_c_303_n 0.00107336f $X=1.235 $Y=2.32 $X2=0
+ $Y2=0
cc_157 N_A_193_47#_c_177_n N_VPWR_c_305_n 0.00564095f $X=1.84 $Y=1.325 $X2=0
+ $Y2=0
cc_158 N_A_193_47#_c_179_n N_VPWR_c_305_n 0.0235612f $X=1.235 $Y=2.32 $X2=0
+ $Y2=0
cc_159 N_A_193_47#_M1007_d N_VPWR_c_301_n 0.00209344f $X=0.965 $Y=2.065 $X2=0
+ $Y2=0
cc_160 N_A_193_47#_c_177_n N_VPWR_c_301_n 0.0108804f $X=1.84 $Y=1.325 $X2=0
+ $Y2=0
cc_161 N_A_193_47#_c_179_n N_VPWR_c_301_n 0.0142974f $X=1.235 $Y=2.32 $X2=0
+ $Y2=0
cc_162 N_A_193_47#_c_170_n N_VGND_c_362_n 0.00621929f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_193_47#_c_170_n N_VGND_c_364_n 0.00439206f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_193_47#_c_174_n N_VGND_c_364_n 0.0235928f $X=1.235 $Y=0.4 $X2=0 $Y2=0
cc_165 N_A_193_47#_M1004_d N_VGND_c_366_n 0.00209344f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_166 N_A_193_47#_c_170_n N_VGND_c_366_n 0.00745018f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_193_47#_c_174_n N_VGND_c_366_n 0.0143018f $X=1.235 $Y=0.4 $X2=0 $Y2=0
cc_168 N_A_299_93#_c_241_n N_VPWR_M1005_d 0.00463289f $X=2.07 $Y=1.66 $X2=0
+ $Y2=0
cc_169 N_A_299_93#_c_244_n N_VPWR_M1005_d 0.00135845f $X=2.155 $Y=1.575 $X2=0
+ $Y2=0
cc_170 N_A_299_93#_M1003_g N_VPWR_c_303_n 0.0165601f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_299_93#_c_240_n N_VPWR_c_303_n 0.031518f $X=1.627 $Y=1.745 $X2=0
+ $Y2=0
cc_172 N_A_299_93#_c_241_n N_VPWR_c_303_n 0.0183424f $X=2.07 $Y=1.66 $X2=0 $Y2=0
cc_173 N_A_299_93#_c_235_n N_VPWR_c_303_n 8.12398e-19 $X=2.155 $Y=1.325 $X2=0
+ $Y2=0
cc_174 N_A_299_93#_c_237_n N_VPWR_c_303_n 2.5512e-19 $X=2.275 $Y=1.16 $X2=0
+ $Y2=0
cc_175 N_A_299_93#_c_240_n N_VPWR_c_305_n 0.0130885f $X=1.627 $Y=1.745 $X2=0
+ $Y2=0
cc_176 N_A_299_93#_M1003_g N_VPWR_c_306_n 0.0046653f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_299_93#_M1003_g N_VPWR_c_301_n 0.00934473f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_299_93#_c_240_n N_VPWR_c_301_n 0.00844061f $X=1.627 $Y=1.745 $X2=0
+ $Y2=0
cc_179 N_A_299_93#_M1003_g N_X_c_345_n 0.0035877f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_299_93#_c_235_n N_X_c_345_n 0.0331607f $X=2.155 $Y=1.325 $X2=0 $Y2=0
cc_181 N_A_299_93#_c_244_n N_X_c_345_n 0.00846694f $X=2.155 $Y=1.575 $X2=0 $Y2=0
cc_182 N_A_299_93#_c_237_n N_X_c_345_n 0.00797237f $X=2.275 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_299_93#_c_238_n N_X_c_345_n 0.00358577f $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_299_93#_c_234_n N_VGND_M1000_d 0.00111119f $X=2.07 $Y=0.82 $X2=0
+ $Y2=0
cc_185 N_A_299_93#_c_235_n N_VGND_M1000_d 0.00165553f $X=2.155 $Y=1.325 $X2=0
+ $Y2=0
cc_186 N_A_299_93#_c_234_n N_VGND_c_362_n 0.00844092f $X=2.07 $Y=0.82 $X2=0
+ $Y2=0
cc_187 N_A_299_93#_c_235_n N_VGND_c_362_n 0.00979705f $X=2.155 $Y=1.325 $X2=0
+ $Y2=0
cc_188 N_A_299_93#_c_236_n N_VGND_c_362_n 0.0169004f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_299_93#_c_237_n N_VGND_c_362_n 3.34849e-19 $X=2.275 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_299_93#_c_238_n N_VGND_c_362_n 0.00323779f $X=2.29 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_299_93#_c_234_n N_VGND_c_364_n 0.002104f $X=2.07 $Y=0.82 $X2=0 $Y2=0
cc_192 N_A_299_93#_c_236_n N_VGND_c_364_n 0.0159334f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_299_93#_c_238_n N_VGND_c_365_n 0.00583607f $X=2.29 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_299_93#_c_234_n N_VGND_c_366_n 0.00432679f $X=2.07 $Y=0.82 $X2=0
+ $Y2=0
cc_195 N_A_299_93#_c_235_n N_VGND_c_366_n 7.18353e-19 $X=2.155 $Y=1.325 $X2=0
+ $Y2=0
cc_196 N_A_299_93#_c_236_n N_VGND_c_366_n 0.00857794f $X=1.62 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_A_299_93#_c_238_n N_VGND_c_366_n 0.0120361f $X=2.29 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_301_n N_X_M1003_d 0.00387172f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_306_n X 0.018001f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_c_301_n X 0.00993603f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_201 X N_VGND_c_365_n 0.0189908f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_202 N_X_M1001_d N_VGND_c_366_n 0.00283025f $X=2.39 $Y=0.235 $X2=0 $Y2=0
cc_203 X N_VGND_c_366_n 0.0110704f $X=2.465 $Y=0.425 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o31ai_2.pxi.spice
* Created: Thu Aug 27 14:40:27 2020
* 
x_PM_SKY130_FD_SC_HD__O31AI_2%A1 N_A1_M1003_g N_A1_M1001_g N_A1_M1005_g
+ N_A1_M1013_g A1 A1 A1 N_A1_c_79_n PM_SKY130_FD_SC_HD__O31AI_2%A1
x_PM_SKY130_FD_SC_HD__O31AI_2%A2 N_A2_M1002_g N_A2_M1006_g N_A2_M1008_g
+ N_A2_M1009_g A2 A2 N_A2_c_131_n PM_SKY130_FD_SC_HD__O31AI_2%A2
x_PM_SKY130_FD_SC_HD__O31AI_2%A3 N_A3_M1014_g N_A3_M1007_g N_A3_M1015_g
+ N_A3_M1011_g A3 A3 N_A3_c_177_n PM_SKY130_FD_SC_HD__O31AI_2%A3
x_PM_SKY130_FD_SC_HD__O31AI_2%B1 N_B1_c_224_n N_B1_M1004_g N_B1_M1000_g
+ N_B1_c_225_n N_B1_c_226_n N_B1_M1010_g N_B1_M1012_g N_B1_c_227_n B1 B1
+ N_B1_c_229_n PM_SKY130_FD_SC_HD__O31AI_2%B1
x_PM_SKY130_FD_SC_HD__O31AI_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1013_s
+ N_A_27_297#_M1008_d N_A_27_297#_c_273_n N_A_27_297#_c_279_n
+ N_A_27_297#_c_274_n N_A_27_297#_c_286_n N_A_27_297#_c_275_n
+ N_A_27_297#_c_276_n N_A_27_297#_c_288_n PM_SKY130_FD_SC_HD__O31AI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__O31AI_2%VPWR N_VPWR_M1001_d N_VPWR_M1000_d N_VPWR_c_318_n
+ N_VPWR_c_319_n VPWR N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_317_n
+ N_VPWR_c_323_n N_VPWR_c_324_n VPWR PM_SKY130_FD_SC_HD__O31AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O31AI_2%A_281_297# N_A_281_297#_M1006_s
+ N_A_281_297#_M1007_s N_A_281_297#_c_374_n N_A_281_297#_c_370_n
+ N_A_281_297#_c_382_n N_A_281_297#_c_387_p
+ PM_SKY130_FD_SC_HD__O31AI_2%A_281_297#
x_PM_SKY130_FD_SC_HD__O31AI_2%Y N_Y_M1004_s N_Y_M1007_d N_Y_M1011_d N_Y_M1012_s
+ N_Y_c_395_n N_Y_c_390_n N_Y_c_402_n Y Y Y Y Y Y N_Y_c_391_n N_Y_c_389_n
+ N_Y_c_393_n N_Y_c_394_n PM_SKY130_FD_SC_HD__O31AI_2%Y
x_PM_SKY130_FD_SC_HD__O31AI_2%A_27_47# N_A_27_47#_M1003_d N_A_27_47#_M1005_d
+ N_A_27_47#_M1009_s N_A_27_47#_M1015_d N_A_27_47#_M1010_d N_A_27_47#_c_445_n
+ N_A_27_47#_c_453_n N_A_27_47#_c_446_n N_A_27_47#_c_460_n N_A_27_47#_c_465_n
+ N_A_27_47#_c_503_p N_A_27_47#_c_447_n N_A_27_47#_c_474_n N_A_27_47#_c_475_n
+ N_A_27_47#_c_483_n N_A_27_47#_c_448_n N_A_27_47#_c_449_n N_A_27_47#_c_450_n
+ PM_SKY130_FD_SC_HD__O31AI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O31AI_2%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_M1014_s
+ N_VGND_c_526_n N_VGND_c_527_n VGND N_VGND_c_528_n N_VGND_c_529_n
+ N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n N_VGND_c_534_n
+ VGND PM_SKY130_FD_SC_HD__O31AI_2%VGND
cc_1 VNB N_A1_M1003_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_2 VNB N_A1_M1001_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_3 VNB N_A1_M1005_g 0.0177503f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_4 VNB N_A1_M1013_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_5 VNB A1 0.0170331f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_6 VNB N_A1_c_79_n 0.04127f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_7 VNB N_A2_M1002_g 0.0206889f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_8 VNB N_A2_M1006_g 4.60057e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_9 VNB N_A2_M1008_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_10 VNB N_A2_M1009_g 0.0218491f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_11 VNB A2 0.00221811f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_12 VNB N_A2_c_131_n 0.0588816f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_13 VNB N_A3_M1014_g 0.019522f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_14 VNB N_A3_M1007_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_15 VNB N_A3_M1015_g 0.0185906f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_16 VNB N_A3_M1011_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_17 VNB A3 0.00524541f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_18 VNB N_A3_c_177_n 0.0376298f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_19 VNB N_B1_c_224_n 0.0172537f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.025
cc_20 VNB N_B1_c_225_n 0.0187688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B1_c_226_n 0.0201789f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_22 VNB N_B1_c_227_n 0.0109834f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_23 VNB B1 0.022182f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_24 VNB N_B1_c_229_n 0.0340798f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_25 VNB N_VPWR_c_317_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_26 VNB N_Y_c_389_n 0.00170777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_445_n 0.0183269f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_28 VNB N_A_27_47#_c_446_n 0.00956771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_447_n 0.00257277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_448_n 0.001463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_449_n 0.00647876f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.19
cc_32 VNB N_A_27_47#_c_450_n 0.0147282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_526_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_34 VNB N_VGND_c_527_n 0.00275589f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_35 VNB N_VGND_c_528_n 0.0166708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_529_n 0.016968f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_37 VNB N_VGND_c_530_n 0.0392591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_531_n 0.238151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_532_n 0.0208501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_533_n 0.0158606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_534_n 0.00507255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_A1_M1001_g 0.0272353f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_43 VPB N_A1_M1013_g 0.0197334f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_44 VPB A1 0.00880193f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_45 VPB N_A2_M1006_g 0.0199119f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_46 VPB N_A2_M1008_g 0.0272353f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_47 VPB A2 0.00892571f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_48 VPB N_A3_M1007_g 0.0272353f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_49 VPB N_A3_M1011_g 0.019707f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_50 VPB A3 0.00508588f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_51 VPB N_B1_M1000_g 0.0200645f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_52 VPB N_B1_c_225_n 0.00682721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_B1_M1012_g 0.0272092f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_54 VPB N_B1_c_227_n 6.88461e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_55 VPB B1 0.00391252f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_56 VPB N_B1_c_229_n 0.0109753f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_57 VPB N_A_27_297#_c_273_n 0.0316657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_297#_c_274_n 0.00762919f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_59 VPB N_A_27_297#_c_275_n 0.00183174f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_60 VPB N_A_27_297#_c_276_n 0.00456453f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_61 VPB N_VPWR_c_318_n 0.0046277f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_62 VPB N_VPWR_c_319_n 0.00557203f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_63 VPB N_VPWR_c_320_n 0.0704177f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_64 VPB N_VPWR_c_321_n 0.0178976f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_65 VPB N_VPWR_c_317_n 0.0467765f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_66 VPB N_VPWR_c_323_n 0.0214916f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_67 VPB N_VPWR_c_324_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.19
cc_68 VPB N_A_281_297#_c_370_n 0.0114154f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_69 VPB N_Y_c_390_n 0.00177653f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_70 VPB N_Y_c_391_n 0.00405913f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.19
cc_71 VPB N_Y_c_389_n 0.00312037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_Y_c_393_n 0.00821962f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_Y_c_394_n 0.0334076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_A1_M1005_g N_A2_M1002_g 0.0146046f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_75 N_A1_M1013_g N_A2_M1006_g 0.0146046f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_76 A1 A2 0.0240198f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_77 A1 N_A2_c_131_n 0.00276376f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A1_c_79_n N_A2_c_131_n 0.0146046f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A1_M1001_g N_A_27_297#_c_273_n 0.00975139f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A1_M1013_g N_A_27_297#_c_273_n 6.18904e-19 $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A1_M1001_g N_A_27_297#_c_279_n 0.0107189f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A1_M1013_g N_A_27_297#_c_279_n 0.0107189f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_83 A1 N_A_27_297#_c_279_n 0.033369f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A1_c_79_n N_A_27_297#_c_279_n 5.85705e-19 $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A1_M1001_g N_A_27_297#_c_274_n 8.84614e-19 $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_86 A1 N_A_27_297#_c_274_n 0.0276077f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A1_c_79_n N_A_27_297#_c_274_n 5.68867e-19 $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A1_M1001_g N_A_27_297#_c_286_n 6.1949e-19 $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A1_M1013_g N_A_27_297#_c_286_n 0.00975139f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A1_M1013_g N_A_27_297#_c_288_n 8.84614e-19 $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_91 A1 N_A_27_297#_c_288_n 0.0196623f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A1_M1001_g N_VPWR_c_318_n 0.00268723f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A1_M1013_g N_VPWR_c_318_n 0.00268723f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A1_M1013_g N_VPWR_c_320_n 0.00541359f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A1_M1001_g N_VPWR_c_317_n 0.0104744f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A1_M1013_g N_VPWR_c_317_n 0.00952874f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A1_M1001_g N_VPWR_c_323_n 0.00541359f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A1_M1003_g N_A_27_47#_c_445_n 0.00620543f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_99 N_A1_M1005_g N_A_27_47#_c_445_n 5.18879e-19 $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A1_M1003_g N_A_27_47#_c_453_n 0.00844123f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_101 N_A1_M1005_g N_A_27_47#_c_453_n 0.00844123f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_102 A1 N_A_27_47#_c_453_n 0.0322881f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A1_c_79_n N_A_27_47#_c_453_n 0.0020061f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A1_M1003_g N_A_27_47#_c_446_n 8.68782e-19 $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_105 A1 N_A_27_47#_c_446_n 0.027058f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A1_c_79_n N_A_27_47#_c_446_n 0.00213315f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_M1003_g N_A_27_47#_c_460_n 5.19281e-19 $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A1_M1005_g N_A_27_47#_c_460_n 0.00620543f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A1_M1005_g N_A_27_47#_c_448_n 8.68782e-19 $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_110 A1 N_A_27_47#_c_448_n 0.0195698f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_111 N_A1_M1003_g N_VGND_c_526_n 0.00268723f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A1_M1005_g N_VGND_c_526_n 0.00146448f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A1_M1005_g N_VGND_c_528_n 0.00422241f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_114 N_A1_M1003_g N_VGND_c_531_n 0.00666944f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A1_M1005_g N_VGND_c_531_n 0.00572376f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A1_M1003_g N_VGND_c_532_n 0.00422241f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_117 N_A2_M1009_g N_A3_M1014_g 0.0173521f $X=2.09 $Y=0.56 $X2=0 $Y2=0
cc_118 A2 A3 0.0251062f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_119 N_A2_c_131_n A3 8.83086e-19 $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_120 A2 N_A3_c_177_n 7.21518e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A2_c_131_n N_A3_c_177_n 0.00907257f $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A2_M1006_g N_A_27_297#_c_286_n 0.00973197f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A2_M1008_g N_A_27_297#_c_286_n 7.44598e-19 $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A2_M1006_g N_A_27_297#_c_275_n 0.0123658f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A2_M1008_g N_A_27_297#_c_275_n 0.00965515f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_126 A2 N_A_27_297#_c_275_n 0.0500927f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A2_c_131_n N_A_27_297#_c_275_n 0.00257719f $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_M1006_g N_A_27_297#_c_276_n 5.83663e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A2_M1008_g N_A_27_297#_c_276_n 0.00636413f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A2_M1006_g N_A_27_297#_c_288_n 0.0013142f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A2_M1006_g N_VPWR_c_320_n 0.00541359f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A2_M1008_g N_VPWR_c_320_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A2_M1006_g N_VPWR_c_317_n 0.00972738f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A2_M1008_g N_VPWR_c_317_n 0.00664112f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A2_M1008_g N_A_281_297#_c_370_n 0.012606f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A2_M1002_g N_A_27_47#_c_460_n 0.0108215f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_137 N_A2_M1002_g N_A_27_47#_c_465_n 0.0114995f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_138 N_A2_M1009_g N_A_27_47#_c_465_n 0.0114904f $X=2.09 $Y=0.56 $X2=0 $Y2=0
cc_139 A2 N_A_27_47#_c_465_n 0.0509375f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A2_c_131_n N_A_27_47#_c_465_n 0.0107859f $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_M1002_g N_A_27_47#_c_448_n 0.00128201f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A2_M1009_g N_VGND_c_527_n 9.94421e-19 $X=2.09 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A2_M1002_g N_VGND_c_528_n 0.00422241f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A2_M1009_g N_VGND_c_529_n 0.00436487f $X=2.09 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A2_M1002_g N_VGND_c_531_n 0.00638873f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_146 N_A2_M1009_g N_VGND_c_531_n 0.00682101f $X=2.09 $Y=0.56 $X2=0 $Y2=0
cc_147 N_A2_M1002_g N_VGND_c_533_n 0.00205456f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A2_M1009_g N_VGND_c_533_n 0.00345545f $X=2.09 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A3_M1015_g N_B1_c_224_n 0.0143974f $X=3.13 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_150 N_A3_M1011_g N_B1_M1000_g 0.0143974f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_151 A3 N_B1_c_227_n 0.00129971f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A3_c_177_n N_B1_c_227_n 0.0143974f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A3_M1007_g N_VPWR_c_320_n 0.00357877f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A3_M1011_g N_VPWR_c_320_n 0.00541359f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A3_M1007_g N_VPWR_c_317_n 0.00664112f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A3_M1011_g N_VPWR_c_317_n 0.00972738f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A3_M1007_g N_A_281_297#_c_370_n 0.012606f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A3_M1007_g N_Y_c_395_n 0.00878637f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A3_M1011_g N_Y_c_395_n 0.0107189f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_160 A3 N_Y_c_395_n 0.0354434f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A3_c_177_n N_Y_c_395_n 5.85705e-19 $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A3_M1007_g N_Y_c_390_n 8.68782e-19 $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_163 A3 N_Y_c_390_n 0.0205842f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A3_c_177_n N_Y_c_390_n 5.56519e-19 $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A3_M1007_g N_Y_c_402_n 7.45387e-19 $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A3_M1011_g N_Y_c_402_n 0.00983765f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A3_M1007_g N_Y_c_391_n 0.00636413f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A3_M1011_g N_Y_c_391_n 5.83663e-19 $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A3_M1015_g N_Y_c_389_n 2.8218e-19 $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_170 A3 N_Y_c_389_n 0.00931709f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A3_c_177_n N_Y_c_389_n 2.56337e-19 $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A3_M1011_g N_Y_c_393_n 9.43996e-19 $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A3_M1014_g N_A_27_47#_c_447_n 0.0127565f $X=2.63 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A3_M1015_g N_A_27_47#_c_447_n 0.00978016f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_175 A3 N_A_27_47#_c_447_n 0.0444901f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A3_c_177_n N_A_27_47#_c_447_n 0.00418969f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A3_M1015_g N_A_27_47#_c_474_n 0.0020512f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A3_M1014_g N_A_27_47#_c_475_n 5.14406e-19 $X=2.63 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A3_M1015_g N_A_27_47#_c_475_n 0.00468939f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_180 A3 N_A_27_47#_c_449_n 0.00945682f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A3_M1014_g N_VGND_c_527_n 0.00881296f $X=2.63 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A3_M1015_g N_VGND_c_527_n 0.00459089f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A3_M1014_g N_VGND_c_529_n 0.00348405f $X=2.63 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A3_M1015_g N_VGND_c_530_n 0.00420723f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A3_M1014_g N_VGND_c_531_n 0.00445075f $X=2.63 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A3_M1015_g N_VGND_c_531_n 0.00598199f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_187 N_B1_M1000_g N_VPWR_c_319_n 0.00672121f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B1_M1012_g N_VPWR_c_319_n 0.00329913f $X=4.09 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B1_M1000_g N_VPWR_c_320_n 0.00541359f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B1_M1012_g N_VPWR_c_321_n 0.00585385f $X=4.09 $Y=1.985 $X2=0 $Y2=0
cc_191 N_B1_M1000_g N_VPWR_c_317_n 0.0099008f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B1_M1012_g N_VPWR_c_317_n 0.0118266f $X=4.09 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B1_M1000_g N_Y_c_402_n 0.0105083f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B1_M1012_g N_Y_c_402_n 6.50333e-19 $X=4.09 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_c_224_n N_Y_c_389_n 0.00476543f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B1_M1000_g N_Y_c_389_n 0.00461631f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_c_225_n N_Y_c_389_n 0.0284534f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B1_c_226_n N_Y_c_389_n 0.00105744f $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_M1012_g N_Y_c_389_n 0.00486325f $X=4.09 $Y=1.985 $X2=0 $Y2=0
cc_200 B1 N_Y_c_389_n 0.0339117f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_201 N_B1_M1000_g N_Y_c_393_n 0.0164958f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B1_c_225_n N_Y_c_393_n 0.00102504f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B1_M1012_g N_Y_c_393_n 0.0197254f $X=4.09 $Y=1.985 $X2=0 $Y2=0
cc_204 B1 N_Y_c_393_n 0.024713f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_205 N_B1_c_229_n N_Y_c_393_n 0.00214841f $X=4.36 $Y=1.16 $X2=0 $Y2=0
cc_206 B1 N_A_27_47#_M1010_d 0.00286201f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_207 N_B1_c_224_n N_A_27_47#_c_447_n 0.00266006f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B1_c_224_n N_A_27_47#_c_474_n 7.12665e-19 $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B1_c_224_n N_A_27_47#_c_475_n 0.00473198f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B1_c_226_n N_A_27_47#_c_475_n 4.93308e-19 $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B1_c_224_n N_A_27_47#_c_483_n 0.0106974f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_225_n N_A_27_47#_c_483_n 6.46342e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B1_c_226_n N_A_27_47#_c_483_n 0.0128241f $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_214 B1 N_A_27_47#_c_450_n 0.0240906f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_215 N_B1_c_229_n N_A_27_47#_c_450_n 0.00129995f $X=4.36 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B1_c_224_n N_VGND_c_530_n 0.00357835f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_226_n N_VGND_c_530_n 0.00357877f $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_224_n N_VGND_c_531_n 0.00554875f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_226_n N_VGND_c_531_n 0.00651204f $X=4.09 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_27_297#_c_279_n N_VPWR_M1001_d 0.00312283f $X=0.955 $Y=1.58 $X2=-0.19
+ $Y2=1.305
cc_221 N_A_27_297#_c_279_n N_VPWR_c_318_n 0.0126919f $X=0.955 $Y=1.58 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_c_286_n N_VPWR_c_320_n 0.0189039f $X=1.12 $Y=1.68 $X2=0 $Y2=0
cc_223 N_A_27_297#_M1001_s N_VPWR_c_317_n 0.00225715f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_224 N_A_27_297#_M1013_s N_VPWR_c_317_n 0.00215201f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_A_27_297#_M1008_d N_VPWR_c_317_n 0.00210147f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_226 N_A_27_297#_c_273_n N_VPWR_c_317_n 0.0133896f $X=0.28 $Y=1.68 $X2=0 $Y2=0
cc_227 N_A_27_297#_c_286_n N_VPWR_c_317_n 0.0122217f $X=1.12 $Y=1.68 $X2=0 $Y2=0
cc_228 N_A_27_297#_c_273_n N_VPWR_c_323_n 0.022803f $X=0.28 $Y=1.68 $X2=0 $Y2=0
cc_229 N_A_27_297#_c_275_n N_A_281_297#_M1006_s 0.00312283f $X=1.795 $Y=1.58
+ $X2=-0.19 $Y2=1.305
cc_230 N_A_27_297#_c_275_n N_A_281_297#_c_374_n 0.0126131f $X=1.795 $Y=1.58
+ $X2=0 $Y2=0
cc_231 N_A_27_297#_M1008_d N_A_281_297#_c_370_n 0.00480843f $X=1.825 $Y=1.485
+ $X2=0 $Y2=0
cc_232 N_A_27_297#_c_275_n N_A_281_297#_c_370_n 0.00271653f $X=1.795 $Y=1.58
+ $X2=0 $Y2=0
cc_233 N_A_27_297#_c_276_n N_A_281_297#_c_370_n 0.0204623f $X=1.96 $Y=1.68 $X2=0
+ $Y2=0
cc_234 N_A_27_297#_c_275_n N_Y_c_390_n 0.0137126f $X=1.795 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A_27_297#_c_276_n N_Y_c_391_n 0.0329599f $X=1.96 $Y=1.68 $X2=0 $Y2=0
cc_236 N_A_27_297#_c_275_n N_A_27_47#_c_465_n 0.00279929f $X=1.795 $Y=1.58 $X2=0
+ $Y2=0
cc_237 N_A_27_297#_c_288_n N_A_27_47#_c_448_n 8.4176e-19 $X=1.12 $Y=1.58 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_317_n N_A_281_297#_M1006_s 0.0039039f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_239 N_VPWR_c_317_n N_A_281_297#_M1007_s 0.0039039f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_320_n N_A_281_297#_c_370_n 0.0818081f $X=3.675 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_317_n N_A_281_297#_c_370_n 0.0502236f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_320_n N_A_281_297#_c_382_n 0.0114055f $X=3.675 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_317_n N_A_281_297#_c_382_n 0.00652883f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_317_n N_Y_M1007_d 0.00226545f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_245 N_VPWR_c_317_n N_Y_M1011_d 0.00215201f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_246 N_VPWR_c_317_n N_Y_M1012_s 0.00248309f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_247 N_VPWR_c_320_n N_Y_c_402_n 0.0189039f $X=3.675 $Y=2.72 $X2=0 $Y2=0
cc_248 N_VPWR_c_317_n N_Y_c_402_n 0.0122217f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_M1000_d N_Y_c_389_n 8.16106e-19 $X=3.625 $Y=1.485 $X2=0 $Y2=0
cc_250 N_VPWR_M1000_d N_Y_c_393_n 0.00390073f $X=3.625 $Y=1.485 $X2=0 $Y2=0
cc_251 N_VPWR_c_319_n N_Y_c_393_n 0.022455f $X=3.84 $Y=2.02 $X2=0 $Y2=0
cc_252 N_VPWR_c_321_n N_Y_c_394_n 0.0222881f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_253 N_VPWR_c_317_n N_Y_c_394_n 0.013017f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_254 N_A_281_297#_c_370_n N_Y_M1007_d 0.00539485f $X=2.835 $Y=2.38 $X2=0 $Y2=0
cc_255 N_A_281_297#_M1007_s N_Y_c_395_n 0.00312283f $X=2.785 $Y=1.485 $X2=0
+ $Y2=0
cc_256 N_A_281_297#_c_370_n N_Y_c_395_n 0.00271653f $X=2.835 $Y=2.38 $X2=0 $Y2=0
cc_257 N_A_281_297#_c_387_p N_Y_c_395_n 0.0126131f $X=2.92 $Y=2.135 $X2=0 $Y2=0
cc_258 N_A_281_297#_c_370_n N_Y_c_391_n 0.0204048f $X=2.835 $Y=2.38 $X2=0 $Y2=0
cc_259 N_Y_c_393_n N_A_27_47#_c_447_n 0.00559305f $X=4.345 $Y=1.665 $X2=0 $Y2=0
cc_260 N_Y_M1004_s N_A_27_47#_c_483_n 0.00559824f $X=3.625 $Y=0.235 $X2=0 $Y2=0
cc_261 N_Y_c_389_n N_A_27_47#_c_483_n 0.0210299f $X=3.84 $Y=0.755 $X2=0 $Y2=0
cc_262 N_Y_c_390_n N_A_27_47#_c_449_n 0.0019114f $X=2.665 $Y=1.58 $X2=0 $Y2=0
cc_263 N_Y_M1004_s N_VGND_c_531_n 0.00313203f $X=3.625 $Y=0.235 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_453_n N_VGND_M1003_s 0.00306532f $X=0.955 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_265 N_A_27_47#_c_465_n N_VGND_M1002_d 0.0116198f $X=2.175 $Y=0.8 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_447_n N_VGND_M1014_s 0.0045572f $X=3.175 $Y=0.8 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_453_n N_VGND_c_526_n 0.012179f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_447_n N_VGND_c_527_n 0.0205027f $X=3.175 $Y=0.8 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_453_n N_VGND_c_528_n 0.0020257f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_460_n N_VGND_c_528_n 0.0188215f $X=1.12 $Y=0.36 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_465_n N_VGND_c_528_n 0.00203365f $X=2.175 $Y=0.8 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_465_n N_VGND_c_529_n 0.00252361f $X=2.175 $Y=0.8 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_503_p N_VGND_c_529_n 0.0211452f $X=2.34 $Y=0.36 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_447_n N_VGND_c_529_n 0.00203142f $X=3.175 $Y=0.8 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_447_n N_VGND_c_530_n 0.0020257f $X=3.175 $Y=0.8 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_474_n N_VGND_c_530_n 0.0189571f $X=3.34 $Y=0.425 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_483_n N_VGND_c_530_n 0.0384264f $X=4.175 $Y=0.34 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_450_n N_VGND_c_530_n 0.021237f $X=4.345 $Y=0.34 $X2=0 $Y2=0
cc_279 N_A_27_47#_M1003_d N_VGND_c_531_n 0.00225715f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1005_d N_VGND_c_531_n 0.00215201f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_M1009_s N_VGND_c_531_n 0.0033921f $X=2.165 $Y=0.235 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1015_d N_VGND_c_531_n 0.00215201f $X=3.205 $Y=0.235 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1010_d N_VGND_c_531_n 0.00208517f $X=4.165 $Y=0.235 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_445_n N_VGND_c_531_n 0.0133626f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_453_n N_VGND_c_531_n 0.00841425f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_460_n N_VGND_c_531_n 0.0121968f $X=1.12 $Y=0.36 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_465_n N_VGND_c_531_n 0.0105952f $X=2.175 $Y=0.8 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_503_p N_VGND_c_531_n 0.0126066f $X=2.34 $Y=0.36 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_447_n N_VGND_c_531_n 0.0091336f $X=3.175 $Y=0.8 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_474_n N_VGND_c_531_n 0.0122645f $X=3.34 $Y=0.425 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_483_n N_VGND_c_531_n 0.0236533f $X=4.175 $Y=0.34 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_450_n N_VGND_c_531_n 0.0127852f $X=4.345 $Y=0.34 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_445_n N_VGND_c_532_n 0.0226868f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_453_n N_VGND_c_532_n 0.0020257f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_465_n N_VGND_c_533_n 0.0387231f $X=2.175 $Y=0.8 $X2=0 $Y2=0

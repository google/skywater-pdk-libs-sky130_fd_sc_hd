* File: sky130_fd_sc_hd__dfrtp_1.pxi.spice
* Created: Thu Aug 27 14:14:41 2020
* 
x_PM_SKY130_FD_SC_HD__DFRTP_1%CLK N_CLK_c_193_n N_CLK_c_197_n N_CLK_c_194_n
+ N_CLK_M1023_g N_CLK_c_198_n N_CLK_M1011_g N_CLK_c_199_n CLK CLK
+ PM_SKY130_FD_SC_HD__DFRTP_1%CLK
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_27_47# N_A_27_47#_M1023_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1012_g N_A_27_47#_M1000_g N_A_27_47#_M1008_g N_A_27_47#_c_235_n
+ N_A_27_47#_c_236_n N_A_27_47#_c_237_n N_A_27_47#_M1006_g N_A_27_47#_c_238_n
+ N_A_27_47#_M1021_g N_A_27_47#_M1018_g N_A_27_47#_c_240_n N_A_27_47#_c_241_n
+ N_A_27_47#_c_242_n N_A_27_47#_c_259_n N_A_27_47#_c_260_n N_A_27_47#_c_243_n
+ N_A_27_47#_c_244_n N_A_27_47#_c_245_n N_A_27_47#_c_246_n N_A_27_47#_c_247_n
+ N_A_27_47#_c_248_n N_A_27_47#_c_249_n N_A_27_47#_c_250_n N_A_27_47#_c_251_n
+ N_A_27_47#_c_252_n PM_SKY130_FD_SC_HD__DFRTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DFRTP_1%D N_D_M1025_g N_D_M1024_g N_D_c_470_n N_D_c_474_n
+ D N_D_c_471_n PM_SKY130_FD_SC_HD__DFRTP_1%D
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_193_47# N_A_193_47#_M1012_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1026_g N_A_193_47#_M1017_g N_A_193_47#_c_523_n
+ N_A_193_47#_M1020_g N_A_193_47#_M1010_g N_A_193_47#_c_524_n
+ N_A_193_47#_c_525_n N_A_193_47#_c_526_n N_A_193_47#_c_534_n
+ N_A_193_47#_c_535_n N_A_193_47#_c_527_n N_A_193_47#_c_528_n
+ N_A_193_47#_c_536_n N_A_193_47#_c_537_n N_A_193_47#_c_538_n
+ N_A_193_47#_c_539_n N_A_193_47#_c_540_n N_A_193_47#_c_541_n
+ N_A_193_47#_c_542_n N_A_193_47#_c_543_n N_A_193_47#_c_544_n
+ N_A_193_47#_c_529_n PM_SKY130_FD_SC_HD__DFRTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_761_289# N_A_761_289#_M1019_d
+ N_A_761_289#_M1014_d N_A_761_289#_M1009_g N_A_761_289#_M1002_g
+ N_A_761_289#_c_738_n N_A_761_289#_c_739_n N_A_761_289#_c_760_n
+ N_A_761_289#_c_735_n N_A_761_289#_c_762_n N_A_761_289#_c_747_n
+ N_A_761_289#_c_767_n N_A_761_289#_c_749_n N_A_761_289#_c_785_p
+ N_A_761_289#_c_750_n N_A_761_289#_c_751_n
+ PM_SKY130_FD_SC_HD__DFRTP_1%A_761_289#
x_PM_SKY130_FD_SC_HD__DFRTP_1%RESET_B N_RESET_B_M1003_g N_RESET_B_M1027_g
+ N_RESET_B_M1004_g N_RESET_B_M1016_g RESET_B RESET_B N_RESET_B_c_847_n
+ N_RESET_B_c_848_n N_RESET_B_c_849_n N_RESET_B_c_850_n N_RESET_B_c_851_n
+ N_RESET_B_c_852_n N_RESET_B_c_853_n N_RESET_B_c_854_n N_RESET_B_c_855_n
+ N_RESET_B_c_856_n PM_SKY130_FD_SC_HD__DFRTP_1%RESET_B
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_543_47# N_A_543_47#_M1008_d N_A_543_47#_M1026_d
+ N_A_543_47#_M1019_g N_A_543_47#_c_1003_n N_A_543_47#_c_1004_n
+ N_A_543_47#_M1014_g N_A_543_47#_c_1012_n N_A_543_47#_c_1033_n
+ N_A_543_47#_c_1005_n N_A_543_47#_c_998_n N_A_543_47#_c_999_n
+ N_A_543_47#_c_1000_n N_A_543_47#_c_1001_n N_A_543_47#_c_1002_n
+ PM_SKY130_FD_SC_HD__DFRTP_1%A_543_47#
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_1283_21# N_A_1283_21#_M1001_d
+ N_A_1283_21#_M1016_d N_A_1283_21#_M1022_g N_A_1283_21#_M1007_g
+ N_A_1283_21#_M1005_g N_A_1283_21#_M1015_g N_A_1283_21#_c_1125_n
+ N_A_1283_21#_c_1126_n N_A_1283_21#_c_1166_n N_A_1283_21#_c_1171_n
+ N_A_1283_21#_c_1230_p N_A_1283_21#_c_1137_n N_A_1283_21#_c_1138_n
+ N_A_1283_21#_c_1127_n N_A_1283_21#_c_1128_n N_A_1283_21#_c_1139_n
+ N_A_1283_21#_c_1129_n N_A_1283_21#_c_1130_n N_A_1283_21#_c_1131_n
+ N_A_1283_21#_c_1132_n N_A_1283_21#_c_1133_n N_A_1283_21#_c_1134_n
+ PM_SKY130_FD_SC_HD__DFRTP_1%A_1283_21#
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_1108_47# N_A_1108_47#_M1020_d
+ N_A_1108_47#_M1021_d N_A_1108_47#_M1013_g N_A_1108_47#_M1001_g
+ N_A_1108_47#_c_1277_n N_A_1108_47#_c_1280_n N_A_1108_47#_c_1270_n
+ N_A_1108_47#_c_1273_n N_A_1108_47#_c_1274_n N_A_1108_47#_c_1275_n
+ N_A_1108_47#_c_1276_n PM_SKY130_FD_SC_HD__DFRTP_1%A_1108_47#
x_PM_SKY130_FD_SC_HD__DFRTP_1%VPWR N_VPWR_M1011_d N_VPWR_M1024_s N_VPWR_M1009_d
+ N_VPWR_M1014_s N_VPWR_M1007_d N_VPWR_M1013_d N_VPWR_M1015_s N_VPWR_c_1373_n
+ N_VPWR_c_1374_n N_VPWR_c_1375_n N_VPWR_c_1376_n N_VPWR_c_1377_n
+ N_VPWR_c_1378_n N_VPWR_c_1379_n N_VPWR_c_1380_n N_VPWR_c_1381_n
+ N_VPWR_c_1382_n N_VPWR_c_1383_n N_VPWR_c_1384_n N_VPWR_c_1385_n VPWR
+ N_VPWR_c_1386_n N_VPWR_c_1387_n N_VPWR_c_1388_n N_VPWR_c_1389_n
+ N_VPWR_c_1390_n N_VPWR_c_1372_n N_VPWR_c_1392_n N_VPWR_c_1393_n
+ N_VPWR_c_1394_n N_VPWR_c_1395_n PM_SKY130_FD_SC_HD__DFRTP_1%VPWR
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_448_47# N_A_448_47#_M1025_d N_A_448_47#_M1024_d
+ N_A_448_47#_c_1520_n N_A_448_47#_c_1537_n N_A_448_47#_c_1528_n
+ PM_SKY130_FD_SC_HD__DFRTP_1%A_448_47#
x_PM_SKY130_FD_SC_HD__DFRTP_1%A_651_413# N_A_651_413#_M1006_d
+ N_A_651_413#_M1027_d N_A_651_413#_c_1554_n N_A_651_413#_c_1555_n
+ N_A_651_413#_c_1556_n N_A_651_413#_c_1557_n
+ PM_SKY130_FD_SC_HD__DFRTP_1%A_651_413#
x_PM_SKY130_FD_SC_HD__DFRTP_1%Q N_Q_M1005_d N_Q_M1015_d N_Q_c_1592_n Q Q Q Q Q
+ PM_SKY130_FD_SC_HD__DFRTP_1%Q
x_PM_SKY130_FD_SC_HD__DFRTP_1%VGND N_VGND_M1023_d N_VGND_M1025_s N_VGND_M1003_d
+ N_VGND_M1022_d N_VGND_M1005_s N_VGND_c_1605_n N_VGND_c_1606_n N_VGND_c_1607_n
+ N_VGND_c_1608_n N_VGND_c_1609_n N_VGND_c_1610_n N_VGND_c_1611_n
+ N_VGND_c_1612_n N_VGND_c_1613_n N_VGND_c_1614_n VGND N_VGND_c_1615_n
+ N_VGND_c_1616_n N_VGND_c_1617_n N_VGND_c_1618_n N_VGND_c_1619_n
+ N_VGND_c_1620_n N_VGND_c_1621_n PM_SKY130_FD_SC_HD__DFRTP_1%VGND
cc_1 VNB N_CLK_c_193_n 0.0577303f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.325
cc_2 VNB N_CLK_c_194_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0158337f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_27_47#_M1012_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_5 VNB N_A_27_47#_M1008_g 0.0209769f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_6 VNB N_A_27_47#_c_235_n 0.00890826f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_7 VNB N_A_27_47#_c_236_n 0.0150251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_237_n 0.00188961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_238_n 0.0380394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1018_g 0.0280213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_240_n 0.0111414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_241_n 7.34103e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_242_n 0.00783792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_243_n 0.0271377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_244_n 0.00215116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_245_n 0.0264033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_246_n 6.62431e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_247_n 0.0023967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_248_n 0.00191399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_249_n 0.0231886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_250_n 0.0236925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_251_n 0.00799011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_252_n 0.00574157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D_M1025_g 0.0533319f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_25 VNB N_D_c_470_n 0.0139927f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_26 VNB N_D_c_471_n 0.0188284f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_27 VNB N_A_193_47#_M1017_g 0.0237069f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_A_193_47#_c_523_n 0.0181872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_c_524_n 0.00292129f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_30 VNB N_A_193_47#_c_525_n 0.00474375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_526_n 0.0376939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_527_n 0.00318417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_528_n 0.027804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_529_n 0.0131434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_761_289#_M1002_g 0.0470937f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_36 VNB N_A_761_289#_c_735_n 0.00648449f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_37 VNB N_RESET_B_M1027_g 0.00906477f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_38 VNB N_RESET_B_M1004_g 0.0270317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_M1016_g 9.0366e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_40 VNB RESET_B 0.00278754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_847_n 0.00606631f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_42 VNB N_RESET_B_c_848_n 0.010211f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_43 VNB N_RESET_B_c_849_n 0.0158918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_RESET_B_c_850_n 6.54108e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_851_n 0.0012119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_852_n 0.0033021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_853_n 0.0257225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_854_n 0.0174472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_855_n 0.0250293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_856_n 0.00240216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_543_47#_M1019_g 0.0193117f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_52 VNB N_A_543_47#_c_998_n 0.0116433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_543_47#_c_999_n 0.00578907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_543_47#_c_1000_n 0.00317656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_543_47#_c_1001_n 0.00141599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_543_47#_c_1002_n 0.0285537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1283_21#_M1022_g 0.02143f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_58 VNB N_A_1283_21#_M1007_g 0.00982494f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_59 VNB N_A_1283_21#_c_1125_n 0.00209314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1283_21#_c_1126_n 6.41492e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1283_21#_c_1127_n 0.00297294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1283_21#_c_1128_n 0.00801962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1283_21#_c_1129_n 0.011929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1283_21#_c_1130_n 0.029969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1283_21#_c_1131_n 0.0073052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1283_21#_c_1132_n 0.0142842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1283_21#_c_1133_n 0.0464685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1283_21#_c_1134_n 0.022252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1108_47#_M1001_g 0.0455697f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_70 VNB N_A_1108_47#_c_1270_n 0.00617495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VPWR_c_1372_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_448_47#_c_1520_n 0.0051081f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_73 VNB N_Q_c_1592_n 0.00479254f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_74 VNB Q 0.0154962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB Q 0.0240401f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_76 VNB N_VGND_c_1605_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_77 VNB N_VGND_c_1606_n 0.0192467f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_78 VNB N_VGND_c_1607_n 0.00858778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1608_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1609_n 0.00480551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1610_n 0.00267922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1611_n 0.0711727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1612_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1613_n 0.0475682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1614_n 0.00362291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1615_n 0.0147253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1616_n 0.0372264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1617_n 0.0151507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1618_n 0.445672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1619_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1620_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1621_n 0.00459558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VPB N_CLK_c_193_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.325
cc_94 VPB N_CLK_c_197_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_95 VPB N_CLK_c_198_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_96 VPB N_CLK_c_199_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_97 VPB CLK 0.0152002f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_98 VPB N_A_27_47#_M1000_g 0.0393762f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_99 VPB N_A_27_47#_c_236_n 0.0162228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_c_237_n 0.00553413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_47#_M1006_g 0.0491475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_c_238_n 0.0112552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_47#_M1021_g 0.0463897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_47#_c_259_n 0.00118305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_c_260_n 0.0297336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_47#_c_244_n 4.26143e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_47#_c_247_n 0.00320885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_c_248_n 3.60888e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_c_249_n 0.012023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_c_251_n 0.00283708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_252_n 9.66093e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_D_M1024_g 0.0392567f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_113 VPB N_D_c_470_n 0.0355299f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_114 VPB N_D_c_474_n 0.0197975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB D 0.0281043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_D_c_471_n 0.00129394f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_117 VPB N_A_193_47#_M1026_g 0.0211021f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_118 VPB N_A_193_47#_M1010_g 0.0185283f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_119 VPB N_A_193_47#_c_524_n 0.00403367f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_120 VPB N_A_193_47#_c_525_n 0.00387694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_193_47#_c_534_n 0.00222651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_193_47#_c_535_n 0.00160169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_193_47#_c_536_n 0.012684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_193_47#_c_537_n 0.00221097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_193_47#_c_538_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_193_47#_c_539_n 0.00178929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_193_47#_c_540_n 0.005939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_193_47#_c_541_n 0.00225318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_193_47#_c_542_n 0.0267174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_193_47#_c_543_n 0.0305358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_193_47#_c_544_n 0.00788798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_193_47#_c_529_n 0.0113511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_761_289#_M1009_g 0.0280169f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_134 VPB N_A_761_289#_M1002_g 0.00821552f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_135 VPB N_A_761_289#_c_738_n 0.0139674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_761_289#_c_739_n 0.0282266f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_137 VPB N_A_761_289#_c_735_n 0.00172612f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_138 VPB N_RESET_B_M1027_g 0.0573733f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_139 VPB N_RESET_B_M1016_g 0.0509764f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_140 VPB N_RESET_B_c_856_n 0.00388678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_543_47#_c_1003_n 0.0276965f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_142 VPB N_A_543_47#_c_1004_n 0.0174138f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_143 VPB N_A_543_47#_c_1005_n 0.00704944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_543_47#_c_999_n 0.00782024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_543_47#_c_1000_n 0.00346469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_543_47#_c_1001_n 0.00113493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_543_47#_c_1002_n 0.0226938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_1283_21#_M1007_g 0.0502048f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_149 VPB N_A_1283_21#_M1015_g 0.0254791f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_150 VPB N_A_1283_21#_c_1137_n 0.00810586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_1283_21#_c_1138_n 0.00304108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_1283_21#_c_1139_n 0.0141175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_1283_21#_c_1129_n 0.00951421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_1283_21#_c_1130_n 0.00513292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_1283_21#_c_1132_n 2.87059e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_1108_47#_M1013_g 0.0262097f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_157 VPB N_A_1108_47#_M1001_g 0.0106007f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_158 VPB N_A_1108_47#_c_1273_n 0.0110964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_1108_47#_c_1274_n 0.00205899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_1108_47#_c_1275_n 0.0232558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1108_47#_c_1276_n 0.0289902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1373_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1374_n 0.00927346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1375_n 0.00273179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1376_n 0.00650484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1377_n 0.00223179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1378_n 0.00425084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1379_n 0.0050535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1380_n 0.0475825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1381_n 0.00507461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1382_n 0.0394977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1383_n 0.0035344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1384_n 0.0122568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1385_n 0.00513086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1386_n 0.0146985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1387_n 0.0265368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1388_n 0.0170787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1389_n 0.0102261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1390_n 0.0156754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1372_n 0.0667768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1392_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1393_n 0.00477715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1394_n 0.00572697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1395_n 0.00459796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_448_47#_c_1520_n 0.00778159f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_186 VPB N_A_651_413#_c_1554_n 4.85478e-19 $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_187 VPB N_A_651_413#_c_1555_n 0.00848337f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.665
cc_188 VPB N_A_651_413#_c_1556_n 0.00246665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_651_413#_c_1557_n 7.0682e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB Q 0.0420037f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_191 N_CLK_c_193_n N_A_27_47#_M1012_g 0.00510767f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_192 N_CLK_c_194_n N_A_27_47#_M1012_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_193 CLK N_A_27_47#_M1012_g 3.09846e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_194 N_CLK_c_197_n N_A_27_47#_M1000_g 0.00531917f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_195 N_CLK_c_199_n N_A_27_47#_M1000_g 0.0275602f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_196 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_197 N_CLK_c_193_n N_A_27_47#_c_241_n 0.00787672f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_198 N_CLK_c_194_n N_A_27_47#_c_241_n 0.00695273f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_199 CLK N_A_27_47#_c_241_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_200 N_CLK_c_193_n N_A_27_47#_c_242_n 0.0070116f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_201 CLK N_A_27_47#_c_242_n 0.0220292f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_202 N_CLK_c_198_n N_A_27_47#_c_259_n 0.0128403f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_203 N_CLK_c_199_n N_A_27_47#_c_259_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_204 CLK N_A_27_47#_c_259_n 0.00728212f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_205 N_CLK_c_193_n N_A_27_47#_c_260_n 4.93713e-19 $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_206 N_CLK_c_198_n N_A_27_47#_c_260_n 2.20356e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_207 N_CLK_c_199_n N_A_27_47#_c_260_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_208 CLK N_A_27_47#_c_260_n 0.0231715f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_209 CLK N_A_27_47#_c_244_n 0.00784263f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_210 N_CLK_c_193_n N_A_27_47#_c_247_n 0.00475399f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_211 N_CLK_c_197_n N_A_27_47#_c_247_n 7.09762e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_212 N_CLK_c_199_n N_A_27_47#_c_247_n 0.00454961f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_213 CLK N_A_27_47#_c_247_n 0.048988f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_214 N_CLK_c_193_n N_A_27_47#_c_249_n 0.0179788f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_215 CLK N_A_27_47#_c_249_n 0.00143822f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_216 N_CLK_c_198_n N_VPWR_c_1373_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_217 N_CLK_c_198_n N_VPWR_c_1386_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_218 N_CLK_c_198_n N_VPWR_c_1372_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_219 N_CLK_c_194_n N_VGND_c_1605_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_220 N_CLK_c_193_n N_VGND_c_1615_n 4.74473e-19 $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_221 N_CLK_c_194_n N_VGND_c_1615_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_222 N_CLK_c_194_n N_VGND_c_1618_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_223 N_A_27_47#_M1008_g N_D_M1025_g 0.0124137f $X=2.64 $Y=0.415 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_235_n N_D_M1025_g 0.00561622f $X=2.642 $Y=1.245 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_243_n N_D_M1025_g 0.00237886f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_246_n N_D_M1025_g 0.00141197f $X=2.675 $Y=1.19 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_250_n N_D_M1025_g 0.0194268f $X=2.585 $Y=0.93 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_251_n N_D_M1025_g 0.00359265f $X=2.585 $Y=0.93 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_243_n N_D_c_470_n 0.00328759f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_249_n N_D_c_470_n 0.00307512f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_237_n N_D_c_474_n 0.00561622f $X=2.72 $Y=1.32 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_243_n N_D_c_474_n 0.00121575f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_243_n D 0.00176122f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_243_n N_D_c_471_n 0.0454089f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_235 N_A_27_47#_M1006_g N_A_193_47#_M1026_g 0.0202456f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_M1008_g N_A_193_47#_M1017_g 0.0132876f $X=2.64 $Y=0.415 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1018_g N_A_193_47#_c_523_n 0.0127456f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1021_g N_A_193_47#_M1010_g 0.0170357f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_236_n N_A_193_47#_c_524_n 0.0110546f $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1006_g N_A_193_47#_c_524_n 0.00405215f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_245_n N_A_193_47#_c_524_n 0.0110887f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_246_n N_A_193_47#_c_524_n 5.58797e-19 $X=2.675 $Y=1.19 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_250_n N_A_193_47#_c_524_n 0.00150746f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_251_n N_A_193_47#_c_524_n 0.0290824f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_238_n N_A_193_47#_c_525_n 0.00866804f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_246 N_A_27_47#_M1018_g N_A_193_47#_c_525_n 3.88889e-19 $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_245_n N_A_193_47#_c_525_n 0.0145489f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_248_n N_A_193_47#_c_525_n 5.12182e-19 $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_252_n N_A_193_47#_c_525_n 0.045569f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1018_g N_A_193_47#_c_526_n 0.021218f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_245_n N_A_193_47#_c_526_n 0.00188252f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_252_n N_A_193_47#_c_526_n 0.00185788f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_238_n N_A_193_47#_c_534_n 0.00133124f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_254 N_A_27_47#_M1021_g N_A_193_47#_c_534_n 0.0109104f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_245_n N_A_193_47#_c_534_n 0.00491458f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_252_n N_A_193_47#_c_534_n 0.00841432f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_236_n N_A_193_47#_c_527_n 0.00114671f $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_245_n N_A_193_47#_c_527_n 0.00894827f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_250_n N_A_193_47#_c_527_n 7.0175e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_251_n N_A_193_47#_c_527_n 0.0184123f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_236_n N_A_193_47#_c_528_n 0.0226065f $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_245_n N_A_193_47#_c_528_n 0.00261571f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_250_n N_A_193_47#_c_528_n 0.0175107f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_251_n N_A_193_47#_c_528_n 8.36786e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_243_n N_A_193_47#_c_536_n 0.0494564f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_245_n N_A_193_47#_c_536_n 0.00684111f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_246_n N_A_193_47#_c_536_n 0.0133153f $X=2.675 $Y=1.19 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_251_n N_A_193_47#_c_536_n 0.00548636f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1000_g N_A_193_47#_c_537_n 0.00307706f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_259_n N_A_193_47#_c_537_n 0.00527405f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_260_n N_A_193_47#_c_537_n 3.65662e-19 $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_243_n N_A_193_47#_c_537_n 0.0136396f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_247_n N_A_193_47#_c_537_n 0.00104863f $X=0.695 $Y=1.19 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1006_g N_A_193_47#_c_538_n 0.00283709f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1021_g N_A_193_47#_c_538_n 0.00608452f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_276 N_A_27_47#_c_245_n N_A_193_47#_c_538_n 0.121215f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_236_n N_A_193_47#_c_539_n 3.78985e-19 $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1006_g N_A_193_47#_c_539_n 0.00277626f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_245_n N_A_193_47#_c_539_n 0.0129897f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_236_n N_A_193_47#_c_540_n 8.09221e-19 $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_237_n N_A_193_47#_c_540_n 0.00542966f $X=2.72 $Y=1.32 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1006_g N_A_193_47#_c_540_n 0.00325095f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_245_n N_A_193_47#_c_540_n 0.00524922f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_246_n N_A_193_47#_c_540_n 2.72172e-19 $X=2.675 $Y=1.19 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_251_n N_A_193_47#_c_540_n 0.00817823f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1021_g N_A_193_47#_c_541_n 0.00147605f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_248_n N_A_193_47#_c_541_n 0.0139913f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_252_n N_A_193_47#_c_541_n 7.23087e-19 $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_237_n N_A_193_47#_c_542_n 0.0187505f $X=2.72 $Y=1.32 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1006_g N_A_193_47#_c_542_n 0.0138904f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_250_n N_A_193_47#_c_542_n 6.13774e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_251_n N_A_193_47#_c_542_n 0.00142642f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_238_n N_A_193_47#_c_543_n 0.00311561f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_294 N_A_27_47#_M1021_g N_A_193_47#_c_543_n 0.0207208f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_248_n N_A_193_47#_c_543_n 0.00104369f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_252_n N_A_193_47#_c_543_n 4.78088e-19 $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_238_n N_A_193_47#_c_544_n 0.00367588f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_298 N_A_27_47#_M1021_g N_A_193_47#_c_544_n 0.00525218f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_299 N_A_27_47#_c_248_n N_A_193_47#_c_544_n 0.00244943f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_252_n N_A_193_47#_c_544_n 0.0147695f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1012_g N_A_193_47#_c_529_n 0.0227708f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_241_n N_A_193_47#_c_529_n 0.01251f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_259_n N_A_193_47#_c_529_n 0.00874344f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_243_n N_A_193_47#_c_529_n 0.0193882f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_244_n N_A_193_47#_c_529_n 0.0021977f $X=0.84 $Y=1.19 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_247_n N_A_193_47#_c_529_n 0.0685829f $X=0.695 $Y=1.19 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_236_n N_A_761_289#_M1002_g 0.00256582f $X=3.105 $Y=1.32
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_245_n N_A_761_289#_M1002_g 0.0022411f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1006_g N_A_761_289#_c_738_n 6.41799e-19 $X=3.18 $Y=2.275
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_c_245_n N_A_761_289#_c_738_n 0.00791634f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_M1006_g N_A_761_289#_c_739_n 0.01719f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_245_n N_A_761_289#_c_735_n 0.0128787f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_M1021_g N_A_761_289#_c_747_n 0.00242771f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_c_245_n N_A_761_289#_c_747_n 0.00205194f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_315 N_A_27_47#_M1021_g N_A_761_289#_c_749_n 0.00383854f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_245_n N_A_761_289#_c_750_n 7.74909e-19 $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_M1021_g N_A_761_289#_c_751_n 2.31682e-19 $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_c_245_n N_RESET_B_M1027_g 0.00162058f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_245_n N_RESET_B_c_847_n 0.0589913f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_245_n N_RESET_B_c_848_n 0.00492178f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_238_n N_RESET_B_c_849_n 5.35574e-19 $X=5.845 $Y=1.395 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_245_n N_RESET_B_c_849_n 0.12382f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_248_n N_RESET_B_c_849_n 0.0255775f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_252_n N_RESET_B_c_849_n 0.0184793f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_245_n N_RESET_B_c_853_n 0.00221649f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_M1021_g N_A_543_47#_c_1003_n 0.0268099f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_245_n N_A_543_47#_c_1003_n 0.00359773f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_M1006_g N_A_543_47#_c_1012_n 0.0169036f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_236_n N_A_543_47#_c_1005_n 0.00114222f $X=3.105 $Y=1.32
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_M1006_g N_A_543_47#_c_1005_n 0.0167379f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_245_n N_A_543_47#_c_1005_n 4.47512e-19 $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_245_n N_A_543_47#_c_998_n 0.0135671f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_245_n N_A_543_47#_c_999_n 0.0379321f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_236_n N_A_543_47#_c_1000_n 0.00382694f $X=3.105 $Y=1.32
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_245_n N_A_543_47#_c_1000_n 0.0134122f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_245_n N_A_543_47#_c_1001_n 0.0100049f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_245_n N_A_543_47#_c_1002_n 0.00476255f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_M1018_g N_A_1283_21#_M1022_g 0.0308149f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_252_n N_A_1283_21#_M1022_g 6.8514e-19 $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_238_n N_A_1283_21#_M1007_g 0.00175162f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_M1021_g N_A_1283_21#_M1007_g 0.00178563f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_238_n N_A_1283_21#_c_1133_n 0.0089256f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_238_n N_A_1108_47#_c_1277_n 8.21465e-19 $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_M1018_g N_A_1108_47#_c_1277_n 0.0109079f $X=6.01 $Y=0.415
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_252_n N_A_1108_47#_c_1277_n 0.0215171f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_M1021_g N_A_1108_47#_c_1280_n 0.00464335f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_238_n N_A_1108_47#_c_1270_n 0.00235645f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_M1018_g N_A_1108_47#_c_1270_n 0.00182809f $X=6.01 $Y=0.415
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_248_n N_A_1108_47#_c_1270_n 0.00772758f $X=6.11 $Y=1.19
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_252_n N_A_1108_47#_c_1270_n 0.0429822f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_238_n N_A_1108_47#_c_1273_n 0.00164867f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_M1021_g N_A_1108_47#_c_1273_n 0.00219772f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_252_n N_A_1108_47#_c_1273_n 8.53289e-19 $X=6.07 $Y=1.11
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_259_n N_VPWR_M1011_d 0.00167655f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_355 N_A_27_47#_M1000_g N_VPWR_c_1373_n 0.00939211f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_259_n N_VPWR_c_1373_n 0.0175536f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_260_n N_VPWR_c_1373_n 0.0127425f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_358 N_A_27_47#_M1021_g N_VPWR_c_1376_n 0.00111281f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1006_g N_VPWR_c_1380_n 0.00357863f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_M1021_g N_VPWR_c_1382_n 0.0055505f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_259_n N_VPWR_c_1386_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_362 N_A_27_47#_c_260_n N_VPWR_c_1386_n 0.0181185f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_363 N_A_27_47#_M1000_g N_VPWR_c_1387_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_M1000_g N_VPWR_c_1372_n 0.00859122f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_M1006_g N_VPWR_c_1372_n 0.00600164f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_M1021_g N_VPWR_c_1372_n 0.00644128f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_259_n N_VPWR_c_1372_n 0.00507261f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_260_n N_VPWR_c_1372_n 0.00973967f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_M1008_g N_A_448_47#_c_1520_n 0.00138047f $X=2.64 $Y=0.415
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_235_n N_A_448_47#_c_1520_n 3.20092e-19 $X=2.642 $Y=1.245
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_243_n N_A_448_47#_c_1520_n 0.0205223f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_246_n N_A_448_47#_c_1520_n 0.00258354f $X=2.675 $Y=1.19
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_250_n N_A_448_47#_c_1520_n 3.50691e-19 $X=2.585 $Y=0.93
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_251_n N_A_448_47#_c_1520_n 0.0463537f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_246_n N_A_448_47#_c_1528_n 6.44071e-19 $X=2.675 $Y=1.19
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_250_n N_A_448_47#_c_1528_n 4.7648e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_251_n N_A_448_47#_c_1528_n 0.0060732f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_M1006_g N_A_651_413#_c_1554_n 8.91651e-19 $X=3.18 $Y=2.275
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_245_n N_A_651_413#_c_1555_n 2.79618e-19 $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_M1006_g N_A_651_413#_c_1556_n 4.86622e-19 $X=3.18 $Y=2.275
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_241_n N_VGND_M1023_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_27_47#_M1012_g N_VGND_c_1605_n 0.0111875f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_241_n N_VGND_c_1605_n 0.0166634f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_244_n N_VGND_c_1605_n 9.27814e-19 $X=0.84 $Y=1.19 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_249_n N_VGND_c_1605_n 5.7379e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_M1012_g N_VGND_c_1606_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_M1012_g N_VGND_c_1607_n 0.00430756f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1008_g N_VGND_c_1611_n 0.00585385f $X=2.64 $Y=0.415 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_250_n N_VGND_c_1611_n 2.72564e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1018_g N_VGND_c_1613_n 0.00357877f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_240_n N_VGND_c_1615_n 0.0108577f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_392 N_A_27_47#_c_241_n N_VGND_c_1615_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_M1023_s N_VGND_c_1618_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_M1012_g N_VGND_c_1618_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_M1008_g N_VGND_c_1618_n 0.00642996f $X=2.64 $Y=0.415 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1018_g N_VGND_c_1618_n 0.00565064f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_240_n N_VGND_c_1618_n 0.00916732f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_241_n N_VGND_c_1618_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_251_n N_VGND_c_1618_n 0.00714893f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_400 N_D_M1024_g N_A_193_47#_M1026_g 0.014327f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_401 N_D_c_474_n N_A_193_47#_c_524_n 0.00459927f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_402 N_D_M1024_g N_A_193_47#_c_536_n 0.00135182f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_403 N_D_c_470_n N_A_193_47#_c_536_n 0.00295589f $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_404 D N_A_193_47#_c_536_n 0.0339847f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_405 D N_A_193_47#_c_537_n 0.00279509f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_406 N_D_c_474_n N_A_193_47#_c_540_n 0.00143055f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_407 N_D_c_474_n N_A_193_47#_c_542_n 0.0151527f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_408 N_D_c_470_n N_A_193_47#_c_529_n 8.20589e-19 $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_409 D N_A_193_47#_c_529_n 0.0745399f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_410 N_D_c_471_n N_A_193_47#_c_529_n 0.0518322f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_411 N_D_M1024_g N_VPWR_c_1374_n 0.0044954f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_412 N_D_c_470_n N_VPWR_c_1374_n 0.00536585f $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_413 D N_VPWR_c_1374_n 0.0228549f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_414 N_D_M1024_g N_VPWR_c_1380_n 0.00420613f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_415 D N_VPWR_c_1387_n 0.0211539f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_416 N_D_M1024_g N_VPWR_c_1372_n 0.00685455f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_417 D N_VPWR_c_1372_n 0.00588351f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_418 N_D_M1025_g N_A_448_47#_c_1520_n 0.0279651f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_419 N_D_M1024_g N_A_448_47#_c_1520_n 0.0259313f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_420 N_D_c_470_n N_A_448_47#_c_1520_n 0.00781441f $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_421 N_D_c_474_n N_A_448_47#_c_1520_n 0.0131062f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_422 D N_A_448_47#_c_1520_n 0.0365307f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_423 N_D_c_471_n N_A_448_47#_c_1520_n 0.0623934f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_424 N_D_M1025_g N_A_448_47#_c_1537_n 0.00588428f $X=2.165 $Y=0.445 $X2=0
+ $Y2=0
cc_425 N_D_M1025_g N_A_448_47#_c_1528_n 0.00163056f $X=2.165 $Y=0.445 $X2=0
+ $Y2=0
cc_426 N_D_c_471_n N_VGND_M1025_s 0.00431154f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_427 N_D_c_471_n N_VGND_c_1606_n 0.00272126f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_428 N_D_M1025_g N_VGND_c_1607_n 0.00675175f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_429 N_D_c_471_n N_VGND_c_1607_n 0.0275242f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_430 N_D_M1025_g N_VGND_c_1611_n 0.00367956f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_431 N_D_M1025_g N_VGND_c_1618_n 0.00677951f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_432 N_D_c_471_n N_VGND_c_1618_n 0.005702f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_433 N_A_193_47#_c_534_n N_A_761_289#_M1014_d 2.38738e-19 $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_434 N_A_193_47#_c_535_n N_A_761_289#_M1014_d 0.00203554f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_435 N_A_193_47#_c_538_n N_A_761_289#_M1014_d 0.00257222f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_436 N_A_193_47#_c_538_n N_A_761_289#_M1009_g 0.0023317f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_437 N_A_193_47#_M1017_g N_A_761_289#_M1002_g 0.00811432f $X=3.12 $Y=0.415
+ $X2=0 $Y2=0
cc_438 N_A_193_47#_c_528_n N_A_761_289#_M1002_g 0.00345535f $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_439 N_A_193_47#_c_538_n N_A_761_289#_c_738_n 0.0223886f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_440 N_A_193_47#_c_538_n N_A_761_289#_c_739_n 0.00270169f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_441 N_A_193_47#_c_523_n N_A_761_289#_c_760_n 0.00348356f $X=5.465 $Y=0.705
+ $X2=0 $Y2=0
cc_442 N_A_193_47#_c_535_n N_A_761_289#_c_735_n 0.00219387f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_443 N_A_193_47#_c_538_n N_A_761_289#_c_762_n 0.00749812f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_444 N_A_193_47#_c_535_n N_A_761_289#_c_747_n 0.0134011f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_445 N_A_193_47#_c_538_n N_A_761_289#_c_747_n 0.0181068f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_446 N_A_193_47#_c_541_n N_A_761_289#_c_747_n 0.00186336f $X=6.11 $Y=1.87
+ $X2=0 $Y2=0
cc_447 N_A_193_47#_c_544_n N_A_761_289#_c_747_n 0.00477525f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_448 N_A_193_47#_c_538_n N_A_761_289#_c_767_n 0.00696518f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_449 N_A_193_47#_c_525_n N_A_761_289#_c_750_n 0.0522946f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_450 N_A_193_47#_c_526_n N_A_761_289#_c_750_n 0.00348356f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_451 N_A_193_47#_c_535_n N_A_761_289#_c_751_n 0.0105163f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_452 N_A_193_47#_c_538_n N_RESET_B_M1027_g 0.00286324f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_453 N_A_193_47#_c_525_n N_RESET_B_c_849_n 0.0127742f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_454 N_A_193_47#_c_526_n N_RESET_B_c_849_n 0.00393129f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_455 N_A_193_47#_c_523_n N_A_543_47#_M1019_g 0.0103966f $X=5.465 $Y=0.705
+ $X2=0 $Y2=0
cc_456 N_A_193_47#_c_525_n N_A_543_47#_c_1003_n 7.67033e-19 $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_457 N_A_193_47#_c_526_n N_A_543_47#_c_1003_n 0.00138652f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_458 N_A_193_47#_c_535_n N_A_543_47#_c_1003_n 0.0016569f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_459 N_A_193_47#_c_538_n N_A_543_47#_c_1004_n 0.0027309f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_460 N_A_193_47#_M1026_g N_A_543_47#_c_1012_n 0.00421429f $X=2.685 $Y=2.275
+ $X2=0 $Y2=0
cc_461 N_A_193_47#_c_536_n N_A_543_47#_c_1012_n 4.97575e-19 $X=2.845 $Y=1.87
+ $X2=0 $Y2=0
cc_462 N_A_193_47#_c_538_n N_A_543_47#_c_1012_n 0.00304089f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_463 N_A_193_47#_c_539_n N_A_543_47#_c_1012_n 0.0046344f $X=3.135 $Y=1.87
+ $X2=0 $Y2=0
cc_464 N_A_193_47#_c_540_n N_A_543_47#_c_1012_n 0.0208127f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_465 N_A_193_47#_c_542_n N_A_543_47#_c_1012_n 4.68077e-19 $X=2.695 $Y=1.74
+ $X2=0 $Y2=0
cc_466 N_A_193_47#_M1017_g N_A_543_47#_c_1033_n 0.00973778f $X=3.12 $Y=0.415
+ $X2=0 $Y2=0
cc_467 N_A_193_47#_c_527_n N_A_543_47#_c_1033_n 0.0121475f $X=3.095 $Y=0.9 $X2=0
+ $Y2=0
cc_468 N_A_193_47#_c_528_n N_A_543_47#_c_1033_n 0.00324607f $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_469 N_A_193_47#_M1026_g N_A_543_47#_c_1005_n 8.68564e-19 $X=2.685 $Y=2.275
+ $X2=0 $Y2=0
cc_470 N_A_193_47#_c_524_n N_A_543_47#_c_1005_n 0.0155497f $X=2.99 $Y=1.575
+ $X2=0 $Y2=0
cc_471 N_A_193_47#_c_538_n N_A_543_47#_c_1005_n 0.0157004f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_472 N_A_193_47#_c_539_n N_A_543_47#_c_1005_n 0.00273426f $X=3.135 $Y=1.87
+ $X2=0 $Y2=0
cc_473 N_A_193_47#_c_540_n N_A_543_47#_c_1005_n 0.0280664f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_474 N_A_193_47#_c_542_n N_A_543_47#_c_1005_n 2.1939e-19 $X=2.695 $Y=1.74
+ $X2=0 $Y2=0
cc_475 N_A_193_47#_M1017_g N_A_543_47#_c_998_n 0.00647277f $X=3.12 $Y=0.415
+ $X2=0 $Y2=0
cc_476 N_A_193_47#_c_524_n N_A_543_47#_c_998_n 0.00810958f $X=2.99 $Y=1.575
+ $X2=0 $Y2=0
cc_477 N_A_193_47#_c_527_n N_A_543_47#_c_998_n 0.0159961f $X=3.095 $Y=0.9 $X2=0
+ $Y2=0
cc_478 N_A_193_47#_c_528_n N_A_543_47#_c_998_n 0.00150777f $X=3.095 $Y=0.9 $X2=0
+ $Y2=0
cc_479 N_A_193_47#_c_524_n N_A_543_47#_c_1000_n 0.0123239f $X=2.99 $Y=1.575
+ $X2=0 $Y2=0
cc_480 N_A_193_47#_c_527_n N_A_543_47#_c_1000_n 7.96251e-19 $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_481 N_A_193_47#_c_538_n N_A_543_47#_c_1000_n 0.00748451f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_482 N_A_193_47#_c_526_n N_A_543_47#_c_1002_n 0.0103966f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_483 N_A_193_47#_M1010_g N_A_1283_21#_M1007_g 0.0335217f $X=6.275 $Y=2.275
+ $X2=0 $Y2=0
cc_484 N_A_193_47#_c_543_n N_A_1283_21#_M1007_g 0.0198765f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_485 N_A_193_47#_c_544_n N_A_1283_21#_M1007_g 0.00149229f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_486 N_A_193_47#_c_525_n N_A_1108_47#_c_1277_n 0.0060004f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_487 N_A_193_47#_c_526_n N_A_1108_47#_c_1277_n 0.00264523f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_488 N_A_193_47#_M1010_g N_A_1108_47#_c_1280_n 0.0120896f $X=6.275 $Y=2.275
+ $X2=0 $Y2=0
cc_489 N_A_193_47#_c_534_n N_A_1108_47#_c_1280_n 7.08603e-19 $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_490 N_A_193_47#_c_538_n N_A_1108_47#_c_1280_n 9.42387e-19 $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_491 N_A_193_47#_c_541_n N_A_1108_47#_c_1280_n 0.00337735f $X=6.11 $Y=1.87
+ $X2=0 $Y2=0
cc_492 N_A_193_47#_c_543_n N_A_1108_47#_c_1280_n 3.21714e-19 $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_493 N_A_193_47#_c_544_n N_A_1108_47#_c_1280_n 0.02818f $X=6.265 $Y=1.74 $X2=0
+ $Y2=0
cc_494 N_A_193_47#_c_543_n N_A_1108_47#_c_1273_n 0.00200126f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_495 N_A_193_47#_c_544_n N_A_1108_47#_c_1273_n 0.0205187f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_496 N_A_193_47#_M1010_g N_A_1108_47#_c_1274_n 0.00233339f $X=6.275 $Y=2.275
+ $X2=0 $Y2=0
cc_497 N_A_193_47#_c_541_n N_A_1108_47#_c_1274_n 0.00209221f $X=6.11 $Y=1.87
+ $X2=0 $Y2=0
cc_498 N_A_193_47#_c_543_n N_A_1108_47#_c_1274_n 4.36865e-19 $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_499 N_A_193_47#_c_544_n N_A_1108_47#_c_1274_n 0.0162391f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_500 N_A_193_47#_c_538_n N_VPWR_M1014_s 0.00127798f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_501 N_A_193_47#_c_529_n N_VPWR_c_1373_n 0.012721f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_502 N_A_193_47#_c_536_n N_VPWR_c_1374_n 0.00656454f $X=2.845 $Y=1.87 $X2=0
+ $Y2=0
cc_503 N_A_193_47#_c_529_n N_VPWR_c_1374_n 4.4131e-19 $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_504 N_A_193_47#_c_538_n N_VPWR_c_1375_n 0.00139202f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_505 N_A_193_47#_c_538_n N_VPWR_c_1376_n 0.00326091f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_506 N_A_193_47#_M1026_g N_VPWR_c_1380_n 0.00427876f $X=2.685 $Y=2.275 $X2=0
+ $Y2=0
cc_507 N_A_193_47#_c_540_n N_VPWR_c_1380_n 0.00166184f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_508 N_A_193_47#_M1010_g N_VPWR_c_1382_n 0.00357877f $X=6.275 $Y=2.275 $X2=0
+ $Y2=0
cc_509 N_A_193_47#_c_529_n N_VPWR_c_1387_n 0.0120448f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_510 N_A_193_47#_M1026_g N_VPWR_c_1372_n 0.0059104f $X=2.685 $Y=2.275 $X2=0
+ $Y2=0
cc_511 N_A_193_47#_M1010_g N_VPWR_c_1372_n 0.00526867f $X=6.275 $Y=2.275 $X2=0
+ $Y2=0
cc_512 N_A_193_47#_c_536_n N_VPWR_c_1372_n 0.0759296f $X=2.845 $Y=1.87 $X2=0
+ $Y2=0
cc_513 N_A_193_47#_c_537_n N_VPWR_c_1372_n 0.0154052f $X=1.245 $Y=1.87 $X2=0
+ $Y2=0
cc_514 N_A_193_47#_c_538_n N_VPWR_c_1372_n 0.131729f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_515 N_A_193_47#_c_539_n N_VPWR_c_1372_n 0.0159609f $X=3.135 $Y=1.87 $X2=0
+ $Y2=0
cc_516 N_A_193_47#_c_540_n N_VPWR_c_1372_n 0.00140124f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_517 N_A_193_47#_c_541_n N_VPWR_c_1372_n 0.0158397f $X=6.11 $Y=1.87 $X2=0
+ $Y2=0
cc_518 N_A_193_47#_c_542_n N_VPWR_c_1372_n 4.39969e-19 $X=2.695 $Y=1.74 $X2=0
+ $Y2=0
cc_519 N_A_193_47#_c_529_n N_VPWR_c_1372_n 0.0029375f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_520 N_A_193_47#_M1026_g N_A_448_47#_c_1520_n 0.00392609f $X=2.685 $Y=2.275
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_c_536_n N_A_448_47#_c_1520_n 0.0288873f $X=2.845 $Y=1.87
+ $X2=0 $Y2=0
cc_522 N_A_193_47#_c_539_n N_A_448_47#_c_1520_n 0.00100139f $X=3.135 $Y=1.87
+ $X2=0 $Y2=0
cc_523 N_A_193_47#_c_540_n N_A_448_47#_c_1520_n 0.0185011f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_524 N_A_193_47#_c_542_n N_A_448_47#_c_1520_n 9.81315e-19 $X=2.695 $Y=1.74
+ $X2=0 $Y2=0
cc_525 N_A_193_47#_c_538_n N_A_651_413#_c_1555_n 0.0297495f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_526 N_A_193_47#_c_538_n N_A_651_413#_c_1556_n 0.00857493f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_527 N_A_193_47#_c_529_n N_VGND_c_1606_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_528 N_A_193_47#_c_529_n N_VGND_c_1607_n 0.00457032f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_M1017_g N_VGND_c_1611_n 0.00368123f $X=3.12 $Y=0.415 $X2=0
+ $Y2=0
cc_530 N_A_193_47#_c_523_n N_VGND_c_1613_n 0.0051118f $X=5.465 $Y=0.705 $X2=0
+ $Y2=0
cc_531 N_A_193_47#_c_525_n N_VGND_c_1613_n 0.00183172f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_532 N_A_193_47#_c_526_n N_VGND_c_1613_n 2.13253e-19 $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_533 N_A_193_47#_M1012_d N_VGND_c_1618_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_534 N_A_193_47#_M1017_g N_VGND_c_1618_n 0.00618454f $X=3.12 $Y=0.415 $X2=0
+ $Y2=0
cc_535 N_A_193_47#_c_523_n N_VGND_c_1618_n 0.00654107f $X=5.465 $Y=0.705 $X2=0
+ $Y2=0
cc_536 N_A_193_47#_c_525_n N_VGND_c_1618_n 0.00150843f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_537 N_A_193_47#_c_529_n N_VGND_c_1618_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_538 N_A_761_289#_M1009_g N_RESET_B_M1027_g 0.0224927f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_539 N_A_761_289#_M1002_g N_RESET_B_M1027_g 0.0177106f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_540 N_A_761_289#_c_738_n N_RESET_B_M1027_g 0.0115545f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_541 N_A_761_289#_c_739_n N_RESET_B_M1027_g 0.0220442f $X=3.94 $Y=1.61 $X2=0
+ $Y2=0
cc_542 N_A_761_289#_c_735_n N_RESET_B_M1027_g 4.12396e-19 $X=5.19 $Y=1.525 $X2=0
+ $Y2=0
cc_543 N_A_761_289#_c_762_n N_RESET_B_M1027_g 0.00253836f $X=5.19 $Y=1.835 $X2=0
+ $Y2=0
cc_544 N_A_761_289#_c_767_n N_RESET_B_M1027_g 9.1253e-19 $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_545 N_A_761_289#_M1002_g N_RESET_B_c_847_n 0.00269192f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_546 N_A_761_289#_M1002_g N_RESET_B_c_848_n 0.0139529f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_547 N_A_761_289#_c_735_n N_RESET_B_c_848_n 0.0051548f $X=5.19 $Y=1.525 $X2=0
+ $Y2=0
cc_548 N_A_761_289#_c_750_n N_RESET_B_c_848_n 0.00197464f $X=5.145 $Y=0.835
+ $X2=0 $Y2=0
cc_549 N_A_761_289#_M1019_d N_RESET_B_c_849_n 3.28012e-19 $X=5.045 $Y=0.235
+ $X2=0 $Y2=0
cc_550 N_A_761_289#_c_738_n N_RESET_B_c_849_n 2.43406e-19 $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_551 N_A_761_289#_c_735_n N_RESET_B_c_849_n 0.00696464f $X=5.19 $Y=1.525 $X2=0
+ $Y2=0
cc_552 N_A_761_289#_c_785_p N_RESET_B_c_849_n 0.00227253f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_553 N_A_761_289#_c_750_n N_RESET_B_c_849_n 0.0121464f $X=5.145 $Y=0.835 $X2=0
+ $Y2=0
cc_554 N_A_761_289#_M1002_g N_RESET_B_c_854_n 0.0635296f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_555 N_A_761_289#_c_785_p N_RESET_B_c_854_n 9.82944e-19 $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_556 N_A_761_289#_c_760_n N_A_543_47#_M1019_g 0.0061779f $X=5.145 $Y=0.705
+ $X2=0 $Y2=0
cc_557 N_A_761_289#_c_735_n N_A_543_47#_M1019_g 0.0120311f $X=5.19 $Y=1.525
+ $X2=0 $Y2=0
cc_558 N_A_761_289#_c_785_p N_A_543_47#_M1019_g 0.00225962f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_559 N_A_761_289#_c_750_n N_A_543_47#_M1019_g 0.00423512f $X=5.145 $Y=0.835
+ $X2=0 $Y2=0
cc_560 N_A_761_289#_c_738_n N_A_543_47#_c_1003_n 0.00207011f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_561 N_A_761_289#_c_735_n N_A_543_47#_c_1003_n 0.00860889f $X=5.19 $Y=1.525
+ $X2=0 $Y2=0
cc_562 N_A_761_289#_c_750_n N_A_543_47#_c_1003_n 8.88512e-19 $X=5.145 $Y=0.835
+ $X2=0 $Y2=0
cc_563 N_A_761_289#_c_751_n N_A_543_47#_c_1003_n 0.00482334f $X=5.19 $Y=1.61
+ $X2=0 $Y2=0
cc_564 N_A_761_289#_c_762_n N_A_543_47#_c_1004_n 0.00308571f $X=5.19 $Y=1.835
+ $X2=0 $Y2=0
cc_565 N_A_761_289#_c_747_n N_A_543_47#_c_1004_n 0.0106757f $X=5.495 $Y=1.92
+ $X2=0 $Y2=0
cc_566 N_A_761_289#_c_767_n N_A_543_47#_c_1004_n 0.00298755f $X=5.275 $Y=1.92
+ $X2=0 $Y2=0
cc_567 N_A_761_289#_c_749_n N_A_543_47#_c_1004_n 0.00453769f $X=5.58 $Y=2.3
+ $X2=0 $Y2=0
cc_568 N_A_761_289#_c_751_n N_A_543_47#_c_1004_n 0.00385118f $X=5.19 $Y=1.61
+ $X2=0 $Y2=0
cc_569 N_A_761_289#_M1009_g N_A_543_47#_c_1012_n 0.00124715f $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_570 N_A_761_289#_M1002_g N_A_543_47#_c_1033_n 0.00466363f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_571 N_A_761_289#_M1009_g N_A_543_47#_c_1005_n 4.99336e-19 $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_572 N_A_761_289#_M1002_g N_A_543_47#_c_1005_n 0.00150033f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_573 N_A_761_289#_c_738_n N_A_543_47#_c_1005_n 0.00842454f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_574 N_A_761_289#_c_739_n N_A_543_47#_c_1005_n 0.0048158f $X=3.94 $Y=1.61
+ $X2=0 $Y2=0
cc_575 N_A_761_289#_M1002_g N_A_543_47#_c_998_n 0.0114869f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_576 N_A_761_289#_M1002_g N_A_543_47#_c_999_n 0.0109334f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_577 N_A_761_289#_c_738_n N_A_543_47#_c_999_n 0.063308f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_578 N_A_761_289#_c_739_n N_A_543_47#_c_999_n 0.00338177f $X=3.94 $Y=1.61
+ $X2=0 $Y2=0
cc_579 N_A_761_289#_c_738_n N_A_543_47#_c_1001_n 0.0116159f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_580 N_A_761_289#_c_735_n N_A_543_47#_c_1001_n 0.0244986f $X=5.19 $Y=1.525
+ $X2=0 $Y2=0
cc_581 N_A_761_289#_c_738_n N_A_543_47#_c_1002_n 0.00751143f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_582 N_A_761_289#_c_749_n N_A_1108_47#_c_1280_n 0.0206716f $X=5.58 $Y=2.3
+ $X2=0 $Y2=0
cc_583 N_A_761_289#_c_738_n N_VPWR_M1014_s 0.00130684f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_584 N_A_761_289#_c_762_n N_VPWR_M1014_s 0.00241466f $X=5.19 $Y=1.835 $X2=0
+ $Y2=0
cc_585 N_A_761_289#_c_767_n N_VPWR_M1014_s 0.00353974f $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_586 N_A_761_289#_M1009_g N_VPWR_c_1375_n 0.0044935f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_587 N_A_761_289#_c_738_n N_VPWR_c_1376_n 0.00261535f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_588 N_A_761_289#_c_747_n N_VPWR_c_1376_n 0.003184f $X=5.495 $Y=1.92 $X2=0
+ $Y2=0
cc_589 N_A_761_289#_c_767_n N_VPWR_c_1376_n 0.008938f $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_590 N_A_761_289#_c_749_n N_VPWR_c_1376_n 0.0216047f $X=5.58 $Y=2.3 $X2=0
+ $Y2=0
cc_591 N_A_761_289#_M1009_g N_VPWR_c_1380_n 0.00432313f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_592 N_A_761_289#_c_747_n N_VPWR_c_1382_n 0.00199878f $X=5.495 $Y=1.92 $X2=0
+ $Y2=0
cc_593 N_A_761_289#_c_749_n N_VPWR_c_1382_n 0.0117479f $X=5.58 $Y=2.3 $X2=0
+ $Y2=0
cc_594 N_A_761_289#_M1014_d N_VPWR_c_1372_n 0.00326756f $X=5.425 $Y=1.645 $X2=0
+ $Y2=0
cc_595 N_A_761_289#_M1009_g N_VPWR_c_1372_n 0.00628822f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_596 N_A_761_289#_c_747_n N_VPWR_c_1372_n 0.00181326f $X=5.495 $Y=1.92 $X2=0
+ $Y2=0
cc_597 N_A_761_289#_c_767_n N_VPWR_c_1372_n 4.80263e-19 $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_598 N_A_761_289#_c_749_n N_VPWR_c_1372_n 0.00306902f $X=5.58 $Y=2.3 $X2=0
+ $Y2=0
cc_599 N_A_761_289#_M1009_g N_A_651_413#_c_1554_n 7.77269e-19 $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_600 N_A_761_289#_M1009_g N_A_651_413#_c_1555_n 0.0117327f $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_601 N_A_761_289#_c_738_n N_A_651_413#_c_1555_n 0.0556558f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_602 N_A_761_289#_c_739_n N_A_651_413#_c_1555_n 0.00332707f $X=3.94 $Y=1.61
+ $X2=0 $Y2=0
cc_603 N_A_761_289#_c_767_n N_A_651_413#_c_1555_n 0.00487217f $X=5.275 $Y=1.92
+ $X2=0 $Y2=0
cc_604 N_A_761_289#_c_785_p N_VGND_c_1608_n 0.0177195f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_605 N_A_761_289#_M1002_g N_VGND_c_1611_n 0.00585385f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_606 N_A_761_289#_c_785_p N_VGND_c_1613_n 0.0185505f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_607 N_A_761_289#_M1019_d N_VGND_c_1618_n 0.00246666f $X=5.045 $Y=0.235 $X2=0
+ $Y2=0
cc_608 N_A_761_289#_M1002_g N_VGND_c_1618_n 0.00633204f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_609 N_A_761_289#_c_785_p N_VGND_c_1618_n 0.00609105f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_848_n N_A_543_47#_M1019_g 0.00182794f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_849_n N_A_543_47#_M1019_g 0.00503251f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_850_n N_A_543_47#_M1019_g 4.85534e-19 $X=4.395 $Y=0.85 $X2=0
+ $Y2=0
cc_613 N_RESET_B_c_853_n N_A_543_47#_M1019_g 0.0070799f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_614 N_RESET_B_c_854_n N_A_543_47#_M1019_g 0.0129551f $X=4.37 $Y=0.765 $X2=0
+ $Y2=0
cc_615 N_RESET_B_c_847_n N_A_543_47#_c_998_n 0.00858647f $X=4.28 $Y=0.85 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_848_n N_A_543_47#_c_998_n 0.0146357f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_617 N_RESET_B_M1027_g N_A_543_47#_c_999_n 0.00939437f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_847_n N_A_543_47#_c_999_n 0.00116894f $X=4.28 $Y=0.85 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_848_n N_A_543_47#_c_999_n 0.0505984f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_849_n N_A_543_47#_c_999_n 0.00103298f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_853_n N_A_543_47#_c_999_n 0.00314155f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_622 N_RESET_B_M1027_g N_A_543_47#_c_1001_n 8.07088e-19 $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_623 N_RESET_B_c_848_n N_A_543_47#_c_1001_n 7.26099e-19 $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_624 N_RESET_B_c_849_n N_A_543_47#_c_1001_n 0.00420388f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_853_n N_A_543_47#_c_1001_n 5.16993e-19 $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_626 N_RESET_B_M1027_g N_A_543_47#_c_1002_n 0.0181811f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_849_n N_A_543_47#_c_1002_n 8.21109e-19 $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_628 N_RESET_B_c_853_n N_A_543_47#_c_1002_n 0.00600523f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_629 N_RESET_B_M1004_g N_A_1283_21#_M1022_g 0.0101625f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_630 N_RESET_B_c_849_n N_A_1283_21#_M1022_g 8.78915e-19 $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_631 N_RESET_B_M1016_g N_A_1283_21#_M1007_g 0.0333609f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_852_n N_A_1283_21#_M1007_g 0.00197455f $X=7.19 $Y=1.165 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_855_n N_A_1283_21#_M1007_g 0.00410139f $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_856_n N_A_1283_21#_M1007_g 0.00166565f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_635 N_RESET_B_M1004_g N_A_1283_21#_c_1125_n 3.49601e-19 $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_636 RESET_B N_A_1283_21#_c_1125_n 0.00296317f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_637 N_RESET_B_c_849_n N_A_1283_21#_c_1125_n 0.0109517f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_851_n N_A_1283_21#_c_1125_n 0.00740908f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_639 N_RESET_B_c_855_n N_A_1283_21#_c_1125_n 4.00963e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_856_n N_A_1283_21#_c_1125_n 0.006652f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_641 N_RESET_B_M1004_g N_A_1283_21#_c_1126_n 0.00733777f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_642 RESET_B N_A_1283_21#_c_1126_n 0.0043842f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_643 N_RESET_B_c_851_n N_A_1283_21#_c_1126_n 4.41459e-19 $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_644 N_RESET_B_M1004_g N_A_1283_21#_c_1166_n 0.00588467f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_645 RESET_B N_A_1283_21#_c_1166_n 0.0122946f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_646 N_RESET_B_c_851_n N_A_1283_21#_c_1166_n 0.00297971f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_647 N_RESET_B_c_855_n N_A_1283_21#_c_1166_n 9.38055e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_856_n N_A_1283_21#_c_1166_n 0.00166967f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_649 N_RESET_B_M1004_g N_A_1283_21#_c_1171_n 0.00390919f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_650 N_RESET_B_M1016_g N_A_1283_21#_c_1138_n 0.00230253f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_651 RESET_B N_A_1283_21#_c_1128_n 0.0127158f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_652 N_RESET_B_c_851_n N_A_1283_21#_c_1128_n 6.44878e-19 $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_653 N_RESET_B_c_856_n N_A_1283_21#_c_1139_n 0.0036174f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_654 N_RESET_B_M1004_g N_A_1283_21#_c_1131_n 0.00557763f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_655 RESET_B N_A_1283_21#_c_1131_n 0.0119774f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_656 N_RESET_B_c_849_n N_A_1283_21#_c_1131_n 0.0122086f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_851_n N_A_1283_21#_c_1131_n 0.00988863f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_658 N_RESET_B_c_855_n N_A_1283_21#_c_1131_n 4.8034e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_856_n N_A_1283_21#_c_1131_n 0.00872348f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_660 RESET_B N_A_1283_21#_c_1132_n 0.0155377f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_661 N_RESET_B_c_851_n N_A_1283_21#_c_1132_n 0.00108995f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_852_n N_A_1283_21#_c_1132_n 0.00126581f $X=7.19 $Y=1.165
+ $X2=0 $Y2=0
cc_663 N_RESET_B_c_856_n N_A_1283_21#_c_1132_n 0.0234117f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_664 N_RESET_B_M1004_g N_A_1283_21#_c_1133_n 0.00837678f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_665 N_RESET_B_c_849_n N_A_1283_21#_c_1133_n 0.00336334f $X=7.045 $Y=0.85
+ $X2=0 $Y2=0
cc_666 N_RESET_B_c_851_n N_A_1283_21#_c_1133_n 0.00369633f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_667 N_RESET_B_c_855_n N_A_1283_21#_c_1133_n 0.0123335f $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_668 N_RESET_B_c_856_n N_A_1283_21#_c_1133_n 5.46251e-19 $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_669 N_RESET_B_M1016_g N_A_1108_47#_M1013_g 0.0209796f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_670 N_RESET_B_M1004_g N_A_1108_47#_M1001_g 0.0345821f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_671 N_RESET_B_M1016_g N_A_1108_47#_M1001_g 0.00874253f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_672 RESET_B N_A_1108_47#_M1001_g 0.00845022f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_673 N_RESET_B_c_855_n N_A_1108_47#_M1001_g 0.0210473f $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_674 N_RESET_B_c_856_n N_A_1108_47#_M1001_g 0.00881611f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_675 N_RESET_B_c_849_n N_A_1108_47#_c_1277_n 0.012043f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_676 N_RESET_B_M1004_g N_A_1108_47#_c_1270_n 3.06785e-19 $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_677 N_RESET_B_c_849_n N_A_1108_47#_c_1270_n 0.0190486f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_678 N_RESET_B_c_852_n N_A_1108_47#_c_1270_n 0.00350005f $X=7.19 $Y=1.165
+ $X2=0 $Y2=0
cc_679 N_RESET_B_c_856_n N_A_1108_47#_c_1270_n 0.00372747f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_680 N_RESET_B_M1016_g N_A_1108_47#_c_1273_n 0.00109897f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_681 N_RESET_B_c_849_n N_A_1108_47#_c_1273_n 0.00621195f $X=7.045 $Y=0.85
+ $X2=0 $Y2=0
cc_682 N_RESET_B_c_856_n N_A_1108_47#_c_1273_n 0.00451828f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_683 N_RESET_B_M1016_g N_A_1108_47#_c_1274_n 0.00180441f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_684 N_RESET_B_M1016_g N_A_1108_47#_c_1275_n 0.0144262f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_685 N_RESET_B_c_852_n N_A_1108_47#_c_1275_n 0.00392251f $X=7.19 $Y=1.165
+ $X2=0 $Y2=0
cc_686 N_RESET_B_c_855_n N_A_1108_47#_c_1275_n 6.25544e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_687 N_RESET_B_c_856_n N_A_1108_47#_c_1275_n 0.0397801f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_688 N_RESET_B_M1016_g N_A_1108_47#_c_1276_n 0.0217285f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_856_n N_A_1108_47#_c_1276_n 0.00253996f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_690 N_RESET_B_M1027_g N_VPWR_c_1375_n 0.00862424f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_691 N_RESET_B_M1027_g N_VPWR_c_1376_n 0.00315462f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_692 N_RESET_B_M1016_g N_VPWR_c_1377_n 0.00837873f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_693 N_RESET_B_M1016_g N_VPWR_c_1378_n 7.11879e-19 $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_694 N_RESET_B_M1016_g N_VPWR_c_1384_n 0.0046653f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_695 N_RESET_B_M1027_g N_VPWR_c_1388_n 0.00345093f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_696 N_RESET_B_M1027_g N_VPWR_c_1372_n 0.00519819f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_697 N_RESET_B_M1016_g N_VPWR_c_1372_n 0.00799591f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_698 N_RESET_B_M1027_g N_A_651_413#_c_1555_n 0.0122302f $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_699 N_RESET_B_M1027_g N_A_651_413#_c_1557_n 0.00113125f $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_700 N_RESET_B_c_849_n N_VGND_M1003_d 0.0025426f $X=7.045 $Y=0.85 $X2=0 $Y2=0
cc_701 N_RESET_B_c_848_n N_VGND_c_1608_n 0.0066953f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_702 N_RESET_B_c_849_n N_VGND_c_1608_n 0.00423599f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_703 N_RESET_B_c_853_n N_VGND_c_1608_n 6.55014e-19 $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_704 N_RESET_B_c_854_n N_VGND_c_1608_n 0.0117447f $X=4.37 $Y=0.765 $X2=0 $Y2=0
cc_705 N_RESET_B_M1004_g N_VGND_c_1609_n 0.00402543f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_706 N_RESET_B_c_849_n N_VGND_c_1609_n 8.29415e-19 $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_RESET_B_c_853_n N_VGND_c_1611_n 0.00162298f $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_708 N_RESET_B_c_854_n N_VGND_c_1611_n 0.00585385f $X=4.37 $Y=0.765 $X2=0
+ $Y2=0
cc_709 N_RESET_B_M1004_g N_VGND_c_1616_n 0.0036601f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_710 N_RESET_B_M1004_g N_VGND_c_1618_n 0.00599573f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_711 N_RESET_B_c_847_n N_VGND_c_1618_n 0.0362506f $X=4.28 $Y=0.85 $X2=0 $Y2=0
cc_712 N_RESET_B_c_848_n N_VGND_c_1618_n 0.00772058f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_713 N_RESET_B_c_849_n N_VGND_c_1618_n 0.139055f $X=7.045 $Y=0.85 $X2=0 $Y2=0
cc_714 N_RESET_B_c_851_n N_VGND_c_1618_n 0.0148902f $X=7.19 $Y=0.965 $X2=0 $Y2=0
cc_715 N_RESET_B_c_853_n N_VGND_c_1618_n 0.00136687f $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_716 N_RESET_B_c_854_n N_VGND_c_1618_n 0.00606683f $X=4.37 $Y=0.765 $X2=0
+ $Y2=0
cc_717 RESET_B A_1462_47# 0.00176151f $X=7.405 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_718 N_A_543_47#_c_1004_n N_VPWR_c_1376_n 0.0111275f $X=5.35 $Y=1.57 $X2=0
+ $Y2=0
cc_719 N_A_543_47#_c_1002_n N_VPWR_c_1376_n 0.00129214f $X=4.85 $Y=1.17 $X2=0
+ $Y2=0
cc_720 N_A_543_47#_c_1012_n N_VPWR_c_1380_n 0.0397779f $X=3.245 $Y=2.3 $X2=0
+ $Y2=0
cc_721 N_A_543_47#_c_1004_n N_VPWR_c_1382_n 0.00290206f $X=5.35 $Y=1.57 $X2=0
+ $Y2=0
cc_722 N_A_543_47#_M1026_d N_VPWR_c_1372_n 0.00221211f $X=2.76 $Y=2.065 $X2=0
+ $Y2=0
cc_723 N_A_543_47#_c_1004_n N_VPWR_c_1372_n 0.00346038f $X=5.35 $Y=1.57 $X2=0
+ $Y2=0
cc_724 N_A_543_47#_c_1012_n N_VPWR_c_1372_n 0.0114478f $X=3.245 $Y=2.3 $X2=0
+ $Y2=0
cc_725 N_A_543_47#_c_1012_n N_A_448_47#_c_1520_n 0.0221744f $X=3.245 $Y=2.3
+ $X2=0 $Y2=0
cc_726 N_A_543_47#_c_1012_n N_A_651_413#_M1006_d 0.00470561f $X=3.245 $Y=2.3
+ $X2=-0.19 $Y2=-0.24
cc_727 N_A_543_47#_c_1005_n N_A_651_413#_M1006_d 6.28858e-19 $X=3.33 $Y=2.135
+ $X2=-0.19 $Y2=-0.24
cc_728 N_A_543_47#_c_1012_n N_A_651_413#_c_1554_n 0.019526f $X=3.245 $Y=2.3
+ $X2=0 $Y2=0
cc_729 N_A_543_47#_c_1005_n N_A_651_413#_c_1554_n 0.00726918f $X=3.33 $Y=2.135
+ $X2=0 $Y2=0
cc_730 N_A_543_47#_c_1004_n N_A_651_413#_c_1555_n 0.00137742f $X=5.35 $Y=1.57
+ $X2=0 $Y2=0
cc_731 N_A_543_47#_c_999_n N_A_651_413#_c_1555_n 4.0432e-19 $X=4.765 $Y=1.27
+ $X2=0 $Y2=0
cc_732 N_A_543_47#_c_1005_n N_A_651_413#_c_1556_n 0.0132883f $X=3.33 $Y=2.135
+ $X2=0 $Y2=0
cc_733 N_A_543_47#_c_1000_n N_A_651_413#_c_1556_n 0.0035943f $X=3.6 $Y=1.27
+ $X2=0 $Y2=0
cc_734 N_A_543_47#_c_1004_n N_A_651_413#_c_1557_n 0.00269162f $X=5.35 $Y=1.57
+ $X2=0 $Y2=0
cc_735 N_A_543_47#_M1019_g N_VGND_c_1608_n 0.00677972f $X=4.97 $Y=0.555 $X2=0
+ $Y2=0
cc_736 N_A_543_47#_c_999_n N_VGND_c_1608_n 0.00223331f $X=4.765 $Y=1.27 $X2=0
+ $Y2=0
cc_737 N_A_543_47#_c_1001_n N_VGND_c_1608_n 6.77929e-19 $X=4.85 $Y=1.17 $X2=0
+ $Y2=0
cc_738 N_A_543_47#_c_1002_n N_VGND_c_1608_n 0.001314f $X=4.85 $Y=1.17 $X2=0
+ $Y2=0
cc_739 N_A_543_47#_c_1033_n N_VGND_c_1611_n 0.0387784f $X=3.43 $Y=0.39 $X2=0
+ $Y2=0
cc_740 N_A_543_47#_M1019_g N_VGND_c_1613_n 0.00542163f $X=4.97 $Y=0.555 $X2=0
+ $Y2=0
cc_741 N_A_543_47#_M1008_d N_VGND_c_1618_n 0.00309942f $X=2.715 $Y=0.235 $X2=0
+ $Y2=0
cc_742 N_A_543_47#_M1019_g N_VGND_c_1618_n 0.00686855f $X=4.97 $Y=0.555 $X2=0
+ $Y2=0
cc_743 N_A_543_47#_c_1033_n N_VGND_c_1618_n 0.0303432f $X=3.43 $Y=0.39 $X2=0
+ $Y2=0
cc_744 N_A_543_47#_c_1033_n A_639_47# 0.0148617f $X=3.43 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_745 N_A_543_47#_c_998_n A_639_47# 0.00606072f $X=3.515 $Y=1.185 $X2=-0.19
+ $Y2=-0.24
cc_746 N_A_1283_21#_c_1137_n N_A_1108_47#_M1013_g 0.0125936f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_747 N_A_1283_21#_c_1139_n N_A_1108_47#_M1013_g 0.00276677f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_748 N_A_1283_21#_c_1126_n N_A_1108_47#_M1001_g 6.19895e-19 $X=7.15 $Y=0.695
+ $X2=0 $Y2=0
cc_749 N_A_1283_21#_c_1166_n N_A_1108_47#_M1001_g 0.0116638f $X=7.815 $Y=0.38
+ $X2=0 $Y2=0
cc_750 N_A_1283_21#_c_1128_n N_A_1108_47#_M1001_g 0.0037075f $X=7.975 $Y=0.82
+ $X2=0 $Y2=0
cc_751 N_A_1283_21#_c_1139_n N_A_1108_47#_M1001_g 0.004469f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_752 N_A_1283_21#_c_1132_n N_A_1108_47#_M1001_g 0.0115506f $X=7.815 $Y=0.82
+ $X2=0 $Y2=0
cc_753 N_A_1283_21#_M1022_g N_A_1108_47#_c_1277_n 0.00955366f $X=6.49 $Y=0.445
+ $X2=0 $Y2=0
cc_754 N_A_1283_21#_c_1126_n N_A_1108_47#_c_1277_n 3.21819e-19 $X=7.15 $Y=0.695
+ $X2=0 $Y2=0
cc_755 N_A_1283_21#_M1007_g N_A_1108_47#_c_1280_n 0.0102686f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_756 N_A_1283_21#_M1022_g N_A_1108_47#_c_1270_n 0.00739655f $X=6.49 $Y=0.445
+ $X2=0 $Y2=0
cc_757 N_A_1283_21#_c_1125_n N_A_1108_47#_c_1270_n 0.0190293f $X=6.79 $Y=0.98
+ $X2=0 $Y2=0
cc_758 N_A_1283_21#_c_1126_n N_A_1108_47#_c_1270_n 0.00468097f $X=7.15 $Y=0.695
+ $X2=0 $Y2=0
cc_759 N_A_1283_21#_c_1131_n N_A_1108_47#_c_1270_n 0.0122822f $X=7.15 $Y=0.78
+ $X2=0 $Y2=0
cc_760 N_A_1283_21#_c_1133_n N_A_1108_47#_c_1270_n 0.0104269f $X=6.695 $Y=0.98
+ $X2=0 $Y2=0
cc_761 N_A_1283_21#_M1007_g N_A_1108_47#_c_1273_n 0.0164997f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_762 N_A_1283_21#_c_1125_n N_A_1108_47#_c_1273_n 0.00480564f $X=6.79 $Y=0.98
+ $X2=0 $Y2=0
cc_763 N_A_1283_21#_c_1133_n N_A_1108_47#_c_1273_n 0.00270124f $X=6.695 $Y=0.98
+ $X2=0 $Y2=0
cc_764 N_A_1283_21#_M1007_g N_A_1108_47#_c_1274_n 0.0114588f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_765 N_A_1283_21#_c_1138_n N_A_1108_47#_c_1274_n 0.00493675f $X=7.53 $Y=2
+ $X2=0 $Y2=0
cc_766 N_A_1283_21#_c_1125_n N_A_1108_47#_c_1275_n 0.00570594f $X=6.79 $Y=0.98
+ $X2=0 $Y2=0
cc_767 N_A_1283_21#_c_1137_n N_A_1108_47#_c_1275_n 0.0202553f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_768 N_A_1283_21#_c_1138_n N_A_1108_47#_c_1275_n 0.0138731f $X=7.53 $Y=2 $X2=0
+ $Y2=0
cc_769 N_A_1283_21#_c_1139_n N_A_1108_47#_c_1275_n 0.0141871f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_770 N_A_1283_21#_c_1132_n N_A_1108_47#_c_1275_n 2.98117e-19 $X=7.815 $Y=0.82
+ $X2=0 $Y2=0
cc_771 N_A_1283_21#_c_1133_n N_A_1108_47#_c_1275_n 8.76062e-19 $X=6.695 $Y=0.98
+ $X2=0 $Y2=0
cc_772 N_A_1283_21#_c_1137_n N_A_1108_47#_c_1276_n 0.00285904f $X=7.99 $Y=2
+ $X2=0 $Y2=0
cc_773 N_A_1283_21#_c_1138_n N_A_1108_47#_c_1276_n 2.53623e-19 $X=7.53 $Y=2
+ $X2=0 $Y2=0
cc_774 N_A_1283_21#_c_1139_n N_A_1108_47#_c_1276_n 0.00684159f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_775 N_A_1283_21#_c_1137_n N_VPWR_M1013_d 0.00225536f $X=7.99 $Y=2 $X2=0 $Y2=0
cc_776 N_A_1283_21#_M1007_g N_VPWR_c_1377_n 0.00383525f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_777 N_A_1283_21#_M1015_g N_VPWR_c_1378_n 8.95466e-19 $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_778 N_A_1283_21#_c_1137_n N_VPWR_c_1378_n 0.021029f $X=7.99 $Y=2 $X2=0 $Y2=0
cc_779 N_A_1283_21#_M1015_g N_VPWR_c_1379_n 0.0284377f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_780 N_A_1283_21#_c_1137_n N_VPWR_c_1379_n 0.0122029f $X=7.99 $Y=2 $X2=0 $Y2=0
cc_781 N_A_1283_21#_c_1139_n N_VPWR_c_1379_n 0.0274877f $X=8.075 $Y=1.915 $X2=0
+ $Y2=0
cc_782 N_A_1283_21#_c_1129_n N_VPWR_c_1379_n 0.0229566f $X=8.645 $Y=1.16 $X2=0
+ $Y2=0
cc_783 N_A_1283_21#_c_1130_n N_VPWR_c_1379_n 0.00320419f $X=8.645 $Y=1.16 $X2=0
+ $Y2=0
cc_784 N_A_1283_21#_M1007_g N_VPWR_c_1382_n 0.00357668f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_785 N_A_1283_21#_c_1230_p N_VPWR_c_1384_n 0.00701792f $X=7.445 $Y=2.21 $X2=0
+ $Y2=0
cc_786 N_A_1283_21#_c_1137_n N_VPWR_c_1384_n 0.00260015f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_787 N_A_1283_21#_c_1137_n N_VPWR_c_1389_n 0.00242671f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_788 N_A_1283_21#_M1015_g N_VPWR_c_1390_n 0.0046653f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_789 N_A_1283_21#_M1016_d N_VPWR_c_1372_n 0.00416801f $X=7.31 $Y=2.065 $X2=0
+ $Y2=0
cc_790 N_A_1283_21#_M1007_g N_VPWR_c_1372_n 0.00559732f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_791 N_A_1283_21#_M1015_g N_VPWR_c_1372_n 0.00895857f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_792 N_A_1283_21#_c_1230_p N_VPWR_c_1372_n 0.00608739f $X=7.445 $Y=2.21 $X2=0
+ $Y2=0
cc_793 N_A_1283_21#_c_1137_n N_VPWR_c_1372_n 0.00960349f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_794 N_A_1283_21#_M1015_g Q 0.00431325f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_795 N_A_1283_21#_c_1129_n Q 0.0266145f $X=8.645 $Y=1.16 $X2=0 $Y2=0
cc_796 N_A_1283_21#_c_1134_n Q 0.0195346f $X=8.657 $Y=0.995 $X2=0 $Y2=0
cc_797 N_A_1283_21#_c_1126_n N_VGND_M1022_d 0.00259202f $X=7.15 $Y=0.695 $X2=0
+ $Y2=0
cc_798 N_A_1283_21#_c_1171_n N_VGND_M1022_d 0.0020638f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_799 N_A_1283_21#_M1022_g N_VGND_c_1609_n 0.00552213f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_800 N_A_1283_21#_c_1126_n N_VGND_c_1609_n 0.0043583f $X=7.15 $Y=0.695 $X2=0
+ $Y2=0
cc_801 N_A_1283_21#_c_1171_n N_VGND_c_1609_n 0.0139352f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_802 N_A_1283_21#_c_1131_n N_VGND_c_1609_n 0.0135486f $X=7.15 $Y=0.78 $X2=0
+ $Y2=0
cc_803 N_A_1283_21#_c_1133_n N_VGND_c_1609_n 0.00108751f $X=6.695 $Y=0.98 $X2=0
+ $Y2=0
cc_804 N_A_1283_21#_c_1127_n N_VGND_c_1610_n 0.0113008f $X=7.975 $Y=0.465 $X2=0
+ $Y2=0
cc_805 N_A_1283_21#_c_1128_n N_VGND_c_1610_n 0.00495943f $X=7.975 $Y=0.82 $X2=0
+ $Y2=0
cc_806 N_A_1283_21#_c_1129_n N_VGND_c_1610_n 0.0109281f $X=8.645 $Y=1.16 $X2=0
+ $Y2=0
cc_807 N_A_1283_21#_c_1130_n N_VGND_c_1610_n 0.00255976f $X=8.645 $Y=1.16 $X2=0
+ $Y2=0
cc_808 N_A_1283_21#_c_1134_n N_VGND_c_1610_n 0.0108863f $X=8.657 $Y=0.995 $X2=0
+ $Y2=0
cc_809 N_A_1283_21#_M1022_g N_VGND_c_1613_n 0.00403211f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_810 N_A_1283_21#_c_1166_n N_VGND_c_1616_n 0.0253037f $X=7.815 $Y=0.38 $X2=0
+ $Y2=0
cc_811 N_A_1283_21#_c_1171_n N_VGND_c_1616_n 0.00758764f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_812 N_A_1283_21#_c_1127_n N_VGND_c_1616_n 0.0178412f $X=7.975 $Y=0.465 $X2=0
+ $Y2=0
cc_813 N_A_1283_21#_c_1131_n N_VGND_c_1616_n 0.00275249f $X=7.15 $Y=0.78 $X2=0
+ $Y2=0
cc_814 N_A_1283_21#_c_1134_n N_VGND_c_1617_n 0.0046653f $X=8.657 $Y=0.995 $X2=0
+ $Y2=0
cc_815 N_A_1283_21#_M1001_d N_VGND_c_1618_n 0.00212393f $X=7.765 $Y=0.235 $X2=0
+ $Y2=0
cc_816 N_A_1283_21#_M1022_g N_VGND_c_1618_n 0.00628912f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_817 N_A_1283_21#_c_1166_n N_VGND_c_1618_n 0.012114f $X=7.815 $Y=0.38 $X2=0
+ $Y2=0
cc_818 N_A_1283_21#_c_1171_n N_VGND_c_1618_n 0.00279545f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_819 N_A_1283_21#_c_1127_n N_VGND_c_1618_n 0.0120802f $X=7.975 $Y=0.465 $X2=0
+ $Y2=0
cc_820 N_A_1283_21#_c_1131_n N_VGND_c_1618_n 0.00245528f $X=7.15 $Y=0.78 $X2=0
+ $Y2=0
cc_821 N_A_1283_21#_c_1133_n N_VGND_c_1618_n 8.11688e-19 $X=6.695 $Y=0.98 $X2=0
+ $Y2=0
cc_822 N_A_1283_21#_c_1134_n N_VGND_c_1618_n 0.00895857f $X=8.657 $Y=0.995 $X2=0
+ $Y2=0
cc_823 N_A_1283_21#_c_1166_n A_1462_47# 0.00399694f $X=7.815 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_824 N_A_1108_47#_M1013_g N_VPWR_c_1377_n 7.45342e-19 $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_825 N_A_1108_47#_c_1280_n N_VPWR_c_1377_n 0.0234228f $X=6.6 $Y=2.295 $X2=0
+ $Y2=0
cc_826 N_A_1108_47#_c_1275_n N_VPWR_c_1377_n 0.00898242f $X=7.655 $Y=1.66 $X2=0
+ $Y2=0
cc_827 N_A_1108_47#_M1013_g N_VPWR_c_1378_n 0.0078865f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_828 N_A_1108_47#_M1013_g N_VPWR_c_1379_n 0.00418219f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_829 N_A_1108_47#_c_1280_n N_VPWR_c_1382_n 0.0505746f $X=6.6 $Y=2.295 $X2=0
+ $Y2=0
cc_830 N_A_1108_47#_M1013_g N_VPWR_c_1384_n 0.00367706f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_831 N_A_1108_47#_M1021_d N_VPWR_c_1372_n 0.00178215f $X=5.92 $Y=2.065 $X2=0
+ $Y2=0
cc_832 N_A_1108_47#_M1013_g N_VPWR_c_1372_n 0.00430058f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_833 N_A_1108_47#_c_1280_n N_VPWR_c_1372_n 0.0242715f $X=6.6 $Y=2.295 $X2=0
+ $Y2=0
cc_834 N_A_1108_47#_c_1280_n A_1270_413# 0.00433468f $X=6.6 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_835 N_A_1108_47#_c_1277_n N_VGND_c_1609_n 0.0213874f $X=6.365 $Y=0.395 $X2=0
+ $Y2=0
cc_836 N_A_1108_47#_M1001_g N_VGND_c_1610_n 0.00268936f $X=7.69 $Y=0.445 $X2=0
+ $Y2=0
cc_837 N_A_1108_47#_c_1277_n N_VGND_c_1613_n 0.0567494f $X=6.365 $Y=0.395 $X2=0
+ $Y2=0
cc_838 N_A_1108_47#_M1001_g N_VGND_c_1616_n 0.00366111f $X=7.69 $Y=0.445 $X2=0
+ $Y2=0
cc_839 N_A_1108_47#_M1020_d N_VGND_c_1618_n 0.00272411f $X=5.54 $Y=0.235 $X2=0
+ $Y2=0
cc_840 N_A_1108_47#_M1001_g N_VGND_c_1618_n 0.00675738f $X=7.69 $Y=0.445 $X2=0
+ $Y2=0
cc_841 N_A_1108_47#_c_1277_n N_VGND_c_1618_n 0.0161501f $X=6.365 $Y=0.395 $X2=0
+ $Y2=0
cc_842 N_A_1108_47#_c_1277_n A_1217_47# 0.00484766f $X=6.365 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_843 N_VPWR_c_1372_n N_A_448_47#_M1024_d 0.00255917f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_844 N_VPWR_c_1374_n N_A_448_47#_c_1520_n 0.00413503f $X=2.015 $Y=2.34 $X2=0
+ $Y2=0
cc_845 N_VPWR_c_1380_n N_A_448_47#_c_1520_n 0.0177638f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_846 N_VPWR_c_1372_n N_A_448_47#_c_1520_n 0.00643929f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_847 N_VPWR_c_1372_n N_A_651_413#_M1006_d 0.00515242f $X=8.97 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_848 N_VPWR_c_1372_n N_A_651_413#_M1027_d 0.00220707f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_849 N_VPWR_c_1380_n N_A_651_413#_c_1554_n 0.0071865f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_850 N_VPWR_c_1372_n N_A_651_413#_c_1554_n 0.00287341f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_851 N_VPWR_c_1375_n N_A_651_413#_c_1555_n 0.0205079f $X=4.155 $Y=2.29 $X2=0
+ $Y2=0
cc_852 N_VPWR_c_1380_n N_A_651_413#_c_1555_n 0.00357601f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_853 N_VPWR_c_1388_n N_A_651_413#_c_1555_n 0.00256078f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_854 N_VPWR_c_1372_n N_A_651_413#_c_1555_n 0.00495172f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_855 N_VPWR_c_1376_n N_A_651_413#_c_1557_n 0.0106232f $X=5.14 $Y=2.34 $X2=0
+ $Y2=0
cc_856 N_VPWR_c_1388_n N_A_651_413#_c_1557_n 0.0071865f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_857 N_VPWR_c_1372_n N_A_651_413#_c_1557_n 0.00287341f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_858 N_VPWR_c_1372_n A_1270_413# 0.00216831f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_859 N_VPWR_c_1372_n N_Q_M1015_d 0.00401809f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_860 N_VPWR_c_1390_n Q 0.00923202f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_861 N_VPWR_c_1372_n Q 0.00900352f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_862 N_A_448_47#_c_1537_n N_VGND_c_1611_n 0.00763796f $X=2.215 $Y=0.39 $X2=0
+ $Y2=0
cc_863 N_A_448_47#_c_1528_n N_VGND_c_1611_n 0.0137117f $X=2.375 $Y=0.39 $X2=0
+ $Y2=0
cc_864 N_A_448_47#_M1025_d N_VGND_c_1618_n 0.00276506f $X=2.24 $Y=0.235 $X2=0
+ $Y2=0
cc_865 N_A_448_47#_c_1537_n N_VGND_c_1618_n 0.00579413f $X=2.215 $Y=0.39 $X2=0
+ $Y2=0
cc_866 N_A_448_47#_c_1528_n N_VGND_c_1618_n 0.0115463f $X=2.375 $Y=0.39 $X2=0
+ $Y2=0
cc_867 Q N_VGND_c_1617_n 0.0165374f $X=8.88 $Y=0.425 $X2=0 $Y2=0
cc_868 N_Q_M1005_d N_VGND_c_1618_n 0.00387432f $X=8.805 $Y=0.235 $X2=0 $Y2=0
cc_869 Q N_VGND_c_1618_n 0.00968619f $X=8.88 $Y=0.425 $X2=0 $Y2=0
cc_870 N_VGND_c_1618_n A_639_47# 0.0110359f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_871 N_VGND_c_1618_n A_805_47# 0.00196925f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_872 N_VGND_c_1618_n A_1217_47# 0.00217995f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_873 N_VGND_c_1618_n A_1462_47# 0.00196947f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__sdlclkp_4.spice
* Created: Thu Aug 27 14:47:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdlclkp_4.pex.spice"
.subckt sky130_fd_sc_hd__sdlclkp_4  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1027 N_VGND_M1027_d N_SCE_M1027_g N_A_27_47#_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1011 N_A_27_47#_M1011_d N_GATE_M1011_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0733385 AS=0.0567 PD=0.813077 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_287_413#_M1007_d N_A_257_147#_M1007_g N_A_27_47#_M1011_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0675 AS=0.0628615 PD=0.735 PS=0.696923 NRD=14.988
+ NRS=19.992 M=1 R=2.4 SA=75001.1 SB=75001.9 A=0.054 P=1.02 MULT=1
MM1022 A_395_47# N_A_257_243#_M1022_g N_A_287_413#_M1007_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0833538 AS=0.0675 PD=0.812308 PS=0.735 NRD=58.836 NRS=16.656 M=1
+ R=2.4 SA=75001.6 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1016 N_VGND_M1016_d N_A_465_315#_M1016_g A_395_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.108042 AS=0.0972462 PD=0.863551 PS=0.947692 NRD=25.704 NRS=50.436 M=1
+ R=2.8 SA=75001.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_465_315#_M1008_d N_A_287_413#_M1008_g N_VGND_M1016_d VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.167208 PD=1.82 PS=1.33645 NRD=0 NRS=14.76 M=1
+ R=4.33333 SA=75001.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A_257_147#_M1020_g N_A_257_243#_M1020_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_257_147#_M1025_d N_CLK_M1025_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_1127_47# N_A_465_315#_M1017_g N_A_1045_47#_M1017_s VNB NSHORT L=0.15
+ W=0.65 AD=0.06825 AS=0.169 PD=0.86 PS=1.82 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_CLK_M1019_g A_1127_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.125125 AS=0.06825 PD=1.035 PS=0.86 NRD=5.532 NRS=9.228 M=1 R=4.33333
+ SA=75000.5 SB=75002 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1019_d N_A_1045_47#_M1003_g N_GCLK_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.125125 AS=0.08775 PD=1.035 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_1045_47#_M1004_g N_GCLK_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1004_d N_A_1045_47#_M1009_g N_GCLK_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_1045_47#_M1015_g N_GCLK_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 A_109_369# N_SCE_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1664 PD=0.85 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_27_47#_M1005_d N_GATE_M1005_g A_109_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.136875 AS=0.0672 PD=1.2317 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667
+ SA=75000.5 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1026 N_A_287_413#_M1026_d N_A_257_243#_M1026_g N_A_27_47#_M1005_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0693 AS=0.0898245 PD=0.75 PS=0.808302 NRD=11.7215
+ NRS=23.443 M=1 R=2.8 SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1010 A_383_413# N_A_257_147#_M1010_g N_A_287_413#_M1026_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.0693 PD=0.86 PS=0.75 NRD=77.3816 NRS=11.7215 M=1 R=2.8
+ SA=75001.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_465_315#_M1023_g A_383_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.108727 AS=0.0924 PD=0.90507 PS=0.86 NRD=70.3487 NRS=77.3816 M=1 R=2.8
+ SA=75002.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1000 N_A_465_315#_M1000_d N_A_287_413#_M1000_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.258873 PD=2.52 PS=2.15493 NRD=0 NRS=19.7 M=1 R=6.66667
+ SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A_257_147#_M1012_g N_A_257_243#_M1012_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.16925 AS=0.1664 PD=1.37 PS=1.8 NRD=64.4584 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_257_147#_M1002_d N_CLK_M1002_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.16925 PD=1.8 PS=1.37 NRD=0 NRS=64.4584 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_A_1045_47#_M1013_d N_A_465_315#_M1013_g N_VPWR_M1013_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_1045_47#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1625 AS=0.135 PD=1.325 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_GCLK_M1001_d N_A_1045_47#_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1625 PD=1.27 PS=1.325 NRD=0 NRS=3.9203 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1018 N_GCLK_M1001_d N_A_1045_47#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1021 N_GCLK_M1021_d N_A_1045_47#_M1021_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1024 N_GCLK_M1021_d N_A_1045_47#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.31 PD=1.27 PS=2.62 NRD=0 NRS=8.8453 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.8993 P=20.53
c_89 VNB 0 5.96947e-20 $X=0.15 $Y=-0.085
c_162 VPB 0 1.88295e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__sdlclkp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o32a_1.pxi.spice
* Created: Tue Sep  1 19:25:42 2020
* 
x_PM_SKY130_FD_SC_HD__O32A_1%A_77_199# N_A_77_199#_M1011_d N_A_77_199#_M1000_d
+ N_A_77_199#_M1009_g N_A_77_199#_M1002_g N_A_77_199#_c_67_n N_A_77_199#_c_73_p
+ N_A_77_199#_c_111_p N_A_77_199#_c_82_p N_A_77_199#_c_83_p N_A_77_199#_c_128_p
+ N_A_77_199#_c_89_p N_A_77_199#_c_129_p N_A_77_199#_c_93_p N_A_77_199#_c_62_n
+ N_A_77_199#_c_63_n N_A_77_199#_c_64_n N_A_77_199#_c_97_p N_A_77_199#_c_65_n
+ PM_SKY130_FD_SC_HD__O32A_1%A_77_199#
x_PM_SKY130_FD_SC_HD__O32A_1%A1 N_A1_M1005_g N_A1_M1010_g A1 N_A1_c_154_n
+ N_A1_c_155_n PM_SKY130_FD_SC_HD__O32A_1%A1
x_PM_SKY130_FD_SC_HD__O32A_1%A2 N_A2_M1008_g N_A2_M1003_g A2 A2 A2 N_A2_c_187_n
+ N_A2_c_188_n PM_SKY130_FD_SC_HD__O32A_1%A2
x_PM_SKY130_FD_SC_HD__O32A_1%A3 N_A3_M1001_g N_A3_M1000_g A3 A3 N_A3_c_224_n
+ N_A3_c_225_n N_A3_c_226_n PM_SKY130_FD_SC_HD__O32A_1%A3
x_PM_SKY130_FD_SC_HD__O32A_1%B2 N_B2_M1011_g N_B2_M1007_g B2 B2 N_B2_c_261_n
+ N_B2_c_262_n N_B2_c_263_n PM_SKY130_FD_SC_HD__O32A_1%B2
x_PM_SKY130_FD_SC_HD__O32A_1%B1 N_B1_c_299_n N_B1_M1006_g N_B1_M1004_g B1
+ N_B1_c_301_n PM_SKY130_FD_SC_HD__O32A_1%B1
x_PM_SKY130_FD_SC_HD__O32A_1%X N_X_M1009_s N_X_M1002_s N_X_c_328_n N_X_c_326_n X
+ X X N_X_c_330_n N_X_c_327_n PM_SKY130_FD_SC_HD__O32A_1%X
x_PM_SKY130_FD_SC_HD__O32A_1%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_352_n
+ N_VPWR_c_353_n N_VPWR_c_354_n VPWR N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_351_n VPWR PM_SKY130_FD_SC_HD__O32A_1%VPWR
x_PM_SKY130_FD_SC_HD__O32A_1%VGND N_VGND_M1009_d N_VGND_M1008_d N_VGND_c_407_n
+ N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n
+ VGND N_VGND_c_413_n N_VGND_c_414_n VGND PM_SKY130_FD_SC_HD__O32A_1%VGND
x_PM_SKY130_FD_SC_HD__O32A_1%A_227_47# N_A_227_47#_M1005_d N_A_227_47#_M1001_d
+ N_A_227_47#_M1006_d N_A_227_47#_c_457_n N_A_227_47#_c_458_n
+ N_A_227_47#_c_452_n N_A_227_47#_c_482_n N_A_227_47#_c_464_n
+ N_A_227_47#_c_451_n PM_SKY130_FD_SC_HD__O32A_1%A_227_47#
cc_1 VNB N_A_77_199#_c_62_n 0.00295064f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=1.835
cc_2 VNB N_A_77_199#_c_63_n 0.00518274f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.16
cc_3 VNB N_A_77_199#_c_64_n 0.026729f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.16
cc_4 VNB N_A_77_199#_c_65_n 0.0197563f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_5 VNB A1 0.00202231f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=0.56
cc_6 VNB N_A1_c_154_n 0.0255876f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.985
cc_7 VNB N_A1_c_155_n 0.0170368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB A2 0.00372928f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=0.56
cc_9 VNB N_A2_c_187_n 0.0243067f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.495
cc_10 VNB N_A2_c_188_n 0.0180721f $X=-0.19 $Y=-0.24 $X2=0.81 $Y2=1.58
cc_11 VNB N_A3_c_224_n 0.023926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A3_c_225_n 0.00304477f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.325
cc_13 VNB N_A3_c_226_n 0.0185641f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.495
cc_14 VNB N_B2_c_261_n 0.0241597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B2_c_262_n 0.00391049f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.325
cc_16 VNB N_B2_c_263_n 0.0186732f $X=-0.19 $Y=-0.24 $X2=0.725 $Y2=1.495
cc_17 VNB N_B1_c_299_n 0.0227545f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=0.235
cc_18 VNB B1 0.0115433f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=0.56
cc_19 VNB N_B1_c_301_n 0.0359229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_326_n 0.0230492f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.325
cc_21 VNB N_X_c_327_n 0.0292838f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=1.96
cc_22 VNB N_VPWR_c_351_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=2.38
cc_23 VNB N_VGND_c_407_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=0.56
cc_24 VNB N_VGND_c_408_n 0.00559947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_409_n 0.0215822f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=1.58
cc_26 VNB N_VGND_c_410_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0.81 $Y2=1.58
cc_27 VNB N_VGND_c_411_n 0.0185558f $X=-0.19 $Y=-0.24 $X2=1.23 $Y2=2.295
cc_28 VNB N_VGND_c_412_n 0.00631415f $X=-0.19 $Y=-0.24 $X2=2.18 $Y2=2.38
cc_29 VNB N_VGND_c_413_n 0.0420839f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=2.38
cc_30 VNB N_VGND_c_414_n 0.201011f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=2.34
cc_31 VNB N_A_227_47#_c_451_n 0.0201726f $X=-0.19 $Y=-0.24 $X2=1.23 $Y2=1.665
cc_32 VPB N_A_77_199#_M1002_g 0.0223975f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.985
cc_33 VPB N_A_77_199#_c_67_n 0.00158251f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.495
cc_34 VPB N_A_77_199#_c_62_n 0.00112837f $X=-0.19 $Y=1.305 $X2=3.05 $Y2=1.835
cc_35 VPB N_A_77_199#_c_63_n 0.00392641f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.16
cc_36 VPB N_A_77_199#_c_64_n 0.00625607f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.16
cc_37 VPB N_A1_M1010_g 0.0197583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB A1 0.00123896f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=0.56
cc_39 VPB N_A1_c_154_n 0.00611554f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.985
cc_40 VPB N_A2_M1003_g 0.0201163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB A2 9.7737e-19 $X=-0.19 $Y=1.305 $X2=0.64 $Y2=0.56
cc_42 VPB N_A2_c_187_n 0.00638193f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.495
cc_43 VPB N_A3_M1000_g 0.0197733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A3_c_224_n 0.00655966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A3_c_225_n 0.00225006f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.325
cc_46 VPB N_B2_M1007_g 0.0199501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_B2_c_261_n 0.00656017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_B2_c_262_n 0.00222996f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.325
cc_49 VPB N_B1_M1004_g 0.0267991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB B1 9.15652e-19 $X=-0.19 $Y=1.305 $X2=0.64 $Y2=0.56
cc_51 VPB N_B1_c_301_n 0.0107316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_328_n 0.00831449f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=0.56
cc_53 VPB N_X_c_326_n 0.00917028f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.325
cc_54 VPB N_X_c_330_n 0.034282f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=1.665
cc_55 VPB N_VPWR_c_352_n 0.00258113f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.985
cc_56 VPB N_VPWR_c_353_n 0.0104645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_354_n 0.0437601f $X=-0.19 $Y=1.305 $X2=0.725 $Y2=1.495
cc_58 VPB N_VPWR_c_355_n 0.0581678f $X=-0.19 $Y=1.305 $X2=1.315 $Y2=2.38
cc_59 VPB N_VPWR_c_356_n 0.0236706f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.16
cc_60 VPB N_VPWR_c_351_n 0.0439941f $X=-0.19 $Y=1.305 $X2=2.345 $Y2=2.38
cc_61 N_A_77_199#_M1002_g N_A1_M1010_g 0.0277968f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_77_199#_c_67_n N_A1_M1010_g 0.00173273f $X=0.725 $Y=1.495 $X2=0 $Y2=0
cc_63 N_A_77_199#_c_73_p N_A1_M1010_g 0.015118f $X=1.145 $Y=1.58 $X2=0 $Y2=0
cc_64 N_A_77_199#_c_73_p A1 0.0165948f $X=1.145 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_77_199#_c_63_n A1 0.0207441f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_77_199#_c_64_n A1 4.93181e-19 $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_77_199#_c_73_p N_A1_c_154_n 0.00199381f $X=1.145 $Y=1.58 $X2=0 $Y2=0
cc_68 N_A_77_199#_c_63_n N_A1_c_154_n 0.00194569f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_77_199#_c_64_n N_A1_c_154_n 0.0205298f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_77_199#_c_65_n N_A1_c_155_n 0.0258937f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_77_199#_c_73_p N_A2_M1003_g 0.00121534f $X=1.145 $Y=1.58 $X2=0 $Y2=0
cc_72 N_A_77_199#_c_82_p N_A2_M1003_g 0.00657261f $X=1.23 $Y=2.295 $X2=0 $Y2=0
cc_73 N_A_77_199#_c_83_p N_A2_M1003_g 0.0108688f $X=2.18 $Y=2.38 $X2=0 $Y2=0
cc_74 N_A_77_199#_c_67_n A2 0.00435198f $X=0.725 $Y=1.495 $X2=0 $Y2=0
cc_75 N_A_77_199#_c_73_p A2 0.0140153f $X=1.145 $Y=1.58 $X2=0 $Y2=0
cc_76 N_A_77_199#_c_82_p A2 0.0338885f $X=1.23 $Y=2.295 $X2=0 $Y2=0
cc_77 N_A_77_199#_c_83_p A2 0.0196403f $X=2.18 $Y=2.38 $X2=0 $Y2=0
cc_78 N_A_77_199#_c_83_p N_A3_M1000_g 0.0103511f $X=2.18 $Y=2.38 $X2=0 $Y2=0
cc_79 N_A_77_199#_c_89_p N_A3_c_224_n 0.0027136f $X=2.345 $Y=2.085 $X2=0 $Y2=0
cc_80 N_A_77_199#_M1000_d N_A3_c_225_n 0.00207764f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_81 N_A_77_199#_c_83_p N_A3_c_225_n 0.00378901f $X=2.18 $Y=2.38 $X2=0 $Y2=0
cc_82 N_A_77_199#_c_89_p N_A3_c_225_n 0.003678f $X=2.345 $Y=2.085 $X2=0 $Y2=0
cc_83 N_A_77_199#_c_93_p N_B2_M1007_g 0.0162959f $X=2.965 $Y=1.96 $X2=0 $Y2=0
cc_84 N_A_77_199#_c_62_n N_B2_M1007_g 0.00430806f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_85 N_A_77_199#_c_93_p N_B2_c_261_n 0.00249924f $X=2.965 $Y=1.96 $X2=0 $Y2=0
cc_86 N_A_77_199#_c_62_n N_B2_c_261_n 0.0021494f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_87 N_A_77_199#_c_97_p N_B2_c_261_n 0.00358227f $X=3.05 $Y=0.73 $X2=0 $Y2=0
cc_88 N_A_77_199#_M1000_d N_B2_c_262_n 0.00214305f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_89 N_A_77_199#_c_89_p N_B2_c_262_n 0.00411586f $X=2.345 $Y=2.085 $X2=0 $Y2=0
cc_90 N_A_77_199#_c_93_p N_B2_c_262_n 0.0148725f $X=2.965 $Y=1.96 $X2=0 $Y2=0
cc_91 N_A_77_199#_c_62_n N_B2_c_262_n 0.0511464f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_92 N_A_77_199#_c_97_p N_B2_c_262_n 0.00508417f $X=3.05 $Y=0.73 $X2=0 $Y2=0
cc_93 N_A_77_199#_c_62_n N_B2_c_263_n 0.00306945f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_94 N_A_77_199#_c_62_n N_B1_c_299_n 0.00863988f $X=3.05 $Y=1.835 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_77_199#_c_97_p N_B1_c_299_n 0.00833006f $X=3.05 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_77_199#_c_93_p N_B1_M1004_g 0.00733449f $X=2.965 $Y=1.96 $X2=0 $Y2=0
cc_97 N_A_77_199#_c_62_n N_B1_M1004_g 0.0156338f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_98 N_A_77_199#_c_62_n B1 0.0216779f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_99 N_A_77_199#_c_62_n N_B1_c_301_n 0.00753027f $X=3.05 $Y=1.835 $X2=0 $Y2=0
cc_100 N_A_77_199#_M1002_g N_X_c_328_n 0.00841572f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_77_199#_c_111_p N_X_c_328_n 0.0141598f $X=0.81 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_77_199#_c_63_n N_X_c_328_n 0.00199187f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_77_199#_c_64_n N_X_c_328_n 0.00199986f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_77_199#_M1002_g N_X_c_326_n 0.00216353f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_77_199#_c_67_n N_X_c_326_n 0.00471102f $X=0.725 $Y=1.495 $X2=0 $Y2=0
cc_106 N_A_77_199#_c_63_n N_X_c_326_n 0.0233364f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_77_199#_c_64_n N_X_c_326_n 0.00786683f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_77_199#_c_65_n N_X_c_326_n 0.00340798f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_77_199#_c_63_n N_X_c_327_n 0.00956978f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_77_199#_c_64_n N_X_c_327_n 0.00254615f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_77_199#_c_65_n N_X_c_327_n 0.00794233f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_77_199#_c_73_p N_VPWR_M1002_d 0.00559347f $X=1.145 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_77_199#_c_111_p N_VPWR_M1002_d 4.07682e-19 $X=0.81 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_77_199#_M1002_g N_VPWR_c_352_n 0.0137346f $X=0.64 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_77_199#_c_73_p N_VPWR_c_352_n 0.00956383f $X=1.145 $Y=1.58 $X2=0
+ $Y2=0
cc_116 N_A_77_199#_c_111_p N_VPWR_c_352_n 0.00573263f $X=0.81 $Y=1.58 $X2=0
+ $Y2=0
cc_117 N_A_77_199#_c_83_p N_VPWR_c_355_n 0.048705f $X=2.18 $Y=2.38 $X2=0 $Y2=0
cc_118 N_A_77_199#_c_128_p N_VPWR_c_355_n 0.0103171f $X=1.315 $Y=2.38 $X2=0
+ $Y2=0
cc_119 N_A_77_199#_c_129_p N_VPWR_c_355_n 0.0212162f $X=2.345 $Y=2.295 $X2=0
+ $Y2=0
cc_120 N_A_77_199#_c_93_p N_VPWR_c_355_n 0.00991715f $X=2.965 $Y=1.96 $X2=0
+ $Y2=0
cc_121 N_A_77_199#_M1002_g N_VPWR_c_356_n 0.0046653f $X=0.64 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_77_199#_M1000_d N_VPWR_c_351_n 0.00325134f $X=2.155 $Y=1.485 $X2=0
+ $Y2=0
cc_123 N_A_77_199#_M1002_g N_VPWR_c_351_n 0.00897386f $X=0.64 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_77_199#_c_83_p N_VPWR_c_351_n 0.0307752f $X=2.18 $Y=2.38 $X2=0 $Y2=0
cc_125 N_A_77_199#_c_128_p N_VPWR_c_351_n 0.006547f $X=1.315 $Y=2.38 $X2=0 $Y2=0
cc_126 N_A_77_199#_c_129_p N_VPWR_c_351_n 0.0126835f $X=2.345 $Y=2.295 $X2=0
+ $Y2=0
cc_127 N_A_77_199#_c_93_p N_VPWR_c_351_n 0.0172698f $X=2.965 $Y=1.96 $X2=0 $Y2=0
cc_128 N_A_77_199#_c_73_p A_227_297# 0.0033478f $X=1.145 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A_77_199#_c_82_p A_227_297# 0.00838463f $X=1.23 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_77_199#_c_83_p A_227_297# 0.00437438f $X=2.18 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_77_199#_c_128_p A_227_297# 0.00207796f $X=1.315 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A_77_199#_c_83_p A_323_297# 0.00963114f $X=2.18 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_77_199#_c_93_p A_539_297# 0.0112172f $X=2.965 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_77_199#_c_62_n A_539_297# 0.00370082f $X=3.05 $Y=1.835 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_77_199#_c_63_n N_VGND_c_407_n 0.00191725f $X=0.55 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_77_199#_c_65_n N_VGND_c_407_n 0.00297551f $X=0.55 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_A_77_199#_c_65_n N_VGND_c_409_n 0.00541359f $X=0.55 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_77_199#_M1011_d N_VGND_c_414_n 0.00330106f $X=2.695 $Y=0.235 $X2=0
+ $Y2=0
cc_139 N_A_77_199#_c_65_n N_VGND_c_414_n 0.0106108f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_77_199#_c_73_p N_A_227_47#_c_452_n 0.00188857f $X=1.145 $Y=1.58 $X2=0
+ $Y2=0
cc_141 N_A_77_199#_M1011_d N_A_227_47#_c_451_n 0.00641276f $X=2.695 $Y=0.235
+ $X2=0 $Y2=0
cc_142 N_A_77_199#_c_97_p N_A_227_47#_c_451_n 0.0228904f $X=3.05 $Y=0.73 $X2=0
+ $Y2=0
cc_143 N_A1_M1010_g N_A2_M1003_g 0.0404118f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_144 A1 A2 0.0193908f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A1_c_154_n A2 6.11112e-19 $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A1_M1010_g A2 9.70262e-19 $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_147 A1 N_A2_c_187_n 0.00112156f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A1_c_154_n N_A2_c_187_n 0.0206718f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A1_c_155_n N_A2_c_188_n 0.0102221f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A1_c_155_n N_X_c_327_n 6.48273e-19 $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_M1010_g N_VPWR_c_352_n 0.00306721f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1010_g N_VPWR_c_355_n 0.00585385f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A1_M1010_g N_VPWR_c_351_n 0.0107141f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A1_c_154_n N_VGND_c_407_n 2.1041e-19 $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A1_c_155_n N_VGND_c_407_n 0.00297551f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A1_c_155_n N_VGND_c_411_n 0.00585385f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A1_c_155_n N_VGND_c_414_n 0.0107321f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_158 A1 N_A_227_47#_c_452_n 0.00420581f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A1_c_154_n N_A_227_47#_c_452_n 0.00187805f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_M1003_g N_A3_M1000_g 0.0365515f $X=1.54 $Y=1.985 $X2=0 $Y2=0
cc_161 A2 N_A3_M1000_g 0.0079345f $X=1.52 $Y=1.445 $X2=0 $Y2=0
cc_162 A2 N_A3_c_224_n 0.00111813f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A2_c_187_n N_A3_c_224_n 0.0214125f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A2_M1003_g N_A3_c_225_n 4.96581e-19 $X=1.54 $Y=1.985 $X2=0 $Y2=0
cc_165 A2 N_A3_c_225_n 0.0472313f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A2_c_187_n N_A3_c_225_n 0.00101459f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A2_c_188_n N_A3_c_226_n 0.0179959f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VPWR_c_355_n 0.00357877f $X=1.54 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A2_M1003_g N_VPWR_c_351_n 0.00574349f $X=1.54 $Y=1.985 $X2=0 $Y2=0
cc_170 A2 A_323_297# 0.00912089f $X=1.52 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_171 N_A2_c_188_n N_VGND_c_408_n 0.00317203f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_188_n N_VGND_c_411_n 0.00427194f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_188_n N_VGND_c_414_n 0.0060737f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_c_188_n N_A_227_47#_c_457_n 0.00518889f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_175 A2 N_A_227_47#_c_458_n 0.0241781f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A2_c_187_n N_A_227_47#_c_458_n 0.00114453f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A2_c_188_n N_A_227_47#_c_458_n 0.0101481f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A3_M1000_g N_B2_M1007_g 0.028111f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A3_c_225_n N_B2_M1007_g 9.88057e-19 $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A3_c_224_n N_B2_c_261_n 0.0204569f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A3_c_225_n N_B2_c_261_n 2.99585e-19 $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A3_M1000_g N_B2_c_262_n 0.00104212f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A3_c_224_n N_B2_c_262_n 0.00221537f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A3_c_225_n N_B2_c_262_n 0.0498586f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A3_c_226_n N_B2_c_263_n 0.0167992f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A3_M1000_g N_VPWR_c_355_n 0.00357877f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A3_M1000_g N_VPWR_c_351_n 0.00582422f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A3_c_226_n N_VGND_c_408_n 0.00317203f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A3_c_226_n N_VGND_c_413_n 0.00428022f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A3_c_226_n N_VGND_c_414_n 0.00630832f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A3_c_226_n N_A_227_47#_c_457_n 5.97614e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A3_c_225_n N_A_227_47#_c_458_n 0.0148298f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A3_c_226_n N_A_227_47#_c_458_n 0.0128054f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A3_c_224_n N_A_227_47#_c_464_n 0.00383363f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A3_c_225_n N_A_227_47#_c_464_n 0.00370042f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B2_c_263_n N_B1_c_299_n 0.0195459f $X=2.71 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_197 N_B2_M1007_g N_B1_M1004_g 0.034815f $X=2.62 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B2_c_262_n N_B1_M1004_g 9.43742e-19 $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B2_c_261_n N_B1_c_301_n 0.0182038f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B2_c_262_n N_B1_c_301_n 2.82126e-19 $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B2_M1007_g N_VPWR_c_355_n 0.00425094f $X=2.62 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B2_M1007_g N_VPWR_c_351_n 0.00652788f $X=2.62 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B2_c_262_n A_539_297# 0.00205228f $X=2.71 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_204 N_B2_c_263_n N_VGND_c_413_n 0.00357877f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B2_c_263_n N_VGND_c_414_n 0.00586478f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B2_c_262_n N_A_227_47#_c_464_n 0.00668657f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B2_c_262_n N_A_227_47#_c_451_n 0.0048873f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B2_c_263_n N_A_227_47#_c_451_n 0.0112784f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B1_M1004_g N_VPWR_c_354_n 0.0045387f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_210 B1 N_VPWR_c_354_n 0.022812f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_211 N_B1_c_301_n N_VPWR_c_354_n 0.00630094f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B1_M1004_g N_VPWR_c_355_n 0.00553297f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1004_g N_VPWR_c_351_n 0.0109531f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_c_299_n N_VGND_c_413_n 0.00357877f $X=3.18 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_299_n N_VGND_c_414_n 0.00654364f $X=3.18 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_299_n N_A_227_47#_c_451_n 0.0132315f $X=3.18 $Y=0.995 $X2=0 $Y2=0
cc_217 B1 N_A_227_47#_c_451_n 0.016123f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_218 N_B1_c_301_n N_A_227_47#_c_451_n 0.00589395f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_219 N_X_c_330_n N_VPWR_c_352_n 0.0402863f $X=0.385 $Y=1.76 $X2=0 $Y2=0
cc_220 N_X_c_330_n N_VPWR_c_356_n 0.0255041f $X=0.385 $Y=1.76 $X2=0 $Y2=0
cc_221 N_X_M1002_s N_VPWR_c_351_n 0.00600901f $X=0.23 $Y=1.485 $X2=0 $Y2=0
cc_222 N_X_c_330_n N_VPWR_c_351_n 0.0146803f $X=0.385 $Y=1.76 $X2=0 $Y2=0
cc_223 N_X_c_327_n N_VGND_c_409_n 0.0336937f $X=0.43 $Y=0.38 $X2=0 $Y2=0
cc_224 N_X_M1009_s N_VGND_c_414_n 0.00209319f $X=0.305 $Y=0.235 $X2=0 $Y2=0
cc_225 N_X_c_327_n N_VGND_c_414_n 0.0193004f $X=0.43 $Y=0.38 $X2=0 $Y2=0
cc_226 N_VPWR_c_351_n A_227_297# 0.00299717f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_227 N_VPWR_c_351_n A_323_297# 0.00313203f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_228 N_VPWR_c_351_n A_539_297# 0.00479441f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_229 N_VGND_c_414_n N_A_227_47#_M1005_d 0.00280738f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_230 N_VGND_c_414_n N_A_227_47#_M1001_d 0.0033081f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_c_414_n N_A_227_47#_M1006_d 0.00233918f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_411_n N_A_227_47#_c_457_n 0.0190643f $X=1.645 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_414_n N_A_227_47#_c_457_n 0.0124836f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_M1008_d N_A_227_47#_c_458_n 0.00957641f $X=1.615 $Y=0.235 $X2=0
+ $Y2=0
cc_235 N_VGND_c_408_n N_A_227_47#_c_458_n 0.0211878f $X=1.81 $Y=0.38 $X2=0 $Y2=0
cc_236 N_VGND_c_411_n N_A_227_47#_c_458_n 0.00252892f $X=1.645 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_413_n N_A_227_47#_c_458_n 0.00312413f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_414_n N_A_227_47#_c_458_n 0.0112698f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_413_n N_A_227_47#_c_482_n 0.0210761f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_414_n N_A_227_47#_c_482_n 0.0126406f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_413_n N_A_227_47#_c_451_n 0.0633699f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_414_n N_A_227_47#_c_451_n 0.0381765f $X=3.45 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__and3b_4.spice.SKY130_FD_SC_HD__AND3B_4.pxi
* Created: Thu Aug 27 14:08:13 2020
* 
x_PM_SKY130_FD_SC_HD__AND3B_4%A_98_199# N_A_98_199#_M1002_d N_A_98_199#_M1009_d
+ N_A_98_199#_M1010_g N_A_98_199#_M1007_g N_A_98_199#_c_80_n N_A_98_199#_c_87_p
+ N_A_98_199#_c_112_p N_A_98_199#_c_81_n N_A_98_199#_c_75_n N_A_98_199#_c_76_n
+ N_A_98_199#_c_77_n N_A_98_199#_c_78_n PM_SKY130_FD_SC_HD__AND3B_4%A_98_199#
x_PM_SKY130_FD_SC_HD__AND3B_4%B N_B_M1001_g N_B_M1000_g B B N_B_c_157_n
+ N_B_c_158_n PM_SKY130_FD_SC_HD__AND3B_4%B
x_PM_SKY130_FD_SC_HD__AND3B_4%C N_C_M1011_g N_C_M1006_g C N_C_c_198_n
+ N_C_c_199_n PM_SKY130_FD_SC_HD__AND3B_4%C
x_PM_SKY130_FD_SC_HD__AND3B_4%A_56_297# N_A_56_297#_M1010_s N_A_56_297#_M1007_s
+ N_A_56_297#_M1000_d N_A_56_297#_c_237_n N_A_56_297#_M1004_g
+ N_A_56_297#_M1003_g N_A_56_297#_c_238_n N_A_56_297#_M1005_g
+ N_A_56_297#_M1008_g N_A_56_297#_c_239_n N_A_56_297#_M1012_g
+ N_A_56_297#_M1013_g N_A_56_297#_c_240_n N_A_56_297#_M1014_g
+ N_A_56_297#_M1015_g N_A_56_297#_c_261_n N_A_56_297#_c_263_n
+ N_A_56_297#_c_294_n N_A_56_297#_c_241_n N_A_56_297#_c_250_n
+ N_A_56_297#_c_251_n N_A_56_297#_c_242_n N_A_56_297#_c_252_n
+ N_A_56_297#_c_243_n N_A_56_297#_c_286_n N_A_56_297#_c_244_n
+ N_A_56_297#_c_245_n PM_SKY130_FD_SC_HD__AND3B_4%A_56_297#
x_PM_SKY130_FD_SC_HD__AND3B_4%A_N N_A_N_M1002_g N_A_N_M1009_g A_N A_N
+ N_A_N_c_384_n N_A_N_c_385_n N_A_N_c_388_n PM_SKY130_FD_SC_HD__AND3B_4%A_N
x_PM_SKY130_FD_SC_HD__AND3B_4%VPWR N_VPWR_M1007_d N_VPWR_M1006_d N_VPWR_M1008_s
+ N_VPWR_M1015_s N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_418_n
+ N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ N_VPWR_c_424_n N_VPWR_c_425_n VPWR N_VPWR_c_426_n N_VPWR_c_414_n
+ PM_SKY130_FD_SC_HD__AND3B_4%VPWR
x_PM_SKY130_FD_SC_HD__AND3B_4%X N_X_M1004_s N_X_M1012_s N_X_M1003_d N_X_M1013_d
+ N_X_c_490_n N_X_c_497_n N_X_c_523_p N_X_c_500_n X X
+ PM_SKY130_FD_SC_HD__AND3B_4%X
x_PM_SKY130_FD_SC_HD__AND3B_4%VGND N_VGND_M1011_d N_VGND_M1005_d N_VGND_M1014_d
+ N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n N_VGND_c_540_n N_VGND_c_541_n
+ N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n N_VGND_c_545_n VGND
+ N_VGND_c_546_n N_VGND_c_547_n PM_SKY130_FD_SC_HD__AND3B_4%VGND
cc_1 VNB N_A_98_199#_c_75_n 0.043058f $X=-0.19 $Y=-0.24 $X2=4.25 $Y2=0.59
cc_2 VNB N_A_98_199#_c_76_n 0.0221176f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_3 VNB N_A_98_199#_c_77_n 0.00309103f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=1.16
cc_4 VNB N_A_98_199#_c_78_n 0.0205132f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=0.995
cc_5 VNB B 0.00113869f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.56
cc_6 VNB N_B_c_157_n 0.0253802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_158_n 0.0163589f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=1.875
cc_8 VNB C 4.72612e-19 $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.56
cc_9 VNB N_C_c_198_n 0.0236109f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.985
cc_10 VNB N_C_c_199_n 0.01733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_56_297#_c_237_n 0.0167541f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.325
cc_12 VNB N_A_56_297#_c_238_n 0.0159963f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=1.99
cc_13 VNB N_A_56_297#_c_239_n 0.01598f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_14 VNB N_A_56_297#_c_240_n 0.0161419f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=0.995
cc_15 VNB N_A_56_297#_c_241_n 0.00133518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_56_297#_c_242_n 0.0257406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_56_297#_c_243_n 0.0245998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_56_297#_c_244_n 0.00188394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_56_297#_c_245_n 0.0627956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB A_N 0.00260728f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.995
cc_21 VNB N_A_N_c_384_n 0.0233327f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.985
cc_22 VNB N_A_N_c_385_n 0.0359603f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=1.325
cc_23 VNB N_VPWR_c_414_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB X 0.00382293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_537_n 0.00278435f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.985
cc_26 VNB N_VGND_c_538_n 3.10008e-19 $X=-0.19 $Y=-0.24 $X2=4.165 $Y2=1.99
cc_27 VNB N_VGND_c_539_n 0.00507182f $X=-0.19 $Y=-0.24 $X2=4.25 $Y2=0.59
cc_28 VNB N_VGND_c_540_n 0.0458115f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_29 VNB N_VGND_c_541_n 0.00512961f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_30 VNB N_VGND_c_542_n 0.0129643f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=1.16
cc_31 VNB N_VGND_c_543_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_544_n 0.01135f $X=-0.19 $Y=-0.24 $X2=4.18 $Y2=2.02
cc_33 VNB N_VGND_c_545_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_34 VNB N_VGND_c_546_n 0.0238808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_547_n 0.251677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_98_199#_M1007_g 0.023375f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.985
cc_37 VPB N_A_98_199#_c_80_n 0.00187533f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.875
cc_38 VPB N_A_98_199#_c_81_n 0.0119273f $X=-0.19 $Y=1.305 $X2=4.305 $Y2=1.875
cc_39 VPB N_A_98_199#_c_75_n 0.0281636f $X=-0.19 $Y=1.305 $X2=4.25 $Y2=0.59
cc_40 VPB N_A_98_199#_c_76_n 0.00684183f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_41 VPB N_A_98_199#_c_77_n 3.66935e-19 $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.16
cc_42 VPB N_B_M1000_g 0.0201191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB B 0.00185118f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.56
cc_44 VPB N_B_c_157_n 0.00618893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_C_M1006_g 0.02026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB C 6.75502e-19 $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.56
cc_47 VPB N_C_c_198_n 0.00451012f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.985
cc_48 VPB N_A_56_297#_M1003_g 0.0196305f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.875
cc_49 VPB N_A_56_297#_M1008_g 0.01823f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_50 VPB N_A_56_297#_M1013_g 0.0181342f $X=-0.19 $Y=1.305 $X2=4.18 $Y2=2.02
cc_51 VPB N_A_56_297#_M1015_g 0.0180492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_56_297#_c_250_n 0.00237981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_56_297#_c_251_n 0.00548881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_56_297#_c_252_n 0.029929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_56_297#_c_243_n 0.0094258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_56_297#_c_244_n 9.37008e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_56_297#_c_245_n 0.0118258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB A_N 0.00182169f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.995
cc_59 VPB N_A_N_c_384_n 0.00484838f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.985
cc_60 VPB N_A_N_c_388_n 0.064139f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.875
cc_61 VPB N_VPWR_c_415_n 0.00431378f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.875
cc_62 VPB N_VPWR_c_416_n 3.15142e-19 $X=-0.19 $Y=1.305 $X2=4.305 $Y2=0.59
cc_63 VPB N_VPWR_c_417_n 0.00515801f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_64 VPB N_VPWR_c_418_n 0.0065666f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=1.16
cc_65 VPB N_VPWR_c_419_n 0.0222531f $X=-0.19 $Y=1.305 $X2=4.18 $Y2=2.02
cc_66 VPB N_VPWR_c_420_n 0.0142875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_421_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_422_n 0.0144022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_423_n 0.00442675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_424_n 0.0121314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_425_n 0.00510002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_426_n 0.0236527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_414_n 0.0546906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB X 0.00271146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 N_A_98_199#_M1007_g N_B_M1000_g 0.0336723f $X=0.685 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_98_199#_c_80_n N_B_M1000_g 0.00818788f $X=0.765 $Y=1.875 $X2=0 $Y2=0
cc_77 N_A_98_199#_c_87_p N_B_M1000_g 0.0170691f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_78 N_A_98_199#_c_80_n B 0.0011498f $X=0.765 $Y=1.875 $X2=0 $Y2=0
cc_79 N_A_98_199#_c_87_p B 0.00626283f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_80 N_A_98_199#_c_76_n B 3.17854e-19 $X=0.625 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_98_199#_c_77_n B 0.0251693f $X=0.765 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_98_199#_c_78_n B 0.00301f $X=0.625 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_98_199#_c_87_p N_B_c_157_n 0.00175888f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_84 N_A_98_199#_c_76_n N_B_c_157_n 0.020415f $X=0.625 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_98_199#_c_77_n N_B_c_157_n 0.00201929f $X=0.765 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_98_199#_c_78_n N_B_c_158_n 0.0274219f $X=0.625 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_98_199#_c_87_p N_C_M1006_g 0.0147309f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_88 N_A_98_199#_c_87_p N_A_56_297#_M1000_d 0.005195f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_89 N_A_98_199#_c_87_p N_A_56_297#_M1003_g 0.0162473f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_90 N_A_98_199#_c_87_p N_A_56_297#_M1008_g 0.0137723f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_91 N_A_98_199#_c_87_p N_A_56_297#_M1013_g 0.0137329f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_92 N_A_98_199#_c_87_p N_A_56_297#_M1015_g 0.0143721f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_93 N_A_98_199#_c_77_n N_A_56_297#_c_261_n 0.0065964f $X=0.765 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_A_98_199#_c_78_n N_A_56_297#_c_261_n 0.010114f $X=0.625 $Y=0.995 $X2=0
+ $Y2=0
cc_95 N_A_98_199#_c_80_n N_A_56_297#_c_263_n 0.00641447f $X=0.765 $Y=1.875 $X2=0
+ $Y2=0
cc_96 N_A_98_199#_c_87_p N_A_56_297#_c_263_n 0.0417797f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_97 N_A_98_199#_c_87_p N_A_56_297#_c_251_n 0.00320895f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_98 N_A_98_199#_c_76_n N_A_56_297#_c_242_n 0.00353092f $X=0.625 $Y=1.16 $X2=0
+ $Y2=0
cc_99 N_A_98_199#_c_77_n N_A_56_297#_c_242_n 0.00461803f $X=0.765 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_98_199#_c_78_n N_A_56_297#_c_242_n 0.00851654f $X=0.625 $Y=0.995
+ $X2=0 $Y2=0
cc_101 N_A_98_199#_c_80_n N_A_56_297#_c_252_n 0.0282418f $X=0.765 $Y=1.875 $X2=0
+ $Y2=0
cc_102 N_A_98_199#_c_112_p N_A_56_297#_c_252_n 0.0190738f $X=0.85 $Y=1.99 $X2=0
+ $Y2=0
cc_103 N_A_98_199#_c_76_n N_A_56_297#_c_252_n 8.36899e-19 $X=0.625 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_98_199#_M1007_g N_A_56_297#_c_243_n 0.00228542f $X=0.685 $Y=1.985
+ $X2=0 $Y2=0
cc_105 N_A_98_199#_c_80_n N_A_56_297#_c_243_n 0.00558849f $X=0.765 $Y=1.875
+ $X2=0 $Y2=0
cc_106 N_A_98_199#_c_76_n N_A_56_297#_c_243_n 0.00758799f $X=0.625 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_98_199#_c_77_n N_A_56_297#_c_243_n 0.0251492f $X=0.765 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_98_199#_c_78_n N_A_56_297#_c_243_n 0.00261927f $X=0.625 $Y=0.995
+ $X2=0 $Y2=0
cc_109 N_A_98_199#_c_87_p N_A_56_297#_c_244_n 0.00152815f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_110 N_A_98_199#_c_87_p A_N 0.0204984f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_111 N_A_98_199#_c_75_n A_N 0.0836589f $X=4.25 $Y=0.59 $X2=0 $Y2=0
cc_112 N_A_98_199#_c_87_p N_A_N_c_384_n 3.40975e-19 $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_113 N_A_98_199#_c_75_n N_A_N_c_385_n 0.0356302f $X=4.25 $Y=0.59 $X2=0 $Y2=0
cc_114 N_A_98_199#_c_87_p N_A_N_c_388_n 0.0132599f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_115 N_A_98_199#_c_80_n N_VPWR_M1007_d 0.00497821f $X=0.765 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_98_199#_c_87_p N_VPWR_M1007_d 0.0090055f $X=4.165 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_117 N_A_98_199#_c_112_p N_VPWR_M1007_d 3.39327e-19 $X=0.85 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_98_199#_c_87_p N_VPWR_M1006_d 0.00511822f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_119 N_A_98_199#_c_87_p N_VPWR_M1008_s 0.00318728f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_120 N_A_98_199#_c_87_p N_VPWR_M1015_s 0.00881898f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_121 N_A_98_199#_c_87_p N_VPWR_c_415_n 0.0186333f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_122 N_A_98_199#_c_87_p N_VPWR_c_416_n 0.016541f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_123 N_A_98_199#_c_87_p N_VPWR_c_417_n 0.020792f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_124 N_A_98_199#_M1007_g N_VPWR_c_418_n 0.0181782f $X=0.685 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_98_199#_c_87_p N_VPWR_c_418_n 0.0207388f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_126 N_A_98_199#_c_112_p N_VPWR_c_418_n 0.00500121f $X=0.85 $Y=1.99 $X2=0
+ $Y2=0
cc_127 N_A_98_199#_M1007_g N_VPWR_c_419_n 0.00413833f $X=0.685 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_98_199#_c_112_p N_VPWR_c_419_n 9.32307e-19 $X=0.85 $Y=1.99 $X2=0
+ $Y2=0
cc_129 N_A_98_199#_c_87_p N_VPWR_c_420_n 0.0091985f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_130 N_A_98_199#_c_87_p N_VPWR_c_422_n 0.00922778f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_131 N_A_98_199#_c_87_p N_VPWR_c_424_n 0.00853679f $X=4.165 $Y=1.99 $X2=0
+ $Y2=0
cc_132 N_A_98_199#_c_87_p N_VPWR_c_426_n 0.0050207f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_133 N_A_98_199#_c_81_n N_VPWR_c_426_n 0.00575061f $X=4.305 $Y=1.875 $X2=0
+ $Y2=0
cc_134 N_A_98_199#_M1007_g N_VPWR_c_414_n 0.00742155f $X=0.685 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_98_199#_c_87_p N_VPWR_c_414_n 0.0595978f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_136 N_A_98_199#_c_112_p N_VPWR_c_414_n 0.00191171f $X=0.85 $Y=1.99 $X2=0
+ $Y2=0
cc_137 N_A_98_199#_c_81_n N_VPWR_c_414_n 0.00853444f $X=4.305 $Y=1.875 $X2=0
+ $Y2=0
cc_138 N_A_98_199#_c_87_p N_X_M1003_d 0.00480695f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_139 N_A_98_199#_c_87_p N_X_M1013_d 0.00452678f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_140 N_A_98_199#_c_87_p N_X_c_490_n 0.0707751f $X=4.165 $Y=1.99 $X2=0 $Y2=0
cc_141 N_A_98_199#_c_75_n N_VGND_c_539_n 0.00103608f $X=4.25 $Y=0.59 $X2=0 $Y2=0
cc_142 N_A_98_199#_c_78_n N_VGND_c_540_n 0.00376052f $X=0.625 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_98_199#_c_75_n N_VGND_c_546_n 0.00953624f $X=4.25 $Y=0.59 $X2=0 $Y2=0
cc_144 N_A_98_199#_c_75_n N_VGND_c_547_n 0.0097021f $X=4.25 $Y=0.59 $X2=0 $Y2=0
cc_145 N_A_98_199#_c_78_n N_VGND_c_547_n 0.00665195f $X=0.625 $Y=0.995 $X2=0
+ $Y2=0
cc_146 N_B_M1000_g N_C_M1006_g 0.0418145f $X=1.21 $Y=1.985 $X2=0 $Y2=0
cc_147 B C 0.0157056f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_148 N_B_c_157_n C 0.00113253f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_149 B N_C_c_198_n 0.00105289f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_150 N_B_c_157_n N_C_c_198_n 0.0200227f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_151 B N_C_c_199_n 7.59316e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_152 N_B_c_158_n N_C_c_199_n 0.0493861f $X=1.127 $Y=0.995 $X2=0 $Y2=0
cc_153 B N_A_56_297#_c_261_n 0.0110968f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_154 N_B_c_157_n N_A_56_297#_c_261_n 0.00180755f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B_c_158_n N_A_56_297#_c_261_n 0.0121282f $X=1.127 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B_M1000_g N_A_56_297#_c_263_n 0.00247352f $X=1.21 $Y=1.985 $X2=0 $Y2=0
cc_157 B N_A_56_297#_c_241_n 0.00493317f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_158 B N_A_56_297#_c_242_n 0.00329776f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_159 N_B_c_158_n N_A_56_297#_c_242_n 0.00147233f $X=1.127 $Y=0.995 $X2=0 $Y2=0
cc_160 B N_A_56_297#_c_243_n 0.00420985f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_161 B N_A_56_297#_c_286_n 0.00537848f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_162 N_B_c_158_n N_A_56_297#_c_286_n 0.00447612f $X=1.127 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B_M1000_g N_VPWR_c_418_n 0.00932461f $X=1.21 $Y=1.985 $X2=0 $Y2=0
cc_164 N_B_M1000_g N_VPWR_c_420_n 0.00295479f $X=1.21 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B_M1000_g N_VPWR_c_414_n 0.00362847f $X=1.21 $Y=1.985 $X2=0 $Y2=0
cc_166 B A_152_47# 0.00271229f $X=1.065 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_167 N_B_c_158_n N_VGND_c_540_n 0.00377907f $X=1.127 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B_c_158_n N_VGND_c_547_n 0.0055266f $X=1.127 $Y=0.995 $X2=0 $Y2=0
cc_169 N_C_c_199_n N_A_56_297#_c_237_n 0.017966f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_170 N_C_M1006_g N_A_56_297#_M1003_g 0.0323588f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_171 N_C_c_199_n N_A_56_297#_c_261_n 2.33057e-19 $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_172 N_C_M1006_g N_A_56_297#_c_263_n 0.00923969f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_173 C N_A_56_297#_c_263_n 0.0110588f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_174 N_C_c_198_n N_A_56_297#_c_263_n 0.00142954f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_175 C N_A_56_297#_c_294_n 0.00601829f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_176 N_C_c_198_n N_A_56_297#_c_294_n 0.00183917f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_177 N_C_c_199_n N_A_56_297#_c_294_n 0.0070961f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_178 C N_A_56_297#_c_241_n 0.00180742f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_179 N_C_c_199_n N_A_56_297#_c_241_n 0.00211339f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C_M1006_g N_A_56_297#_c_250_n 0.00370421f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_181 C N_A_56_297#_c_286_n 0.00519792f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_182 N_C_c_199_n N_A_56_297#_c_286_n 0.0122444f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_183 N_C_M1006_g N_A_56_297#_c_244_n 5.42739e-19 $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_184 C N_A_56_297#_c_244_n 0.0259704f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_185 N_C_c_198_n N_A_56_297#_c_244_n 0.00249723f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_186 C N_A_56_297#_c_245_n 2.97304e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_187 N_C_c_198_n N_A_56_297#_c_245_n 0.0113804f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_188 N_C_M1006_g N_VPWR_c_415_n 0.00171766f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_189 N_C_M1006_g N_VPWR_c_418_n 0.00111348f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_190 N_C_M1006_g N_VPWR_c_420_n 0.00422112f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_191 N_C_M1006_g N_VPWR_c_414_n 0.00588844f $X=1.66 $Y=1.985 $X2=0 $Y2=0
cc_192 N_C_c_199_n N_VGND_c_537_n 0.00662989f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_193 N_C_c_199_n N_VGND_c_540_n 0.00398339f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_194 N_C_c_199_n N_VGND_c_547_n 0.00583361f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_56_297#_c_240_n A_N 0.00386664f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_56_297#_c_245_n N_A_N_c_384_n 0.018687f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_56_297#_c_240_n N_A_N_c_385_n 0.0219107f $X=3.455 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_56_297#_M1015_g N_A_N_c_388_n 0.0376211f $X=3.455 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_56_297#_c_263_n N_VPWR_M1006_d 0.00722999f $X=1.885 $Y=1.61 $X2=0
+ $Y2=0
cc_200 N_A_56_297#_c_250_n N_VPWR_M1006_d 4.46631e-19 $X=1.97 $Y=1.525 $X2=0
+ $Y2=0
cc_201 N_A_56_297#_M1003_g N_VPWR_c_415_n 0.00170185f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_A_56_297#_M1003_g N_VPWR_c_416_n 0.00109012f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_56_297#_M1008_g N_VPWR_c_416_n 0.00838688f $X=2.605 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_56_297#_M1013_g N_VPWR_c_416_n 0.00785375f $X=3.025 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_56_297#_M1015_g N_VPWR_c_416_n 0.00105243f $X=3.455 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_56_297#_M1013_g N_VPWR_c_417_n 0.00104065f $X=3.025 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_56_297#_M1015_g N_VPWR_c_417_n 0.0076562f $X=3.455 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_56_297#_c_252_n N_VPWR_c_419_n 0.00843196f $X=0.425 $Y=1.66 $X2=0
+ $Y2=0
cc_209 N_A_56_297#_M1003_g N_VPWR_c_422_n 0.00422112f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_56_297#_M1008_g N_VPWR_c_422_n 0.00322931f $X=2.605 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_56_297#_M1013_g N_VPWR_c_424_n 0.00337001f $X=3.025 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_56_297#_M1015_g N_VPWR_c_424_n 0.00351072f $X=3.455 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_56_297#_M1007_s N_VPWR_c_414_n 0.006758f $X=0.28 $Y=1.485 $X2=0 $Y2=0
cc_214 N_A_56_297#_M1000_d N_VPWR_c_414_n 0.00341753f $X=1.285 $Y=1.485 $X2=0
+ $Y2=0
cc_215 N_A_56_297#_M1003_g N_VPWR_c_414_n 0.00585201f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_56_297#_M1008_g N_VPWR_c_414_n 0.00386154f $X=2.605 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_56_297#_M1013_g N_VPWR_c_414_n 0.00397572f $X=3.025 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_56_297#_M1015_g N_VPWR_c_414_n 0.00411677f $X=3.455 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_56_297#_c_252_n N_VPWR_c_414_n 0.0114138f $X=0.425 $Y=1.66 $X2=0
+ $Y2=0
cc_220 N_A_56_297#_M1003_g N_X_c_490_n 0.00208318f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_56_297#_M1008_g N_X_c_490_n 0.00844125f $X=2.605 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A_56_297#_M1013_g N_X_c_490_n 0.00844125f $X=3.025 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_56_297#_M1015_g N_X_c_490_n 0.00534716f $X=3.455 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_56_297#_c_251_n N_X_c_490_n 0.0554173f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_56_297#_c_245_n N_X_c_490_n 0.00414616f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_56_297#_c_238_n N_X_c_497_n 0.011111f $X=2.595 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_56_297#_c_239_n N_X_c_497_n 0.0110478f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_56_297#_c_245_n N_X_c_497_n 0.00235864f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_56_297#_c_251_n N_X_c_500_n 0.0529713f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_56_297#_c_245_n N_X_c_500_n 0.00234013f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_56_297#_c_240_n X 0.00741445f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_56_297#_c_245_n X 0.00354528f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_56_297#_c_239_n X 0.00322576f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_56_297#_M1013_g X 0.00399219f $X=3.025 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_56_297#_c_240_n X 0.00346564f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_56_297#_M1015_g X 0.00491067f $X=3.455 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_56_297#_c_251_n X 0.0262398f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_56_297#_c_245_n X 0.0149733f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_56_297#_c_261_n A_152_47# 0.00967848f $X=1.42 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_240 N_A_56_297#_c_261_n A_257_47# 0.00436202f $X=1.42 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_241 N_A_56_297#_c_286_n A_257_47# 0.00523052f $X=1.51 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_242 N_A_56_297#_c_294_n N_VGND_M1011_d 0.00939743f $X=1.885 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_56_297#_c_241_n N_VGND_M1011_d 0.00126621f $X=2 $Y=1.02 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_56_297#_c_237_n N_VGND_c_537_n 0.0075957f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_56_297#_c_238_n N_VGND_c_537_n 0.00103561f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_56_297#_c_294_n N_VGND_c_537_n 0.0217515f $X=1.885 $Y=0.71 $X2=0
+ $Y2=0
cc_247 N_A_56_297#_c_286_n N_VGND_c_537_n 0.00639825f $X=1.51 $Y=0.45 $X2=0
+ $Y2=0
cc_248 N_A_56_297#_c_237_n N_VGND_c_538_n 0.00104703f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_56_297#_c_238_n N_VGND_c_538_n 0.0076774f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_56_297#_c_239_n N_VGND_c_538_n 0.00625485f $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_56_297#_c_240_n N_VGND_c_538_n 4.98572e-19 $X=3.455 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_56_297#_c_239_n N_VGND_c_539_n 4.98572e-19 $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A_56_297#_c_240_n N_VGND_c_539_n 0.00652699f $X=3.455 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A_56_297#_c_261_n N_VGND_c_540_n 0.0273292f $X=1.42 $Y=0.45 $X2=0 $Y2=0
cc_255 N_A_56_297#_c_294_n N_VGND_c_540_n 0.00276954f $X=1.885 $Y=0.71 $X2=0
+ $Y2=0
cc_256 N_A_56_297#_c_242_n N_VGND_c_540_n 0.0318852f $X=0.47 $Y=0.38 $X2=0 $Y2=0
cc_257 N_A_56_297#_c_286_n N_VGND_c_540_n 0.00615001f $X=1.51 $Y=0.45 $X2=0
+ $Y2=0
cc_258 N_A_56_297#_c_237_n N_VGND_c_542_n 0.00501198f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_56_297#_c_238_n N_VGND_c_542_n 0.00351072f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_56_297#_c_239_n N_VGND_c_544_n 0.00351072f $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_56_297#_c_240_n N_VGND_c_544_n 0.00350947f $X=3.455 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_56_297#_M1010_s N_VGND_c_547_n 0.0024621f $X=0.305 $Y=0.235 $X2=0
+ $Y2=0
cc_263 N_A_56_297#_c_237_n N_VGND_c_547_n 0.00840993f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_56_297#_c_238_n N_VGND_c_547_n 0.00411677f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_56_297#_c_239_n N_VGND_c_547_n 0.0040731f $X=3.025 $Y=0.995 $X2=0
+ $Y2=0
cc_266 N_A_56_297#_c_240_n N_VGND_c_547_n 0.00407112f $X=3.455 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_56_297#_c_261_n N_VGND_c_547_n 0.0261818f $X=1.42 $Y=0.45 $X2=0 $Y2=0
cc_268 N_A_56_297#_c_294_n N_VGND_c_547_n 0.00673056f $X=1.885 $Y=0.71 $X2=0
+ $Y2=0
cc_269 N_A_56_297#_c_242_n N_VGND_c_547_n 0.0183637f $X=0.47 $Y=0.38 $X2=0 $Y2=0
cc_270 N_A_56_297#_c_286_n N_VGND_c_547_n 0.00600073f $X=1.51 $Y=0.45 $X2=0
+ $Y2=0
cc_271 A_N N_VPWR_M1015_s 0.00299822f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_272 N_A_N_c_388_n N_VPWR_c_417_n 0.00882316f $X=3.902 $Y=1.325 $X2=0 $Y2=0
cc_273 N_A_N_c_388_n N_VPWR_c_426_n 0.00422112f $X=3.902 $Y=1.325 $X2=0 $Y2=0
cc_274 N_A_N_c_388_n N_VPWR_c_414_n 0.00708071f $X=3.902 $Y=1.325 $X2=0 $Y2=0
cc_275 A_N X 0.0498985f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_276 N_A_N_c_384_n X 9.66564e-19 $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_N_c_385_n X 2.93679e-19 $X=3.902 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_N_c_388_n X 4.22939e-19 $X=3.902 $Y=1.325 $X2=0 $Y2=0
cc_279 A_N N_VGND_M1014_d 0.003576f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_280 A_N N_VGND_c_539_n 0.00987137f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_281 N_A_N_c_384_n N_VGND_c_539_n 2.41939e-19 $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_N_c_385_n N_VGND_c_539_n 0.00780265f $X=3.902 $Y=0.995 $X2=0 $Y2=0
cc_283 A_N N_VGND_c_546_n 0.00251532f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_284 N_A_N_c_385_n N_VGND_c_546_n 0.00446012f $X=3.902 $Y=0.995 $X2=0 $Y2=0
cc_285 A_N N_VGND_c_547_n 0.0049869f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_286 N_A_N_c_385_n N_VGND_c_547_n 0.00798639f $X=3.902 $Y=0.995 $X2=0 $Y2=0
cc_287 N_VPWR_c_414_n N_X_M1003_d 0.00330361f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_414_n N_X_M1013_d 0.00318969f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_M1008_s N_X_c_490_n 0.00316343f $X=2.68 $Y=1.485 $X2=0 $Y2=0
cc_290 N_X_c_497_n N_VGND_M1005_d 0.00327388f $X=3.145 $Y=0.73 $X2=0 $Y2=0
cc_291 N_X_c_497_n N_VGND_c_538_n 0.0162283f $X=3.145 $Y=0.73 $X2=0 $Y2=0
cc_292 X N_VGND_c_539_n 0.00184492f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_293 N_X_c_497_n N_VGND_c_542_n 0.00263122f $X=3.145 $Y=0.73 $X2=0 $Y2=0
cc_294 N_X_c_500_n N_VGND_c_542_n 0.00436709f $X=2.475 $Y=0.68 $X2=0 $Y2=0
cc_295 N_X_c_497_n N_VGND_c_544_n 0.00263122f $X=3.145 $Y=0.73 $X2=0 $Y2=0
cc_296 N_X_c_523_p N_VGND_c_544_n 0.0123718f $X=3.24 $Y=0.42 $X2=0 $Y2=0
cc_297 X N_VGND_c_544_n 0.00279855f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_298 N_X_M1004_s N_VGND_c_547_n 0.00434391f $X=2.24 $Y=0.235 $X2=0 $Y2=0
cc_299 N_X_M1012_s N_VGND_c_547_n 0.00251147f $X=3.1 $Y=0.235 $X2=0 $Y2=0
cc_300 N_X_c_497_n N_VGND_c_547_n 0.0101713f $X=3.145 $Y=0.73 $X2=0 $Y2=0
cc_301 N_X_c_523_p N_VGND_c_547_n 0.00722256f $X=3.24 $Y=0.42 $X2=0 $Y2=0
cc_302 N_X_c_500_n N_VGND_c_547_n 0.00604783f $X=2.475 $Y=0.68 $X2=0 $Y2=0
cc_303 X N_VGND_c_547_n 0.00467557f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_304 A_152_47# N_VGND_c_547_n 0.00316087f $X=0.76 $Y=0.235 $X2=0 $Y2=0
cc_305 A_257_47# N_VGND_c_547_n 0.00192961f $X=1.285 $Y=0.235 $X2=1.885 $Y2=0.71

* File: sky130_fd_sc_hd__xnor2_1.spice
* Created: Thu Aug 27 14:48:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__xnor2_1.spice.pex"
.subckt sky130_fd_sc_hd__xnor2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1005 A_129_47# N_B_M1005_g N_A_47_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.169 PD=0.86 PS=1.82 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g A_129_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.06825 PD=0.92 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.5 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1001 N_A_285_47#_M1001_d N_A_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_285_47#_M1006_d N_B_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1009_d N_A_47_47#_M1009_g N_A_285_47#_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.195 AS=0.08775 PD=1.9 PS=0.92 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_47_47#_M1008_d N_B_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.3 PD=1.27 PS=2.6 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.4
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_47_47#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.365 AS=0.135 PD=1.73 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1002 A_377_297# N_A_M1002_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.365 PD=1.21 PS=1.73 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g A_377_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.105 PD=1.33 PS=1.21 NRD=10.8153 NRS=9.8303 M=1 R=6.66667 SA=75001.9
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_47_47#_M1000_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.36 AS=0.165 PD=2.72 PS=1.33 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__xnor2_1.spice.SKY130_FD_SC_HD__XNOR2_1.pxi"
*
.ends
*
*

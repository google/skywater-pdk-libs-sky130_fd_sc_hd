* File: sky130_fd_sc_hd__o221a_2.spice
* Created: Thu Aug 27 14:36:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o221a_2.spice.pex"
.subckt sky130_fd_sc_hd__o221a_2  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1006 N_A_141_47#_M1006_d N_C1_M1006_g N_A_38_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.23725 PD=0.92 PS=2.03 NRD=0 NRS=14.76 M=1 R=4.33333
+ SA=75000.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1003 N_A_225_47#_M1003_d N_B1_M1003_g N_A_141_47#_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_141_47#_M1007_d N_B2_M1007_g N_A_225_47#_M1003_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_225_47#_M1001_d N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A1_M1013_g N_A_225_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1004_d N_A_38_47#_M1004_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1004_d N_A_38_47#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_C1_M1011_g N_A_38_47#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.325 PD=1.33 PS=2.65 NRD=5.8903 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1005 A_237_297# N_B1_M1005_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1 AD=0.1125
+ AS=0.165 PD=1.225 PS=1.33 NRD=11.3078 NRS=3.9203 M=1 R=6.66667 SA=75000.7
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_38_47#_M1009_d N_B2_M1009_g A_237_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.3875 AS=0.1125 PD=1.775 PS=1.225 NRD=0 NRS=11.3078 M=1 R=6.66667
+ SA=75001.1 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 A_497_297# N_A2_M1010_g N_A_38_47#_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.3875 PD=1.21 PS=1.775 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75002
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g A_497_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.105 PD=1.33 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.4 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1012_d N_A_38_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_38_47#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_40 VNB 0 1.90646e-19 $X=0.12 $Y=-0.085
*
.include "sky130_fd_sc_hd__o221a_2.spice.SKY130_FD_SC_HD__O221A_2.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__o2bb2ai_4.pex.spice
* Created: Tue Sep  1 19:24:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%A2_N 1 3 6 8 10 13 15 17 20 22 24 27 29 40
+ 41
c62 22 0 1.79953e-19 $X=1.75 $Y=0.995
r63 39 41 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.75 $Y2=1.16
r64 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r65 37 39 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.61 $Y2=1.16
r66 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r67 34 36 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=0.59 $Y=1.16
+ $X2=0.91 $Y2=1.16
r68 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r69 31 34 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.59
+ $Y2=1.16
r70 29 40 24.8225 $w=2.08e-07 $l=4.7e-07 $layer=LI1_cond $X=1.14 $Y=1.18
+ $X2=1.61 $Y2=1.18
r71 29 35 29.0476 $w=2.08e-07 $l=5.5e-07 $layer=LI1_cond $X=1.14 $Y=1.18
+ $X2=0.59 $Y2=1.18
r72 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r73 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r74 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r75 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r76 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r77 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r78 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r79 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r80 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r81 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r82 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r83 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r84 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r85 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r86 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r87 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%A1_N 1 3 6 8 10 13 15 17 20 22 24 27 29 40
+ 41
c78 1 0 8.27827e-20 $X=2.17 $Y=0.995
r79 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.28 $Y=1.16
+ $X2=3.43 $Y2=1.16
r80 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.28
+ $Y=1.16 $X2=3.28 $Y2=1.16
r81 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.28 $Y2=1.16
r82 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=3.01 $Y2=1.16
r83 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.59 $Y2=1.16
r84 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r85 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.17 $Y=1.16 $X2=2.26
+ $Y2=1.16
r86 29 40 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=2.98 $Y=1.18 $X2=3.28
+ $Y2=1.18
r87 29 35 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=2.98 $Y=1.18 $X2=2.26
+ $Y2=1.18
r88 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r89 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.985
r90 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r92 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r93 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.985
r94 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.16
r95 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r96 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.16
r97 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.985
r98 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r99 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r100 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r101 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r102 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%A_113_47# 1 2 3 4 5 6 21 23 25 28 30 32 35
+ 37 39 42 44 46 48 49 53 55 56 59 61 65 67 71 73 77 79 82 83 88 92 94 96 98 109
c156 53 0 8.27827e-20 $X=1.54 $Y=0.73
r157 108 109 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.6 $Y=1.16
+ $X2=5.63 $Y2=1.16
r158 105 106 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.18 $Y=1.16
+ $X2=5.21 $Y2=1.16
r159 104 105 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=5.18 $Y2=1.16
r160 103 104 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.76 $Y=1.16
+ $X2=4.79 $Y2=1.16
r161 99 101 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.34 $Y=1.16
+ $X2=4.37 $Y2=1.16
r162 89 108 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.48 $Y=1.16
+ $X2=5.6 $Y2=1.16
r163 89 106 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.48 $Y=1.16
+ $X2=5.21 $Y2=1.16
r164 88 89 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.48
+ $Y=1.16 $X2=5.48 $Y2=1.16
r165 86 103 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.76 $Y2=1.16
r166 86 101 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.37 $Y2=1.16
r167 85 88 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=4.46 $Y=1.18
+ $X2=5.48 $Y2=1.18
r168 85 86 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r169 83 85 28.7836 $w=2.08e-07 $l=5.45e-07 $layer=LI1_cond $X=3.915 $Y=1.18
+ $X2=4.46 $Y2=1.18
r170 81 83 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.83 $Y=1.285
+ $X2=3.915 $Y2=1.18
r171 81 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.83 $Y=1.285
+ $X2=3.83 $Y2=1.455
r172 80 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=1.54
+ $X2=3.22 $Y2=1.54
r173 79 82 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.745 $Y=1.54
+ $X2=3.83 $Y2=1.455
r174 79 80 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.745 $Y=1.54
+ $X2=3.345 $Y2=1.54
r175 75 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.625
+ $X2=3.22 $Y2=1.54
r176 75 77 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.22 $Y=1.625
+ $X2=3.22 $Y2=2.3
r177 74 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=1.54
+ $X2=2.38 $Y2=1.54
r178 73 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=1.54
+ $X2=3.22 $Y2=1.54
r179 73 74 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.095 $Y=1.54
+ $X2=2.505 $Y2=1.54
r180 69 96 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=1.625
+ $X2=2.38 $Y2=1.54
r181 69 71 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.38 $Y=1.625
+ $X2=2.38 $Y2=2.3
r182 68 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=1.54
+ $X2=1.54 $Y2=1.54
r183 67 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=1.54
+ $X2=2.38 $Y2=1.54
r184 67 68 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.255 $Y=1.54
+ $X2=1.665 $Y2=1.54
r185 63 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.625
+ $X2=1.54 $Y2=1.54
r186 63 65 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.54 $Y=1.625
+ $X2=1.54 $Y2=2.3
r187 62 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=1.54
+ $X2=0.7 $Y2=1.54
r188 61 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=1.54
+ $X2=1.54 $Y2=1.54
r189 61 62 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.415 $Y=1.54
+ $X2=0.825 $Y2=1.54
r190 57 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.625
+ $X2=0.7 $Y2=1.54
r191 57 59 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=1.625
+ $X2=0.7 $Y2=2.3
r192 55 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=1.54
+ $X2=0.7 $Y2=1.54
r193 55 56 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.575 $Y=1.54
+ $X2=0.255 $Y2=1.54
r194 51 53 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=0.7 $Y=0.775
+ $X2=1.54 $Y2=0.775
r195 49 51 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=0.255 $Y=0.775
+ $X2=0.7 $Y2=0.775
r196 48 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.255 $Y2=1.54
r197 47 49 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.255 $Y2=0.775
r198 47 48 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.17 $Y2=1.455
r199 44 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=1.16
r200 44 46 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=0.56
r201 40 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.6 $Y=1.325
+ $X2=5.6 $Y2=1.16
r202 40 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.6 $Y=1.325
+ $X2=5.6 $Y2=1.985
r203 37 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=1.16
r204 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=0.56
r205 33 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.18 $Y=1.325
+ $X2=5.18 $Y2=1.16
r206 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.18 $Y=1.325
+ $X2=5.18 $Y2=1.985
r207 30 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=1.16
r208 30 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=0.56
r209 26 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.76 $Y=1.325
+ $X2=4.76 $Y2=1.16
r210 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.76 $Y=1.325
+ $X2=4.76 $Y2=1.985
r211 23 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=1.16
r212 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=0.56
r213 19 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.34 $Y=1.325
+ $X2=4.34 $Y2=1.16
r214 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.34 $Y=1.325
+ $X2=4.34 $Y2=1.985
r215 6 98 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.62
r216 6 77 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=2.3
r217 5 96 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.62
r218 5 71 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=2.3
r219 4 94 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.62
r220 4 65 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2.3
r221 3 92 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.62
r222 3 59 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2.3
r223 2 53 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.73
r224 1 51 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 35
+ 41
c81 1 0 2.9244e-20 $X=6.54 $Y=0.995
r82 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.65 $Y=1.16 $X2=7.8
+ $Y2=1.16
r83 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.38 $Y=1.16
+ $X2=7.65 $Y2=1.16
r84 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.96 $Y=1.16
+ $X2=7.38 $Y2=1.16
r85 35 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.65
+ $Y=1.16 $X2=7.65 $Y2=1.16
r86 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.63 $Y=1.16
+ $X2=6.96 $Y2=1.16
r87 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.63
+ $Y=1.16 $X2=6.63 $Y2=1.16
r88 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.54 $Y=1.16 $X2=6.63
+ $Y2=1.16
r89 29 35 0.259574 $w=1.408e-06 $l=3e-08 $layer=LI1_cond $X=7.17 $Y=1.19
+ $X2=7.17 $Y2=1.16
r90 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.8 $Y=1.325
+ $X2=7.8 $Y2=1.16
r91 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.8 $Y=1.325 $X2=7.8
+ $Y2=1.985
r92 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.8 $Y=0.995
+ $X2=7.8 $Y2=1.16
r93 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.8 $Y=0.995 $X2=7.8
+ $Y2=0.56
r94 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.38 $Y=1.325
+ $X2=7.38 $Y2=1.16
r95 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.38 $Y=1.325
+ $X2=7.38 $Y2=1.985
r96 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.38 $Y=0.995
+ $X2=7.38 $Y2=1.16
r97 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.38 $Y=0.995
+ $X2=7.38 $Y2=0.56
r98 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.96 $Y=1.325
+ $X2=6.96 $Y2=1.16
r99 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.96 $Y=1.325
+ $X2=6.96 $Y2=1.985
r100 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.96 $Y=0.995
+ $X2=6.96 $Y2=1.16
r101 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.96 $Y=0.995
+ $X2=6.96 $Y2=0.56
r102 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.54 $Y=1.325
+ $X2=6.54 $Y2=1.16
r103 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.54 $Y=1.325
+ $X2=6.54 $Y2=1.985
r104 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.54 $Y=0.995
+ $X2=6.54 $Y2=1.16
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.54 $Y=0.995
+ $X2=6.54 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 40
+ 41
r75 39 41 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=9.3 $Y=1.16 $X2=9.48
+ $Y2=1.16
r76 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.3 $Y=1.16
+ $X2=9.3 $Y2=1.16
r77 37 39 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=9.06 $Y=1.16 $X2=9.3
+ $Y2=1.16
r78 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.64 $Y=1.16
+ $X2=9.06 $Y2=1.16
r79 34 36 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=8.28 $Y=1.16
+ $X2=8.64 $Y2=1.16
r80 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.28
+ $Y=1.16 $X2=8.28 $Y2=1.16
r81 31 34 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.22 $Y=1.16 $X2=8.28
+ $Y2=1.16
r82 29 40 17.4286 $w=2.08e-07 $l=3.3e-07 $layer=LI1_cond $X=8.97 $Y=1.18 $X2=9.3
+ $Y2=1.18
r83 29 35 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=8.97 $Y=1.18
+ $X2=8.28 $Y2=1.18
r84 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.48 $Y=1.325
+ $X2=9.48 $Y2=1.16
r85 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.48 $Y=1.325
+ $X2=9.48 $Y2=1.985
r86 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.48 $Y=0.995
+ $X2=9.48 $Y2=1.16
r87 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.48 $Y=0.995
+ $X2=9.48 $Y2=0.56
r88 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.325
+ $X2=9.06 $Y2=1.16
r89 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.06 $Y=1.325
+ $X2=9.06 $Y2=1.985
r90 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=0.995
+ $X2=9.06 $Y2=1.16
r91 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.06 $Y=0.995
+ $X2=9.06 $Y2=0.56
r92 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.64 $Y=1.325
+ $X2=8.64 $Y2=1.16
r93 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.64 $Y=1.325
+ $X2=8.64 $Y2=1.985
r94 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.64 $Y=0.995
+ $X2=8.64 $Y2=1.16
r95 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.64 $Y=0.995
+ $X2=8.64 $Y2=0.56
r96 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.22 $Y=1.325
+ $X2=8.22 $Y2=1.16
r97 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.22 $Y=1.325 $X2=8.22
+ $Y2=1.985
r98 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.22 $Y=0.995
+ $X2=8.22 $Y2=1.16
r99 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.22 $Y=0.995 $X2=8.22
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46
+ 50 52 56 60 64 67 68 70 71 72 73 75 76 78 79 80 82 94 113 114 120 123 126 131
r150 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r151 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r152 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r153 117 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r154 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r155 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r156 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r157 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r158 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r159 105 108 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=8.05 $Y2=2.72
r160 105 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r161 104 107 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=8.05 $Y2=2.72
r162 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r163 102 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.935 $Y=2.72
+ $X2=5.81 $Y2=2.72
r164 102 104 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.935 $Y=2.72
+ $X2=6.21 $Y2=2.72
r165 101 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r166 101 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r167 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 98 123 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=3.885 $Y2=2.72
r169 98 100 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=4.83 $Y2=2.72
r170 97 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r171 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r172 94 123 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.885 $Y2=2.72
r173 94 96 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.45 $Y2=2.72
r174 93 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r175 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r176 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 90 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r178 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r179 87 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.12 $Y2=2.72
r180 87 89 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.61 $Y2=2.72
r181 86 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r182 86 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r183 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 83 117 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r185 83 85 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.69 $Y2=2.72
r186 82 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=1.12 $Y2=2.72
r187 82 85 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=0.69 $Y2=2.72
r188 80 131 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=2.72
+ $X2=0.23 $Y2=2.72
r189 78 110 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=8.97 $Y2=2.72
r190 78 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=9.27 $Y2=2.72
r191 77 113 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.395 $Y=2.72
+ $X2=9.89 $Y2=2.72
r192 77 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.395 $Y=2.72
+ $X2=9.27 $Y2=2.72
r193 75 107 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.305 $Y=2.72
+ $X2=8.05 $Y2=2.72
r194 75 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.305 $Y=2.72
+ $X2=8.43 $Y2=2.72
r195 74 110 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.555 $Y=2.72
+ $X2=8.97 $Y2=2.72
r196 74 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.555 $Y=2.72
+ $X2=8.43 $Y2=2.72
r197 72 100 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.845 $Y=2.72
+ $X2=4.83 $Y2=2.72
r198 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.845 $Y=2.72
+ $X2=4.97 $Y2=2.72
r199 70 92 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.675 $Y=2.72
+ $X2=2.53 $Y2=2.72
r200 70 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.675 $Y=2.72
+ $X2=2.8 $Y2=2.72
r201 69 96 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.925 $Y=2.72
+ $X2=3.45 $Y2=2.72
r202 69 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.925 $Y=2.72
+ $X2=2.8 $Y2=2.72
r203 67 89 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.61 $Y2=2.72
r204 67 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.96 $Y2=2.72
r205 66 92 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.085 $Y=2.72
+ $X2=2.53 $Y2=2.72
r206 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=2.72
+ $X2=1.96 $Y2=2.72
r207 62 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=2.635
+ $X2=9.27 $Y2=2.72
r208 62 64 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=9.27 $Y=2.635
+ $X2=9.27 $Y2=1.96
r209 58 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=2.635
+ $X2=8.43 $Y2=2.72
r210 58 60 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.43 $Y=2.635
+ $X2=8.43 $Y2=1.96
r211 54 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.81 $Y=2.635
+ $X2=5.81 $Y2=2.72
r212 54 56 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.81 $Y=2.635
+ $X2=5.81 $Y2=1.96
r213 53 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=4.97 $Y2=2.72
r214 52 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.685 $Y=2.72
+ $X2=5.81 $Y2=2.72
r215 52 53 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.685 $Y=2.72
+ $X2=5.095 $Y2=2.72
r216 48 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=2.635
+ $X2=4.97 $Y2=2.72
r217 48 50 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.97 $Y=2.635
+ $X2=4.97 $Y2=1.96
r218 44 123 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=2.635
+ $X2=3.885 $Y2=2.72
r219 44 46 10.9102 $w=7.38e-07 $l=6.75e-07 $layer=LI1_cond $X=3.885 $Y=2.635
+ $X2=3.885 $Y2=1.96
r220 40 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=2.635
+ $X2=2.8 $Y2=2.72
r221 40 42 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.8 $Y=2.635
+ $X2=2.8 $Y2=1.96
r222 36 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.635
+ $X2=1.96 $Y2=2.72
r223 36 38 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.96 $Y=2.635
+ $X2=1.96 $Y2=1.96
r224 32 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r225 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=1.96
r226 28 117 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.202 $Y2=2.72
r227 28 30 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.28 $Y2=1.96
r228 9 64 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.135
+ $Y=1.485 $X2=9.27 $Y2=1.96
r229 8 60 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=1.485 $X2=8.43 $Y2=1.96
r230 7 56 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.675
+ $Y=1.485 $X2=5.81 $Y2=1.96
r231 6 50 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.835
+ $Y=1.485 $X2=4.97 $Y2=1.96
r232 5 46 150 $w=1.7e-07 $l=8.29156e-07 $layer=licon1_PDIFF $count=4 $X=3.505
+ $Y=1.485 $X2=4.13 $Y2=1.96
r233 4 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=1.96
r234 3 38 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.96
r235 2 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.96
r236 1 30 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%Y 1 2 3 4 5 6 19 25 27 29 33 35 38 39 43
+ 48 49 51 52 55
r86 52 55 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=7.59 $Y=1.625
+ $X2=7.59 $Y2=1.87
r87 52 54 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=1.625
+ $X2=7.59 $Y2=1.54
r88 44 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.875 $Y=1.54
+ $X2=6.75 $Y2=1.54
r89 43 54 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.465 $Y=1.54
+ $X2=7.59 $Y2=1.54
r90 43 44 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.465 $Y=1.54
+ $X2=6.875 $Y2=1.54
r91 40 49 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.155 $Y=1.54
+ $X2=6.015 $Y2=1.54
r92 39 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.625 $Y=1.54
+ $X2=6.75 $Y2=1.54
r93 39 40 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.625 $Y=1.54
+ $X2=6.155 $Y2=1.54
r94 38 49 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=1.455
+ $X2=6.015 $Y2=1.54
r95 37 38 22.6373 $w=2.78e-07 $l=5.5e-07 $layer=LI1_cond $X=6.015 $Y=0.905
+ $X2=6.015 $Y2=1.455
r96 36 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.515 $Y=1.54
+ $X2=5.39 $Y2=1.54
r97 35 49 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.875 $Y=1.54
+ $X2=6.015 $Y2=1.54
r98 35 36 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.875 $Y=1.54
+ $X2=5.515 $Y2=1.54
r99 31 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.39 $Y=1.625
+ $X2=5.39 $Y2=1.54
r100 31 33 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.39 $Y=1.625
+ $X2=5.39 $Y2=2.3
r101 30 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.675 $Y=1.54
+ $X2=4.55 $Y2=1.54
r102 29 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.265 $Y=1.54
+ $X2=5.39 $Y2=1.54
r103 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.265 $Y=1.54
+ $X2=4.675 $Y2=1.54
r104 25 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=1.625
+ $X2=4.55 $Y2=1.54
r105 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.55 $Y=1.625
+ $X2=4.55 $Y2=2.3
r106 21 24 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=4.58 $Y=0.775
+ $X2=5.42 $Y2=0.775
r107 19 37 6.82866 $w=2.6e-07 $l=1.94422e-07 $layer=LI1_cond $X=5.875 $Y=0.775
+ $X2=6.015 $Y2=0.905
r108 19 24 20.1678 $w=2.58e-07 $l=4.55e-07 $layer=LI1_cond $X=5.875 $Y=0.775
+ $X2=5.42 $Y2=0.775
r109 6 54 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=7.455
+ $Y=1.485 $X2=7.59 $Y2=1.62
r110 5 51 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.615
+ $Y=1.485 $X2=6.75 $Y2=1.62
r111 4 48 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.255
+ $Y=1.485 $X2=5.39 $Y2=1.62
r112 4 33 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.255
+ $Y=1.485 $X2=5.39 $Y2=2.3
r113 3 46 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.485 $X2=4.55 $Y2=1.62
r114 3 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.485 $X2=4.55 $Y2=2.3
r115 2 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.235 $X2=5.42 $Y2=0.73
r116 1 21 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%A_1241_297# 1 2 3 4 5 18 20 21 24 26 28 29
+ 30 34 36 38 40 42 48
r63 38 50 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.72 $Y=1.625
+ $X2=9.72 $Y2=1.54
r64 38 40 25.0935 $w=3.08e-07 $l=6.75e-07 $layer=LI1_cond $X=9.72 $Y=1.625
+ $X2=9.72 $Y2=2.3
r65 37 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.975 $Y=1.54
+ $X2=8.85 $Y2=1.54
r66 36 50 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.565 $Y=1.54
+ $X2=9.72 $Y2=1.54
r67 36 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.565 $Y=1.54
+ $X2=8.975 $Y2=1.54
r68 32 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.625
+ $X2=8.85 $Y2=1.54
r69 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.85 $Y=1.625
+ $X2=8.85 $Y2=2.3
r70 31 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.135 $Y=1.54
+ $X2=8.01 $Y2=1.54
r71 30 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.725 $Y=1.54
+ $X2=8.85 $Y2=1.54
r72 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.725 $Y=1.54
+ $X2=8.135 $Y2=1.54
r73 29 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.01 $Y=2.295
+ $X2=8.01 $Y2=2.38
r74 28 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.01 $Y=1.625
+ $X2=8.01 $Y2=1.54
r75 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=8.01 $Y=1.625
+ $X2=8.01 $Y2=2.295
r76 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=2.38
+ $X2=7.17 $Y2=2.38
r77 26 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.885 $Y=2.38
+ $X2=8.01 $Y2=2.38
r78 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.885 $Y=2.38
+ $X2=7.295 $Y2=2.38
r79 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=2.295
+ $X2=7.17 $Y2=2.38
r80 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.17 $Y=2.295
+ $X2=7.17 $Y2=1.96
r81 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.045 $Y=2.38
+ $X2=7.17 $Y2=2.38
r82 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.045 $Y=2.38
+ $X2=6.455 $Y2=2.38
r83 16 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.315 $Y=2.295
+ $X2=6.455 $Y2=2.38
r84 16 18 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.315 $Y=2.295
+ $X2=6.315 $Y2=1.96
r85 5 50 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.555
+ $Y=1.485 $X2=9.69 $Y2=1.62
r86 5 40 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.555
+ $Y=1.485 $X2=9.69 $Y2=2.3
r87 4 48 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.485 $X2=8.85 $Y2=1.62
r88 4 34 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.485 $X2=8.85 $Y2=2.3
r89 3 46 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.01 $Y2=2.3
r90 3 44 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.01 $Y2=1.62
r91 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.035
+ $Y=1.485 $X2=7.17 $Y2=1.96
r92 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=6.205
+ $Y=1.485 $X2=6.33 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%A_27_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
c73 23 0 1.79953e-19 $X=2 $Y=0.725
r74 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.64 $Y=0.725
+ $X2=3.64 $Y2=0.39
r75 31 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.815
+ $X2=2.8 $Y2=0.815
r76 30 32 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.475 $Y=0.815
+ $X2=3.64 $Y2=0.725
r77 30 31 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.475 $Y=0.815
+ $X2=2.965 $Y2=0.815
r78 26 40 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.8 $Y=0.725 $X2=2.8
+ $Y2=0.815
r79 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.8 $Y=0.725 $X2=2.8
+ $Y2=0.39
r80 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0.815 $X2=2
+ $Y2=0.815
r81 24 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=0.815
+ $X2=2.8 $Y2=0.815
r82 24 25 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.635 $Y=0.815
+ $X2=2.125 $Y2=0.815
r83 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2 $Y=0.725 $X2=2
+ $Y2=0.815
r84 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2 $Y=0.475 $X2=2
+ $Y2=0.365
r85 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2 $Y=0.475 $X2=2
+ $Y2=0.725
r86 18 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=0.28 $Y=0.365
+ $X2=1.12 $Y2=0.365
r87 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=0.365 $X2=2
+ $Y2=0.365
r88 16 21 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=1.875 $Y=0.365
+ $X2=1.12 $Y2=0.365
r89 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.39
r90 4 28 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.39
r91 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.73
r92 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r93 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r94 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 55 67 71 84 85 88 91 96
r142 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r143 88 89 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r144 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r145 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r146 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r147 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r148 79 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=7.59
+ $Y2=0
r149 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r150 76 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=0 $X2=7.59
+ $Y2=0
r151 76 78 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.675 $Y=0
+ $X2=8.05 $Y2=0
r152 75 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r153 75 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=6.67
+ $Y2=0
r154 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r155 72 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=0 $X2=6.75
+ $Y2=0
r156 72 74 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.835 $Y=0 $X2=7.13
+ $Y2=0
r157 71 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=0 $X2=7.59
+ $Y2=0
r158 71 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.505 $Y=0
+ $X2=7.13 $Y2=0
r159 70 89 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=6.67 $Y2=0
r160 69 70 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r161 67 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.75
+ $Y2=0
r162 67 69 209.749 $w=1.68e-07 $l=3.215e-06 $layer=LI1_cond $X=6.665 $Y=0
+ $X2=3.45 $Y2=0
r163 66 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r164 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r165 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r166 63 96 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=0.23 $Y2=0
r167 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r168 58 62 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r169 58 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r170 55 96 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=0 $X2=0.23
+ $Y2=0
r171 53 81 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.185 $Y=0
+ $X2=8.97 $Y2=0
r172 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.185 $Y=0 $X2=9.27
+ $Y2=0
r173 52 84 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=9.355 $Y=0
+ $X2=9.89 $Y2=0
r174 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=0 $X2=9.27
+ $Y2=0
r175 50 78 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.345 $Y=0 $X2=8.05
+ $Y2=0
r176 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.345 $Y=0 $X2=8.43
+ $Y2=0
r177 49 81 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.515 $Y=0
+ $X2=8.97 $Y2=0
r178 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.515 $Y=0 $X2=8.43
+ $Y2=0
r179 47 65 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=0
+ $X2=2.99 $Y2=0
r180 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.22
+ $Y2=0
r181 46 69 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.305 $Y=0
+ $X2=3.45 $Y2=0
r182 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.22
+ $Y2=0
r183 44 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=0
+ $X2=2.07 $Y2=0
r184 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.38
+ $Y2=0
r185 43 65 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=2.99 $Y2=0
r186 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.38
+ $Y2=0
r187 39 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=0.085
+ $X2=9.27 $Y2=0
r188 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.27 $Y=0.085
+ $X2=9.27 $Y2=0.39
r189 35 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0
r190 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0.39
r191 31 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=0.085
+ $X2=7.59 $Y2=0
r192 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.59 $Y=0.085
+ $X2=7.59 $Y2=0.39
r193 27 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0
r194 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0.39
r195 23 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0
r196 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0.39
r197 19 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0
r198 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0.39
r199 6 41 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.135
+ $Y=0.235 $X2=9.27 $Y2=0.39
r200 5 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.235 $X2=8.43 $Y2=0.39
r201 4 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.455
+ $Y=0.235 $X2=7.59 $Y2=0.39
r202 3 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.615
+ $Y=0.235 $X2=6.75 $Y2=0.39
r203 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.39
r204 1 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_4%A_807_47# 1 2 3 4 5 6 7 24 26 27 30 31 32
+ 33 36 38 42 44 48 50 54 58 59 60
c117 58 0 2.9244e-20 $X=7.17 $Y=0.815
r118 52 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.69 $Y=0.725
+ $X2=9.69 $Y2=0.39
r119 51 60 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=0.815
+ $X2=8.85 $Y2=0.815
r120 50 52 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=9.525 $Y=0.815
+ $X2=9.69 $Y2=0.725
r121 50 51 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=9.525 $Y=0.815
+ $X2=9.015 $Y2=0.815
r122 46 60 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.85 $Y=0.725
+ $X2=8.85 $Y2=0.815
r123 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.85 $Y=0.725
+ $X2=8.85 $Y2=0.39
r124 45 59 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=0.815
+ $X2=8.01 $Y2=0.815
r125 44 60 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=0.815
+ $X2=8.85 $Y2=0.815
r126 44 45 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=8.685 $Y=0.815
+ $X2=8.175 $Y2=0.815
r127 40 59 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.01 $Y=0.725
+ $X2=8.01 $Y2=0.815
r128 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.01 $Y=0.725
+ $X2=8.01 $Y2=0.39
r129 39 58 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0.815
+ $X2=7.17 $Y2=0.815
r130 38 59 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.845 $Y=0.815
+ $X2=8.01 $Y2=0.815
r131 38 39 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.845 $Y=0.815
+ $X2=7.335 $Y2=0.815
r132 34 58 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.17 $Y=0.725
+ $X2=7.17 $Y2=0.815
r133 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.17 $Y=0.725
+ $X2=7.17 $Y2=0.39
r134 32 58 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=7.005 $Y=0.82
+ $X2=7.17 $Y2=0.815
r135 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.005 $Y=0.82
+ $X2=6.495 $Y2=0.82
r136 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.41 $Y=0.735
+ $X2=6.495 $Y2=0.82
r137 30 57 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.41 $Y=0.475
+ $X2=6.41 $Y2=0.365
r138 30 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.41 $Y=0.475
+ $X2=6.41 $Y2=0.735
r139 27 29 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=4.245 $Y=0.365
+ $X2=5 $Y2=0.365
r140 26 57 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=0.365
+ $X2=6.41 $Y2=0.365
r141 26 29 69.4085 $w=2.18e-07 $l=1.325e-06 $layer=LI1_cond $X=6.325 $Y=0.365
+ $X2=5 $Y2=0.365
r142 22 27 6.88292 $w=2.2e-07 $l=1.49432e-07 $layer=LI1_cond $X=4.152 $Y=0.475
+ $X2=4.245 $Y2=0.365
r143 22 24 6.29484 $w=1.83e-07 $l=1.05e-07 $layer=LI1_cond $X=4.152 $Y=0.475
+ $X2=4.152 $Y2=0.58
r144 7 54 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.555
+ $Y=0.235 $X2=9.69 $Y2=0.39
r145 6 48 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.715
+ $Y=0.235 $X2=8.85 $Y2=0.39
r146 5 42 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.875
+ $Y=0.235 $X2=8.01 $Y2=0.39
r147 4 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.035
+ $Y=0.235 $X2=7.17 $Y2=0.39
r148 3 57 91 $w=1.7e-07 $l=6.98212e-07 $layer=licon1_NDIFF $count=2 $X=5.705
+ $Y=0.235 $X2=6.33 $Y2=0.39
r149 2 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.39
r150 1 24 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.235 $X2=4.16 $Y2=0.58
.ends


* File: sky130_fd_sc_hd__clkdlybuf4s15_1.spice.SKY130_FD_SC_HD__CLKDLYBUF4S15_1.pxi
* Created: Thu Aug 27 14:11:15 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A N_A_M1002_g N_A_M1004_g A N_A_c_68_n
+ N_A_c_69_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_27_47# N_A_27_47#_M1002_s
+ N_A_27_47#_M1004_s N_A_27_47#_c_98_n N_A_27_47#_M1007_g N_A_27_47#_M1001_g
+ N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_102_n N_A_27_47#_c_107_n
+ N_A_27_47#_c_103_n N_A_27_47#_c_104_n N_A_27_47#_c_108_n N_A_27_47#_c_109_n
+ N_A_27_47#_c_105_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_282_47# N_A_282_47#_M1007_d
+ N_A_282_47#_M1001_d N_A_282_47#_c_163_n N_A_282_47#_M1005_g
+ N_A_282_47#_M1000_g N_A_282_47#_c_164_n N_A_282_47#_c_165_n
+ N_A_282_47#_c_166_n N_A_282_47#_c_167_n N_A_282_47#_c_168_n
+ N_A_282_47#_c_169_n N_A_282_47#_c_175_n N_A_282_47#_c_170_n
+ N_A_282_47#_c_171_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_282_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_394_47# N_A_394_47#_M1005_s
+ N_A_394_47#_M1000_s N_A_394_47#_M1003_g N_A_394_47#_M1006_g
+ N_A_394_47#_c_228_n N_A_394_47#_c_234_n N_A_394_47#_c_229_n
+ N_A_394_47#_c_230_n N_A_394_47#_c_235_n N_A_394_47#_c_236_n
+ N_A_394_47#_c_231_n N_A_394_47#_c_232_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_394_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%VPWR N_VPWR_M1004_d N_VPWR_M1000_d
+ N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n VPWR
+ N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_292_n N_VPWR_c_300_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%X N_X_M1003_d N_X_M1006_d X X X X X X
+ N_X_c_334_n X PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%VGND N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n VGND
+ N_VGND_c_353_n N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%VGND
cc_1 VNB N_A_M1002_g 0.043536f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_c_68_n 0.025392f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_3 VNB N_A_c_69_n 0.0126988f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_4 VNB N_A_27_47#_c_98_n 0.0222651f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_5 VNB N_A_27_47#_M1001_g 6.60529e-19 $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_6 VNB N_A_27_47#_c_100_n 0.0494468f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.025
cc_7 VNB N_A_27_47#_c_101_n 0.0135496f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.325
cc_8 VNB N_A_27_47#_c_102_n 0.0185426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_103_n 0.0019047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_104_n 0.0101074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_105_n 0.00431793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_282_47#_c_163_n 0.02332f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_13 VNB N_A_282_47#_c_164_n 0.0247086f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.325
cc_14 VNB N_A_282_47#_c_165_n 0.00453903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_282_47#_c_166_n 0.00498788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_282_47#_c_167_n 0.0138999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_282_47#_c_168_n 0.024662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_282_47#_c_169_n 0.00192115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_282_47#_c_170_n 0.00131782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_282_47#_c_171_n 0.00281555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_394_47#_M1003_g 0.0365036f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_22 VNB N_A_394_47#_c_228_n 0.00430508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_394_47#_c_229_n 0.0012699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_394_47#_c_230_n 0.003261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_394_47#_c_231_n 0.00383365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_394_47#_c_232_n 0.02422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_292_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB X 0.0368703f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_29 VNB N_X_c_334_n 0.0114984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_349_n 0.0055024f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_31 VNB N_VGND_c_350_n 0.00558775f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_32 VNB N_VGND_c_351_n 0.0474987f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_33 VNB N_VGND_c_352_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_353_n 0.0171204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_354_n 0.0185118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_355_n 0.208271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_356_n 0.00602727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_M1004_g 0.0296455f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_39 VPB N_A_c_68_n 0.0057428f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_40 VPB N_A_c_69_n 0.00232387f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_41 VPB N_A_27_47#_M1001_g 0.0394294f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_42 VPB N_A_27_47#_c_107_n 0.0316915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_108_n 0.0016672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_109_n 0.00769094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_105_n 0.0035471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_282_47#_M1000_g 0.0381846f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_47 VPB N_A_282_47#_c_164_n 0.00684497f $X=-0.19 $Y=1.305 $X2=0.39 $Y2=1.325
cc_48 VPB N_A_282_47#_c_168_n 0.00947587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_282_47#_c_175_n 0.00707847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_282_47#_c_170_n 0.00993186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_394_47#_M1006_g 0.0242977f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_52 VPB N_A_394_47#_c_234_n 0.00945826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_394_47#_c_235_n 0.00856849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_394_47#_c_236_n 0.00426045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_394_47#_c_231_n 0.0014633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_394_47#_c_232_n 0.00592207f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_293_n 0.00558649f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_58 VPB N_VPWR_c_294_n 0.00597825f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_59 VPB N_VPWR_c_295_n 0.0462082f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_60 VPB N_VPWR_c_296_n 0.00766468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_297_n 0.0177606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_298_n 0.0187787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_292_n 0.0523513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_300_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB X 0.0195614f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_66 VPB X 0.0295358f $X=-0.19 $Y=1.305 $X2=0.39 $Y2=1.16
cc_67 N_A_M1002_g N_A_27_47#_c_98_n 0.00905157f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_68_n N_A_27_47#_M1001_g 0.014263f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_M1002_g N_A_27_47#_c_100_n 0.0192598f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_c_69_n N_A_27_47#_c_100_n 7.78656e-19 $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_A_27_47#_c_102_n 0.0134754f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_M1004_g N_A_27_47#_c_107_n 0.0163822f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_A_27_47#_c_103_n 0.0102222f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_c_69_n N_A_27_47#_c_103_n 0.00953108f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_M1002_g N_A_27_47#_c_104_n 0.00420722f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_A_27_47#_c_104_n 0.00401319f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_69_n N_A_27_47#_c_104_n 0.0285757f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_A_27_47#_c_108_n 0.0125955f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_c_69_n N_A_27_47#_c_108_n 0.00915457f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_M1004_g N_A_27_47#_c_109_n 0.00422287f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_c_68_n N_A_27_47#_c_109_n 0.00371254f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_69_n N_A_27_47#_c_109_n 0.0257309f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_A_27_47#_c_105_n 0.00465755f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_c_68_n N_A_27_47#_c_105_n 0.00587612f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_c_69_n N_A_27_47#_c_105_n 0.023714f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VPWR_c_293_n 0.00938211f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_VPWR_c_297_n 0.0054895f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_VPWR_c_292_n 0.0115145f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1002_g N_VGND_c_349_n 0.00344941f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VGND_c_353_n 0.00424868f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_VGND_c_355_n 0.00744605f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_101_n N_A_282_47#_c_164_n 0.00454252f $X=1.335 $Y=1.145 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_c_98_n N_A_282_47#_c_165_n 0.00953719f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_98_n N_A_282_47#_c_166_n 0.00341603f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_105_n N_A_282_47#_c_166_n 0.00770619f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_98_n N_A_282_47#_c_169_n 0.00572408f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_M1001_g N_A_282_47#_c_175_n 0.0126518f $X=1.335 $Y=2.075 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_101_n N_A_282_47#_c_170_n 0.0132526f $X=1.335 $Y=1.145 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_108_n N_A_282_47#_c_170_n 0.00825752f $X=0.73 $Y=1.58 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_105_n N_A_282_47#_c_170_n 0.011307f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_101_n N_A_282_47#_c_171_n 0.00290025f $X=1.335 $Y=1.145
+ $X2=0 $Y2=0
cc_102 N_A_27_47#_c_105_n N_A_282_47#_c_171_n 0.00935483f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_108_n N_VPWR_M1004_d 0.0229122f $X=0.73 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_27_47#_c_105_n N_VPWR_M1004_d 3.3297e-19 $X=0.925 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_27_47#_M1001_g N_VPWR_c_293_n 0.00862604f $X=1.335 $Y=2.075 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_100_n N_VPWR_c_293_n 6.02664e-19 $X=1.26 $Y=1.145 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_108_n N_VPWR_c_293_n 0.0274169f $X=0.73 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1001_g N_VPWR_c_295_n 0.0054895f $X=1.335 $Y=2.075 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_107_n N_VPWR_c_297_n 0.0217658f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_110 N_A_27_47#_M1004_s N_VPWR_c_292_n 0.00213418f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1001_g N_VPWR_c_292_n 0.0120171f $X=1.335 $Y=2.075 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_107_n N_VPWR_c_292_n 0.0128348f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_103_n N_VGND_M1002_d 0.0134372f $X=0.73 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_27_47#_c_98_n N_VGND_c_349_n 0.00511159f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_100_n N_VGND_c_349_n 6.32636e-19 $X=1.26 $Y=1.145 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_103_n N_VGND_c_349_n 0.0254149f $X=0.73 $Y=0.8 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_98_n N_VGND_c_351_n 0.0054895f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_103_n N_VGND_c_351_n 0.00488709f $X=0.73 $Y=0.8 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_102_n N_VGND_c_353_n 0.0216552f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_103_n N_VGND_c_353_n 0.00239555f $X=0.73 $Y=0.8 $X2=0 $Y2=0
cc_121 N_A_27_47#_M1002_s N_VGND_c_355_n 0.00213418f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_c_98_n N_VGND_c_355_n 0.0120171f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_102_n N_VGND_c_355_n 0.0128089f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_103_n N_VGND_c_355_n 0.0138547f $X=0.73 $Y=0.8 $X2=0 $Y2=0
cc_125 N_A_282_47#_c_163_n N_A_394_47#_M1003_g 0.0109525f $X=2.31 $Y=1 $X2=0
+ $Y2=0
cc_126 N_A_282_47#_M1000_g N_A_394_47#_M1006_g 0.012465f $X=2.31 $Y=2.075 $X2=0
+ $Y2=0
cc_127 N_A_282_47#_c_163_n N_A_394_47#_c_228_n 0.0154705f $X=2.31 $Y=1 $X2=0
+ $Y2=0
cc_128 N_A_282_47#_c_165_n N_A_394_47#_c_228_n 0.0385933f $X=1.55 $Y=0.38 $X2=0
+ $Y2=0
cc_129 N_A_282_47#_M1000_g N_A_394_47#_c_234_n 0.0270821f $X=2.31 $Y=2.075 $X2=0
+ $Y2=0
cc_130 N_A_282_47#_c_170_n N_A_394_47#_c_234_n 0.0743939f $X=1.572 $Y=1.835
+ $X2=0 $Y2=0
cc_131 N_A_282_47#_c_163_n N_A_394_47#_c_229_n 0.0102603f $X=2.31 $Y=1 $X2=0
+ $Y2=0
cc_132 N_A_282_47#_c_167_n N_A_394_47#_c_229_n 0.0277028f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_282_47#_c_168_n N_A_394_47#_c_229_n 0.00842051f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_282_47#_c_163_n N_A_394_47#_c_230_n 0.00418154f $X=2.31 $Y=1 $X2=0
+ $Y2=0
cc_135 N_A_282_47#_c_164_n N_A_394_47#_c_230_n 0.00526724f $X=2.2 $Y=1.165 $X2=0
+ $Y2=0
cc_136 N_A_282_47#_c_167_n N_A_394_47#_c_230_n 0.0239185f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_282_47#_c_169_n N_A_394_47#_c_230_n 0.0148501f $X=1.572 $Y=0.825
+ $X2=0 $Y2=0
cc_138 N_A_282_47#_c_167_n N_A_394_47#_c_235_n 0.0198283f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_282_47#_c_168_n N_A_394_47#_c_235_n 0.0082263f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_282_47#_M1000_g N_A_394_47#_c_236_n 0.0115419f $X=2.31 $Y=2.075 $X2=0
+ $Y2=0
cc_141 N_A_282_47#_c_164_n N_A_394_47#_c_236_n 0.0056487f $X=2.2 $Y=1.165 $X2=0
+ $Y2=0
cc_142 N_A_282_47#_c_167_n N_A_394_47#_c_236_n 0.0386906f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_282_47#_c_168_n N_A_394_47#_c_236_n 6.19808e-19 $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_282_47#_c_170_n N_A_394_47#_c_236_n 0.014358f $X=1.572 $Y=1.835 $X2=0
+ $Y2=0
cc_145 N_A_282_47#_c_163_n N_A_394_47#_c_231_n 0.00218389f $X=2.31 $Y=1 $X2=0
+ $Y2=0
cc_146 N_A_282_47#_M1000_g N_A_394_47#_c_231_n 0.00170496f $X=2.31 $Y=2.075
+ $X2=0 $Y2=0
cc_147 N_A_282_47#_c_167_n N_A_394_47#_c_231_n 0.0162311f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_148 N_A_282_47#_c_168_n N_A_394_47#_c_231_n 0.00483008f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_282_47#_c_168_n N_A_394_47#_c_232_n 0.0217057f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_282_47#_c_175_n N_VPWR_c_293_n 0.0228386f $X=1.55 $Y=2 $X2=0 $Y2=0
cc_151 N_A_282_47#_M1000_g N_VPWR_c_294_n 0.00597906f $X=2.31 $Y=2.075 $X2=0
+ $Y2=0
cc_152 N_A_282_47#_M1000_g N_VPWR_c_295_n 0.00357668f $X=2.31 $Y=2.075 $X2=0
+ $Y2=0
cc_153 N_A_282_47#_c_175_n N_VPWR_c_295_n 0.0242182f $X=1.55 $Y=2 $X2=0 $Y2=0
cc_154 N_A_282_47#_M1001_d N_VPWR_c_292_n 0.00213418f $X=1.41 $Y=1.665 $X2=0
+ $Y2=0
cc_155 N_A_282_47#_M1000_g N_VPWR_c_292_n 0.00735699f $X=2.31 $Y=2.075 $X2=0
+ $Y2=0
cc_156 N_A_282_47#_c_175_n N_VPWR_c_292_n 0.0141671f $X=1.55 $Y=2 $X2=0 $Y2=0
cc_157 N_A_282_47#_c_165_n N_VGND_c_349_n 0.0102136f $X=1.55 $Y=0.38 $X2=0 $Y2=0
cc_158 N_A_282_47#_c_163_n N_VGND_c_350_n 0.00530768f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_159 N_A_282_47#_c_163_n N_VGND_c_351_n 0.00424868f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_160 N_A_282_47#_c_165_n N_VGND_c_351_n 0.0241445f $X=1.55 $Y=0.38 $X2=0 $Y2=0
cc_161 N_A_282_47#_M1007_d N_VGND_c_355_n 0.00213418f $X=1.41 $Y=0.235 $X2=0
+ $Y2=0
cc_162 N_A_282_47#_c_163_n N_VGND_c_355_n 0.00802257f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_163 N_A_282_47#_c_165_n N_VGND_c_355_n 0.0141471f $X=1.55 $Y=0.38 $X2=0 $Y2=0
cc_164 N_A_394_47#_c_235_n N_VPWR_M1000_d 0.00975842f $X=2.855 $Y=1.505 $X2=0
+ $Y2=0
cc_165 N_A_394_47#_M1006_g N_VPWR_c_294_n 0.00993071f $X=3.17 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_394_47#_c_235_n N_VPWR_c_294_n 0.0338738f $X=2.855 $Y=1.505 $X2=0
+ $Y2=0
cc_167 N_A_394_47#_c_232_n N_VPWR_c_294_n 4.16759e-19 $X=3.11 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_394_47#_c_234_n N_VPWR_c_295_n 0.0304911f $X=2.095 $Y=2 $X2=0 $Y2=0
cc_169 N_A_394_47#_M1006_g N_VPWR_c_298_n 0.00533769f $X=3.17 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_394_47#_M1000_s N_VPWR_c_292_n 0.00213418f $X=1.97 $Y=1.665 $X2=0
+ $Y2=0
cc_171 N_A_394_47#_M1006_g N_VPWR_c_292_n 0.0112012f $X=3.17 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_394_47#_c_234_n N_VPWR_c_292_n 0.0176502f $X=2.095 $Y=2 $X2=0 $Y2=0
cc_173 N_A_394_47#_M1003_g X 0.0310376f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A_394_47#_c_229_n X 0.0138867f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_175 N_A_394_47#_c_235_n X 0.0137399f $X=2.855 $Y=1.505 $X2=0 $Y2=0
cc_176 N_A_394_47#_c_231_n X 0.0410932f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_394_47#_M1006_g X 0.0109775f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_394_47#_M1003_g N_X_c_334_n 0.00485391f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A_394_47#_c_229_n N_VGND_M1005_d 0.015296f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_180 N_A_394_47#_M1003_g N_VGND_c_350_n 0.00616133f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_394_47#_c_228_n N_VGND_c_350_n 0.0106109f $X=2.095 $Y=0.38 $X2=0
+ $Y2=0
cc_182 N_A_394_47#_c_229_n N_VGND_c_350_n 0.0271231f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_183 N_A_394_47#_c_232_n N_VGND_c_350_n 3.93243e-19 $X=3.11 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_394_47#_c_228_n N_VGND_c_351_n 0.0209424f $X=2.095 $Y=0.38 $X2=0
+ $Y2=0
cc_185 N_A_394_47#_c_229_n N_VGND_c_351_n 0.00610976f $X=2.855 $Y=0.8 $X2=0
+ $Y2=0
cc_186 N_A_394_47#_M1003_g N_VGND_c_354_n 0.0043439f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_187 N_A_394_47#_c_229_n N_VGND_c_354_n 0.0024529f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_188 N_A_394_47#_M1005_s N_VGND_c_355_n 0.00213418f $X=1.97 $Y=0.235 $X2=0
+ $Y2=0
cc_189 N_A_394_47#_M1003_g N_VGND_c_355_n 0.00800603f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_190 N_A_394_47#_c_228_n N_VGND_c_355_n 0.0124245f $X=2.095 $Y=0.38 $X2=0
+ $Y2=0
cc_191 N_A_394_47#_c_229_n N_VGND_c_355_n 0.0166411f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_192 N_VPWR_c_292_n N_X_M1006_d 0.00213418f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_298_n X 0.0249747f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_c_292_n X 0.0145277f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_195 N_X_c_334_n N_VGND_c_354_n 0.0196893f $X=3.48 $Y=0.415 $X2=0 $Y2=0
cc_196 N_X_M1003_d N_VGND_c_355_n 0.00214967f $X=3.245 $Y=0.235 $X2=0 $Y2=0
cc_197 N_X_c_334_n N_VGND_c_355_n 0.0139935f $X=3.48 $Y=0.415 $X2=0 $Y2=0

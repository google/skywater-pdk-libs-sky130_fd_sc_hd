* File: sky130_fd_sc_hd__maj3_4.spice.pex
* Created: Thu Aug 27 14:27:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MAJ3_4%C 3 6 10 13 15 16 17 18 21 22 24 25 27 28 30
+ 34 36 39 41 45
c105 28 0 1.93111e-19 $X=2.78 $Y=1.16
c106 27 0 1.67168e-19 $X=2.78 $Y=1.16
c107 25 0 3.16076e-20 $X=2.63 $Y=1.16
c108 16 0 1.11508e-19 $X=0.805 $Y=1.915
r109 41 45 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.18 $X2=0.69
+ $Y2=1.18
r110 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.16
+ $X2=0.59 $Y2=1.325
r111 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.16
+ $X2=0.59 $Y2=0.995
r112 30 41 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.72 $Y2=1.18
r113 30 45 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.59 $Y=1.18 $X2=0.69
+ $Y2=1.18
r114 30 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r115 28 40 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.782 $Y=1.16
+ $X2=2.782 $Y2=1.325
r116 28 39 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.782 $Y=1.16
+ $X2=2.782 $Y2=0.995
r117 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.16 $X2=2.78 $Y2=1.16
r118 25 27 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.63 $Y=1.16
+ $X2=2.78 $Y2=1.16
r119 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.545 $Y=1.245
+ $X2=2.63 $Y2=1.16
r120 23 24 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.545 $Y=1.245
+ $X2=2.545 $Y2=2.225
r121 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=2.31
+ $X2=2.545 $Y2=2.225
r122 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.46 $Y=2.31
+ $X2=1.79 $Y2=2.31
r123 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=2.225
+ $X2=1.79 $Y2=2.31
r124 19 20 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.705 $Y=2.085
+ $X2=1.705 $Y2=2.225
r125 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=2
+ $X2=1.705 $Y2=2.085
r126 17 18 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.62 $Y=2 $X2=0.89
+ $Y2=2
r127 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=1.915
+ $X2=0.89 $Y2=2
r128 15 30 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=1.285
+ $X2=0.805 $Y2=1.18
r129 15 16 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.805 $Y=1.285
+ $X2=0.805 $Y2=1.915
r130 13 40 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.695 $Y=1.985
+ $X2=2.695 $Y2=1.325
r131 10 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.695 $Y=0.56
+ $X2=2.695 $Y2=0.995
r132 6 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.68 $Y=1.985
+ $X2=0.68 $Y2=1.325
r133 3 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.68 $Y=0.56
+ $X2=0.68 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_4%A 1 3 6 8 10 13 15 16 23 24
c43 23 0 6.74376e-20 $X=1.285 $Y=1.16
r44 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.285 $Y=1.16
+ $X2=1.495 $Y2=1.16
r45 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.285
+ $Y=1.16 $X2=1.285 $Y2=1.16
r46 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.075 $Y=1.16
+ $X2=1.285 $Y2=1.16
r47 15 16 10.0469 $w=3.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.255 $Y=1.19
+ $X2=1.255 $Y2=1.53
r48 15 23 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.255 $Y=1.19
+ $X2=1.255 $Y2=1.16
r49 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.325
+ $X2=1.495 $Y2=1.16
r50 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.495 $Y=1.325
+ $X2=1.495 $Y2=1.985
r51 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=1.16
r52 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r53 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.325
+ $X2=1.075 $Y2=1.16
r54 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.075 $Y=1.325
+ $X2=1.075 $Y2=1.985
r55 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=0.995
+ $X2=1.075 $Y2=1.16
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.075 $Y=0.995
+ $X2=1.075 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_4%B 1 3 6 8 10 13 15 22
c40 15 0 1.93111e-19 $X=2.065 $Y=1.19
c41 6 0 6.74376e-20 $X=1.915 $Y=1.985
r42 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.125 $Y=1.16
+ $X2=2.335 $Y2=1.16
r43 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.915 $Y=1.16
+ $X2=2.125 $Y2=1.16
r44 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.16 $X2=2.125 $Y2=1.16
r45 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.325
+ $X2=2.335 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.335 $Y=1.325
+ $X2=2.335 $Y2=1.985
r47 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=0.995
+ $X2=2.335 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.335 $Y=0.995
+ $X2=2.335 $Y2=0.56
r49 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.325
+ $X2=1.915 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.915 $Y=1.325
+ $X2=1.915 $Y2=1.985
r51 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_4%A_47_297# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 45 47 50 53 55 58 59 64 68 73 74 77 87
c168 87 0 1.67168e-19 $X=4.59 $Y=1.16
c169 50 0 1.32843e-19 $X=1.705 $Y=1.545
c170 13 0 1.56657e-19 $X=3.33 $Y=0.995
r171 84 85 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.75 $Y=1.16
+ $X2=4.17 $Y2=1.16
r172 73 74 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=1.62
+ $X2=0.275 $Y2=1.455
r173 71 74 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.17 $Y=0.885
+ $X2=0.17 $Y2=1.455
r174 70 71 8.70114 $w=5.48e-07 $l=1.13e-07 $layer=LI1_cond $X=0.36 $Y=0.772
+ $X2=0.36 $Y2=0.885
r175 68 70 8.52478 $w=5.48e-07 $l=3.92e-07 $layer=LI1_cond $X=0.36 $Y=0.38
+ $X2=0.36 $Y2=0.772
r176 65 87 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.38 $Y=1.16
+ $X2=4.59 $Y2=1.16
r177 65 85 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.38 $Y=1.16
+ $X2=4.17 $Y2=1.16
r178 64 65 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.38
+ $Y=1.16 $X2=4.38 $Y2=1.16
r179 62 84 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.54 $Y=1.16
+ $X2=3.75 $Y2=1.16
r180 62 81 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.54 $Y=1.16
+ $X2=3.33 $Y2=1.16
r181 61 64 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=3.54 $Y=1.18
+ $X2=4.38 $Y2=1.18
r182 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.16 $X2=3.54 $Y2=1.16
r183 59 61 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=3.285 $Y=1.18
+ $X2=3.54 $Y2=1.18
r184 58 59 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.2 $Y=1.075
+ $X2=3.285 $Y2=1.18
r185 57 58 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.2 $Y=0.885
+ $X2=3.2 $Y2=1.075
r186 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=0.8
+ $X2=3.2 $Y2=0.885
r187 55 77 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.115 $Y=0.8
+ $X2=2.29 $Y2=0.8
r188 51 77 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0.772
+ $X2=2.29 $Y2=0.772
r189 51 75 21.5123 $w=2.23e-07 $l=4.2e-07 $layer=LI1_cond $X=2.125 $Y=0.772
+ $X2=1.705 $Y2=0.772
r190 51 53 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.125 $Y=0.66
+ $X2=2.125 $Y2=0.38
r191 50 80 14.5568 $w=3.52e-07 $l=5.70526e-07 $layer=LI1_cond $X=1.705 $Y=1.545
+ $X2=2.125 $Y2=1.9
r192 49 75 2.38091 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.705 $Y=0.885
+ $X2=1.705 $Y2=0.772
r193 49 50 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.705 $Y=0.885
+ $X2=1.705 $Y2=1.545
r194 48 70 6.02202 $w=2.25e-07 $l=2.75e-07 $layer=LI1_cond $X=0.635 $Y=0.772
+ $X2=0.36 $Y2=0.772
r195 47 75 4.35367 $w=2.23e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.772
+ $X2=1.705 $Y2=0.772
r196 47 48 50.4514 $w=2.23e-07 $l=9.85e-07 $layer=LI1_cond $X=1.62 $Y=0.772
+ $X2=0.635 $Y2=0.772
r197 43 73 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.275 $Y=1.645
+ $X2=0.275 $Y2=1.62
r198 43 45 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=0.275 $Y=1.645
+ $X2=0.275 $Y2=2.3
r199 37 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.16
r200 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.985
r201 34 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=1.16
r202 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=0.56
r203 30 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.325
+ $X2=4.17 $Y2=1.16
r204 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.17 $Y=1.325
+ $X2=4.17 $Y2=1.985
r205 27 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=0.995
+ $X2=4.17 $Y2=1.16
r206 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.17 $Y=0.995
+ $X2=4.17 $Y2=0.56
r207 23 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.75 $Y=1.325
+ $X2=3.75 $Y2=1.16
r208 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.75 $Y=1.325
+ $X2=3.75 $Y2=1.985
r209 20 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.75 $Y=0.995
+ $X2=3.75 $Y2=1.16
r210 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.75 $Y=0.995
+ $X2=3.75 $Y2=0.56
r211 16 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.325
+ $X2=3.33 $Y2=1.16
r212 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.33 $Y=1.325
+ $X2=3.33 $Y2=1.985
r213 13 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=0.995
+ $X2=3.33 $Y2=1.16
r214 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.33 $Y=0.995
+ $X2=3.33 $Y2=0.56
r215 4 80 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.99
+ $Y=1.485 $X2=2.125 $Y2=1.63
r216 3 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.485 $X2=0.38 $Y2=1.62
r217 3 45 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.485 $X2=0.38 $Y2=2.3
r218 2 53 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.235 $X2=2.125 $Y2=0.38
r219 1 68 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.325
+ $Y=0.235 $X2=0.47 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_4%VPWR 1 2 3 4 15 19 23 27 29 31 33 35 40 48 54
+ 57 60 64 68
r81 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r82 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r83 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r84 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r85 55 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.23 $Y2=2.72
r86 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 52 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r88 52 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r89 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r90 49 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=2.72
+ $X2=3.96 $Y2=2.72
r91 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.045 $Y=2.72
+ $X2=4.37 $Y2=2.72
r92 48 63 3.67103 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.887 $Y2=2.72
r93 48 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.37 $Y2=2.72
r94 47 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r95 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r96 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r97 44 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 43 46 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r99 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r100 41 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.285 $Y2=2.72
r101 41 43 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.61 $Y2=2.72
r102 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=3.01 $Y2=2.72
r103 40 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.53 $Y2=2.72
r104 37 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r105 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=2.72
+ $X2=1.285 $Y2=2.72
r106 35 37 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.12 $Y=2.72
+ $X2=0.23 $Y2=2.72
r107 33 68 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r108 29 63 3.24416 $w=2.1e-07 $l=1.13666e-07 $layer=LI1_cond $X=4.82 $Y=2.635
+ $X2=4.887 $Y2=2.72
r109 29 31 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=4.82 $Y=2.635
+ $X2=4.82 $Y2=1.96
r110 25 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=2.635
+ $X2=3.96 $Y2=2.72
r111 25 27 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.96 $Y=2.635
+ $X2=3.96 $Y2=1.96
r112 24 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=2.72
+ $X2=3.01 $Y2=2.72
r113 23 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=2.72
+ $X2=3.96 $Y2=2.72
r114 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.875 $Y=2.72
+ $X2=3.175 $Y2=2.72
r115 19 22 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=3.01 $Y=1.62
+ $X2=3.01 $Y2=2.34
r116 17 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=2.635
+ $X2=3.01 $Y2=2.72
r117 17 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.01 $Y=2.635
+ $X2=3.01 $Y2=2.34
r118 13 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.72
r119 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.34
r120 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=1.485 $X2=4.8 $Y2=1.96
r121 3 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.825
+ $Y=1.485 $X2=3.96 $Y2=1.96
r122 2 22 400 $w=1.7e-07 $l=9.67587e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.485 $X2=3.01 $Y2=2.34
r123 2 19 400 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=2.77 $Y=1.485
+ $X2=3.01 $Y2=1.62
r124 1 15 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.485 $X2=1.285 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_4%X 1 2 3 4 13 15 18 19 21 25 29 32 39 40 41 47
+ 48
c72 18 0 1.56657e-19 $X=3.58 $Y=0.715
r73 41 48 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.825 $Y=1.54
+ $X2=4.845 $Y2=1.54
r74 41 59 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.825 $Y=1.54
+ $X2=4.38 $Y2=1.54
r75 41 48 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=4.845 $Y=1.45
+ $X2=4.845 $Y2=1.455
r76 40 41 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=4.845 $Y=1.19
+ $X2=4.845 $Y2=1.45
r77 39 47 1.16746 $w=1.88e-07 $l=2e-08 $layer=LI1_cond $X=4.825 $Y=0.81
+ $X2=4.845 $Y2=0.81
r78 39 40 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=4.845 $Y=0.92
+ $X2=4.845 $Y2=1.19
r79 39 47 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=4.845 $Y=0.92
+ $X2=4.845 $Y2=0.905
r80 32 34 3.84769 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=0.4 $X2=3.54
+ $Y2=0.49
r81 29 59 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=4.38 $Y=2.34
+ $X2=4.38 $Y2=1.625
r82 23 39 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=4.38 $Y=0.81
+ $X2=4.825 $Y2=0.81
r83 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.38 $Y=0.715
+ $X2=4.38 $Y2=0.4
r84 22 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=1.54
+ $X2=3.54 $Y2=1.54
r85 21 59 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=1.54
+ $X2=4.38 $Y2=1.54
r86 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.215 $Y=1.54
+ $X2=3.705 $Y2=1.54
r87 20 38 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.705 $Y=0.81
+ $X2=3.58 $Y2=0.81
r88 19 23 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=0.81
+ $X2=4.38 $Y2=0.81
r89 19 20 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=4.215 $Y=0.81
+ $X2=3.705 $Y2=0.81
r90 18 38 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=3.58 $Y=0.715
+ $X2=3.58 $Y2=0.81
r91 18 34 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.58 $Y=0.715
+ $X2=3.58 $Y2=0.49
r92 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=1.625 $X2=3.54
+ $Y2=1.54
r93 13 15 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=3.54 $Y=1.625
+ $X2=3.54 $Y2=2.34
r94 4 59 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.485 $X2=4.38 $Y2=1.62
r95 4 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.485 $X2=4.38 $Y2=2.34
r96 3 36 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.54 $Y2=1.62
r97 3 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.54 $Y2=2.34
r98 2 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.245
+ $Y=0.235 $X2=4.38 $Y2=0.4
r99 1 38 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.235 $X2=3.54 $Y2=0.74
r100 1 32 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.235 $X2=3.54 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_4%VGND 1 2 3 4 15 19 21 25 27 29 31 33 38 46 52
+ 55 58 62 66
r79 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r80 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r81 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r82 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r83 53 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.23
+ $Y2=0
r84 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r85 50 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r86 50 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r87 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r88 47 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=0 $X2=3.96
+ $Y2=0
r89 47 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.045 $Y=0 $X2=4.37
+ $Y2=0
r90 46 61 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.887
+ $Y2=0
r91 46 49 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.37
+ $Y2=0
r92 45 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r93 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r94 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r95 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r96 41 44 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r97 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r98 39 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.285
+ $Y2=0
r99 39 41 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.61
+ $Y2=0
r100 38 55 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=3.032
+ $Y2=0
r101 38 44 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.53
+ $Y2=0
r102 35 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r103 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.285
+ $Y2=0
r104 33 35 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.23
+ $Y2=0
r105 31 66 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0
+ $X2=0.23 $Y2=0
r106 27 61 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.8 $Y=0.085
+ $X2=4.887 $Y2=0
r107 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.8 $Y=0.085
+ $X2=4.8 $Y2=0.38
r108 23 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0
r109 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0.38
r110 22 55 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.205 $Y=0
+ $X2=3.032 $Y2=0
r111 21 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.96
+ $Y2=0
r112 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.875 $Y=0
+ $X2=3.205 $Y2=0
r113 17 55 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.032 $Y=0.085
+ $X2=3.032 $Y2=0
r114 17 19 9.85422 $w=3.43e-07 $l=2.95e-07 $layer=LI1_cond $X=3.032 $Y=0.085
+ $X2=3.032 $Y2=0.38
r115 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.085
+ $X2=1.285 $Y2=0
r116 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.285 $Y=0.085
+ $X2=1.285 $Y2=0.38
r117 4 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.665
+ $Y=0.235 $X2=4.8 $Y2=0.38
r118 3 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.825
+ $Y=0.235 $X2=3.96 $Y2=0.38
r119 2 19 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.235 $X2=3.025 $Y2=0.38
r120 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.235 $X2=1.285 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_16.spice
* Created: Thu Aug 27 14:23:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_16.spice.pex"
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_16  VNB VPB A KAPWR X VGND VPWR
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_A_110_47#_M1012_d N_A_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75008.4
+ A=0.063 P=1.14 MULT=1
MM1022 N_A_110_47#_M1012_d N_A_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75007.9
+ A=0.063 P=1.14 MULT=1
MM1026 N_A_110_47#_M1026_d N_A_M1026_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75007.5
+ A=0.063 P=1.14 MULT=1
MM1039 N_A_110_47#_M1026_d N_A_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75007.1
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1039_s N_A_110_47#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75006.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_110_47#_M1003_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75006.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1003_d N_A_110_47#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75005.8
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_110_47#_M1007_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75005.3
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1007_d N_A_110_47#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.6 SB=75004.9
+ A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_110_47#_M1015_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.1 SB=75004.5
+ A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1015_d N_A_110_47#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.5 SB=75004.1
+ A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_110_47#_M1018_g N_X_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.0588 PD=0.695 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.9
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1018_d N_A_110_47#_M1020_g N_X_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.0588 PD=0.695 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.3
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_110_47#_M1023_g N_X_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.8 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1023_d N_A_110_47#_M1029_g N_X_M1029_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_110_47#_M1031_g N_X_M1029_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1031_d N_A_110_47#_M1032_g N_X_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.1 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_A_110_47#_M1033_g N_X_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.5 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1033_d N_A_110_47#_M1036_g N_X_M1036_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.9 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_110_47#_M1037_g N_X_M1036_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75008.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_KAPWR_M1009_d N_A_M1009_g N_A_110_47#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75008.4 A=0.15 P=2.3 MULT=1
MM1019 N_KAPWR_M1019_d N_A_M1019_g N_A_110_47#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75007.9 A=0.15 P=2.3 MULT=1
MM1021 N_KAPWR_M1019_d N_A_M1021_g N_A_110_47#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75007.5
+ A=0.15 P=2.3 MULT=1
MM1038 N_KAPWR_M1038_d N_A_M1038_g N_A_110_47#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75007.1 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_110_47#_M1000_g N_KAPWR_M1038_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1000_d N_A_110_47#_M1001_g N_KAPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75006.2 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_110_47#_M1005_g N_KAPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75005.8 A=0.15 P=2.3 MULT=1
MM1006 N_X_M1005_d N_A_110_47#_M1006_g N_KAPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1010_d N_A_110_47#_M1010_g N_KAPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1010_d N_A_110_47#_M1011_g N_KAPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1013_d N_A_110_47#_M1013_g N_KAPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1014 N_X_M1013_d N_A_110_47#_M1014_g N_KAPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1375 PD=1.28 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.9
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1016 N_X_M1016_d N_A_110_47#_M1016_g N_KAPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1375 PD=1.28 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.3
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1024 N_X_M1016_d N_A_110_47#_M1024_g N_KAPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.8
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1025 N_X_M1025_d N_A_110_47#_M1025_g N_KAPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1027 N_X_M1025_d N_A_110_47#_M1027_g N_KAPWR_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1028 N_X_M1028_d N_A_110_47#_M1028_g N_KAPWR_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1030 N_X_M1028_d N_A_110_47#_M1030_g N_KAPWR_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.5 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1034 N_X_M1034_d N_A_110_47#_M1034_g N_KAPWR_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1035 N_X_M1034_d N_A_110_47#_M1035_g N_KAPWR_M1035_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=15.3759 P=22.37
*
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_16.spice.SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__o31a_2.spice.pex
* Created: Thu Aug 27 14:39:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O31A_2%A_108_21# 1 2 7 9 12 14 16 18 21 23 26 27 29
+ 30 32 33 34 35 36 37 40 44
c108 40 0 1.67512e-19 $X=3.51 $Y=1.495
c109 27 0 2.02454e-20 $X=1.115 $Y=1.16
c110 26 0 8.42142e-20 $X=1.115 $Y=1.16
r111 44 46 16.8246 $w=4.83e-07 $l=4.65e-07 $layer=LI1_cond $X=3.352 $Y=0.36
+ $X2=3.352 $Y2=0.825
r112 40 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.51 $Y=1.495
+ $X2=3.51 $Y2=0.825
r113 38 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.08 $Y=1.58
+ $X2=2.955 $Y2=1.58
r114 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=1.58
+ $X2=3.51 $Y2=1.495
r115 37 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.425 $Y=1.58
+ $X2=3.08 $Y2=1.58
r116 35 42 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=1.665
+ $X2=2.955 $Y2=1.58
r117 35 36 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=2.955 $Y=1.665
+ $X2=2.955 $Y2=2.295
r118 33 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.83 $Y=2.38
+ $X2=2.955 $Y2=2.295
r119 33 34 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.83 $Y=2.38
+ $X2=1.82 $Y2=2.38
r120 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.735 $Y=2.295
+ $X2=1.82 $Y2=2.38
r121 31 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.735 $Y=1.615
+ $X2=1.735 $Y2=2.295
r122 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.65 $Y=1.53
+ $X2=1.735 $Y2=1.615
r123 29 30 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.65 $Y=1.53
+ $X2=1.2 $Y2=1.53
r124 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.16 $X2=1.115 $Y2=1.16
r125 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=1.445
+ $X2=1.2 $Y2=1.53
r126 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.115 $Y=1.445
+ $X2=1.115 $Y2=1.16
r127 19 27 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=1.115 $Y=1.325
+ $X2=1.145 $Y2=1.16
r128 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.115 $Y=1.325
+ $X2=1.115 $Y2=1.985
r129 16 27 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=1.115 $Y=0.995
+ $X2=1.145 $Y2=1.16
r130 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.115 $Y=0.995
+ $X2=1.115 $Y2=0.56
r131 15 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.69 $Y=1.16
+ $X2=0.615 $Y2=1.16
r132 14 27 5.03009 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.04 $Y=1.16
+ $X2=1.145 $Y2=1.16
r133 14 15 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.04 $Y=1.16
+ $X2=0.69 $Y2=1.16
r134 10 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.325
+ $X2=0.615 $Y2=1.16
r135 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.615 $Y=1.325
+ $X2=0.615 $Y2=1.985
r136 7 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=1.16
r137 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=0.56
r138 2 42 300 $w=1.7e-07 $l=3.62077e-07 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=1.485 $X2=2.915 $Y2=1.66
r139 1 44 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=3.11
+ $Y=0.235 $X2=3.275 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%A1 3 6 8 11 13
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.16
+ $X2=1.595 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.16
+ $X2=1.595 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.16 $X2=1.595 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.655 $Y=1.985
+ $X2=1.655 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.655 $Y=0.56
+ $X2=1.655 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%A2 1 3 6 8 9 10 15
c36 15 0 1.90303e-19 $X=2.075 $Y=1.16
r37 9 10 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.09 $Y=1.53 $X2=2.09
+ $Y2=1.87
r38 9 26 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=2.09 $Y=1.53
+ $X2=2.09 $Y2=1.325
r39 8 26 8.18414 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.067 $Y=1.16
+ $X2=2.067 $Y2=1.325
r40 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.16 $X2=2.075 $Y2=1.16
r41 4 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.325
+ $X2=2.075 $Y2=1.16
r42 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.075 $Y=1.325
+ $X2=2.075 $Y2=1.985
r43 1 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=0.995
+ $X2=2.075 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.075 $Y=0.995
+ $X2=2.075 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%A3 1 3 6 8 11
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.555
+ $Y=1.16 $X2=2.555 $Y2=1.16
r36 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=1.16
r37 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=1.985
r38 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=0.995
+ $X2=2.555 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.555 $Y=0.995
+ $X2=2.555 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%B1 3 6 8 11 13
r33 11 14 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.052 $Y=1.16
+ $X2=3.052 $Y2=1.325
r34 11 13 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.052 $Y=1.16
+ $X2=3.052 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=1.16 $X2=3.035 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.13 $Y=1.985
+ $X2=3.13 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.035 $Y=0.56
+ $X2=3.035 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%VPWR 1 2 3 10 12 18 20 22 25 26 27 33 45
c47 18 0 2.02454e-20 $X=1.385 $Y=1.96
c48 3 0 1.67512e-19 $X=3.205 $Y=1.485
r49 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 36 39 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 35 38 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 33 44 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=3.467 $Y2=2.72
r56 33 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 32 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r58 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 29 41 4.4818 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=2.72 $X2=0.19
+ $Y2=2.72
r60 29 31 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.38 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 27 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 27 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 25 31 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 25 26 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.322 $Y2=2.72
r65 24 35 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.48 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 24 26 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.48 $Y=2.72
+ $X2=1.322 $Y2=2.72
r67 20 44 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.422 $Y=2.635
+ $X2=3.467 $Y2=2.72
r68 20 22 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=3.422 $Y=2.635
+ $X2=3.422 $Y2=1.96
r69 16 26 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.322 $Y=2.635
+ $X2=1.322 $Y2=2.72
r70 16 18 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=1.322 $Y=2.635
+ $X2=1.322 $Y2=1.96
r71 12 15 27.7368 $w=2.93e-07 $l=7.1e-07 $layer=LI1_cond $X=0.232 $Y=1.63
+ $X2=0.232 $Y2=2.34
r72 10 41 2.99573 $w=2.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.232 $Y=2.635
+ $X2=0.19 $Y2=2.72
r73 10 15 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.232 $Y=2.635
+ $X2=0.232 $Y2=2.34
r74 3 22 300 $w=1.7e-07 $l=5.72495e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=1.485 $X2=3.42 $Y2=1.96
r75 2 18 300 $w=1.7e-07 $l=5.64137e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=1.485 $X2=1.385 $Y2=1.96
r76 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r77 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%X 1 2 7 8 9 10 11 12 13 23 30 38 47
r33 47 48 1.93707 $w=4.38e-07 $l=3.5e-08 $layer=LI1_cond $X=0.77 $Y=1.87
+ $X2=0.77 $Y2=1.835
r34 30 43 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.705 $Y=0.85
+ $X2=0.705 $Y2=0.825
r35 13 51 6.54797 $w=4.38e-07 $l=2.5e-07 $layer=LI1_cond $X=0.77 $Y=2.21
+ $X2=0.77 $Y2=1.96
r36 12 51 1.70247 $w=4.38e-07 $l=6.5e-08 $layer=LI1_cond $X=0.77 $Y=1.895
+ $X2=0.77 $Y2=1.96
r37 12 47 0.654797 $w=4.38e-07 $l=2.5e-08 $layer=LI1_cond $X=0.77 $Y=1.895
+ $X2=0.77 $Y2=1.87
r38 12 48 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.705 $Y=1.81
+ $X2=0.705 $Y2=1.835
r39 11 12 10.4092 $w=3.08e-07 $l=2.8e-07 $layer=LI1_cond $X=0.705 $Y=1.53
+ $X2=0.705 $Y2=1.81
r40 11 32 8.73626 $w=3.08e-07 $l=2.35e-07 $layer=LI1_cond $X=0.705 $Y=1.53
+ $X2=0.705 $Y2=1.295
r41 10 23 2.602 $w=2.2e-07 $l=1.55e-07 $layer=LI1_cond $X=0.705 $Y=1.185
+ $X2=0.55 $Y2=1.185
r42 10 28 3.84985 $w=3.1e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=1.185
+ $X2=0.705 $Y2=1.075
r43 10 32 3.84985 $w=3.1e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=1.185
+ $X2=0.705 $Y2=1.295
r44 9 43 1.80611 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=0.77 $Y=0.795 $X2=0.77
+ $Y2=0.825
r45 9 28 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=0.705 $Y=0.88
+ $X2=0.705 $Y2=1.075
r46 9 30 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=0.705 $Y=0.88 $X2=0.705
+ $Y2=0.85
r47 8 9 7.46469 $w=4.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.77 $Y=0.51 $X2=0.77
+ $Y2=0.795
r48 8 38 3.92878 $w=4.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.77 $Y=0.51 $X2=0.77
+ $Y2=0.36
r49 7 23 16.5009 $w=2.18e-07 $l=3.15e-07 $layer=LI1_cond $X=0.235 $Y=1.185
+ $X2=0.55 $Y2=1.185
r50 2 51 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=1.485 $X2=0.825 $Y2=1.96
r51 1 38 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=0.69
+ $Y=0.235 $X2=0.825 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%VGND 1 2 3 10 12 16 19 20 21 27 33 34 41
r55 41 44 9.87808 $w=4.18e-07 $l=3.6e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.33
+ $Y2=0.36
r56 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r57 34 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r58 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r59 31 41 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.33
+ $Y2=0
r60 31 33 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=3.45
+ $Y2=0
r61 30 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r62 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 27 41 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.33
+ $Y2=0
r64 27 29 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.07
+ $Y2=0
r65 26 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r66 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 23 37 4.4818 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r68 23 25 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=1.15
+ $Y2=0
r69 21 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r70 21 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 19 25 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.15
+ $Y2=0
r72 19 20 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.385
+ $Y2=0
r73 18 29 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r74 18 20 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.385
+ $Y2=0
r75 14 20 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=0.085
+ $X2=1.385 $Y2=0
r76 14 16 7.30937 $w=4.48e-07 $l=2.75e-07 $layer=LI1_cond $X=1.385 $Y=0.085
+ $X2=1.385 $Y2=0.36
r77 10 37 2.99573 $w=2.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.232 $Y=0.085
+ $X2=0.19 $Y2=0
r78 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.232 $Y=0.085
+ $X2=0.232 $Y2=0.38
r79 3 44 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.235 $X2=2.315 $Y2=0.36
r80 2 16 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=1.19
+ $Y=0.235 $X2=1.385 $Y2=0.36
r81 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_2%A_346_47# 1 2 7 10 11 12
c23 11 0 1.90303e-19 $X=1.95 $Y=0.74
r24 12 14 5.03913 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.825 $Y=0.655
+ $X2=2.825 $Y2=0.56
r25 10 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.71 $Y=0.74
+ $X2=2.825 $Y2=0.655
r26 10 11 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.71 $Y=0.74
+ $X2=1.95 $Y2=0.74
r27 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=0.655
+ $X2=1.95 $Y2=0.74
r28 7 9 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.865 $Y=0.655
+ $X2=1.865 $Y2=0.56
r29 2 14 182 $w=1.7e-07 $l=3.99061e-07 $layer=licon1_NDIFF $count=1 $X=2.63
+ $Y=0.235 $X2=2.795 $Y2=0.56
r30 1 9 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.73
+ $Y=0.235 $X2=1.865 $Y2=0.56
.ends


* NGSPICE file created from sky130_fd_sc_hd__nand3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
M1000 a_218_47# B a_408_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=5.135e+11p ps=5.48e+06u
M1001 VPWR B Y VPB phighvt w=1e+06u l=150000u
+  ad=1.4015e+12p pd=1.289e+07u as=8.1e+11p ps=7.62e+06u
M1002 a_408_47# B a_218_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 VGND C a_218_47# VNB nshort w=650000u l=150000u
+  ad=4.085e+11p pd=3.91e+06u as=0p ps=0u
M1006 a_408_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1007 VPWR C Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_218_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_47# a_408_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_47# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends


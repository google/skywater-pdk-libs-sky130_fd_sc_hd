* File: sky130_fd_sc_hd__a311o_2.spice.SKY130_FD_SC_HD__A311O_2.pxi
* Created: Thu Aug 27 14:04:01 2020
* 
x_PM_SKY130_FD_SC_HD__A311O_2%A_79_21# N_A_79_21#_M1001_d N_A_79_21#_M1006_d
+ N_A_79_21#_M1000_d N_A_79_21#_c_58_n N_A_79_21#_M1007_g N_A_79_21#_M1004_g
+ N_A_79_21#_c_59_n N_A_79_21#_M1012_g N_A_79_21#_M1010_g N_A_79_21#_c_60_n
+ N_A_79_21#_c_61_n N_A_79_21#_c_71_p N_A_79_21#_c_141_p N_A_79_21#_c_68_p
+ N_A_79_21#_c_114_p N_A_79_21#_c_82_p N_A_79_21#_c_73_p N_A_79_21#_c_83_p
+ N_A_79_21#_c_98_p N_A_79_21#_c_102_p N_A_79_21#_c_99_p N_A_79_21#_c_158_p
+ N_A_79_21#_c_122_p PM_SKY130_FD_SC_HD__A311O_2%A_79_21#
x_PM_SKY130_FD_SC_HD__A311O_2%A3 N_A3_M1002_g N_A3_M1011_g A3 N_A3_c_174_n
+ N_A3_c_175_n PM_SKY130_FD_SC_HD__A311O_2%A3
x_PM_SKY130_FD_SC_HD__A311O_2%A2 N_A2_M1009_g N_A2_M1005_g A2 N_A2_c_214_n
+ N_A2_c_215_n PM_SKY130_FD_SC_HD__A311O_2%A2
x_PM_SKY130_FD_SC_HD__A311O_2%A1 N_A1_M1001_g N_A1_M1013_g A1 N_A1_c_250_n
+ N_A1_c_251_n PM_SKY130_FD_SC_HD__A311O_2%A1
x_PM_SKY130_FD_SC_HD__A311O_2%B1 N_B1_M1008_g N_B1_M1003_g B1 N_B1_c_285_n
+ N_B1_c_286_n N_B1_c_287_n PM_SKY130_FD_SC_HD__A311O_2%B1
x_PM_SKY130_FD_SC_HD__A311O_2%C1 N_C1_M1006_g N_C1_M1000_g C1 N_C1_c_317_n
+ N_C1_c_318_n PM_SKY130_FD_SC_HD__A311O_2%C1
x_PM_SKY130_FD_SC_HD__A311O_2%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1005_d
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n VPWR N_VPWR_c_348_n
+ N_VPWR_c_339_n PM_SKY130_FD_SC_HD__A311O_2%VPWR
x_PM_SKY130_FD_SC_HD__A311O_2%X N_X_M1007_s N_X_M1004_s X X X X X X N_X_c_397_n
+ PM_SKY130_FD_SC_HD__A311O_2%X
x_PM_SKY130_FD_SC_HD__A311O_2%A_319_297# N_A_319_297#_M1011_d
+ N_A_319_297#_M1013_d N_A_319_297#_c_414_n N_A_319_297#_c_418_n
+ N_A_319_297#_c_415_n N_A_319_297#_c_416_n N_A_319_297#_c_421_n
+ PM_SKY130_FD_SC_HD__A311O_2%A_319_297#
x_PM_SKY130_FD_SC_HD__A311O_2%VGND N_VGND_M1007_d N_VGND_M1012_d N_VGND_M1008_d
+ N_VGND_c_438_n N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n VGND
+ N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n
+ N_VGND_c_447_n PM_SKY130_FD_SC_HD__A311O_2%VGND
cc_1 VNB N_A_79_21#_c_58_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_59_n 0.0173524f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_60_n 0.0017627f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.16
cc_4 VNB N_A_79_21#_c_61_n 0.0612097f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.16
cc_5 VNB N_A3_c_174_n 0.0223052f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_6 VNB N_A3_c_175_n 0.0187184f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_7 VNB A2 0.00398814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_214_n 0.0213583f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_9 VNB N_A2_c_215_n 0.0166976f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_10 VNB A1 0.00522468f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB N_A1_c_250_n 0.0222552f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_12 VNB N_A1_c_251_n 0.0172419f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_13 VNB N_B1_c_285_n 0.0223968f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_14 VNB N_B1_c_286_n 0.00314824f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB N_B1_c_287_n 0.0189953f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_16 VNB C1 0.0133916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C1_c_317_n 0.0298364f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_18 VNB N_C1_c_318_n 0.0235626f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_19 VNB N_VPWR_c_339_n 0.17485f $X=-0.19 $Y=-0.24 $X2=3.88 $Y2=0.42
cc_20 VNB N_VGND_c_438_n 0.00997672f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_21 VNB N_VGND_c_439_n 0.0331381f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_22 VNB N_VGND_c_440_n 0.00506574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_441_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_24 VNB N_VGND_c_442_n 0.0184034f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=0.825
cc_25 VNB N_VGND_c_443_n 0.0438139f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.74
cc_26 VNB N_VGND_c_444_n 0.0182832f $X=-0.19 $Y=-0.24 $X2=2.875 $Y2=0.57
cc_27 VNB N_VGND_c_445_n 0.219751f $X=-0.19 $Y=-0.24 $X2=2.875 $Y2=0.57
cc_28 VNB N_VGND_c_446_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_447_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=3.88 $Y2=1.96
cc_30 VPB N_A_79_21#_M1004_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_31 VPB N_A_79_21#_M1010_g 0.0200354f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_32 VPB N_A_79_21#_c_60_n 0.00256655f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_33 VPB N_A_79_21#_c_61_n 0.0143985f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_34 VPB N_A3_M1011_g 0.0218732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A3_c_174_n 0.00414182f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_36 VPB N_A2_M1005_g 0.0209847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A2 0.00122755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A2_c_214_n 0.00436976f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_39 VPB N_A1_M1013_g 0.0217366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB A1 9.1039e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_41 VPB N_A1_c_250_n 0.00439161f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_42 VPB N_B1_M1003_g 0.022223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B1_c_285_n 0.00414456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_44 VPB N_B1_c_286_n 0.00124017f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_45 VPB N_C1_M1000_g 0.0278425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB C1 0.0026577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_C1_c_317_n 0.00572067f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_48 VPB N_VPWR_c_340_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_49 VPB N_VPWR_c_341_n 0.0431432f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_50 VPB N_VPWR_c_342_n 0.00502493f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_51 VPB N_VPWR_c_343_n 0.00561515f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_52 VPB N_VPWR_c_344_n 0.0230176f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.495
cc_53 VPB N_VPWR_c_345_n 0.00420575f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_54 VPB N_VPWR_c_346_n 0.0200876f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_55 VPB N_VPWR_c_347_n 0.00631443f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.74
cc_56 VPB N_VPWR_c_348_n 0.0502786f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=0.655
cc_57 VPB N_VPWR_c_339_n 0.044982f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=0.42
cc_58 N_A_79_21#_M1010_g N_A3_M1011_g 0.0240362f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_60_n N_A3_M1011_g 0.00342104f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_79_21#_c_68_p N_A3_M1011_g 0.0166179f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_60_n A3 0.0140465f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_61_n A3 0.00126615f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_71_p A3 0.0132681f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_68_p A3 0.0135626f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_73_p A3 4.14162e-19 $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_60_n N_A3_c_174_n 0.00107425f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_61_n N_A3_c_174_n 0.0214547f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_71_p N_A3_c_174_n 0.00214908f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_68_p N_A3_c_174_n 0.00264114f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_73_p N_A3_c_174_n 3.68129e-19 $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_59_n N_A3_c_175_n 0.01685f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_60_n N_A3_c_175_n 0.00342104f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_71_p N_A3_c_175_n 0.0109942f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_82_p N_A3_c_175_n 0.00662151f $X=1.61 $Y=0.655 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_83_p N_A3_c_175_n 0.00525832f $X=1.695 $Y=0.34 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_68_p N_A2_M1005_g 0.0111977f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_68_p A2 0.017476f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_73_p A2 0.0118015f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_68_p N_A2_c_214_n 0.00197275f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_73_p N_A2_c_214_n 0.00119993f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_71_p N_A2_c_215_n 6.70141e-19 $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_82_p N_A2_c_215_n 0.00365704f $X=1.61 $Y=0.655 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_73_p N_A2_c_215_n 0.0104978f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_68_p N_A1_M1013_g 0.0115635f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_68_p A1 0.0152527f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_73_p A1 0.0111258f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_68_p N_A1_c_250_n 0.00227792f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_73_p N_A1_c_250_n 0.00141243f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_73_p N_A1_c_251_n 0.0105433f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_98_p N_A1_c_251_n 0.00403733f $X=2.875 $Y=0.57 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_99_p N_A1_c_251_n 7.22281e-19 $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_68_p N_B1_M1003_g 0.0163705f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_68_p N_B1_c_285_n 0.00258743f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_102_p N_B1_c_285_n 0.00285103f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_68_p N_B1_c_286_n 0.0210947f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_102_p N_B1_c_286_n 0.0161005f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_99_p N_B1_c_286_n 0.0054721f $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_102_p N_B1_c_287_n 0.0112997f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_68_p N_C1_M1000_g 0.018342f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_68_p C1 0.0193768f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_102_p C1 0.019189f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_68_p N_C1_c_317_n 0.00277415f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_102_p N_C1_c_317_n 0.00275628f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_102_p N_C1_c_318_n 0.0152672f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_68_p N_VPWR_M1010_d 0.00684331f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_114_p N_VPWR_M1010_d 0.00795071f $X=1.185 $Y=1.58 $X2=0
+ $Y2=0
cc_107 N_A_79_21#_c_68_p N_VPWR_M1005_d 0.0108392f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_79_21#_M1004_g N_VPWR_c_341_n 0.00450113f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_79_21#_M1010_g N_VPWR_c_342_n 0.0088938f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_68_p N_VPWR_c_342_n 0.0157471f $X=3.795 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_114_p N_VPWR_c_342_n 0.0021188f $X=1.185 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A_79_21#_M1004_g N_VPWR_c_344_n 0.00542953f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_79_21#_M1010_g N_VPWR_c_344_n 0.00542953f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_79_21#_c_122_p N_VPWR_c_348_n 0.0116048f $X=3.88 $Y=1.96 $X2=0 $Y2=0
cc_115 N_A_79_21#_M1000_d N_VPWR_c_339_n 0.00525232f $X=3.745 $Y=1.485 $X2=0
+ $Y2=0
cc_116 N_A_79_21#_M1004_g N_VPWR_c_339_n 0.0104585f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_79_21#_M1010_g N_VPWR_c_339_n 0.0101795f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_122_p N_VPWR_c_339_n 0.00646998f $X=3.88 $Y=1.96 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_58_n N_X_c_397_n 0.0128056f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_79_21#_M1004_g N_X_c_397_n 0.0197519f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_59_n N_X_c_397_n 0.0110976f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_79_21#_M1010_g N_X_c_397_n 0.0178012f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_60_n N_X_c_397_n 0.0463319f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_61_n N_X_c_397_n 0.0325857f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_68_p N_A_319_297#_M1011_d 0.00916616f $X=3.795 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_126 N_A_79_21#_c_68_p N_A_319_297#_M1013_d 0.00983405f $X=3.795 $Y=1.58 $X2=0
+ $Y2=0
cc_127 N_A_79_21#_c_68_p N_A_319_297#_c_414_n 0.0155382f $X=3.795 $Y=1.58 $X2=0
+ $Y2=0
cc_128 N_A_79_21#_c_68_p N_A_319_297#_c_415_n 0.0454313f $X=3.795 $Y=1.58 $X2=0
+ $Y2=0
cc_129 N_A_79_21#_c_68_p N_A_319_297#_c_416_n 0.0204563f $X=3.795 $Y=1.58 $X2=0
+ $Y2=0
cc_130 N_A_79_21#_c_68_p A_635_297# 0.0179778f $X=3.795 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_79_21#_c_60_n N_VGND_M1012_d 7.32946e-19 $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_71_p N_VGND_M1012_d 0.00691221f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_141_p N_VGND_M1012_d 0.0032487f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_102_p N_VGND_M1008_d 0.00974295f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_79_21#_c_58_n N_VGND_c_439_n 0.00321527f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_59_n N_VGND_c_440_n 0.00337722f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_61_n N_VGND_c_440_n 7.26766e-19 $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_71_p N_VGND_c_440_n 0.011029f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_141_p N_VGND_c_440_n 0.0125012f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_82_p N_VGND_c_440_n 0.00279984f $X=1.61 $Y=0.655 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_83_p N_VGND_c_440_n 0.0133992f $X=1.695 $Y=0.34 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_102_p N_VGND_c_441_n 0.0242585f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_58_n N_VGND_c_442_n 0.00542953f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_59_n N_VGND_c_442_n 0.00542953f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_71_p N_VGND_c_443_n 0.00248434f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_73_p N_VGND_c_443_n 0.0741173f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_83_p N_VGND_c_443_n 0.00971947f $X=1.695 $Y=0.34 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_102_p N_VGND_c_443_n 0.00334994f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_79_21#_c_102_p N_VGND_c_444_n 0.00321699f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_79_21#_c_158_p N_VGND_c_444_n 0.011459f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_151 N_A_79_21#_M1001_d N_VGND_c_445_n 0.00351743f $X=2.605 $Y=0.235 $X2=0
+ $Y2=0
cc_152 N_A_79_21#_M1006_d N_VGND_c_445_n 0.00370147f $X=3.745 $Y=0.235 $X2=0
+ $Y2=0
cc_153 N_A_79_21#_c_58_n N_VGND_c_445_n 0.0104585f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_59_n N_VGND_c_445_n 0.0100565f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_71_p N_VGND_c_445_n 0.00536968f $X=1.525 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_141_p N_VGND_c_445_n 8.6794e-19 $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_73_p N_VGND_c_445_n 0.0459185f $X=2.79 $Y=0.34 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_83_p N_VGND_c_445_n 0.00619703f $X=1.695 $Y=0.34 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_102_p N_VGND_c_445_n 0.0139244f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_79_21#_c_158_p N_VGND_c_445_n 0.00644035f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_71_p A_319_47# 0.00199183f $X=1.525 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_79_21#_c_82_p A_319_47# 0.00263527f $X=1.61 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_79_21#_c_73_p A_319_47# 0.00824289f $X=2.79 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_164 N_A_79_21#_c_83_p A_319_47# 4.1826e-19 $X=1.695 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_165 N_A_79_21#_c_73_p A_417_47# 0.0107491f $X=2.79 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A3_M1011_g N_A2_M1005_g 0.0209777f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_167 A3 A2 0.0233553f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A3_c_174_n A2 0.00187555f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A3_c_175_n A2 0.00235477f $X=1.58 $Y=0.995 $X2=0 $Y2=0
cc_170 A3 N_A2_c_214_n 3.82878e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A3_c_174_n N_A2_c_214_n 0.0191719f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A3_c_175_n N_A2_c_215_n 0.0307705f $X=1.58 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A3_M1011_g N_VPWR_c_342_n 0.00974622f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A3_M1011_g N_VPWR_c_346_n 0.00579312f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A3_M1011_g N_VPWR_c_339_n 0.0111786f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A3_M1011_g N_X_c_397_n 0.00104911f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A3_c_175_n N_X_c_397_n 0.0011072f $X=1.58 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A3_M1011_g N_A_319_297#_c_414_n 0.00170398f $X=1.52 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A3_M1011_g N_A_319_297#_c_418_n 0.00458013f $X=1.52 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A3_c_175_n N_VGND_c_440_n 0.00529004f $X=1.58 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A3_c_175_n N_VGND_c_443_n 0.0039519f $X=1.58 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A3_c_175_n N_VGND_c_445_n 0.00629046f $X=1.58 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_M1005_g N_A1_M1013_g 0.0374809f $X=2.01 $Y=1.985 $X2=0 $Y2=0
cc_184 A2 A1 0.0312731f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_185 N_A2_c_214_n A1 0.00206857f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_c_215_n A1 5.23002e-19 $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_187 A2 N_A1_c_250_n 3.90049e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A2_c_214_n N_A1_c_250_n 0.0164411f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_189 A2 N_A1_c_251_n 0.00148821f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A2_c_215_n N_A1_c_251_n 0.0300119f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_M1005_g N_VPWR_c_343_n 0.00434844f $X=2.01 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A2_M1005_g N_VPWR_c_346_n 0.00436487f $X=2.01 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A2_M1005_g N_VPWR_c_339_n 0.00633402f $X=2.01 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A2_M1005_g N_A_319_297#_c_415_n 0.0105704f $X=2.01 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A2_c_215_n N_VGND_c_443_n 0.00357877f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_215_n N_VGND_c_445_n 0.00572424f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_197 A2 A_417_47# 0.00326828f $X=1.99 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_198 N_A1_M1013_g N_B1_M1003_g 0.0254459f $X=2.53 $Y=1.985 $X2=0 $Y2=0
cc_199 A1 N_B1_c_285_n 3.23806e-19 $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_200 N_A1_c_250_n N_B1_c_285_n 0.0133736f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_201 A1 N_B1_c_286_n 0.0210328f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A1_c_250_n N_B1_c_286_n 0.0023628f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_203 A1 N_B1_c_287_n 0.00202093f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_204 N_A1_c_251_n N_B1_c_287_n 0.0181509f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A1_M1013_g N_VPWR_c_343_n 0.00329367f $X=2.53 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A1_M1013_g N_VPWR_c_348_n 0.00435702f $X=2.53 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A1_M1013_g N_VPWR_c_339_n 0.00639196f $X=2.53 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A1_M1013_g N_A_319_297#_c_415_n 0.0132799f $X=2.53 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A1_M1013_g N_A_319_297#_c_421_n 0.00862402f $X=2.53 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A1_c_251_n N_VGND_c_443_n 0.00357877f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A1_c_251_n N_VGND_c_445_n 0.00587291f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_M1003_g N_C1_M1000_g 0.0365368f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_c_285_n C1 0.00110765f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B1_c_286_n C1 0.0109995f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_215 N_B1_c_285_n N_C1_c_317_n 0.0127802f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B1_c_286_n N_C1_c_317_n 0.00125938f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B1_c_287_n N_C1_c_318_n 0.0229775f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_M1003_g N_VPWR_c_348_n 0.00585385f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B1_M1003_g N_VPWR_c_339_n 0.0114532f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B1_c_287_n N_VGND_c_441_n 0.00458634f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_287_n N_VGND_c_443_n 0.00428022f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_287_n N_VGND_c_445_n 0.00654566f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_223 N_C1_M1000_g N_VPWR_c_348_n 0.00585385f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_224 N_C1_M1000_g N_VPWR_c_339_n 0.0120554f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_225 N_C1_c_318_n N_VGND_c_441_n 0.00467817f $X=3.755 $Y=0.995 $X2=0 $Y2=0
cc_226 N_C1_c_318_n N_VGND_c_444_n 0.00428022f $X=3.755 $Y=0.995 $X2=0 $Y2=0
cc_227 N_C1_c_318_n N_VGND_c_445_n 0.00708574f $X=3.755 $Y=0.995 $X2=0 $Y2=0
cc_228 N_VPWR_c_339_n N_X_M1004_s 0.00217524f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_342_n N_X_c_397_n 0.0276609f $X=1.245 $Y=2 $X2=0 $Y2=0
cc_230 N_VPWR_c_344_n N_X_c_397_n 0.0150775f $X=1.16 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_339_n N_X_c_397_n 0.0119688f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_339_n N_A_319_297#_M1011_d 0.00315939f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_233 N_VPWR_c_339_n N_A_319_297#_M1013_d 0.00389706f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_342_n N_A_319_297#_c_414_n 0.0115483f $X=1.245 $Y=2 $X2=0 $Y2=0
cc_235 N_VPWR_c_342_n N_A_319_297#_c_418_n 0.0287862f $X=1.245 $Y=2 $X2=0 $Y2=0
cc_236 N_VPWR_c_346_n N_A_319_297#_c_418_n 0.0153379f $X=2.125 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_339_n N_A_319_297#_c_418_n 0.00944122f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_M1005_d N_A_319_297#_c_415_n 0.00587854f $X=2.085 $Y=1.485 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_343_n N_A_319_297#_c_415_n 0.0141687f $X=2.29 $Y=2.34 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_346_n N_A_319_297#_c_415_n 0.00336467f $X=2.125 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_348_n N_A_319_297#_c_415_n 0.00327382f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_339_n N_A_319_297#_c_415_n 0.0144643f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_343_n N_A_319_297#_c_421_n 0.0125922f $X=2.29 $Y=2.34 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_348_n N_A_319_297#_c_421_n 0.0196089f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_339_n N_A_319_297#_c_421_n 0.0118379f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_339_n A_635_297# 0.0179632f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_247 N_VPWR_c_341_n N_VGND_c_439_n 0.0086775f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_248 N_X_c_397_n N_VGND_c_442_n 0.0150775f $X=0.68 $Y=0.38 $X2=1.1 $Y2=0.825
cc_249 N_X_M1007_s N_VGND_c_445_n 0.00217524f $X=0.545 $Y=0.235 $X2=2.875
+ $Y2=0.57
cc_250 N_X_c_397_n N_VGND_c_445_n 0.0119688f $X=0.68 $Y=0.38 $X2=2.875 $Y2=0.57
cc_251 N_VGND_c_445_n A_319_47# 0.00273039f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_252 N_VGND_c_445_n A_417_47# 0.00297142f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

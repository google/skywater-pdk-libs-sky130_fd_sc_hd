* File: sky130_fd_sc_hd__a32o_2.pex.spice
* Created: Thu Aug 27 14:05:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A32O_2%A_21_199# 1 2 7 9 12 14 16 19 23 26 27 29 30
+ 33 34 35 38 44 50
r96 44 45 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.03
+ $X2=2.04 $Y2=1.945
r97 36 38 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.42 $Y=0.615
+ $X2=2.42 $Y2=0.36
r98 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.255 $Y=0.7
+ $X2=2.42 $Y2=0.615
r99 34 35 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.255 $Y=0.7
+ $X2=1.89 $Y2=0.7
r100 33 45 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=2 $Y=1.63 $X2=2
+ $Y2=1.945
r101 30 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2 $Y=1.53
+ $X2=1.795 $Y2=1.53
r102 30 33 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2 $Y=1.615 $X2=2
+ $Y2=1.63
r103 29 40 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=1.445
+ $X2=1.795 $Y2=1.53
r104 28 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.795 $Y=0.785
+ $X2=1.89 $Y2=0.7
r105 28 29 38.5263 $w=1.88e-07 $l=6.6e-07 $layer=LI1_cond $X=1.795 $Y=0.785
+ $X2=1.795 $Y2=1.445
r106 26 40 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.7 $Y=1.53
+ $X2=1.795 $Y2=1.53
r107 26 27 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=1.7 $Y=1.53
+ $X2=0.705 $Y2=1.53
r108 24 50 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.62 $Y=1.16
+ $X2=0.89 $Y2=1.16
r109 24 47 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.62 $Y=1.16
+ $X2=0.47 $Y2=1.16
r110 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r111 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=1.445
+ $X2=0.705 $Y2=1.53
r112 21 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.62 $Y=1.445
+ $X2=0.62 $Y2=1.16
r113 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r114 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r115 14 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r116 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r117 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r118 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r119 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r120 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r121 2 44 600 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2.03
r122 2 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.63
r123 1 38 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.235 $X2=2.42 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%B2 3 6 9 10 12 13
r40 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.365
+ $Y=1.16 $X2=1.365 $Y2=1.16
r41 13 18 0.833091 $w=4.13e-07 $l=3e-08 $layer=LI1_cond $X=1.322 $Y=1.19
+ $X2=1.322 $Y2=1.16
r42 12 18 8.60861 $w=4.13e-07 $l=3.1e-07 $layer=LI1_cond $X=1.322 $Y=0.85
+ $X2=1.322 $Y2=1.16
r43 9 17 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.365 $Y2=1.16
r44 9 11 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.757 $Y=1.16
+ $X2=1.757 $Y2=1.325
r45 9 10 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.757 $Y=1.16
+ $X2=1.757 $Y2=0.995
r46 6 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.985
+ $X2=1.83 $Y2=1.325
r47 3 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.685 $Y=0.56
+ $X2=1.685 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%B1 3 6 10 12 15 19
c45 19 0 1.98392e-19 $X=2.25 $Y=0.995
c46 10 0 2.94838e-20 $X=2.25 $Y=1.16
r47 13 15 8.37803 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.43 $Y=1.245 $X2=2.43
+ $Y2=1.445
r48 12 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=1.16
+ $X2=2.43 $Y2=1.245
r49 10 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.25 $Y2=0.995
r50 9 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=1.16 $X2=2.43
+ $Y2=1.16
r51 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r52 4 10 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.325
+ $X2=2.25 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.325 $X2=2.25
+ $Y2=1.985
r54 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.19 $Y=0.56 $X2=2.19
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%A1 3 6 11 12 13 15 18
c40 18 0 1.97052e-19 $X=2.75 $Y=0.995
c41 11 0 1.98392e-19 $X=2.77 $Y=1.16
r42 12 19 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.75 $Y2=1.325
r43 12 18 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.75 $Y2=0.995
r44 11 13 8.5315 $w=2.98e-07 $l=2.05e-07 $layer=LI1_cond $X=2.835 $Y=1.16
+ $X2=2.835 $Y2=0.955
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.16 $X2=2.77 $Y2=1.16
r46 8 15 6.82517 $w=1.93e-07 $l=1.2e-07 $layer=LI1_cond $X=2.87 $Y=0.512
+ $X2=2.99 $Y2=0.512
r47 8 13 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.87 $Y=0.61
+ $X2=2.87 $Y2=0.955
r48 6 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.985
+ $X2=2.67 $Y2=1.325
r49 3 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.56 $X2=2.67
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%A2 1 3 6 8 9 10 11 17
c44 17 0 2.91989e-20 $X=3.25 $Y=1.16
c45 8 0 1.97052e-19 $X=3.45 $Y=0.51
r46 25 31 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=1.325
+ $X2=3.425 $Y2=1.16
r47 19 31 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=1.16
r48 18 31 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=3.25 $Y=1.16
+ $X2=3.425 $Y2=1.16
r49 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.16 $X2=3.25 $Y2=1.16
r50 11 25 9.84378 $w=2.38e-07 $l=2.05e-07 $layer=LI1_cond $X=3.425 $Y=1.53
+ $X2=3.425 $Y2=1.325
r51 10 31 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=3.425 $Y2=1.16
r52 9 19 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=3.425 $Y=0.85
+ $X2=3.425 $Y2=0.995
r53 8 9 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=3.425 $Y=0.51
+ $X2=3.425 $Y2=0.85
r54 4 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.25 $Y=1.325 $X2=3.25
+ $Y2=1.985
r56 1 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.25 $Y=0.995 $X2=3.25
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%A3 1 3 6 8 9 15
r26 12 15 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.67 $Y=1.16 $X2=3.9
+ $Y2=1.16
r27 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.935 $Y=1.16
+ $X2=3.935 $Y2=1.53
r28 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9 $Y=1.16
+ $X2=3.9 $Y2=1.16
r29 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.325 $X2=3.67
+ $Y2=1.985
r31 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.995 $X2=3.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%X 1 2 3 12 14 19 20 21 22 23 24 33 36
r41 33 36 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=0.825
+ $X2=0.24 $Y2=0.85
r42 23 24 10.0225 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=1.955
+ $X2=0.24 $Y2=2.21
r43 22 23 10.0225 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=1.53
+ $X2=0.24 $Y2=1.785
r44 21 22 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=0.24 $Y=1.19
+ $X2=0.24 $Y2=1.53
r45 20 33 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.74 $X2=0.24
+ $Y2=0.825
r46 20 21 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.24 $Y=0.88
+ $X2=0.24 $Y2=1.19
r47 20 36 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.88 $X2=0.24
+ $Y2=0.85
r48 15 23 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.24 $Y2=1.87
r49 14 19 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=1.87 $X2=1.1
+ $Y2=1.87
r50 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=1.87
+ $X2=0.345 $Y2=1.87
r51 10 20 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.24 $Y2=0.74
r52 10 12 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.68 $Y2=0.74
r53 3 19 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.95
r54 2 23 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
r55 1 12 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%VPWR 1 2 3 12 16 18 20 23 24 25 27 39 44 48
r61 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 39 47 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.927 $Y2=2.72
r66 39 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r74 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r76 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r79 23 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=2.72
+ $X2=2.88 $Y2=2.72
r81 22 41 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.45 $Y2=2.72
r82 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.88 $Y2=2.72
r83 18 47 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.882 $Y=2.635
+ $X2=3.927 $Y2=2.72
r84 18 20 21.8448 $w=3.33e-07 $l=6.35e-07 $layer=LI1_cond $X=3.882 $Y=2.635
+ $X2=3.882 $Y2=2
r85 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2.72
r86 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2.225
r87 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r88 10 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.21
r89 3 20 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=2
r90 2 16 600 $w=1.7e-07 $l=8.04674e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2.225
r91 1 12 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%A_299_297# 1 2 3 12 14 15 16 18 25
c33 25 0 2.91989e-20 $X=3.46 $Y=1.96
c34 16 0 2.94838e-20 $X=2.46 $Y=1.965
r35 19 23 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.88
+ $X2=2.46 $Y2=1.88
r36 18 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=1.88
+ $X2=3.46 $Y2=1.88
r37 18 19 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.375 $Y=1.88
+ $X2=2.545 $Y2=1.88
r38 16 23 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.965
+ $X2=2.46 $Y2=1.88
r39 16 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.46 $Y=1.965
+ $X2=2.46 $Y2=2.295
r40 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=2.46 $Y2=2.295
r41 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=1.705 $Y2=2.38
r42 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=2.295
+ $X2=1.705 $Y2=2.38
r43 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.62 $Y=2.295
+ $X2=1.62 $Y2=1.95
r44 3 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=1.96
r45 2 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.96
r46 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_2%VGND 1 2 3 10 12 14 16 18 25 36 42 45
r61 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r62 40 42 6.65775 $w=5.28e-07 $l=3e-08 $layer=LI1_cond $X=1.61 $Y=0.18 $X2=1.64
+ $Y2=0.18
r63 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r64 38 40 3.04661 $w=5.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.475 $Y=0.18
+ $X2=1.61 $Y2=0.18
r65 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r66 34 38 7.33444 $w=5.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.475 $Y2=0.18
r67 34 36 10.8327 $w=5.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=0.935 $Y2=0.18
r68 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 29 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r70 29 41 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=1.61
+ $Y2=0
r71 28 42 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=1.64
+ $Y2=0
r72 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r73 25 44 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.927
+ $Y2=0
r74 25 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.45
+ $Y2=0
r75 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r76 23 36 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=0.935
+ $Y2=0
r77 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r78 21 31 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r79 21 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r80 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r81 18 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r82 14 44 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.882 $Y=0.085
+ $X2=3.927 $Y2=0
r83 14 16 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=3.882 $Y=0.085
+ $X2=3.882 $Y2=0.38
r84 10 31 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r85 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r86 3 16 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.38
r87 2 38 91 $w=1.7e-07 $l=5.69078e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.475 $Y2=0.36
r88 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__dlygate4sd1_1.pex.spice
* Created: Thu Aug 27 14:18:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A 3 7 9 10 14
c33 14 0 5.56024e-20 $X=0.31 $Y=1.16
r34 14 17 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.36 $Y=1.16
+ $X2=0.36 $Y2=1.325
r35 14 16 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.36 $Y=1.16
+ $X2=0.36 $Y2=0.995
r36 9 10 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.16 $X2=0.32
+ $Y2=1.53
r37 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.16 $X2=0.31 $Y2=1.16
r38 7 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r39 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_27_47# 1 2 9 13 17 21 23 24 25 26 27
+ 28 32
c71 32 0 2.77055e-20 $X=0.89 $Y=1.16
c72 27 0 1.90252e-19 $X=0.81 $Y=1.325
c73 25 0 5.56024e-20 $X=0.725 $Y=1.895
r74 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r75 29 31 20.4279 $w=2.15e-07 $l=3.6e-07 $layer=LI1_cond $X=0.852 $Y=0.8
+ $X2=0.852 $Y2=1.16
r76 27 31 9.93147 $w=2.15e-07 $l=1.84811e-07 $layer=LI1_cond $X=0.81 $Y=1.325
+ $X2=0.852 $Y2=1.16
r77 27 28 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.81 $Y=1.325
+ $X2=0.81 $Y2=1.785
r78 25 28 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.725 $Y=1.895
+ $X2=0.81 $Y2=1.785
r79 25 26 18.0724 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=0.725 $Y=1.895
+ $X2=0.38 $Y2=1.895
r80 23 29 2.11506 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.725 $Y=0.8
+ $X2=0.852 $Y2=0.8
r81 23 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.725 $Y=0.8
+ $X2=0.38 $Y2=0.8
r82 19 24 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.237 $Y=0.715
+ $X2=0.38 $Y2=0.8
r83 19 21 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=0.237 $Y=0.715
+ $X2=0.237 $Y2=0.51
r84 15 26 7.00622 $w=2.2e-07 $l=1.95407e-07 $layer=LI1_cond $X=0.232 $Y=2.005
+ $X2=0.38 $Y2=1.895
r85 15 17 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.232 $Y=2.005
+ $X2=0.232 $Y2=2.21
r86 11 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r87 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=2.275
r88 7 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r89 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.445
r90 2 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.21
r91 1 21 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_193_47# 1 2 7 9 10 12 14 16 19 25 30
+ 32 36
c64 36 0 1.90252e-19 $X=1.84 $Y=1.16
r65 35 36 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.83 $Y=1.16 $X2=1.84
+ $Y2=1.16
r66 28 30 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.1 $Y=2.32
+ $X2=1.235 $Y2=2.32
r67 23 25 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.1 $Y=0.4
+ $X2=1.235 $Y2=0.4
r68 20 35 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.63 $Y=1.16 $X2=1.83
+ $Y2=1.16
r69 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.16 $X2=1.63 $Y2=1.16
r70 17 32 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=1.175
+ $X2=1.235 $Y2=1.175
r71 17 19 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=1.32 $Y=1.175
+ $X2=1.63 $Y2=1.175
r72 16 30 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.235 $Y=2.175
+ $X2=1.235 $Y2=2.32
r73 15 32 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.235 $Y=1.275
+ $X2=1.235 $Y2=1.175
r74 15 16 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.235 $Y=1.275
+ $X2=1.235 $Y2=2.175
r75 14 32 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.235 $Y=1.075
+ $X2=1.235 $Y2=1.175
r76 13 25 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.235 $Y=0.545
+ $X2=1.235 $Y2=0.4
r77 13 14 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.235 $Y=0.545
+ $X2=1.235 $Y2=1.075
r78 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.16
r79 10 12 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.915
r80 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r81 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.83 $Y=0.995 $X2=1.83
+ $Y2=0.675
r82 2 28 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=2.065 $X2=1.1 $Y2=2.34
r83 1 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%A_299_93# 1 2 9 12 16 19 21 22 23 24
+ 26 30 32
r67 30 33 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.16 $X2=2.29
+ $Y2=1.325
r68 30 32 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.16 $X2=2.29
+ $Y2=0.995
r69 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=1.16 $X2=2.275 $Y2=1.16
r70 27 29 17.5021 $w=2.37e-07 $l=3.4e-07 $layer=LI1_cond $X=2.215 $Y=0.82
+ $X2=2.215 $Y2=1.16
r71 23 29 9.48765 $w=2.37e-07 $l=1.92678e-07 $layer=LI1_cond $X=2.155 $Y=1.325
+ $X2=2.215 $Y2=1.16
r72 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.155 $Y=1.325
+ $X2=2.155 $Y2=1.575
r73 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.07 $Y=1.66
+ $X2=2.155 $Y2=1.575
r74 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.07 $Y=1.66
+ $X2=1.74 $Y2=1.66
r75 20 26 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.74 $Y=0.82
+ $X2=1.627 $Y2=0.82
r76 19 27 2.684 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.07 $Y=0.82 $X2=2.215
+ $Y2=0.82
r77 19 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.07 $Y=0.82
+ $X2=1.74 $Y2=0.82
r78 16 22 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.627 $Y=1.745
+ $X2=1.74 $Y2=1.66
r79 16 18 5.69333 $w=2.25e-07 $l=1.05e-07 $layer=LI1_cond $X=1.627 $Y=1.745
+ $X2=1.627 $Y2=1.85
r80 12 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=1.985
+ $X2=2.315 $Y2=1.325
r81 9 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.315 $Y=0.56
+ $X2=2.315 $Y2=0.995
r82 2 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.705 $X2=1.63 $Y2=1.85
r83 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.465 $X2=1.62 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%VPWR 1 2 9 13 15 17 22 29 30 33 36 41
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 34 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r45 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 30 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 27 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.27 $Y=2.72 $X2=2.09
+ $Y2=2.72
r49 27 29 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 23 33 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.657 $Y2=2.72
r54 23 25 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 22 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=2.09
+ $Y2=2.72
r56 22 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=1.61
+ $Y2=2.72
r57 19 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 17 33 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.55 $Y=2.72
+ $X2=0.657 $Y2=2.72
r59 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=0.23
+ $Y2=2.72
r60 15 41 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 11 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=2.635
+ $X2=2.09 $Y2=2.72
r62 11 13 20.3278 $w=3.58e-07 $l=6.35e-07 $layer=LI1_cond $X=2.09 $Y=2.635
+ $X2=2.09 $Y2=2
r63 7 33 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.657 $Y=2.635
+ $X2=0.657 $Y2=2.72
r64 7 9 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.657 $Y=2.635
+ $X2=0.657 $Y2=2.34
r65 2 13 600 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.705 $X2=2.105 $Y2=2
r66 1 9 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%X 1 2 10 11 12 13 14 15
r17 14 15 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.57 $Y=1.87
+ $X2=2.57 $Y2=2.21
r18 11 14 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=2.57 $Y=1.625
+ $X2=2.57 $Y2=1.87
r19 11 12 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.57 $Y=1.625
+ $X2=2.57 $Y2=1.495
r20 10 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.615 $Y=0.825
+ $X2=2.615 $Y2=1.495
r21 9 13 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=0.68
+ $X2=2.555 $Y2=0.51
r22 9 10 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.555 $Y=0.68
+ $X2=2.555 $Y2=0.825
r23 2 14 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=2.39
+ $Y=1.485 $X2=2.525 $Y2=1.87
r24 1 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.235 $X2=2.525 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD1_1%VGND 1 2 9 13 15 17 22 29 30 33 36 41
c46 9 0 2.77055e-20 $X=0.68 $Y=0.38
r47 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r48 34 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r49 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r50 30 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r51 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.075
+ $Y2=0
r53 27 29 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.99
+ $Y2=0
r54 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r55 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r56 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r57 23 33 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.657
+ $Y2=0
r58 23 25 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.61
+ $Y2=0
r59 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=2.075
+ $Y2=0
r60 22 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=1.61
+ $Y2=0
r61 19 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 17 33 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.657
+ $Y2=0
r63 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.23
+ $Y2=0
r64 15 41 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r65 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0
r66 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0.38
r67 7 33 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.657 $Y=0.085
+ $X2=0.657 $Y2=0
r68 7 9 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.657 $Y=0.085
+ $X2=0.657 $Y2=0.38
r69 2 13 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.465 $X2=2.105 $Y2=0.38
r70 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


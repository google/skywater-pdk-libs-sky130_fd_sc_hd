* File: sky130_fd_sc_hd__o22a_1.pex.spice
* Created: Tue Sep  1 19:23:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O22A_1%A_78_199# 1 2 7 9 12 17 18 20 21 22 23 25 28
+ 29
c72 28 0 8.9786e-20 $X=1.62 $Y=0.73
c73 20 0 9.14711e-20 $X=0.81 $Y=0.805
c74 17 0 1.46941e-19 $X=0.69 $Y=1.16
r75 33 35 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.49
+ $Y2=1.16
r76 28 29 10.1417 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=1.62 $Y=0.77 $X2=1.42
+ $Y2=0.77
r77 23 32 3.02357 $w=3.85e-07 $l=1.61369e-07 $layer=LI1_cond $X=1.927 $Y=1.805
+ $X2=1.94 $Y2=1.65
r78 23 25 4.63971 $w=3.83e-07 $l=1.55e-07 $layer=LI1_cond $X=1.927 $Y=1.805
+ $X2=1.927 $Y2=1.96
r79 21 32 4.58935 $w=2.1e-07 $l=2.28637e-07 $layer=LI1_cond $X=1.735 $Y=1.6
+ $X2=1.94 $Y2=1.65
r80 21 22 48.8528 $w=2.08e-07 $l=9.25e-07 $layer=LI1_cond $X=1.735 $Y=1.6
+ $X2=0.81 $Y2=1.6
r81 20 29 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=0.81 $Y=0.805
+ $X2=1.42 $Y2=0.805
r82 18 35 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.69 $Y=1.16 $X2=0.49
+ $Y2=1.16
r83 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.16 $X2=0.69 $Y2=1.16
r84 15 22 6.97695 $w=2.1e-07 $l=1.83123e-07 $layer=LI1_cond $X=0.672 $Y=1.495
+ $X2=0.81 $Y2=1.6
r85 15 17 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=0.672 $Y=1.495
+ $X2=0.672 $Y2=1.16
r86 14 20 7.21025 $w=1.8e-07 $l=1.77381e-07 $layer=LI1_cond $X=0.672 $Y=0.895
+ $X2=0.81 $Y2=0.805
r87 14 17 11.1054 $w=2.73e-07 $l=2.65e-07 $layer=LI1_cond $X=0.672 $Y=0.895
+ $X2=0.672 $Y2=1.16
r88 10 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r89 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r90 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r91 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r92 2 32 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.485 $X2=1.98 $Y2=1.62
r93 2 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=1.485 $X2=1.98 $Y2=1.96
r94 1 28 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%B1 3 5 7 8 13
c33 13 0 1.33197e-20 $X=1.385 $Y=1.16
c34 8 0 1.86282e-19 $X=1.15 $Y=1.19
r35 13 14 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.41 $Y2=1.16
r36 11 13 31.4985 $w=3.29e-07 $l=2.15e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.385 $Y2=1.16
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r38 5 14 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r39 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
r40 1 13 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.16
r41 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%B2 3 5 7 8 11 12 15
c36 11 0 1.86282e-19 $X=1.83 $Y=1.16
r37 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=1.83 $Y2=1.325
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.16 $X2=1.83 $Y2=1.16
r39 8 12 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=1.635 $Y=1.2
+ $X2=1.83 $Y2=1.2
r40 8 15 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=1.2 $X2=1.61
+ $Y2=1.2
r41 5 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r42 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.995 $X2=1.83
+ $Y2=0.56
r43 3 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.77 $Y=1.985
+ $X2=1.77 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%A2 3 6 8 11 12 15
c43 15 0 8.9786e-20 $X=2.32 $Y=0.995
c44 8 0 1.33197e-20 $X=2.545 $Y=1.615
r45 11 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.32 $Y2=1.325
r46 11 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.32 $Y2=0.995
r47 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.16 $X2=2.33 $Y2=1.16
r48 8 12 15.555 $w=2e-07 $l=2.55e-07 $layer=LI1_cond $X=2.545 $Y=1.615 $X2=2.545
+ $Y2=1.87
r49 8 10 20.0427 $w=2.96e-07 $l=5.20312e-07 $layer=LI1_cond $X=2.545 $Y=1.615
+ $X2=2.405 $Y2=1.16
r50 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.39 $Y=1.985
+ $X2=2.39 $Y2=1.325
r51 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.33 $Y=0.56 $X2=2.33
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%A1 3 6 8 11 13
r25 11 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.16
+ $X2=2.845 $Y2=1.325
r26 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.16
+ $X2=2.845 $Y2=0.995
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.835
+ $Y=1.16 $X2=2.835 $Y2=1.16
r28 8 12 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=2.99 $Y=1.175
+ $X2=2.835 $Y2=1.175
r29 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.985
+ $X2=2.75 $Y2=1.325
r30 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.56 $X2=2.75
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%X 1 2 7 10
r13 10 13 42.1876 $w=2.78e-07 $l=1.025e-06 $layer=LI1_cond $X=0.225 $Y=0.595
+ $X2=0.225 $Y2=1.62
r14 7 17 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=0.225 $Y=2.21 $X2=0.225
+ $Y2=2.3
r15 7 13 24.2836 $w=2.78e-07 $l=5.9e-07 $layer=LI1_cond $X=0.225 $Y=2.21
+ $X2=0.225 $Y2=1.62
r16 2 17 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r17 2 13 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r18 1 10 182 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%VPWR 1 2 7 9 13 15 20 29 37
c41 1 0 1.46941e-19 $X=0.565 $Y=1.485
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 24 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 24 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 23 26 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 21 23 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.34 $Y=2.72 $X2=1.61
+ $Y2=2.72
r50 20 36 4.71668 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=3.017 $Y2=2.72
r51 20 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.53 $Y2=2.72
r52 15 21 10.0822 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=0.947 $Y=2.72
+ $X2=1.34 $Y2=2.72
r53 15 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 15 29 11.5799 $w=7.83e-07 $l=7.6e-07 $layer=LI1_cond $X=0.947 $Y=2.72
+ $X2=0.947 $Y2=1.96
r55 15 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.555 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 13 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 13 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 9 12 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.975 $Y=1.66
+ $X2=2.975 $Y2=2.34
r59 7 36 2.96544 $w=3.2e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=3.017 $Y2=2.72
r60 7 12 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.34
r61 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=2.34
r62 2 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.66
r63 1 29 150 $w=1.7e-07 $l=8.13542e-07 $layer=licon1_PDIFF $count=4 $X=0.565
+ $Y=1.485 $X2=1.175 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%VGND 1 2 9 11 15 17 19 26 27 30 33
r49 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 31 34 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r51 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 27 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r53 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r54 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.54
+ $Y2=0
r55 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.99
+ $Y2=0
r56 19 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r57 19 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r58 17 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0
r61 13 15 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.36
r62 12 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r63 11 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.54
+ $Y2=0
r64 11 12 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=2.455 $Y=0
+ $X2=0.765 $Y2=0
r65 7 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r66 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0.38
r67 2 15 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.405
+ $Y=0.235 $X2=2.54 $Y2=0.36
r68 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_1%A_215_47# 1 2 3 10 14 15 16 20
r41 18 20 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.965 $Y=0.695
+ $X2=2.965 $Y2=0.39
r42 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0.78
+ $X2=2.12 $Y2=0.78
r43 16 18 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.795 $Y=0.78
+ $X2=2.965 $Y2=0.695
r44 16 17 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.795 $Y=0.78
+ $X2=2.285 $Y2=0.78
r45 15 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.695 $X2=2.12
+ $Y2=0.78
r46 14 23 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.12 $Y=0.475 $X2=2.12
+ $Y2=0.385
r47 14 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.12 $Y=0.475
+ $X2=2.12 $Y2=0.695
r48 10 23 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.385
+ $X2=2.12 $Y2=0.385
r49 10 12 46.5202 $w=1.78e-07 $l=7.55e-07 $layer=LI1_cond $X=1.955 $Y=0.385
+ $X2=1.2 $Y2=0.385
r50 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.39
r51 2 25 182 $w=1.7e-07 $l=5.92832e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.12 $Y2=0.73
r52 2 23 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.12 $Y2=0.39
r53 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.39
.ends


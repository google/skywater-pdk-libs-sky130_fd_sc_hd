* File: sky130_fd_sc_hd__dlrbp_1.spice
* Created: Thu Aug 27 14:16:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlrbp_1.pex.spice"
.subckt sky130_fd_sc_hd__dlrbp_1  VNB VPB GATE D RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_GATE_M1021_g N_A_27_47#_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_193_47#_M1010_d N_A_27_47#_M1010_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g N_A_299_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_465_47# N_A_299_47#_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.0567 PD=0.802308 PS=0.69 NRD=32.628 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1018 N_A_560_47#_M1018_d N_A_193_47#_M1018_g A_465_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0612 AS=0.0609231 PD=0.7 PS=0.687692 NRD=0 NRS=38.076 M=1 R=2.4
+ SA=75001.1 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1011 A_658_47# N_A_27_47#_M1011_g N_A_560_47#_M1018_d VNB NSHORT L=0.15 W=0.36
+ AD=0.0609231 AS=0.0612 PD=0.687692 PS=0.7 NRD=38.076 NRS=21.66 M=1 R=2.4
+ SA=75001.6 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1023 N_VGND_M1023_d N_A_711_307#_M1023_g A_658_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_941_47# N_A_560_47#_M1015_g N_A_711_307#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.095875 AS=0.169 PD=0.945 PS=1.82 NRD=17.076 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_RESET_B_M1020_g A_941_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.23075 AS=0.095875 PD=1.36 PS=0.945 NRD=0 NRS=17.076 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1008 N_Q_M1008_d N_A_711_307#_M1008_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.23075 PD=1.82 PS=1.36 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_711_307#_M1002_g N_A_1308_47#_M1002_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_Q_N_M1019_d N_A_1308_47#_M1019_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_GATE_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_VPWR_M1017_d N_D_M1017_g N_A_299_47#_M1017_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1012 A_465_369# N_A_299_47#_M1012_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116891 AS=0.0864 PD=1.17132 PS=0.91 NRD=39.2818 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_560_47#_M1001_d N_A_27_47#_M1001_g A_465_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0767094 PD=0.69 PS=0.768679 NRD=0 NRS=59.8683 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1022 A_645_413# N_A_193_47#_M1022_g N_A_560_47#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0693 AS=0.0567 PD=0.75 PS=0.69 NRD=51.5943 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_711_307#_M1009_g A_645_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0693 PD=1.36 PS=0.75 NRD=0 NRS=51.5943 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_711_307#_M1013_d N_A_560_47#_M1013_g N_VPWR_M1013_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.155 AS=0.26 PD=1.31 PS=2.52 NRD=6.8753 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_RESET_B_M1005_g N_A_711_307#_M1013_d VPB PHIGHVT L=0.15
+ W=1 AD=0.355 AS=0.155 PD=1.71 PS=1.31 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_Q_M1004_d N_A_711_307#_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.355 PD=2.52 PS=1.71 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_A_711_307#_M1016_g N_A_1308_47#_M1016_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1014 N_Q_N_M1014_d N_A_1308_47#_M1014_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.161 P=19.61
c_149 VPB 0 1.54454e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__dlrbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__or4b_2.spice.pex
* Created: Thu Aug 27 14:44:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4B_2%D_N 3 7 9 15
c28 7 0 3.82892e-19 $X=0.47 $Y=1.695
r29 12 15 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r31 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r32 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r33 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r34 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%A_176_21# 1 2 3 10 12 15 17 19 22 24 26 30 32
+ 36 40 41 43
c110 41 0 2.9293e-19 $X=1.375 $Y=1.16
c111 40 0 2.66826e-20 $X=1.375 $Y=1.16
c112 22 0 1.38646e-19 $X=1.375 $Y=1.985
r113 41 49 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.375 $Y=1.16
+ $X2=0.955 $Y2=1.16
r114 40 42 19.1271 $w=2.36e-07 $l=3.7e-07 $layer=LI1_cond $X=1.477 $Y=1.16
+ $X2=1.477 $Y2=1.53
r115 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.375
+ $Y=1.16 $X2=1.375 $Y2=1.16
r116 34 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.97 $Y=0.735
+ $X2=2.97 $Y2=0.47
r117 33 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.82
+ $X2=2.07 $Y2=0.82
r118 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.885 $Y=0.82
+ $X2=2.97 $Y2=0.735
r119 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.885 $Y=0.82
+ $X2=2.155 $Y2=0.82
r120 28 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.735
+ $X2=2.07 $Y2=0.82
r121 28 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.07 $Y=0.735
+ $X2=2.07 $Y2=0.47
r122 27 42 2.65936 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.665 $Y=1.53
+ $X2=1.477 $Y2=1.53
r123 26 47 4.30016 $w=3.33e-07 $l=1.25e-07 $layer=LI1_cond $X=3.392 $Y=1.53
+ $X2=3.392 $Y2=1.655
r124 26 27 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=3.225 $Y=1.53
+ $X2=1.665 $Y2=1.53
r125 25 40 17.5763 $w=2.36e-07 $l=3.4e-07 $layer=LI1_cond $X=1.477 $Y=0.82
+ $X2=1.477 $Y2=1.16
r126 24 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.82
+ $X2=2.07 $Y2=0.82
r127 24 25 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.985 $Y=0.82
+ $X2=1.585 $Y2=0.82
r128 20 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.16
r129 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.985
r130 17 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=1.16
r131 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=0.56
r132 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.16
r133 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.985
r134 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.16
r135 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r136 3 47 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=1.485 $X2=3.39 $Y2=1.655
r137 2 36 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.265 $X2=2.97 $Y2=0.47
r138 1 30 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.265 $X2=2.07 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%A 3 7 9 12
c37 9 0 1.8796e-19 $X=2.07 $Y=1.19
r38 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.16
+ $X2=1.92 $Y2=1.325
r39 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.16
+ $X2=1.92 $Y2=0.995
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r41 9 13 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=1.92 $Y2=1.175
r42 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.86 $Y=1.695
+ $X2=1.86 $Y2=1.325
r43 3 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.86 $Y=0.475
+ $X2=1.86 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%B 3 6 7 10
c39 10 0 1.10744e-19 $X=2.28 $Y=2.3
r40 10 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.28 $Y=2.3
+ $X2=2.28 $Y2=2.165
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=2.3 $X2=2.28 $Y2=2.3
r42 7 11 9.93485 $w=2.88e-07 $l=2.5e-07 $layer=LI1_cond $X=2.53 $Y=2.27 $X2=2.28
+ $Y2=2.27
r43 6 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.34 $Y=1.695 $X2=2.34
+ $Y2=2.165
r44 3 6 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.34 $Y=0.475
+ $X2=2.34 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%C 3 7 9 10 14
c30 14 0 1.8796e-19 $X=2.76 $Y=1.16
r31 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.16
+ $X2=2.76 $Y2=1.325
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=1.16 $X2=2.76 $Y2=1.16
r33 9 10 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=1.175
+ $X2=3.45 $Y2=1.175
r34 9 15 12.7545 $w=1.98e-07 $l=2.3e-07 $layer=LI1_cond $X=2.99 $Y=1.175
+ $X2=2.76 $Y2=1.175
r35 5 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=0.995
+ $X2=2.76 $Y2=1.16
r36 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.76 $Y=0.995 $X2=2.76
+ $Y2=0.475
r37 3 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.7 $Y=1.695 $X2=2.7
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%A_27_53# 1 2 9 12 15 17 21 22 25 27 30 31 33
+ 37 40 46
c103 40 0 1.51706e-19 $X=1.577 $Y=1.87
c104 37 0 2.66826e-20 $X=0.637 $Y=1.605
c105 30 0 1.10744e-19 $X=2.945 $Y=2.215
c106 27 0 1.38646e-19 $X=2.86 $Y=1.87
c107 25 0 3.75993e-20 $X=1.44 $Y=2.08
r108 34 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=2.3
+ $X2=3.18 $Y2=2.3
r109 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.105
+ $Y=2.3 $X2=3.105 $Y2=2.3
r110 31 33 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.03 $Y=2.3
+ $X2=3.105 $Y2=2.3
r111 30 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=2.215
+ $X2=3.03 $Y2=2.3
r112 29 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.945 $Y=1.955
+ $X2=2.945 $Y2=2.215
r113 28 40 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.715 $Y=1.87
+ $X2=1.577 $Y2=1.87
r114 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.86 $Y=1.87
+ $X2=2.945 $Y2=1.955
r115 27 28 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.86 $Y=1.87
+ $X2=1.715 $Y2=1.87
r116 26 38 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.765 $Y=2.08
+ $X2=0.637 $Y2=2.08
r117 25 40 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=1.577 $Y=2.08
+ $X2=1.577 $Y2=1.87
r118 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.44 $Y=2.08
+ $X2=0.765 $Y2=2.08
r119 23 37 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.68 $Y=0.905
+ $X2=0.68 $Y2=1.605
r120 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.68 $Y2=0.905
r121 21 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.35 $Y2=0.82
r122 17 38 15.0496 $w=2.53e-07 $l=3.33e-07 $layer=LI1_cond $X=0.637 $Y=1.747
+ $X2=0.637 $Y2=2.08
r123 17 37 7.70102 $w=2.53e-07 $l=1.42e-07 $layer=LI1_cond $X=0.637 $Y=1.747
+ $X2=0.637 $Y2=1.605
r124 17 19 10.1091 $w=2.83e-07 $l=2.5e-07 $layer=LI1_cond $X=0.51 $Y=1.747
+ $X2=0.26 $Y2=1.747
r125 13 22 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.217 $Y=0.735
+ $X2=0.35 $Y2=0.82
r126 13 15 10.2198 $w=2.63e-07 $l=2.35e-07 $layer=LI1_cond $X=0.217 $Y=0.735
+ $X2=0.217 $Y2=0.5
r127 9 12 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=3.18 $Y=0.475
+ $X2=3.18 $Y2=1.695
r128 7 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=2.165
+ $X2=3.18 $Y2=2.3
r129 7 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.18 $Y=2.165 $X2=3.18
+ $Y2=1.695
r130 2 19 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.72
r131 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%VPWR 1 2 7 9 14 24 25 28 35
c50 28 0 1.58738e-19 $X=0.68 $Y=2.42
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 28 31 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.68 $Y=2.42 $X2=0.68
+ $Y2=2.72
r53 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 22 25 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 22 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 21 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 18 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 18 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 15 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r63 15 17 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 14 19 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.647 $Y=2.72
+ $X2=1.815 $Y2=2.72
r65 14 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 14 35 10.3204 $w=3.33e-07 $l=3e-07 $layer=LI1_cond $X=1.647 $Y=2.72
+ $X2=1.647 $Y2=2.42
r67 14 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.48 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 9 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r69 9 11 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 7 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 7 11 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r72 2 35 600 $w=1.7e-07 $l=1.03016e-06 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.65 $Y2=2.42
r73 1 28 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=0.535
+ $Y=2.185 $X2=0.68 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%X 1 2 8 9 13 15
c30 13 0 1.86554e-19 $X=1.165 $Y=1.66
r31 10 13 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.02 $Y=1.66
+ $X2=1.165 $Y2=1.66
r32 9 15 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=0.675
+ $X2=1.11 $Y2=0.51
r33 8 10 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=1.495
+ $X2=1.02 $Y2=1.66
r34 7 9 4.52581 $w=3.1e-07 $l=1.53542e-07 $layer=LI1_cond $X=1.02 $Y=0.79
+ $X2=1.11 $Y2=0.675
r35 7 8 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.02 $Y=0.79 $X2=1.02
+ $Y2=1.495
r36 2 13 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.66
r37 1 15 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.165 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_2%VGND 1 2 3 4 17 21 25 27 29 31 33 38 43 49 52
+ 55 59 61
c68 21 0 1.41224e-19 $X=1.6 $Y=0.4
r69 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r70 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r71 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r72 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r73 47 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r74 47 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r75 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r76 44 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.55
+ $Y2=0
r77 44 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.99
+ $Y2=0
r78 43 58 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.452
+ $Y2=0
r79 43 46 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=2.99
+ $Y2=0
r80 42 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r81 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r82 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r83 39 52 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.625
+ $Y2=0
r84 39 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.07
+ $Y2=0
r85 38 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.55
+ $Y2=0
r86 38 41 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.07
+ $Y2=0
r87 37 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r88 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r89 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r90 34 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.715
+ $Y2=0
r91 34 36 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=1.15
+ $Y2=0
r92 33 52 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.625
+ $Y2=0
r93 33 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.15
+ $Y2=0
r94 31 50 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r95 31 61 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r96 27 58 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.452 $Y2=0
r97 27 29 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0.5
r98 23 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=0.085
+ $X2=2.55 $Y2=0
r99 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.55 $Y=0.085
+ $X2=2.55 $Y2=0.4
r100 19 52 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=0.085
+ $X2=1.625 $Y2=0
r101 19 21 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.625 $Y=0.085
+ $X2=1.625 $Y2=0.4
r102 15 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r103 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.4
r104 4 29 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.265 $X2=3.39 $Y2=0.5
r105 3 25 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.265 $X2=2.55 $Y2=0.4
r106 2 21 182 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.6 $Y2=0.4
r107 1 17 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=0.715 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__a221oi_2.pxi.spice
* Created: Thu Aug 27 14:02:05 2020
* 
x_PM_SKY130_FD_SC_HD__A221OI_2%C1 N_C1_c_88_n N_C1_M1001_g N_C1_M1000_g
+ N_C1_c_89_n N_C1_M1018_g N_C1_M1004_g C1 C1 N_C1_c_91_n
+ PM_SKY130_FD_SC_HD__A221OI_2%C1
x_PM_SKY130_FD_SC_HD__A221OI_2%B2 N_B2_c_126_n N_B2_M1008_g N_B2_M1002_g
+ N_B2_c_127_n N_B2_M1019_g N_B2_M1011_g N_B2_c_134_n N_B2_c_128_n N_B2_c_129_n
+ B2 B2 N_B2_c_130_n N_B2_c_131_n PM_SKY130_FD_SC_HD__A221OI_2%B2
x_PM_SKY130_FD_SC_HD__A221OI_2%B1 N_B1_c_207_n N_B1_M1013_g N_B1_M1003_g
+ N_B1_c_208_n N_B1_M1014_g N_B1_M1007_g B1 N_B1_c_210_n
+ PM_SKY130_FD_SC_HD__A221OI_2%B1
x_PM_SKY130_FD_SC_HD__A221OI_2%A2 N_A2_c_250_n N_A2_M1015_g N_A2_M1005_g
+ N_A2_c_251_n N_A2_M1016_g N_A2_M1006_g N_A2_c_252_n N_A2_c_253_n N_A2_c_262_n
+ N_A2_c_263_n N_A2_c_254_n N_A2_c_255_n A2 N_A2_c_257_n A2
+ PM_SKY130_FD_SC_HD__A221OI_2%A2
x_PM_SKY130_FD_SC_HD__A221OI_2%A1 N_A1_c_335_n N_A1_M1009_g N_A1_M1010_g
+ N_A1_c_336_n N_A1_M1012_g N_A1_M1017_g A1 N_A1_c_337_n
+ PM_SKY130_FD_SC_HD__A221OI_2%A1
x_PM_SKY130_FD_SC_HD__A221OI_2%A_27_297# N_A_27_297#_M1000_d N_A_27_297#_M1004_d
+ N_A_27_297#_M1002_s N_A_27_297#_M1007_d N_A_27_297#_c_378_n
+ N_A_27_297#_c_379_n N_A_27_297#_c_380_n N_A_27_297#_c_381_n
+ N_A_27_297#_c_382_n N_A_27_297#_c_383_n N_A_27_297#_c_401_n
+ N_A_27_297#_c_384_n N_A_27_297#_c_402_n N_A_27_297#_c_404_n
+ PM_SKY130_FD_SC_HD__A221OI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__A221OI_2%Y N_Y_M1001_d N_Y_M1013_s N_Y_M1009_s N_Y_M1000_s
+ N_Y_c_433_n N_Y_c_434_n N_Y_c_435_n N_Y_c_436_n Y Y Y Y Y N_Y_c_446_n
+ PM_SKY130_FD_SC_HD__A221OI_2%Y
x_PM_SKY130_FD_SC_HD__A221OI_2%A_301_297# N_A_301_297#_M1002_d
+ N_A_301_297#_M1003_s N_A_301_297#_M1011_d N_A_301_297#_M1010_s
+ N_A_301_297#_M1006_s N_A_301_297#_c_509_n N_A_301_297#_c_510_n
+ N_A_301_297#_c_511_n N_A_301_297#_c_517_n N_A_301_297#_c_550_p
+ N_A_301_297#_c_520_n N_A_301_297#_c_505_n N_A_301_297#_c_551_p
+ N_A_301_297#_c_538_n N_A_301_297#_c_541_n N_A_301_297#_c_526_n
+ PM_SKY130_FD_SC_HD__A221OI_2%A_301_297#
x_PM_SKY130_FD_SC_HD__A221OI_2%VPWR N_VPWR_M1005_d N_VPWR_M1017_d N_VPWR_c_566_n
+ N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n
+ VPWR N_VPWR_c_572_n N_VPWR_c_565_n PM_SKY130_FD_SC_HD__A221OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A221OI_2%VGND N_VGND_M1001_s N_VGND_M1018_s N_VGND_M1019_s
+ N_VGND_M1016_s N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n VGND
+ N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n
+ PM_SKY130_FD_SC_HD__A221OI_2%VGND
x_PM_SKY130_FD_SC_HD__A221OI_2%A_383_47# N_A_383_47#_M1008_d N_A_383_47#_M1014_d
+ N_A_383_47#_c_706_n PM_SKY130_FD_SC_HD__A221OI_2%A_383_47#
x_PM_SKY130_FD_SC_HD__A221OI_2%A_735_47# N_A_735_47#_M1015_d N_A_735_47#_M1012_d
+ N_A_735_47#_c_722_n N_A_735_47#_c_723_n N_A_735_47#_c_721_n
+ PM_SKY130_FD_SC_HD__A221OI_2%A_735_47#
cc_1 VNB N_C1_c_88_n 0.0216908f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_C1_c_89_n 0.0211039f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_3 VNB C1 0.00916578f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_C1_c_91_n 0.0625251f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_5 VNB N_B2_c_126_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_6 VNB N_B2_c_127_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_7 VNB N_B2_c_128_n 0.00349181f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_8 VNB N_B2_c_129_n 0.0193014f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_9 VNB N_B2_c_130_n 0.0259184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B2_c_131_n 0.00702447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B1_c_207_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_12 VNB N_B1_c_208_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_13 VNB B1 0.00141292f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB N_B1_c_210_n 0.0299865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_250_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_16 VNB N_A2_c_251_n 0.0215628f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_17 VNB N_A2_c_252_n 0.00358835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_253_n 0.0192902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_254_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_20 VNB N_A2_c_255_n 0.0018962f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_21 VNB A2 0.0315903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_c_257_n 0.0279975f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.53
cc_23 VNB N_A1_c_335_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_24 VNB N_A1_c_336_n 0.0161471f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_25 VNB N_A1_c_337_n 0.0313079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_433_n 0.0192794f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_27 VNB N_Y_c_434_n 0.00219468f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_28 VNB N_Y_c_435_n 0.00219468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_436_n 0.0137838f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_30 VNB Y 8.46493e-19 $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_31 VNB N_VPWR_c_565_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_635_n 0.010359f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.985
cc_33 VNB N_VGND_c_636_n 0.0306077f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_34 VNB N_VGND_c_637_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_35 VNB N_VGND_c_638_n 0.00705803f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_36 VNB N_VGND_c_639_n 0.0365625f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_37 VNB N_VGND_c_640_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_641_n 0.0368904f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.53
cc_39 VNB N_VGND_c_642_n 0.00326621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_643_n 0.0137583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_644_n 0.28511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_645_n 0.0178184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_646_n 0.0202879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_735_47#_c_721_n 0.00247692f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.985
cc_45 VPB N_C1_M1000_g 0.0229738f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_46 VPB N_C1_M1004_g 0.0223988f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_47 VPB C1 0.0121511f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_48 VPB N_C1_c_91_n 0.0140903f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_49 VPB N_B2_M1002_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_50 VPB N_B2_M1011_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_51 VPB N_B2_c_134_n 0.00732858f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_52 VPB N_B2_c_128_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_53 VPB N_B2_c_129_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_54 VPB N_B2_c_130_n 0.00475082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_B2_c_131_n 0.00397829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_B1_M1003_g 0.0183531f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_57 VPB N_B1_M1007_g 0.0183545f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_58 VPB N_B1_c_210_n 0.00400363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A2_M1005_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_60 VPB N_A2_M1006_g 0.0245822f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_61 VPB N_A2_c_252_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A2_c_253_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A2_c_262_n 0.00788007f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_64 VPB N_A2_c_263_n 2.50157e-19 $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_65 VPB N_A2_c_254_n 0.00130531f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_66 VPB N_A2_c_257_n 0.00538302f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.53
cc_67 VPB N_A1_M1010_g 0.0183373f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_68 VPB N_A1_M1017_g 0.0183337f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_69 VPB N_A1_c_337_n 0.00400351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_297#_c_378_n 0.0198753f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_71 VPB N_A_27_297#_c_379_n 0.00189584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_297#_c_380_n 0.00752692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_297#_c_381_n 0.0042542f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_74 VPB N_A_27_297#_c_382_n 0.00363527f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_75 VPB N_A_27_297#_c_383_n 0.0129913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_297#_c_384_n 2.51509e-19 $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.53
cc_77 VPB Y 9.49571e-19 $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_78 VPB N_A_301_297#_c_505_n 0.00338184f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_566_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_80 VPB N_VPWR_c_567_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_81 VPB N_VPWR_c_568_n 0.0889431f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_82 VPB N_VPWR_c_569_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_570_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_84 VPB N_VPWR_c_571_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_85 VPB N_VPWR_c_572_n 0.0239409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_565_n 0.0561213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 N_C1_c_91_n N_B2_c_131_n 0.00827878f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_88 C1 N_A_27_297#_M1000_d 0.00294588f $X=0.15 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_89 N_C1_M1000_g N_A_27_297#_c_378_n 0.00879529f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_90 N_C1_M1004_g N_A_27_297#_c_378_n 4.50768e-19 $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_91 C1 N_A_27_297#_c_378_n 0.0230229f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_92 N_C1_c_91_n N_A_27_297#_c_378_n 0.00113906f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_93 N_C1_M1000_g N_A_27_297#_c_379_n 0.0101149f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_94 N_C1_M1004_g N_A_27_297#_c_379_n 0.0112878f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_95 N_C1_M1000_g N_A_27_297#_c_380_n 7.04098e-19 $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_96 N_C1_c_89_n N_Y_c_433_n 0.0145972f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_97 N_C1_c_88_n Y 0.00566405f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_98 N_C1_M1000_g Y 0.00118191f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_99 N_C1_c_89_n Y 0.00516881f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_100 N_C1_M1004_g Y 0.0124849f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_101 C1 Y 0.0332756f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_102 N_C1_c_91_n Y 0.0272823f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_103 N_C1_c_88_n N_Y_c_446_n 0.00490933f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_104 N_C1_c_89_n N_Y_c_446_n 0.0104706f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C1_M1000_g N_VPWR_c_568_n 0.00357835f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_106 N_C1_M1004_g N_VPWR_c_568_n 0.00357877f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_107 N_C1_M1000_g N_VPWR_c_565_n 0.00618882f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_108 N_C1_M1004_g N_VPWR_c_565_n 0.00655123f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_109 N_C1_c_88_n N_VGND_c_636_n 0.00344311f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_110 C1 N_VGND_c_636_n 0.0208398f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_111 N_C1_c_91_n N_VGND_c_636_n 0.00623008f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C1_c_88_n N_VGND_c_644_n 0.0104691f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_113 N_C1_c_89_n N_VGND_c_644_n 0.00704379f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_114 N_C1_c_88_n N_VGND_c_645_n 0.00543342f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C1_c_89_n N_VGND_c_645_n 0.00425316f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C1_c_89_n N_VGND_c_646_n 0.00335921f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B2_c_126_n N_B1_c_207_n 0.0268983f $X=1.84 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_118 N_B2_M1002_g N_B1_M1003_g 0.0428045f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B2_c_134_n N_B1_M1003_g 0.00991308f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_120 N_B2_c_127_n N_B1_c_208_n 0.0269138f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B2_M1011_g N_B1_M1007_g 0.0429016f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B2_c_134_n N_B1_M1007_g 0.0102793f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_123 N_B2_c_134_n B1 0.0391837f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_124 N_B2_c_128_n B1 0.0172311f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B2_c_129_n B1 6.66616e-19 $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B2_c_130_n B1 2.07818e-19 $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B2_c_131_n B1 0.0169874f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B2_c_134_n N_B1_c_210_n 0.00214031f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_129 N_B2_c_128_n N_B1_c_210_n 0.00458063f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B2_c_129_n N_B1_c_210_n 0.0223771f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B2_c_130_n N_B1_c_210_n 0.0223106f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B2_c_131_n N_B1_c_210_n 0.00592594f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_133 N_B2_c_127_n N_A2_c_250_n 0.0206567f $X=3.1 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 N_B2_M1011_g N_A2_M1005_g 0.0205948f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B2_c_134_n N_A2_M1005_g 5.77655e-19 $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_136 N_B2_c_128_n N_A2_M1005_g 3.59226e-19 $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_137 N_B2_M1011_g N_A2_c_252_n 3.59226e-19 $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B2_c_128_n N_A2_c_252_n 0.0307171f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B2_c_129_n N_A2_c_252_n 7.80994e-19 $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B2_c_128_n N_A2_c_253_n 7.80994e-19 $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B2_c_129_n N_A2_c_253_n 0.0197715f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B2_M1011_g N_A2_c_263_n 5.77655e-19 $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B2_c_134_n N_A2_c_263_n 0.0154679f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_144 N_B2_c_134_n N_A_27_297#_M1002_s 0.00124334f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_145 N_B2_c_131_n N_A_27_297#_M1002_s 0.00104582f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B2_c_134_n N_A_27_297#_M1007_d 0.00164852f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_147 N_B2_M1002_g N_A_27_297#_c_381_n 0.00483682f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B2_c_131_n N_A_27_297#_c_381_n 0.00801592f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B2_M1002_g N_A_27_297#_c_382_n 0.00284873f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B2_M1002_g N_A_27_297#_c_383_n 0.0113813f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B2_c_131_n N_A_27_297#_c_383_n 0.0273041f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_152 N_B2_c_134_n N_A_27_297#_c_401_n 0.0315971f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_153 N_B2_c_134_n N_A_27_297#_c_402_n 0.00677369f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_154 N_B2_c_131_n N_A_27_297#_c_402_n 0.00564423f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B2_c_134_n N_A_27_297#_c_404_n 0.0122128f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B2_c_126_n N_Y_c_433_n 0.0144101f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B2_c_134_n N_Y_c_433_n 0.0113377f $X=2.935 $Y=1.53 $X2=0 $Y2=0
cc_158 N_B2_c_130_n N_Y_c_433_n 0.00296008f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B2_c_131_n N_Y_c_433_n 0.0425899f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B2_c_126_n N_Y_c_434_n 4.06217e-19 $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_127_n N_Y_c_434_n 3.90908e-19 $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B2_c_127_n N_Y_c_436_n 0.0126004f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B2_c_128_n N_Y_c_436_n 0.0255336f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B2_c_129_n N_Y_c_436_n 0.00296008f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B2_c_131_n Y 0.0122751f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B2_c_131_n N_A_301_297#_M1002_d 0.0042535f $X=1.84 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_167 N_B2_c_134_n N_A_301_297#_M1003_s 0.00166235f $X=2.935 $Y=1.53 $X2=0
+ $Y2=0
cc_168 N_B2_c_134_n N_A_301_297#_M1011_d 0.00151125f $X=2.935 $Y=1.53 $X2=0
+ $Y2=0
cc_169 N_B2_M1002_g N_A_301_297#_c_509_n 0.00851673f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_B2_M1011_g N_A_301_297#_c_510_n 0.0121306f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B2_c_134_n N_A_301_297#_c_511_n 0.00292685f $X=2.935 $Y=1.53 $X2=0
+ $Y2=0
cc_172 N_B2_M1002_g N_VPWR_c_568_n 0.00357877f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B2_M1011_g N_VPWR_c_568_n 0.00357877f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B2_M1002_g N_VPWR_c_565_n 0.00657948f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B2_M1011_g N_VPWR_c_565_n 0.00546478f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B2_c_127_n N_VGND_c_637_n 0.00512705f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B2_c_126_n N_VGND_c_639_n 0.00421857f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B2_c_127_n N_VGND_c_639_n 0.00421857f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B2_c_126_n N_VGND_c_644_n 0.00707621f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B2_c_127_n N_VGND_c_644_n 0.00607688f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B2_c_126_n N_VGND_c_646_n 0.00481673f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B2_c_126_n N_A_383_47#_c_706_n 0.00314362f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B2_c_127_n N_A_383_47#_c_706_n 0.00328545f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_M1003_g N_A_27_297#_c_401_n 0.00924026f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1007_g N_A_27_297#_c_401_n 0.00924026f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_c_207_n N_Y_c_433_n 0.00698837f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_187 B1 N_Y_c_433_n 0.0400369f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_188 N_B1_c_207_n N_Y_c_434_n 0.00400433f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_208_n N_Y_c_434_n 0.00299412f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_210_n N_Y_c_434_n 0.00224214f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B1_c_208_n N_Y_c_436_n 0.00762805f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B1_M1003_g N_A_301_297#_c_509_n 0.00851673f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_B1_M1007_g N_A_301_297#_c_510_n 0.00851673f $X=2.68 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_B1_M1003_g N_VPWR_c_568_n 0.00357877f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_M1007_g N_VPWR_c_568_n 0.00357877f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_M1003_g N_VPWR_c_565_n 0.00525341f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_M1007_g N_VPWR_c_565_n 0.00525341f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B1_c_207_n N_VGND_c_639_n 0.00357877f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_208_n N_VGND_c_639_n 0.00357877f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B1_c_207_n N_VGND_c_644_n 0.00525237f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B1_c_208_n N_VGND_c_644_n 0.00525237f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_207_n N_A_383_47#_c_706_n 0.00924081f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B1_c_208_n N_A_383_47#_c_706_n 0.00930415f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_c_250_n N_A1_c_335_n 0.0269138f $X=3.6 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_205 N_A2_M1005_g N_A1_M1010_g 0.0433395f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A2_c_262_n N_A1_M1010_g 0.0108086f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_207 N_A2_c_251_n N_A1_c_336_n 0.0123204f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A2_M1006_g N_A1_M1017_g 0.042557f $X=4.86 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_c_262_n N_A1_M1017_g 0.0113924f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_210 N_A2_c_252_n A1 0.0133594f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A2_c_253_n A1 2.2122e-19 $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_c_262_n A1 0.0349894f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_213 N_A2_c_255_n A1 0.0172564f $X=4.82 $Y=1.175 $X2=0 $Y2=0
cc_214 N_A2_c_257_n A1 2.00336e-19 $X=4.86 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A2_c_252_n N_A1_c_337_n 0.00527477f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_c_253_n N_A1_c_337_n 0.022397f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A2_c_262_n N_A1_c_337_n 0.00214031f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_218 N_A2_c_254_n N_A1_c_337_n 0.00362491f $X=4.735 $Y=1.445 $X2=0 $Y2=0
cc_219 N_A2_c_255_n N_A1_c_337_n 0.00144374f $X=4.82 $Y=1.175 $X2=0 $Y2=0
cc_220 N_A2_c_257_n N_A1_c_337_n 0.0222902f $X=4.86 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A2_c_250_n N_Y_c_435_n 3.91234e-19 $X=3.6 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_250_n N_Y_c_436_n 0.0126004f $X=3.6 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_252_n N_Y_c_436_n 0.0255336f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A2_c_253_n N_Y_c_436_n 0.00296008f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A2_c_262_n N_Y_c_436_n 0.0071501f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_226 N_A2_c_263_n N_A_301_297#_M1011_d 0.00151125f $X=3.765 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A2_c_262_n N_A_301_297#_M1010_s 0.00165831f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_228 N_A2_c_263_n N_A_301_297#_c_511_n 0.00292685f $X=3.765 $Y=1.53 $X2=0
+ $Y2=0
cc_229 N_A2_M1005_g N_A_301_297#_c_517_n 0.0095558f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A2_c_262_n N_A_301_297#_c_517_n 0.0190307f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_231 N_A2_c_263_n N_A_301_297#_c_517_n 0.013811f $X=3.765 $Y=1.53 $X2=0 $Y2=0
cc_232 N_A2_M1006_g N_A_301_297#_c_520_n 0.01084f $X=4.86 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A2_c_262_n N_A_301_297#_c_520_n 0.0245652f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_234 A2 N_A_301_297#_c_520_n 0.00397033f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_235 N_A2_M1006_g N_A_301_297#_c_505_n 6.58332e-19 $X=4.86 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A2_c_262_n N_A_301_297#_c_505_n 0.00786716f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_237 A2 N_A_301_297#_c_505_n 0.0166332f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_238 N_A2_c_262_n N_A_301_297#_c_526_n 0.0126919f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_239 N_A2_c_262_n N_VPWR_M1005_d 0.00130005f $X=4.65 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_240 N_A2_c_263_n N_VPWR_M1005_d 3.52503e-19 $X=3.765 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_241 N_A2_c_262_n N_VPWR_M1017_d 0.00167975f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_242 N_A2_M1005_g N_VPWR_c_566_n 0.00302074f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A2_M1006_g N_VPWR_c_567_n 0.00302074f $X=4.86 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A2_M1005_g N_VPWR_c_568_n 0.00585385f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A2_M1006_g N_VPWR_c_572_n 0.00585385f $X=4.86 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A2_M1005_g N_VPWR_c_565_n 0.0061234f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A2_M1006_g N_VPWR_c_565_n 0.00700524f $X=4.86 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A2_c_250_n N_VGND_c_637_n 0.00518302f $X=3.6 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A2_c_251_n N_VGND_c_638_n 0.00482486f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_250 A2 N_VGND_c_638_n 0.0143134f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_251 N_A2_c_257_n N_VGND_c_638_n 2.31083e-19 $X=4.86 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A2_c_250_n N_VGND_c_641_n 0.00421857f $X=3.6 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A2_c_251_n N_VGND_c_641_n 0.00539841f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A2_c_250_n N_VGND_c_644_n 0.00605179f $X=3.6 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A2_c_251_n N_VGND_c_644_n 0.010585f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A2_c_250_n N_A_735_47#_c_722_n 0.0032342f $X=3.6 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A2_c_251_n N_A_735_47#_c_723_n 0.00266812f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A2_c_251_n N_A_735_47#_c_721_n 0.00529392f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A2_c_262_n N_A_735_47#_c_721_n 0.00314708f $X=4.65 $Y=1.53 $X2=0 $Y2=0
cc_260 N_A2_c_255_n N_A_735_47#_c_721_n 0.0145302f $X=4.82 $Y=1.175 $X2=0 $Y2=0
cc_261 N_A2_c_257_n N_A_735_47#_c_721_n 0.00153445f $X=4.86 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A1_c_335_n N_Y_c_435_n 0.00298551f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_c_336_n N_Y_c_435_n 0.00373093f $X=4.44 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A1_c_337_n N_Y_c_435_n 0.00224214f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A1_c_335_n N_Y_c_436_n 0.00811447f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_266 A1 N_Y_c_436_n 0.029959f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_267 N_A1_M1010_g N_A_301_297#_c_517_n 0.00956194f $X=4.02 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A1_M1017_g N_A_301_297#_c_520_n 0.00956194f $X=4.44 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A1_M1010_g N_VPWR_c_566_n 0.00157837f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A1_M1017_g N_VPWR_c_567_n 0.00157837f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A1_M1010_g N_VPWR_c_570_n 0.00585385f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A1_M1017_g N_VPWR_c_570_n 0.00585385f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A1_M1010_g N_VPWR_c_565_n 0.00591203f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A1_M1017_g N_VPWR_c_565_n 0.00591203f $X=4.44 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A1_c_335_n N_VGND_c_641_n 0.00357877f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A1_c_336_n N_VGND_c_641_n 0.00357877f $X=4.44 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A1_c_335_n N_VGND_c_644_n 0.00525237f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A1_c_336_n N_VGND_c_644_n 0.00525237f $X=4.44 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A1_c_335_n N_A_735_47#_c_722_n 0.00930415f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A1_c_336_n N_A_735_47#_c_722_n 0.0111772f $X=4.44 $Y=0.995 $X2=0 $Y2=0
cc_281 A1 N_A_735_47#_c_722_n 0.00209698f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_282 N_A_27_297#_c_379_n N_Y_M1000_s 0.00312348f $X=1.025 $Y=2.38 $X2=0 $Y2=0
cc_283 N_A_27_297#_c_381_n N_Y_c_433_n 0.00832345f $X=1.11 $Y=1.66 $X2=0 $Y2=0
cc_284 N_A_27_297#_c_379_n Y 0.0139178f $X=1.025 $Y=2.38 $X2=0 $Y2=0
cc_285 N_A_27_297#_c_383_n N_A_301_297#_M1002_d 0.00496426f $X=1.925 $Y=1.87
+ $X2=-0.19 $Y2=1.305
cc_286 N_A_27_297#_c_401_n N_A_301_297#_M1003_s 0.00317012f $X=2.765 $Y=1.87
+ $X2=0 $Y2=0
cc_287 N_A_27_297#_M1002_s N_A_301_297#_c_509_n 0.00310345f $X=1.915 $Y=1.485
+ $X2=0 $Y2=0
cc_288 N_A_27_297#_c_383_n N_A_301_297#_c_509_n 0.00506389f $X=1.925 $Y=1.87
+ $X2=0 $Y2=0
cc_289 N_A_27_297#_c_401_n N_A_301_297#_c_509_n 0.00506389f $X=2.765 $Y=1.87
+ $X2=0 $Y2=0
cc_290 N_A_27_297#_c_402_n N_A_301_297#_c_509_n 0.0112088f $X=2.05 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_M1007_d N_A_301_297#_c_510_n 0.00312348f $X=2.755 $Y=1.485
+ $X2=0 $Y2=0
cc_292 N_A_27_297#_c_401_n N_A_301_297#_c_510_n 0.00506389f $X=2.765 $Y=1.87
+ $X2=0 $Y2=0
cc_293 N_A_27_297#_c_404_n N_A_301_297#_c_510_n 0.0112811f $X=2.89 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_c_379_n N_A_301_297#_c_538_n 0.011663f $X=1.025 $Y=2.38 $X2=0
+ $Y2=0
cc_295 N_A_27_297#_c_382_n N_A_301_297#_c_538_n 0.0106948f $X=1.15 $Y=2.295
+ $X2=0 $Y2=0
cc_296 N_A_27_297#_c_383_n N_A_301_297#_c_538_n 0.0150802f $X=1.925 $Y=1.87
+ $X2=0 $Y2=0
cc_297 N_A_27_297#_c_401_n N_A_301_297#_c_541_n 0.0116461f $X=2.765 $Y=1.87
+ $X2=0 $Y2=0
cc_298 N_A_27_297#_c_379_n N_VPWR_c_568_n 0.0496214f $X=1.025 $Y=2.38 $X2=0
+ $Y2=0
cc_299 N_A_27_297#_c_380_n N_VPWR_c_568_n 0.0221816f $X=0.435 $Y=2.38 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_M1000_d N_VPWR_c_565_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_301 N_A_27_297#_M1004_d N_VPWR_c_565_n 0.00209324f $X=0.975 $Y=1.485 $X2=0
+ $Y2=0
cc_302 N_A_27_297#_M1002_s N_VPWR_c_565_n 0.00215227f $X=1.915 $Y=1.485 $X2=0
+ $Y2=0
cc_303 N_A_27_297#_M1007_d N_VPWR_c_565_n 0.0021603f $X=2.755 $Y=1.485 $X2=0
+ $Y2=0
cc_304 N_A_27_297#_c_379_n N_VPWR_c_565_n 0.0302976f $X=1.025 $Y=2.38 $X2=0
+ $Y2=0
cc_305 N_A_27_297#_c_380_n N_VPWR_c_565_n 0.0130666f $X=0.435 $Y=2.38 $X2=0
+ $Y2=0
cc_306 N_A_27_297#_c_383_n N_VPWR_c_565_n 0.00927461f $X=1.925 $Y=1.87 $X2=0
+ $Y2=0
cc_307 N_A_27_297#_c_401_n N_VPWR_c_565_n 0.00127799f $X=2.765 $Y=1.87 $X2=0
+ $Y2=0
cc_308 N_Y_M1000_s N_VPWR_c_565_n 0.00216833f $X=0.555 $Y=1.485 $X2=0 $Y2=0
cc_309 N_Y_c_433_n N_VGND_M1018_s 0.0108248f $X=2.285 $Y=0.775 $X2=0 $Y2=0
cc_310 N_Y_c_436_n N_VGND_M1019_s 0.00301529f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_311 Y N_VGND_c_636_n 5.94864e-19 $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_312 N_Y_c_436_n N_VGND_c_637_n 0.0131987f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_313 N_Y_c_433_n N_VGND_c_639_n 0.00199263f $X=2.285 $Y=0.775 $X2=0 $Y2=0
cc_314 N_Y_c_436_n N_VGND_c_639_n 0.00259935f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_315 N_Y_c_436_n N_VGND_c_641_n 0.00245397f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_316 N_Y_M1001_d N_VGND_c_644_n 0.00218509f $X=0.555 $Y=0.235 $X2=0 $Y2=0
cc_317 N_Y_M1013_s N_VGND_c_644_n 0.00216833f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_318 N_Y_M1009_s N_VGND_c_644_n 0.00216833f $X=4.095 $Y=0.235 $X2=0 $Y2=0
cc_319 N_Y_c_433_n N_VGND_c_644_n 0.0112358f $X=2.285 $Y=0.775 $X2=0 $Y2=0
cc_320 N_Y_c_436_n N_VGND_c_644_n 0.0124588f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_321 N_Y_c_446_n N_VGND_c_644_n 0.0118848f $X=0.69 $Y=0.39 $X2=0 $Y2=0
cc_322 N_Y_c_433_n N_VGND_c_645_n 0.00198695f $X=2.285 $Y=0.775 $X2=0 $Y2=0
cc_323 N_Y_c_446_n N_VGND_c_645_n 0.01433f $X=0.69 $Y=0.39 $X2=0 $Y2=0
cc_324 N_Y_c_433_n N_VGND_c_646_n 0.0528344f $X=2.285 $Y=0.775 $X2=0 $Y2=0
cc_325 N_Y_c_433_n N_A_383_47#_M1008_d 0.00191752f $X=2.285 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_326 N_Y_c_436_n N_A_383_47#_M1014_d 0.00191752f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_327 N_Y_M1013_s N_A_383_47#_c_706_n 0.00305026f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_328 N_Y_c_433_n N_A_383_47#_c_706_n 0.0140059f $X=2.285 $Y=0.775 $X2=0 $Y2=0
cc_329 N_Y_c_434_n N_A_383_47#_c_706_n 0.0166948f $X=2.635 $Y=0.775 $X2=0 $Y2=0
cc_330 N_Y_c_436_n N_A_383_47#_c_706_n 0.014941f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_331 N_Y_c_436_n N_A_735_47#_M1015_d 0.00191752f $X=4.065 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_332 N_Y_M1009_s N_A_735_47#_c_722_n 0.00305026f $X=4.095 $Y=0.235 $X2=0 $Y2=0
cc_333 N_Y_c_435_n N_A_735_47#_c_722_n 0.0153374f $X=4.23 $Y=0.73 $X2=0 $Y2=0
cc_334 N_Y_c_436_n N_A_735_47#_c_722_n 0.014941f $X=4.065 $Y=0.775 $X2=0 $Y2=0
cc_335 N_Y_c_435_n N_A_735_47#_c_721_n 0.0112424f $X=4.23 $Y=0.73 $X2=0 $Y2=0
cc_336 N_A_301_297#_c_517_n N_VPWR_M1005_d 0.00325521f $X=4.105 $Y=1.87
+ $X2=-0.19 $Y2=1.305
cc_337 N_A_301_297#_c_520_n N_VPWR_M1017_d 0.00325404f $X=4.99 $Y=1.87 $X2=0
+ $Y2=0
cc_338 N_A_301_297#_c_517_n N_VPWR_c_566_n 0.0123301f $X=4.105 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_301_297#_c_520_n N_VPWR_c_567_n 0.0123301f $X=4.99 $Y=1.87 $X2=0
+ $Y2=0
cc_340 N_A_301_297#_c_509_n N_VPWR_c_568_n 0.0329893f $X=2.345 $Y=2.38 $X2=0
+ $Y2=0
cc_341 N_A_301_297#_c_510_n N_VPWR_c_568_n 0.0515207f $X=3.225 $Y=2.38 $X2=0
+ $Y2=0
cc_342 N_A_301_297#_c_538_n N_VPWR_c_568_n 0.0151494f $X=1.63 $Y=2.3 $X2=0 $Y2=0
cc_343 N_A_301_297#_c_541_n N_VPWR_c_568_n 0.0137033f $X=2.47 $Y=2.3 $X2=0 $Y2=0
cc_344 N_A_301_297#_c_550_p N_VPWR_c_570_n 0.0142343f $X=4.23 $Y=1.96 $X2=0
+ $Y2=0
cc_345 N_A_301_297#_c_551_p N_VPWR_c_572_n 0.0142403f $X=5.075 $Y=1.96 $X2=0
+ $Y2=0
cc_346 N_A_301_297#_M1002_d N_VPWR_c_565_n 0.00207714f $X=1.505 $Y=1.485 $X2=0
+ $Y2=0
cc_347 N_A_301_297#_M1003_s N_VPWR_c_565_n 0.00213597f $X=2.335 $Y=1.485 $X2=0
+ $Y2=0
cc_348 N_A_301_297#_M1011_d N_VPWR_c_565_n 0.00306733f $X=3.175 $Y=1.485 $X2=0
+ $Y2=0
cc_349 N_A_301_297#_M1010_s N_VPWR_c_565_n 0.00223619f $X=4.095 $Y=1.485 $X2=0
+ $Y2=0
cc_350 N_A_301_297#_M1006_s N_VPWR_c_565_n 0.00349344f $X=4.935 $Y=1.485 $X2=0
+ $Y2=0
cc_351 N_A_301_297#_c_509_n N_VPWR_c_565_n 0.0204667f $X=2.345 $Y=2.38 $X2=0
+ $Y2=0
cc_352 N_A_301_297#_c_510_n N_VPWR_c_565_n 0.0315845f $X=3.225 $Y=2.38 $X2=0
+ $Y2=0
cc_353 N_A_301_297#_c_517_n N_VPWR_c_565_n 0.0123955f $X=4.105 $Y=1.87 $X2=0
+ $Y2=0
cc_354 N_A_301_297#_c_550_p N_VPWR_c_565_n 0.00955092f $X=4.23 $Y=1.96 $X2=0
+ $Y2=0
cc_355 N_A_301_297#_c_520_n N_VPWR_c_565_n 0.012579f $X=4.99 $Y=1.87 $X2=0 $Y2=0
cc_356 N_A_301_297#_c_551_p N_VPWR_c_565_n 0.00781266f $X=5.075 $Y=1.96 $X2=0
+ $Y2=0
cc_357 N_A_301_297#_c_538_n N_VPWR_c_565_n 0.00938745f $X=1.63 $Y=2.3 $X2=0
+ $Y2=0
cc_358 N_A_301_297#_c_541_n N_VPWR_c_565_n 0.00938745f $X=2.47 $Y=2.3 $X2=0
+ $Y2=0
cc_359 N_VGND_c_644_n N_A_383_47#_M1008_d 0.00215227f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_360 N_VGND_c_644_n N_A_383_47#_M1014_d 0.00215227f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_637_n N_A_383_47#_c_706_n 0.0142796f $X=3.355 $Y=0.39 $X2=0
+ $Y2=0
cc_362 N_VGND_c_639_n N_A_383_47#_c_706_n 0.0646671f $X=3.27 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_644_n N_A_383_47#_c_706_n 0.0418989f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_644_n N_A_735_47#_M1015_d 0.00215227f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_365 N_VGND_c_644_n N_A_735_47#_M1012_d 0.00215206f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_637_n N_A_735_47#_c_722_n 0.014815f $X=3.355 $Y=0.39 $X2=0 $Y2=0
cc_367 N_VGND_c_641_n N_A_735_47#_c_722_n 0.0504977f $X=4.985 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_644_n N_A_735_47#_c_722_n 0.0327385f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_641_n N_A_735_47#_c_723_n 0.015211f $X=4.985 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_644_n N_A_735_47#_c_723_n 0.00940707f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_638_n N_A_735_47#_c_721_n 0.0161415f $X=5.07 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__probec_p_8.spice.pex
* Created: Thu Aug 27 14:45:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__PROBEC_P_8%A 3 7 11 15 17 19 23 25 26 27
c86 17 0 1.32483e-19 $X=1.31 $Y=1.025
c87 11 0 1.49006e-19 $X=0.89 $Y=0.56
r88 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.16 $X2=0.985 $Y2=1.16
r89 32 34 28.8152 $w=2.76e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.16
+ $X2=0.47 $Y2=1.16
r90 27 38 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=0.985 $Y2=1.175
r91 26 38 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.985 $Y2=1.175
r92 25 26 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r93 25 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r94 17 37 56.7572 $w=2.76e-07 $l=3.25e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=0.985 $Y2=1.16
r95 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r96 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r97 9 37 16.5906 $w=2.76e-07 $l=9.5e-08 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.985 $Y2=1.16
r98 9 34 73.3478 $w=2.76e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.47 $Y2=1.16
r99 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r100 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r101 5 34 17.0164 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r102 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.985
r103 1 34 17.0164 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r104 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__PROBEC_P_8%A_27_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 85 87 88 89 90 93 99 101 104 106 112 116 118 119
+ 130
c315 118 0 1.04918e-19 $X=1.1 $Y=0.82
c316 67 0 1.42978e-20 $X=4.25 $Y=1.985
c317 59 0 4.49167e-20 $X=3.83 $Y=1.985
c318 43 0 8.80506e-20 $X=2.99 $Y=1.985
c319 31 0 1.89403e-19 $X=2.57 $Y=0.56
c320 27 0 1.90765e-19 $X=2.15 $Y=1.985
c321 19 0 1.90765e-19 $X=1.73 $Y=1.985
r322 129 130 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.67 $Y2=1.16
r323 126 127 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.83 $Y2=1.16
r324 125 126 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.41 $Y2=1.16
r325 124 125 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r326 123 124 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r327 113 129 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=3.88 $Y=1.16
+ $X2=4.25 $Y2=1.16
r328 113 127 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=3.88 $Y=1.16
+ $X2=3.83 $Y2=1.16
r329 112 113 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r330 110 123 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=2.15 $Y2=1.16
r331 110 120 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=1.73 $Y2=1.16
r332 109 112 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.84 $Y=1.16
+ $X2=3.88 $Y2=1.16
r333 109 110 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.84
+ $Y=1.16 $X2=1.84 $Y2=1.16
r334 107 119 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.507 $Y2=1.16
r335 107 109 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.84 $Y2=1.16
r336 106 116 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.445
+ $X2=1.507 $Y2=1.53
r337 105 119 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.16
r338 105 106 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.445
r339 104 119 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.075
+ $X2=1.507 $Y2=1.16
r340 103 104 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.507 $Y=0.905
+ $X2=1.507 $Y2=1.075
r341 102 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.82
+ $X2=1.1 $Y2=0.82
r342 101 103 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.42 $Y=0.82
+ $X2=1.507 $Y2=0.905
r343 101 102 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.42 $Y=0.82
+ $X2=1.185 $Y2=0.82
r344 97 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.82
r345 97 99 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.56
r346 93 95 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.1 $Y=1.63 $X2=1.1
+ $Y2=2.31
r347 91 116 26.5529 $w=1.68e-07 $l=4.07e-07 $layer=LI1_cond $X=1.1 $Y=1.53
+ $X2=1.507 $Y2=1.53
r348 91 93 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.1 $Y=1.615
+ $X2=1.1 $Y2=1.63
r349 89 91 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.53
+ $X2=1.1 $Y2=1.53
r350 89 90 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=1.53
+ $X2=0.425 $Y2=1.53
r351 87 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.82
+ $X2=1.1 $Y2=0.82
r352 87 88 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.82
+ $X2=0.345 $Y2=0.82
r353 83 88 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.345 $Y2=0.82
r354 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.56
r355 79 81 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r356 77 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r357 77 79 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r358 73 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.16
r359 73 75 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.985
r360 69 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=1.16
r361 69 71 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=0.56
r362 65 129 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.16
r363 65 67 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.985
r364 61 129 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=1.16
r365 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
r366 57 127 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.16
r367 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.985
r368 53 127 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.16
r369 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
r370 49 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r371 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r372 45 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r373 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r374 41 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r375 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r376 37 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r377 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r378 33 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r379 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r380 29 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r381 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r382 25 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r383 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r384 21 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r385 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r386 17 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r387 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r388 13 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r389 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r390 4 95 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.31
r391 4 93 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.63
r392 3 81 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r393 3 79 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r394 2 99 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.56
r395 1 85 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__PROBEC_P_8%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 43 48
+ 49 51 52 54 55 56 57 58 60 63 64 71 90 97 101 104 106 108 109 111
c138 71 0 1.51059e-19 $X=4.46 $Y=2.875
c139 63 0 1.51706e-19 $X=5.72 $Y=2.72
r140 109 114 0.16865 $w=2.8e-07 $l=3.2e-07 $layer=MET2_cond $X=5.68 $Y=2.72
+ $X2=5.36 $Y2=2.72
r141 108 109 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=5.68 $Y=2.72
+ $X2=5.68 $Y2=2.72
r142 106 108 0.0908117 $w=2.6e-07 $l=1.6e-07 $layer=MET1_cond $X=5.52 $Y=2.72
+ $X2=5.68 $Y2=2.72
r143 105 111 0.128044 $w=4.8e-07 $l=4.5e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.28 $Y2=2.72
r144 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r145 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r146 98 106 0.0939428 $w=4.8e-07 $l=2.3e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.52 $Y2=2.72
r147 98 114 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=5.36 $Y=2.72
+ $X2=5.36 $Y2=2.72
r148 98 111 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.28 $Y2=2.72
r149 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r150 95 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=4.88 $Y2=2.72
r151 95 97 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=5.29 $Y2=2.72
r152 94 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r153 94 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r154 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 91 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.72
+ $X2=4.04 $Y2=2.72
r156 91 93 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.72
+ $X2=4.37 $Y2=2.72
r157 90 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.88 $Y2=2.72
r158 90 93 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.715 $Y=2.72
+ $X2=4.37 $Y2=2.72
r159 89 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r160 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r161 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r162 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r163 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r164 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r165 68 71 0.0160563 $w=1.704e-06 $l=9.6e-07 $layer=MET5_cond $X=5.52 $Y=3.025
+ $X2=4.56 $Y2=3.025
r166 67 68 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=5.52 $Y=3.025
+ $X2=5.52 $Y2=3.025
r167 64 109 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=5.72 $Y=2.72
+ $X2=5.72 $Y2=2.72
r168 63 67 0.0123962 $w=1.18e-06 $l=3.05e-07 $layer=MET4_cond $X=5.52 $Y=2.72
+ $X2=5.52 $Y2=3.025
r169 63 64 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=5.72 $Y=2.72
+ $X2=5.72 $Y2=2.72
r170 60 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r171 58 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r172 56 88 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.99 $Y2=2.72
r173 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.2 $Y2=2.72
r174 54 85 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r175 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.36 $Y2=2.72
r176 53 88 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.99 $Y2=2.72
r177 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.36 $Y2=2.72
r178 51 82 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r179 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.52 $Y2=2.72
r180 50 85 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=2.07 $Y2=2.72
r181 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.52 $Y2=2.72
r182 48 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r183 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r184 47 82 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=1.15 $Y2=2.72
r185 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r186 43 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.88 $Y=1.66
+ $X2=4.88 $Y2=2.34
r187 41 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2.72
r188 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2.34
r189 37 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.635
+ $X2=4.04 $Y2=2.72
r190 37 39 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.04 $Y=2.635
+ $X2=4.04 $Y2=2
r191 36 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.72
+ $X2=3.2 $Y2=2.72
r192 35 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.72
+ $X2=4.04 $Y2=2.72
r193 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=2.72
+ $X2=3.365 $Y2=2.72
r194 31 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635 $X2=3.2
+ $Y2=2.72
r195 31 33 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2
r196 27 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r197 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2
r198 23 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r199 23 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2
r200 19 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r201 19 21 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2
r202 6 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2.34
r203 6 43 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.66
r204 5 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=2
r205 4 33 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2
r206 3 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2
r207 2 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
r208 1 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__PROBEC_P_8%noxref_6 1 2 3 4 5 6 7 8 27 31 33 34 35
+ 36 39 43 45 47 51 55 57 59 62 65 69 71 72 73 74 75 76 80 81 82 84 85 87 89 90
+ 93 95 105
c251 105 0 8.80506e-20 $X=2.475 $Y=1.19
c252 90 0 7.58861e-19 $X=2.05 $Y=1.36
c253 87 0 1.26775e-19 $X=2.53 $Y=1.19
c254 85 0 1.42978e-20 $X=4.75 $Y=1.19
c255 84 0 1.73336e-19 $X=4.75 $Y=1.19
c256 82 0 4.49167e-20 $X=4.36 $Y=1.19
c257 81 0 1.26775e-19 $X=2.66 $Y=1.19
c258 76 0 1.51059e-19 $X=4.417 $Y=1.185
c259 75 0 1.07952e-19 $X=4.417 $Y=0.82
c260 69 0 1.51706e-19 $X=4.46 $Y=1.755
c261 65 0 1.51706e-19 $X=4.46 $Y=0.56
r262 101 105 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=2.5 $Y=1.19 $X2=2.5
+ $Y2=1.19
r263 93 105 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=2.475 $Y=1.19
+ $X2=2.475 $Y2=1.19
r264 90 95 0.0191979 $w=4.93e-06 $l=8.9e-07 $layer=MET5_cond $X=2.05 $Y=1.36
+ $X2=1.16 $Y2=1.36
r265 89 93 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=2.475 $Y=1.19
+ $X2=2.475 $Y2=1.19
r266 89 90 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=2.05 $Y=1.36
+ $X2=2.05 $Y2=1.36
r267 87 101 0.0170272 $w=2.6e-07 $l=3e-08 $layer=MET1_cond $X=2.53 $Y=1.19
+ $X2=2.5 $Y2=1.19
r268 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.75 $Y=1.19
+ $X2=4.75 $Y2=1.19
r269 82 84 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=4.36 $Y=1.19
+ $X2=4.75 $Y2=1.19
r270 81 87 0.089401 $w=2.6e-07 $l=1.3e-07 $layer=MET1_cond $X=2.66 $Y=1.19
+ $X2=2.53 $Y2=1.19
r271 80 82 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.245 $Y=1.19
+ $X2=4.36 $Y2=1.19
r272 80 81 1.96163 $w=1.4e-07 $l=1.585e-06 $layer=MET1_cond $X=4.245 $Y=1.19
+ $X2=2.66 $Y2=1.19
r273 77 85 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=4.545 $Y=1.185
+ $X2=4.75 $Y2=1.185
r274 76 77 0.597719 $w=2.6e-07 $l=1.28e-07 $layer=LI1_cond $X=4.417 $Y=1.185
+ $X2=4.545 $Y2=1.185
r275 69 79 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.46 $Y=1.755
+ $X2=4.46 $Y2=1.615
r276 63 75 4.27425 $w=2.12e-07 $l=1.04307e-07 $layer=LI1_cond $X=4.46 $Y=0.735
+ $X2=4.417 $Y2=0.82
r277 63 65 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.46 $Y=0.735
+ $X2=4.46 $Y2=0.56
r278 62 76 5.8752 $w=2.53e-07 $l=1.3e-07 $layer=LI1_cond $X=4.417 $Y=1.055
+ $X2=4.417 $Y2=1.185
r279 61 75 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=4.417 $Y=0.905
+ $X2=4.417 $Y2=0.82
r280 61 62 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=4.417 $Y=0.905
+ $X2=4.417 $Y2=1.055
r281 60 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=1.53
+ $X2=3.62 $Y2=1.53
r282 59 79 5.12497 $w=2.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.417 $Y=1.53
+ $X2=4.417 $Y2=1.615
r283 59 76 15.5919 $w=2.53e-07 $l=3.45e-07 $layer=LI1_cond $X=4.417 $Y=1.53
+ $X2=4.417 $Y2=1.185
r284 59 60 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.29 $Y=1.53
+ $X2=3.705 $Y2=1.53
r285 58 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0.82
+ $X2=3.62 $Y2=0.82
r286 57 75 2.15711 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.29 $Y=0.82
+ $X2=4.417 $Y2=0.82
r287 57 58 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.29 $Y=0.82
+ $X2=3.705 $Y2=0.82
r288 53 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.615
+ $X2=3.62 $Y2=1.53
r289 53 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.62 $Y=1.615
+ $X2=3.62 $Y2=1.755
r290 49 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.82
r291 49 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.56
r292 48 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.53
+ $X2=2.78 $Y2=1.53
r293 47 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=1.53
+ $X2=3.62 $Y2=1.53
r294 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=1.53
+ $X2=2.865 $Y2=1.53
r295 46 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=2.78 $Y2=0.82
r296 45 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.82
+ $X2=3.62 $Y2=0.82
r297 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=0.82
+ $X2=2.865 $Y2=0.82
r298 41 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=1.615
+ $X2=2.78 $Y2=1.53
r299 41 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=1.615
+ $X2=2.78 $Y2=1.755
r300 37 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.82
r301 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.56
r302 35 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=1.53
+ $X2=2.78 $Y2=1.53
r303 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=1.53
+ $X2=2.025 $Y2=1.53
r304 33 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.82
+ $X2=2.78 $Y2=0.82
r305 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=0.82
+ $X2=2.025 $Y2=0.82
r306 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=2.025 $Y2=1.53
r307 29 31 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=1.94 $Y2=1.755
r308 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=2.025 $Y2=0.82
r309 25 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.56
r310 8 69 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=1.755
r311 7 55 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.755
r312 6 43 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.755
r313 5 31 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.755
r314 4 65 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.56
r315 3 51 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.56
r316 2 39 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.56
r317 1 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__PROBEC_P_8%VGND 1 2 3 4 5 6 21 25 29 33 35 39 43 46
+ 47 49 50 51 52 53 55 58 62 65 70 75 87 94 98 101 104 106 108 109 111
c151 65 0 1.07952e-19 $X=4.46 $Y=-0.455
c152 58 0 1.51706e-19 $X=5.52 $Y=-0.304
r153 109 114 0.16865 $w=2.8e-07 $l=3.2e-07 $layer=MET2_cond $X=5.68 $Y=0
+ $X2=5.36 $Y2=0
r154 108 109 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=5.68 $Y=0 $X2=5.68
+ $Y2=0
r155 106 108 0.0908117 $w=2.6e-07 $l=1.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.68 $Y2=0
r156 105 111 0.128044 $w=4.8e-07 $l=4.5e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.28 $Y2=0
r157 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r158 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r159 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r160 95 106 0.0939428 $w=4.8e-07 $l=2.3e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.52 $Y2=0
r161 95 114 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=5.36 $Y=0 $X2=5.36
+ $Y2=0
r162 95 111 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.28 $Y2=0
r163 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r164 92 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=4.88 $Y2=0
r165 92 94 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.29
+ $Y2=0
r166 91 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r167 91 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r168 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r169 88 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0
+ $X2=4.04 $Y2=0
r170 88 90 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0
+ $X2=4.37 $Y2=0
r171 87 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.88 $Y2=0
r172 87 90 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.37
+ $Y2=0
r173 86 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r174 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r175 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r176 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r177 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r178 80 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r179 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r180 77 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r181 77 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r182 70 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r183 62 109 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=5.72 $Y=0 $X2=5.72
+ $Y2=0
r184 59 65 0.0160563 $w=1.704e-06 $l=9.6e-07 $layer=MET5_cond $X=5.52 $Y=-0.305
+ $X2=4.56 $Y2=-0.305
r185 58 62 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=5.72 $Y=0
+ $X2=5.72 $Y2=0
r186 58 59 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=5.52
+ $Y=-0.304 $X2=5.52 $Y2=-0.304
r187 55 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r188 55 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r189 53 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=0
+ $X2=0.515 $Y2=0
r190 53 75 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r191 51 85 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.99
+ $Y2=0
r192 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.2
+ $Y2=0
r193 49 82 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=0
+ $X2=2.07 $Y2=0
r194 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.36
+ $Y2=0
r195 48 85 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=2.99 $Y2=0
r196 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.36
+ $Y2=0
r197 46 79 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.15 $Y2=0
r198 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r199 45 82 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=0
+ $X2=2.07 $Y2=0
r200 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r201 41 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r202 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.38
r203 37 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r204 37 39 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.4
r205 36 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.2
+ $Y2=0
r206 35 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0
+ $X2=4.04 $Y2=0
r207 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=0
+ $X2=3.365 $Y2=0
r208 31 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.085 $X2=3.2
+ $Y2=0
r209 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0.4
r210 27 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r211 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.4
r212 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r213 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r214 19 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r215 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r216 6 43 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.38
r217 5 39 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.4
r218 4 33 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.4
r219 3 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.4
r220 2 25 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r221 1 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__PROBEC_P_8%X 1 4 8 10
c39 10 0 6.59968e-20 $X=1.06 $Y=1.36
c40 4 0 1.32483e-19 $X=-0.549 $Y=1.36
r41 5 10 0.0302819 $w=1.6e-06 $l=1.609e-06 $layer=MET5_cond $X=-0.549 $Y=1.36
+ $X2=1.06 $Y2=1.36
r42 4 8 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=-0.124 $Y=1.19
+ $X2=-0.124 $Y2=1.19
r43 4 5 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=-0.549 $Y=1.36
+ $X2=-0.549 $Y2=1.36
r44 1 8 0.033007 $w=3.2e-07 $l=2.06e-07 $layer=MET3_cond $X=-0.33 $Y=1.19
+ $X2=-0.124 $Y2=1.19
.ends


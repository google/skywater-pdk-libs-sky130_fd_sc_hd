* File: sky130_fd_sc_hd__or3b_4.spice
* Created: Thu Aug 27 14:43:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or3b_4.pex.spice"
.subckt sky130_fd_sc_hd__or3b_4  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_C_N_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1013_d N_A_176_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_176_21#_M1003_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1003_d N_A_176_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.3
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_176_21#_M1012_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.8
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1009 N_A_176_21#_M1009_d N_A_M1009_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_176_21#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_A_176_21#_M1008_d N_A_27_47#_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VPWR_M1014_d N_C_N_M1014_g N_A_27_47#_M1014_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=70.4866 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1014_d N_A_176_21#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.205282 AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_176_21#_M1007_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1007_d N_A_176_21#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_176_21#_M1015_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1000 A_542_297# N_A_M1000_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75002.1 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1011 A_626_297# N_B_M1011_g A_542_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=15.7403 M=1 R=6.66667 SA=75002.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_A_176_21#_M1001_d N_A_27_47#_M1001_g A_626_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.165 PD=2.52 PS=1.33 NRD=0 NRS=21.6503 M=1 R=6.66667 SA=75003
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__or3b_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o221a_4.pxi.spice
* Created: Tue Sep  1 19:22:39 2020
* 
x_PM_SKY130_FD_SC_HD__O221A_4%C1 N_C1_c_118_n N_C1_M1013_g N_C1_M1003_g
+ N_C1_c_119_n N_C1_M1027_g N_C1_M1019_g C1 N_C1_c_121_n C1
+ PM_SKY130_FD_SC_HD__O221A_4%C1
x_PM_SKY130_FD_SC_HD__O221A_4%B1 N_B1_c_161_n N_B1_M1018_g N_B1_M1001_g
+ N_B1_M1020_g N_B1_M1004_g N_B1_c_169_n N_B1_c_162_n N_B1_c_163_n B1 B1
+ N_B1_c_164_n N_B1_c_165_n N_B1_c_166_n PM_SKY130_FD_SC_HD__O221A_4%B1
x_PM_SKY130_FD_SC_HD__O221A_4%B2 N_B2_c_245_n N_B2_M1016_g N_B2_M1022_g
+ N_B2_c_246_n N_B2_M1024_g N_B2_M1025_g B2 N_B2_c_248_n
+ PM_SKY130_FD_SC_HD__O221A_4%B2
x_PM_SKY130_FD_SC_HD__O221A_4%A1 N_A1_M1008_g N_A1_M1009_g N_A1_c_286_n
+ N_A1_M1021_g N_A1_M1023_g N_A1_c_295_n N_A1_c_287_n N_A1_c_288_n N_A1_c_289_n
+ A1 N_A1_c_291_n N_A1_c_292_n PM_SKY130_FD_SC_HD__O221A_4%A1
x_PM_SKY130_FD_SC_HD__O221A_4%A2 N_A2_c_375_n N_A2_M1007_g N_A2_M1012_g
+ N_A2_c_376_n N_A2_M1014_g N_A2_M1015_g A2 N_A2_c_377_n N_A2_c_378_n
+ PM_SKY130_FD_SC_HD__O221A_4%A2
x_PM_SKY130_FD_SC_HD__O221A_4%A_109_47# N_A_109_47#_M1013_s N_A_109_47#_M1003_s
+ N_A_109_47#_M1022_s N_A_109_47#_M1012_s N_A_109_47#_c_422_n
+ N_A_109_47#_M1006_g N_A_109_47#_M1000_g N_A_109_47#_c_423_n
+ N_A_109_47#_M1010_g N_A_109_47#_M1002_g N_A_109_47#_c_424_n
+ N_A_109_47#_M1011_g N_A_109_47#_M1005_g N_A_109_47#_c_425_n
+ N_A_109_47#_M1017_g N_A_109_47#_M1026_g N_A_109_47#_c_432_n
+ N_A_109_47#_c_439_n N_A_109_47#_c_503_p N_A_109_47#_c_440_n
+ N_A_109_47#_c_456_n N_A_109_47#_c_472_n N_A_109_47#_c_476_n
+ N_A_109_47#_c_433_n N_A_109_47#_c_479_n N_A_109_47#_c_540_p
+ N_A_109_47#_c_441_n N_A_109_47#_c_426_n N_A_109_47#_c_449_n
+ N_A_109_47#_c_462_n N_A_109_47#_c_480_n N_A_109_47#_c_435_n
+ N_A_109_47#_c_427_n PM_SKY130_FD_SC_HD__O221A_4%A_109_47#
x_PM_SKY130_FD_SC_HD__O221A_4%VPWR N_VPWR_M1003_d N_VPWR_M1019_d N_VPWR_M1004_s
+ N_VPWR_M1023_d N_VPWR_M1002_s N_VPWR_M1026_s N_VPWR_c_591_n N_VPWR_c_592_n
+ N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n
+ N_VPWR_c_598_n N_VPWR_c_599_n VPWR N_VPWR_c_600_n N_VPWR_c_601_n
+ N_VPWR_c_602_n N_VPWR_c_590_n N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n
+ N_VPWR_c_607_n N_VPWR_c_608_n PM_SKY130_FD_SC_HD__O221A_4%VPWR
x_PM_SKY130_FD_SC_HD__O221A_4%A_277_297# N_A_277_297#_M1001_d
+ N_A_277_297#_M1025_d N_A_277_297#_c_701_n N_A_277_297#_c_709_n
+ N_A_277_297#_c_710_n PM_SKY130_FD_SC_HD__O221A_4%A_277_297#
x_PM_SKY130_FD_SC_HD__O221A_4%A_717_297# N_A_717_297#_M1009_s
+ N_A_717_297#_M1015_d N_A_717_297#_c_721_n N_A_717_297#_c_729_n
+ N_A_717_297#_c_730_n PM_SKY130_FD_SC_HD__O221A_4%A_717_297#
x_PM_SKY130_FD_SC_HD__O221A_4%X N_X_M1006_d N_X_M1011_d N_X_M1000_d N_X_M1005_d
+ N_X_c_749_n N_X_c_787_n N_X_c_752_n N_X_c_754_n N_X_c_739_n N_X_c_740_n
+ N_X_c_743_n N_X_c_744_n N_X_c_741_n N_X_c_776_n N_X_c_793_n N_X_c_745_n
+ N_X_c_746_n X PM_SKY130_FD_SC_HD__O221A_4%X
x_PM_SKY130_FD_SC_HD__O221A_4%A_27_47# N_A_27_47#_M1013_d N_A_27_47#_M1027_d
+ N_A_27_47#_M1016_d N_A_27_47#_M1020_s N_A_27_47#_c_814_n N_A_27_47#_c_815_n
+ N_A_27_47#_c_821_n N_A_27_47#_c_816_n N_A_27_47#_c_817_n N_A_27_47#_c_847_p
+ PM_SKY130_FD_SC_HD__O221A_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O221A_4%A_277_47# N_A_277_47#_M1018_d N_A_277_47#_M1024_s
+ N_A_277_47#_M1008_d N_A_277_47#_M1014_s N_A_277_47#_c_856_n
+ N_A_277_47#_c_857_n N_A_277_47#_c_877_n N_A_277_47#_c_858_n
+ N_A_277_47#_c_882_n N_A_277_47#_c_859_n N_A_277_47#_c_860_n
+ PM_SKY130_FD_SC_HD__O221A_4%A_277_47#
x_PM_SKY130_FD_SC_HD__O221A_4%VGND N_VGND_M1008_s N_VGND_M1007_d N_VGND_M1021_s
+ N_VGND_M1010_s N_VGND_M1017_s N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n
+ N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n
+ N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n VGND
+ N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n N_VGND_c_938_n
+ PM_SKY130_FD_SC_HD__O221A_4%VGND
cc_1 VNB N_C1_c_118_n 0.0216914f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_C1_c_119_n 0.0157516f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB C1 0.00832616f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_C1_c_121_n 0.0548155f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B1_c_161_n 0.0163525f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B1_c_162_n 0.00406355f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_7 VNB N_B1_c_163_n 0.0229117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B1_c_164_n 0.0193711f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_9 VNB N_B1_c_165_n 0.00498181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_166_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B2_c_245_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_12 VNB N_B2_c_246_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_13 VNB B2 0.00159717f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB N_B2_c_248_n 0.0301299f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_15 VNB N_A1_c_286_n 0.0163539f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_16 VNB N_A1_c_287_n 0.00734966f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_17 VNB N_A1_c_288_n 0.0241564f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_18 VNB N_A1_c_289_n 6.01426e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB A1 0.00643559f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.175
cc_20 VNB N_A1_c_291_n 0.0217006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A1_c_292_n 0.0206213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_c_375_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_23 VNB N_A2_c_376_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_24 VNB N_A2_c_377_n 0.0026962f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_25 VNB N_A2_c_378_n 0.0307879f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_26 VNB N_A_109_47#_c_422_n 0.0161429f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_27 VNB N_A_109_47#_c_423_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_109_47#_c_424_n 0.0157964f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_29 VNB N_A_109_47#_c_425_n 0.0191719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_109_47#_c_426_n 0.00101507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_109_47#_c_427_n 0.065651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_590_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_739_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_740_n 0.00222337f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.175
cc_35 VNB N_X_c_741_n 0.0124437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB X 0.0220587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_814_n 0.00972331f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_38 VNB N_A_27_47#_c_815_n 0.0176737f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_39 VNB N_A_27_47#_c_816_n 0.00212357f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_40 VNB N_A_27_47#_c_817_n 0.00292106f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_41 VNB N_A_277_47#_c_856_n 0.00788475f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_42 VNB N_A_277_47#_c_857_n 0.0186463f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_43 VNB N_A_277_47#_c_858_n 0.00511104f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_44 VNB N_A_277_47#_c_859_n 7.13203e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_277_47#_c_860_n 0.00356355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_922_n 0.00801397f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_47 VNB N_VGND_c_923_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_48 VNB N_VGND_c_924_n 0.00559268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_925_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_926_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_927_n 0.0173887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_928_n 0.0737806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_929_n 0.00458525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_930_n 0.0166557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_931_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_932_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_933_n 0.00326325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_934_n 0.0166796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_935_n 0.0186844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_936_n 0.369769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_937_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_938_n 0.00487447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VPB N_C1_M1003_g 0.0251042f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_64 VPB N_C1_M1019_g 0.0180908f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_65 VPB N_C1_c_121_n 0.0135355f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_66 VPB N_B1_M1001_g 0.0172552f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_B1_M1004_g 0.0223541f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_B1_c_169_n 0.00738794f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_69 VPB N_B1_c_162_n 0.00272228f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_70 VPB N_B1_c_163_n 0.00465795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_B1_c_164_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_72 VPB N_B1_c_165_n 0.00266467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B2_M1022_g 0.0183523f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_74 VPB N_B2_M1025_g 0.0183554f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_75 VPB N_B2_c_248_n 0.00401205f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_76 VPB N_A1_M1009_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_77 VPB N_A1_M1023_g 0.0181634f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_78 VPB N_A1_c_295_n 0.00703656f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_79 VPB N_A1_c_287_n 0.00395225f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_80 VPB N_A1_c_288_n 0.00501007f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_81 VPB N_A1_c_289_n 0.00134466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A1_c_292_n 0.00460764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A2_M1012_g 0.0183623f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_84 VPB N_A2_M1015_g 0.0183486f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_85 VPB N_A2_c_378_n 0.00405299f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_86 VPB N_A_109_47#_M1000_g 0.0178567f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_87 VPB N_A_109_47#_M1002_g 0.0184409f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_88 VPB N_A_109_47#_M1005_g 0.0180964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_109_47#_M1026_g 0.0219226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_109_47#_c_432_n 8.73209e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_109_47#_c_433_n 0.00145536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_109_47#_c_426_n 0.00112774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_109_47#_c_435_n 0.00358247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_109_47#_c_427_n 0.0107251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_591_n 0.0116091f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_96 VPB N_VPWR_c_592_n 0.00760781f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_97 VPB N_VPWR_c_593_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_98 VPB N_VPWR_c_594_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_595_n 0.0167545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_596_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_597_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_598_n 0.0349357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_599_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_600_n 0.0163654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_601_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_602_n 0.0204409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_590_n 0.0650947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_604_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_605_n 0.0349195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_606_n 0.0226617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_607_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_608_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_X_c_743_n 5.78753e-19 $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_114 VPB N_X_c_744_n 0.00162727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_X_c_745_n 7.30684e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_X_c_746_n 0.00204415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB X 0.0210324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 N_C1_c_119_n N_B1_c_161_n 0.0117542f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_119 N_C1_M1019_g N_B1_M1001_g 0.042145f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_120 N_C1_c_121_n N_B1_c_164_n 0.0221541f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C1_c_121_n N_B1_c_165_n 0.00431609f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C1_M1003_g N_A_109_47#_c_432_n 5.02033e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_123 N_C1_M1019_g N_A_109_47#_c_432_n 0.00185021f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_124 N_C1_M1019_g N_A_109_47#_c_439_n 0.00337644f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_125 N_C1_M1019_g N_A_109_47#_c_440_n 0.0116537f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C1_c_118_n N_A_109_47#_c_441_n 0.00407862f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_127 N_C1_c_119_n N_A_109_47#_c_441_n 0.00268818f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C1_c_118_n N_A_109_47#_c_426_n 0.00265667f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_129 N_C1_M1003_g N_A_109_47#_c_426_n 0.00296785f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_130 N_C1_c_119_n N_A_109_47#_c_426_n 0.00290895f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_131 N_C1_M1019_g N_A_109_47#_c_426_n 0.0022611f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_132 C1 N_A_109_47#_c_426_n 0.014625f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_133 N_C1_c_121_n N_A_109_47#_c_426_n 0.0229217f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_134 N_C1_M1019_g N_A_109_47#_c_449_n 0.00117879f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C1_M1003_g N_VPWR_c_592_n 0.00412378f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_136 C1 N_VPWR_c_592_n 0.0193718f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_137 N_C1_c_121_n N_VPWR_c_592_n 0.00610779f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_138 N_C1_M1019_g N_VPWR_c_593_n 0.00153671f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_139 N_C1_M1003_g N_VPWR_c_600_n 0.00583607f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_140 N_C1_M1019_g N_VPWR_c_600_n 0.00585385f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_141 N_C1_M1003_g N_VPWR_c_590_n 0.0113526f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_142 N_C1_M1019_g N_VPWR_c_590_n 0.00593664f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_143 N_C1_c_118_n N_A_27_47#_c_815_n 2.3414e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_144 C1 N_A_27_47#_c_815_n 0.0198144f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_145 N_C1_c_121_n N_A_27_47#_c_815_n 0.00595621f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_146 N_C1_c_118_n N_A_27_47#_c_821_n 0.0119436f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_147 N_C1_c_119_n N_A_27_47#_c_821_n 0.0127333f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_148 C1 N_A_27_47#_c_821_n 0.00170999f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_149 N_C1_c_121_n N_A_27_47#_c_821_n 3.07604e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_150 N_C1_c_118_n N_VGND_c_928_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C1_c_119_n N_VGND_c_928_n 0.00357877f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C1_c_118_n N_VGND_c_936_n 0.00617937f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_153 N_C1_c_119_n N_VGND_c_936_n 0.00525237f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B1_c_161_n N_B2_c_245_n 0.0267413f $X=1.31 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_155 N_B1_M1001_g N_B2_M1022_g 0.0439673f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B1_c_169_n N_B2_M1022_g 0.00999193f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B1_c_166_n N_B2_c_246_n 0.0270078f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B1_M1004_g N_B2_M1025_g 0.0439959f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B1_c_169_n N_B2_M1025_g 0.0102793f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_160 N_B1_c_169_n B2 0.0392598f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_161 N_B1_c_162_n B2 0.0172313f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_162 N_B1_c_163_n B2 6.72338e-19 $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_163 N_B1_c_164_n B2 2.00573e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B1_c_165_n B2 0.0168834f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_169_n N_B2_c_248_n 0.00214031f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_166 N_B1_c_162_n N_B2_c_248_n 0.0045316f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B1_c_163_n N_B2_c_248_n 0.0212121f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_c_164_n N_B2_c_248_n 0.0222883f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B1_c_165_n N_B2_c_248_n 0.00592644f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_169_n N_A1_M1009_g 5.97813e-19 $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_171 N_B1_c_162_n N_A1_M1009_g 3.83263e-19 $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_172 N_B1_M1004_g N_A1_c_287_n 0.00176113f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_c_169_n N_A1_c_287_n 0.0111855f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_174 N_B1_c_162_n N_A1_c_287_n 0.02397f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B1_c_163_n N_A1_c_287_n 0.00115452f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B1_c_162_n N_A1_c_288_n 6.13515e-19 $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B1_c_163_n N_A1_c_288_n 0.00577551f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B1_c_169_n N_A_109_47#_M1022_s 0.00165831f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_179 N_B1_M1001_g N_A_109_47#_c_439_n 8.39534e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1001_g N_A_109_47#_c_440_n 0.0115072f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B1_c_169_n N_A_109_47#_c_440_n 0.0157986f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_182 N_B1_c_164_n N_A_109_47#_c_440_n 3.01349e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B1_c_165_n N_A_109_47#_c_440_n 0.0294941f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B1_M1004_g N_A_109_47#_c_456_n 0.0136543f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_c_169_n N_A_109_47#_c_456_n 0.0362387f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_186 N_B1_c_161_n N_A_109_47#_c_441_n 5.18533e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_M1001_g N_A_109_47#_c_426_n 2.21952e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B1_c_164_n N_A_109_47#_c_426_n 6.28465e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B1_c_165_n N_A_109_47#_c_426_n 0.0411536f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B1_c_169_n N_A_109_47#_c_462_n 0.0120079f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_191 N_B1_c_165_n N_VPWR_M1019_d 0.00295416f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B1_c_169_n N_VPWR_M1004_s 0.00207834f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_193 N_B1_M1001_g N_VPWR_c_593_n 0.00304122f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B1_M1001_g N_VPWR_c_590_n 0.00590802f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_M1004_g N_VPWR_c_590_n 0.00726073f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_M1001_g N_VPWR_c_605_n 0.00583607f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_M1004_g N_VPWR_c_605_n 0.00585385f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B1_M1004_g N_VPWR_c_606_n 0.00509285f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B1_c_169_n N_A_277_297#_M1001_d 0.00113984f $X=2.415 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_200 N_B1_c_165_n N_A_277_297#_M1001_d 0.00115696f $X=1.31 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_201 N_B1_c_169_n N_A_277_297#_M1025_d 0.00164895f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_202 N_B1_c_164_n N_A_27_47#_c_816_n 2.30167e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B1_c_165_n N_A_27_47#_c_816_n 0.0144623f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B1_c_161_n N_A_27_47#_c_817_n 0.0105068f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B1_c_165_n N_A_27_47#_c_817_n 0.00390962f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B1_c_166_n N_A_27_47#_c_817_n 0.00917393f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B1_c_161_n N_A_277_47#_c_856_n 0.00372494f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B1_c_169_n N_A_277_47#_c_856_n 0.0115695f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_209 N_B1_c_164_n N_A_277_47#_c_856_n 0.00149384f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B1_c_165_n N_A_277_47#_c_856_n 0.0134879f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B1_c_163_n N_A_277_47#_c_857_n 0.001729f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B1_c_166_n N_A_277_47#_c_857_n 0.00973721f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_162_n N_A_277_47#_c_859_n 0.0258144f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B1_c_163_n N_A_277_47#_c_859_n 0.00124486f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_215 N_B1_c_166_n N_A_277_47#_c_859_n 0.00532475f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_166_n N_VGND_c_922_n 0.00226541f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_161_n N_VGND_c_928_n 0.00357877f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_166_n N_VGND_c_928_n 0.00357877f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_161_n N_VGND_c_936_n 0.00528062f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B1_c_166_n N_VGND_c_936_n 0.00657948f $X=2.58 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B2_M1022_g N_A_109_47#_c_440_n 0.00924026f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_222 N_B2_M1025_g N_A_109_47#_c_456_n 0.00924026f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B2_M1022_g N_VPWR_c_590_n 0.00525237f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B2_M1025_g N_VPWR_c_590_n 0.00525237f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B2_M1022_g N_VPWR_c_605_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B2_M1025_g N_VPWR_c_605_n 0.00357877f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B2_M1022_g N_A_277_297#_c_701_n 0.00851673f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_B2_M1025_g N_A_277_297#_c_701_n 0.00856088f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_B2_c_245_n N_A_27_47#_c_817_n 0.00886996f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B2_c_246_n N_A_27_47#_c_817_n 0.00886996f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B2_c_245_n N_A_277_47#_c_856_n 0.0113911f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B2_c_246_n N_A_277_47#_c_856_n 0.0109578f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_233 B2 N_A_277_47#_c_856_n 0.0405927f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_234 N_B2_c_248_n N_A_277_47#_c_856_n 0.00224214f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B2_c_245_n N_VGND_c_928_n 0.00357877f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B2_c_246_n N_VGND_c_928_n 0.00357877f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B2_c_245_n N_VGND_c_936_n 0.00525341f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B2_c_246_n N_VGND_c_936_n 0.00525341f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A1_c_291_n N_A2_c_375_n 0.0244283f $X=3.445 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_240 N_A1_M1009_g N_A2_M1012_g 0.0244283f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A1_c_295_n N_A2_M1012_g 0.00998745f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_242 N_A1_c_286_n N_A2_c_376_n 0.0124239f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A1_M1023_g N_A2_M1015_g 0.0433032f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A1_c_295_n N_A2_M1015_g 0.0111274f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_245 N_A1_c_295_n N_A2_c_377_n 0.041432f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_246 N_A1_c_287_n N_A2_c_377_n 0.0180739f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A1_c_288_n N_A2_c_377_n 7.22994e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_248 A1 N_A2_c_377_n 0.0170581f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_249 N_A1_c_295_n N_A2_c_378_n 0.00214031f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_250 N_A1_c_287_n N_A2_c_378_n 0.00480848f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A1_c_288_n N_A2_c_378_n 0.0244283f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A1_c_289_n N_A2_c_378_n 0.00409887f $X=4.65 $Y=1.445 $X2=0 $Y2=0
cc_253 A1 N_A2_c_378_n 0.00143632f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_254 N_A1_c_292_n N_A2_c_378_n 0.022243f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A1_c_295_n N_A_109_47#_M1012_s 0.00165831f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_256 N_A1_c_286_n N_A_109_47#_c_422_n 0.012217f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A1_M1023_g N_A_109_47#_M1000_g 0.0413591f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A1_M1009_g N_A_109_47#_c_456_n 0.0136543f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A1_c_295_n N_A_109_47#_c_456_n 0.021464f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_260 N_A1_c_287_n N_A_109_47#_c_456_n 0.0409127f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_c_288_n N_A_109_47#_c_456_n 4.10999e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A1_M1023_g N_A_109_47#_c_472_n 0.0122904f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_c_295_n N_A_109_47#_c_472_n 0.0276413f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_264 A1 N_A_109_47#_c_472_n 0.00526294f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_265 N_A1_c_292_n N_A_109_47#_c_472_n 0.00105533f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A1_M1023_g N_A_109_47#_c_476_n 0.00365504f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A1_M1023_g N_A_109_47#_c_433_n 3.59092e-19 $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A1_c_289_n N_A_109_47#_c_433_n 0.00554134f $X=4.65 $Y=1.445 $X2=0 $Y2=0
cc_269 A1 N_A_109_47#_c_479_n 0.0172581f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_270 N_A1_c_295_n N_A_109_47#_c_480_n 0.0120079f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_271 N_A1_M1023_g N_A_109_47#_c_435_n 0.00114998f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A1_c_295_n N_A_109_47#_c_435_n 0.0124942f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_273 A1 N_A_109_47#_c_435_n 0.00457456f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_274 N_A1_c_289_n N_A_109_47#_c_427_n 5.4516e-19 $X=4.65 $Y=1.445 $X2=0 $Y2=0
cc_275 A1 N_A_109_47#_c_427_n 0.00154253f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_276 N_A1_c_292_n N_A_109_47#_c_427_n 0.0226678f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A1_c_287_n N_VPWR_M1004_s 0.00719325f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_278 N_A1_M1023_g N_VPWR_c_594_n 0.00302074f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A1_M1009_g N_VPWR_c_598_n 0.00585385f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A1_M1023_g N_VPWR_c_598_n 0.00585385f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A1_M1009_g N_VPWR_c_590_n 0.00723564f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A1_M1023_g N_VPWR_c_590_n 0.00593924f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A1_M1009_g N_VPWR_c_606_n 0.00518337f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A1_c_295_n N_A_717_297#_M1009_s 0.00166235f $X=4.525 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_285 N_A1_c_295_n N_A_717_297#_M1015_d 0.00166402f $X=4.525 $Y=1.53 $X2=0
+ $Y2=0
cc_286 N_A1_c_287_n N_A_277_47#_c_857_n 0.044257f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A1_c_288_n N_A_277_47#_c_857_n 0.003211f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A1_c_291_n N_A_277_47#_c_857_n 0.0112531f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A1_c_291_n N_A_277_47#_c_877_n 0.0108131f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A1_c_286_n N_A_277_47#_c_858_n 0.00252178f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A1_c_295_n N_A_277_47#_c_858_n 0.00567223f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_292 A1 N_A_277_47#_c_858_n 0.016536f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_293 N_A1_c_292_n N_A_277_47#_c_858_n 0.00153559f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A1_c_286_n N_A_277_47#_c_882_n 0.00513121f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A1_c_295_n N_A_277_47#_c_860_n 0.00640335f $X=4.525 $Y=1.53 $X2=0 $Y2=0
cc_296 N_A1_c_287_n N_A_277_47#_c_860_n 0.00423127f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A1_c_291_n N_A_277_47#_c_860_n 0.0011539f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A1_c_291_n N_VGND_c_922_n 0.00320738f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A1_c_286_n N_VGND_c_924_n 0.00159991f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_300 A1 N_VGND_c_924_n 0.0118366f $X=4.76 $Y=1.105 $X2=0 $Y2=0
cc_301 N_A1_c_292_n N_VGND_c_924_n 2.31083e-19 $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A1_c_291_n N_VGND_c_930_n 0.00422241f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A1_c_286_n N_VGND_c_932_n 0.00541359f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A1_c_286_n N_VGND_c_936_n 0.00955595f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A1_c_291_n N_VGND_c_936_n 0.00704983f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A2_M1012_g N_A_109_47#_c_456_n 0.00924026f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A2_M1015_g N_A_109_47#_c_472_n 0.00924026f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A2_M1012_g N_VPWR_c_598_n 0.00357877f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A2_M1015_g N_VPWR_c_598_n 0.00357877f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A2_M1012_g N_VPWR_c_590_n 0.00525237f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A2_M1015_g N_VPWR_c_590_n 0.00525237f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A2_M1012_g N_A_717_297#_c_721_n 0.00851673f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A2_M1015_g N_A_717_297#_c_721_n 0.00851673f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A2_c_375_n N_A_277_47#_c_877_n 0.0061357f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_c_376_n N_A_277_47#_c_877_n 4.92877e-19 $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A2_c_375_n N_A_277_47#_c_858_n 0.00870364f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A2_c_376_n N_A_277_47#_c_858_n 0.0106817f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A2_c_377_n N_A_277_47#_c_858_n 0.0333876f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A2_c_378_n N_A_277_47#_c_858_n 0.00222133f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A2_c_375_n N_A_277_47#_c_882_n 5.22217e-19 $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A2_c_376_n N_A_277_47#_c_882_n 0.00630957f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A2_c_375_n N_A_277_47#_c_860_n 0.0013024f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A2_c_377_n N_A_277_47#_c_860_n 0.00911001f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A2_c_375_n N_VGND_c_923_n 0.00146448f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A2_c_376_n N_VGND_c_923_n 0.00146448f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A2_c_375_n N_VGND_c_930_n 0.00423334f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A2_c_376_n N_VGND_c_932_n 0.00423334f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A2_c_375_n N_VGND_c_936_n 0.0057435f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A2_c_376_n N_VGND_c_936_n 0.0057435f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_109_47#_c_440_n N_VPWR_M1019_d 0.00316782f $X=1.825 $Y=1.87 $X2=0
+ $Y2=0
cc_331 N_A_109_47#_c_456_n N_VPWR_M1004_s 0.0253174f $X=4.015 $Y=1.87 $X2=0
+ $Y2=0
cc_332 N_A_109_47#_c_472_n N_VPWR_M1023_d 0.00288072f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_333 N_A_109_47#_c_476_n N_VPWR_M1023_d 0.00215579f $X=5.06 $Y=1.785 $X2=0
+ $Y2=0
cc_334 N_A_109_47#_c_435_n N_VPWR_M1023_d 0.00140313f $X=5.29 $Y=1.53 $X2=0
+ $Y2=0
cc_335 N_A_109_47#_c_432_n N_VPWR_c_592_n 0.0143011f $X=0.705 $Y=1.585 $X2=0
+ $Y2=0
cc_336 N_A_109_47#_c_440_n N_VPWR_c_593_n 0.0123301f $X=1.825 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_109_47#_M1000_g N_VPWR_c_594_n 0.00157837f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_109_47#_c_472_n N_VPWR_c_594_n 0.0126457f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_109_47#_M1000_g N_VPWR_c_595_n 0.00585385f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_109_47#_M1002_g N_VPWR_c_595_n 0.00585385f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_109_47#_M1002_g N_VPWR_c_596_n 0.00157837f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_109_47#_M1005_g N_VPWR_c_596_n 0.00157837f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_109_47#_M1026_g N_VPWR_c_597_n 0.00338128f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_109_47#_c_503_p N_VPWR_c_600_n 0.0142343f $X=0.68 $Y=2.3 $X2=0 $Y2=0
cc_345 N_A_109_47#_M1005_g N_VPWR_c_601_n 0.00585385f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_109_47#_M1026_g N_VPWR_c_601_n 0.00585385f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_347 N_A_109_47#_M1003_s N_VPWR_c_590_n 0.00284632f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_348 N_A_109_47#_M1022_s N_VPWR_c_590_n 0.00215227f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_349 N_A_109_47#_M1012_s N_VPWR_c_590_n 0.00215227f $X=4.005 $Y=1.485 $X2=0
+ $Y2=0
cc_350 N_A_109_47#_M1000_g N_VPWR_c_590_n 0.00957154f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A_109_47#_M1002_g N_VPWR_c_590_n 0.00588483f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_109_47#_M1005_g N_VPWR_c_590_n 0.0104367f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A_109_47#_M1026_g N_VPWR_c_590_n 0.0117628f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_109_47#_c_503_p N_VPWR_c_590_n 0.00955092f $X=0.68 $Y=2.3 $X2=0 $Y2=0
cc_355 N_A_109_47#_c_440_n N_VPWR_c_590_n 0.0110499f $X=1.825 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_109_47#_c_456_n N_VPWR_c_590_n 0.0145632f $X=4.015 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_109_47#_c_472_n N_VPWR_c_590_n 0.00815405f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_109_47#_c_449_n N_VPWR_c_590_n 9.70401e-19 $X=0.705 $Y=1.87 $X2=0
+ $Y2=0
cc_359 N_A_109_47#_c_456_n N_VPWR_c_606_n 0.0531577f $X=4.015 $Y=1.87 $X2=0
+ $Y2=0
cc_360 N_A_109_47#_c_440_n N_A_277_297#_M1001_d 0.00323299f $X=1.825 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_361 N_A_109_47#_c_456_n N_A_277_297#_M1025_d 0.00328736f $X=4.015 $Y=1.87
+ $X2=0 $Y2=0
cc_362 N_A_109_47#_M1022_s N_A_277_297#_c_701_n 0.00312348f $X=1.805 $Y=1.485
+ $X2=0 $Y2=0
cc_363 N_A_109_47#_c_440_n N_A_277_297#_c_701_n 0.00506389f $X=1.825 $Y=1.87
+ $X2=0 $Y2=0
cc_364 N_A_109_47#_c_456_n N_A_277_297#_c_701_n 0.00506389f $X=4.015 $Y=1.87
+ $X2=0 $Y2=0
cc_365 N_A_109_47#_c_462_n N_A_277_297#_c_701_n 0.0112811f $X=1.95 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_109_47#_c_440_n N_A_277_297#_c_709_n 0.0115714f $X=1.825 $Y=1.87
+ $X2=0 $Y2=0
cc_367 N_A_109_47#_c_456_n N_A_277_297#_c_710_n 0.0116461f $X=4.015 $Y=1.87
+ $X2=0 $Y2=0
cc_368 N_A_109_47#_c_456_n N_A_717_297#_M1009_s 0.00328796f $X=4.015 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_369 N_A_109_47#_c_472_n N_A_717_297#_M1015_d 0.00325314f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_370 N_A_109_47#_M1012_s N_A_717_297#_c_721_n 0.00312348f $X=4.005 $Y=1.485
+ $X2=0 $Y2=0
cc_371 N_A_109_47#_c_456_n N_A_717_297#_c_721_n 0.00506389f $X=4.015 $Y=1.87
+ $X2=0 $Y2=0
cc_372 N_A_109_47#_c_472_n N_A_717_297#_c_721_n 0.00506389f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_373 N_A_109_47#_c_480_n N_A_717_297#_c_721_n 0.0112811f $X=4.14 $Y=1.87 $X2=0
+ $Y2=0
cc_374 N_A_109_47#_c_456_n N_A_717_297#_c_729_n 0.0116461f $X=4.015 $Y=1.87
+ $X2=0 $Y2=0
cc_375 N_A_109_47#_c_472_n N_A_717_297#_c_730_n 0.0116461f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_376 N_A_109_47#_c_435_n N_X_M1000_d 0.00205826f $X=5.29 $Y=1.53 $X2=0 $Y2=0
cc_377 N_A_109_47#_c_422_n N_X_c_749_n 0.00513121f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A_109_47#_c_423_n N_X_c_749_n 0.00630972f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A_109_47#_c_424_n N_X_c_749_n 5.22228e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_109_47#_M1002_g N_X_c_752_n 0.010803f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A_109_47#_c_540_p N_X_c_752_n 0.00496418f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_382 N_A_109_47#_c_540_p N_X_c_754_n 0.0041562f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_109_47#_c_435_n N_X_c_754_n 0.004312f $X=5.29 $Y=1.53 $X2=0 $Y2=0
cc_384 N_A_109_47#_c_427_n N_X_c_754_n 0.00139251f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A_109_47#_c_423_n N_X_c_739_n 0.00870364f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A_109_47#_c_424_n N_X_c_739_n 0.00870364f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A_109_47#_c_540_p N_X_c_739_n 0.036111f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_388 N_A_109_47#_c_427_n N_X_c_739_n 0.00222133f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_109_47#_c_422_n N_X_c_740_n 0.0025255f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_390 N_A_109_47#_c_423_n N_X_c_740_n 0.00113286f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_391 N_A_109_47#_c_479_n N_X_c_740_n 0.0117845f $X=5.375 $Y=1.175 $X2=0 $Y2=0
cc_392 N_A_109_47#_c_540_p N_X_c_740_n 0.0152659f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_393 N_A_109_47#_c_427_n N_X_c_740_n 0.00230301f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_394 N_A_109_47#_M1005_g N_X_c_743_n 0.0129283f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_395 N_A_109_47#_c_540_p N_X_c_743_n 0.0149264f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_396 N_A_109_47#_M1002_g N_X_c_744_n 0.00102397f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A_109_47#_c_540_p N_X_c_744_n 0.0135282f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_398 N_A_109_47#_c_435_n N_X_c_744_n 0.00517831f $X=5.29 $Y=1.53 $X2=0 $Y2=0
cc_399 N_A_109_47#_c_427_n N_X_c_744_n 0.00220442f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_400 N_A_109_47#_c_424_n N_X_c_741_n 0.00113286f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_109_47#_c_425_n N_X_c_741_n 0.0132219f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_109_47#_c_540_p N_X_c_741_n 0.0265405f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_403 N_A_109_47#_c_427_n N_X_c_741_n 0.00230339f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_404 N_A_109_47#_c_423_n N_X_c_776_n 5.22228e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A_109_47#_c_424_n N_X_c_776_n 0.00630972f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A_109_47#_c_425_n N_X_c_776_n 0.0106039f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A_109_47#_M1026_g N_X_c_745_n 0.0164003f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A_109_47#_c_540_p N_X_c_745_n 0.00274549f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_409 N_A_109_47#_c_540_p N_X_c_746_n 0.0203891f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_410 N_A_109_47#_c_427_n N_X_c_746_n 0.00222737f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_411 N_A_109_47#_c_425_n X 0.0216562f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_412 N_A_109_47#_c_540_p X 0.0166688f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_413 N_A_109_47#_c_426_n N_A_27_47#_c_815_n 0.00107689f $X=0.705 $Y=1.445
+ $X2=0 $Y2=0
cc_414 N_A_109_47#_M1013_s N_A_27_47#_c_821_n 0.00304656f $X=0.545 $Y=0.235
+ $X2=0 $Y2=0
cc_415 N_A_109_47#_c_441_n N_A_27_47#_c_821_n 0.0161979f $X=0.68 $Y=0.73 $X2=0
+ $Y2=0
cc_416 N_A_109_47#_c_441_n N_A_27_47#_c_816_n 0.0103589f $X=0.68 $Y=0.73 $X2=0
+ $Y2=0
cc_417 N_A_109_47#_c_422_n N_VGND_c_924_n 0.00159991f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A_109_47#_c_435_n N_VGND_c_924_n 0.00109643f $X=5.29 $Y=1.53 $X2=0
+ $Y2=0
cc_419 N_A_109_47#_c_422_n N_VGND_c_925_n 0.00541359f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A_109_47#_c_423_n N_VGND_c_925_n 0.00423334f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_A_109_47#_c_423_n N_VGND_c_926_n 0.00146448f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_422 N_A_109_47#_c_424_n N_VGND_c_926_n 0.00146448f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_423 N_A_109_47#_c_425_n N_VGND_c_927_n 0.00321527f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_424 N_A_109_47#_c_424_n N_VGND_c_934_n 0.00423334f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_A_109_47#_c_425_n N_VGND_c_934_n 0.00424308f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_426 N_A_109_47#_M1013_s N_VGND_c_936_n 0.00216833f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_427 N_A_109_47#_c_422_n N_VGND_c_936_n 0.00952874f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A_109_47#_c_423_n N_VGND_c_936_n 0.0057163f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_A_109_47#_c_424_n N_VGND_c_936_n 0.0057163f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A_109_47#_c_425_n N_VGND_c_936_n 0.00706016f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_590_n N_A_277_297#_M1001_d 0.00226339f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_432 N_VPWR_c_590_n N_A_277_297#_M1025_d 0.002144f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_433 N_VPWR_c_590_n N_A_277_297#_c_701_n 0.020508f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_434 N_VPWR_c_605_n N_A_277_297#_c_701_n 0.0330174f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_590_n N_A_277_297#_c_709_n 0.00938288f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_605_n N_A_277_297#_c_709_n 0.0136719f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_590_n N_A_277_297#_c_710_n 0.00938745f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_605_n N_A_277_297#_c_710_n 0.0137033f $X=2.665 $Y=2.465 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_590_n N_A_717_297#_M1009_s 0.00219968f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_440 N_VPWR_c_590_n N_A_717_297#_M1015_d 0.00219968f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_598_n N_A_717_297#_c_721_n 0.0330174f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_590_n N_A_717_297#_c_721_n 0.0204707f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_598_n N_A_717_297#_c_729_n 0.0137033f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_590_n N_A_717_297#_c_729_n 0.00938745f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_598_n N_A_717_297#_c_730_n 0.0137033f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_590_n N_A_717_297#_c_730_n 0.00938745f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_590_n N_X_M1000_d 0.00392989f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_448 N_VPWR_c_590_n N_X_M1005_d 0.00284632f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_449 N_VPWR_c_595_n N_X_c_787_n 0.012815f $X=5.695 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_590_n N_X_c_787_n 0.00801045f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_451 N_VPWR_M1002_s N_X_c_752_n 0.00197151f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_452 N_VPWR_c_596_n N_X_c_752_n 0.0133483f $X=5.82 $Y=2.3 $X2=0 $Y2=0
cc_453 N_VPWR_c_590_n N_X_c_752_n 0.00580743f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_M1002_s N_X_c_744_n 2.21014e-19 $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_455 N_VPWR_c_601_n N_X_c_793_n 0.0142343f $X=6.535 $Y=2.72 $X2=0 $Y2=0
cc_456 N_VPWR_c_590_n N_X_c_793_n 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_457 N_VPWR_M1026_s X 0.00286582f $X=6.525 $Y=1.485 $X2=0 $Y2=0
cc_458 N_VPWR_c_597_n X 0.0174458f $X=6.66 $Y=1.96 $X2=0 $Y2=0
cc_459 N_X_c_739_n N_VGND_M1010_s 0.00162089f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_460 N_X_c_741_n N_VGND_M1017_s 0.00285873f $X=6.24 $Y=0.725 $X2=0 $Y2=0
cc_461 N_X_c_740_n N_VGND_c_924_n 0.00830019f $X=5.565 $Y=0.815 $X2=0 $Y2=0
cc_462 N_X_c_749_n N_VGND_c_925_n 0.0188551f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_463 N_X_c_739_n N_VGND_c_925_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_464 N_X_c_739_n N_VGND_c_926_n 0.0122559f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_465 N_X_c_741_n N_VGND_c_927_n 0.0215642f $X=6.24 $Y=0.725 $X2=0 $Y2=0
cc_466 N_X_c_739_n N_VGND_c_934_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_467 N_X_c_741_n N_VGND_c_934_n 0.00194867f $X=6.24 $Y=0.725 $X2=0 $Y2=0
cc_468 N_X_c_776_n N_VGND_c_934_n 0.0188551f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_469 N_X_c_741_n N_VGND_c_935_n 0.00149652f $X=6.24 $Y=0.725 $X2=0 $Y2=0
cc_470 N_X_M1006_d N_VGND_c_936_n 0.00215201f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_471 N_X_M1011_d N_VGND_c_936_n 0.00215201f $X=6.105 $Y=0.235 $X2=0 $Y2=0
cc_472 N_X_c_749_n N_VGND_c_936_n 0.0122069f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_473 N_X_c_739_n N_VGND_c_936_n 0.00835832f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_474 N_X_c_741_n N_VGND_c_936_n 0.00746305f $X=6.24 $Y=0.725 $X2=0 $Y2=0
cc_475 N_X_c_776_n N_VGND_c_936_n 0.0122069f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_817_n N_A_277_47#_M1018_d 0.00312026f $X=2.78 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_477 N_A_27_47#_c_817_n N_A_277_47#_M1024_s 0.00315249f $X=2.78 $Y=0.38 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_M1016_d N_A_277_47#_c_856_n 0.00162317f $X=1.805 $Y=0.235
+ $X2=0 $Y2=0
cc_479 N_A_27_47#_c_816_n N_A_277_47#_c_856_n 0.0115481f $X=1.1 $Y=0.73 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_817_n N_A_277_47#_c_856_n 0.0588671f $X=2.78 $Y=0.38 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_M1020_s N_A_277_47#_c_857_n 0.00319828f $X=2.645 $Y=0.235
+ $X2=0 $Y2=0
cc_482 N_A_27_47#_c_817_n N_A_277_47#_c_857_n 0.018919f $X=2.78 $Y=0.38 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_817_n N_VGND_c_922_n 0.017428f $X=2.78 $Y=0.38 $X2=0 $Y2=0
cc_484 N_A_27_47#_c_814_n N_VGND_c_928_n 0.0180288f $X=0.215 $Y=0.475 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_821_n N_VGND_c_928_n 0.0363282f $X=1.015 $Y=0.365 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_817_n N_VGND_c_928_n 0.0998324f $X=2.78 $Y=0.38 $X2=0 $Y2=0
cc_487 N_A_27_47#_c_847_p N_VGND_c_928_n 0.0114305f $X=1.1 $Y=0.39 $X2=0 $Y2=0
cc_488 N_A_27_47#_M1013_d N_VGND_c_936_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_M1027_d N_VGND_c_936_n 0.0021521f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_M1016_d N_VGND_c_936_n 0.00215227f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_M1020_s N_VGND_c_936_n 0.00209344f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_814_n N_VGND_c_936_n 0.00999725f $X=0.215 $Y=0.475 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_c_821_n N_VGND_c_936_n 0.023578f $X=1.015 $Y=0.365 $X2=0 $Y2=0
cc_494 N_A_27_47#_c_817_n N_VGND_c_936_n 0.0632734f $X=2.78 $Y=0.38 $X2=0 $Y2=0
cc_495 N_A_27_47#_c_847_p N_VGND_c_936_n 0.00653933f $X=1.1 $Y=0.39 $X2=0 $Y2=0
cc_496 N_A_277_47#_c_857_n N_VGND_M1008_s 0.00285834f $X=3.555 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_497 N_A_277_47#_c_858_n N_VGND_M1007_d 0.00162089f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_498 N_A_277_47#_c_857_n N_VGND_c_922_n 0.018331f $X=3.555 $Y=0.81 $X2=0 $Y2=0
cc_499 N_A_277_47#_c_858_n N_VGND_c_923_n 0.0122559f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_500 N_A_277_47#_c_858_n N_VGND_c_924_n 0.00830019f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_501 N_A_277_47#_c_857_n N_VGND_c_928_n 0.00296885f $X=3.555 $Y=0.81 $X2=0
+ $Y2=0
cc_502 N_A_277_47#_c_857_n N_VGND_c_930_n 0.00203746f $X=3.555 $Y=0.81 $X2=0
+ $Y2=0
cc_503 N_A_277_47#_c_877_n N_VGND_c_930_n 0.0188551f $X=3.72 $Y=0.42 $X2=0 $Y2=0
cc_504 N_A_277_47#_c_858_n N_VGND_c_930_n 0.00198695f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_505 N_A_277_47#_c_858_n N_VGND_c_932_n 0.00198695f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_506 N_A_277_47#_c_882_n N_VGND_c_932_n 0.0188551f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_507 N_A_277_47#_M1018_d N_VGND_c_936_n 0.00216833f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_277_47#_M1024_s N_VGND_c_936_n 0.00216833f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_277_47#_M1008_d N_VGND_c_936_n 0.00215201f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_510 N_A_277_47#_M1014_s N_VGND_c_936_n 0.00215201f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_277_47#_c_857_n N_VGND_c_936_n 0.0109066f $X=3.555 $Y=0.81 $X2=0
+ $Y2=0
cc_512 N_A_277_47#_c_877_n N_VGND_c_936_n 0.0122069f $X=3.72 $Y=0.42 $X2=0 $Y2=0
cc_513 N_A_277_47#_c_858_n N_VGND_c_936_n 0.00835832f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_514 N_A_277_47#_c_882_n N_VGND_c_936_n 0.0122069f $X=4.56 $Y=0.39 $X2=0 $Y2=0

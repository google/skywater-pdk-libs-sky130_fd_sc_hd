* File: sky130_fd_sc_hd__a21o_2.pxi.spice
* Created: Tue Sep  1 18:52:07 2020
* 
x_PM_SKY130_FD_SC_HD__A21O_2%A_80_199# N_A_80_199#_M1001_d N_A_80_199#_M1002_s
+ N_A_80_199#_M1004_g N_A_80_199#_c_54_n N_A_80_199#_M1003_g N_A_80_199#_M1009_g
+ N_A_80_199#_c_55_n N_A_80_199#_M1007_g N_A_80_199#_c_56_n N_A_80_199#_c_66_p
+ N_A_80_199#_c_105_p N_A_80_199#_c_63_n N_A_80_199#_c_80_p N_A_80_199#_c_57_n
+ N_A_80_199#_c_58_n N_A_80_199#_c_59_n PM_SKY130_FD_SC_HD__A21O_2%A_80_199#
x_PM_SKY130_FD_SC_HD__A21O_2%B1 N_B1_c_125_n N_B1_M1001_g N_B1_M1002_g B1
+ N_B1_c_127_n PM_SKY130_FD_SC_HD__A21O_2%B1
x_PM_SKY130_FD_SC_HD__A21O_2%A1 N_A1_M1006_g N_A1_M1000_g A1 A1 N_A1_c_161_n
+ N_A1_c_162_n PM_SKY130_FD_SC_HD__A21O_2%A1
x_PM_SKY130_FD_SC_HD__A21O_2%A2 N_A2_c_199_n N_A2_M1005_g N_A2_M1008_g A2
+ N_A2_c_201_n A2 PM_SKY130_FD_SC_HD__A21O_2%A2
x_PM_SKY130_FD_SC_HD__A21O_2%VPWR N_VPWR_M1004_s N_VPWR_M1009_s N_VPWR_M1000_d
+ N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n VPWR
+ N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_227_n N_VPWR_c_236_n
+ N_VPWR_c_237_n PM_SKY130_FD_SC_HD__A21O_2%VPWR
x_PM_SKY130_FD_SC_HD__A21O_2%X N_X_M1003_d N_X_M1004_d N_X_c_287_p N_X_c_275_n X
+ N_X_c_273_n PM_SKY130_FD_SC_HD__A21O_2%X
x_PM_SKY130_FD_SC_HD__A21O_2%A_386_297# N_A_386_297#_M1002_d
+ N_A_386_297#_M1008_d N_A_386_297#_c_292_n N_A_386_297#_c_302_n
+ N_A_386_297#_c_293_n N_A_386_297#_c_298_n N_A_386_297#_c_307_n
+ PM_SKY130_FD_SC_HD__A21O_2%A_386_297#
x_PM_SKY130_FD_SC_HD__A21O_2%VGND N_VGND_M1003_s N_VGND_M1007_s N_VGND_M1005_d
+ N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n
+ N_VGND_c_314_n VGND N_VGND_c_315_n N_VGND_c_316_n N_VGND_c_317_n
+ PM_SKY130_FD_SC_HD__A21O_2%VGND
cc_1 VNB N_A_80_199#_M1004_g 0.0127435f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_2 VNB N_A_80_199#_c_54_n 0.0186908f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.995
cc_3 VNB N_A_80_199#_c_55_n 0.0160705f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=0.995
cc_4 VNB N_A_80_199#_c_56_n 8.53597e-19 $X=-0.19 $Y=-0.24 $X2=1.125 $Y2=1.69
cc_5 VNB N_A_80_199#_c_57_n 0.00103783f $X=-0.19 $Y=-0.24 $X2=1.085 $Y2=1.16
cc_6 VNB N_A_80_199#_c_58_n 0.00106484f $X=-0.19 $Y=-0.24 $X2=1.125 $Y2=0.995
cc_7 VNB N_A_80_199#_c_59_n 0.04927f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=1.235
cc_8 VNB N_B1_c_125_n 0.0188897f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=0.235
cc_9 VNB B1 0.00214757f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_10 VNB N_B1_c_127_n 0.0324598f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_11 VNB A1 0.00253827f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_12 VNB N_A1_c_161_n 0.0237277f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.56
cc_13 VNB N_A1_c_162_n 0.0186174f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_14 VNB N_A2_c_199_n 0.0208749f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=0.235
cc_15 VNB A2 0.0210285f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_16 VNB N_A2_c_201_n 0.0326999f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.995
cc_17 VNB N_VPWR_c_227_n 0.136896f $X=-0.19 $Y=-0.24 $X2=1.125 $Y2=1.805
cc_18 VNB N_X_c_273_n 0.00717477f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=0.56
cc_19 VNB N_VGND_c_309_n 0.0157553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_310_n 0.0130853f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.56
cc_21 VNB N_VGND_c_311_n 0.0121717f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.325
cc_22 VNB N_VGND_c_312_n 0.00274225f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=0.995
cc_23 VNB N_VGND_c_313_n 0.0100784f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=0.56
cc_24 VNB N_VGND_c_314_n 0.0164267f $X=-0.19 $Y=-0.24 $X2=1.125 $Y2=1.69
cc_25 VNB N_VGND_c_315_n 0.0362654f $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=0.74
cc_26 VNB N_VGND_c_316_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_317_n 0.186751f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.145
cc_28 VPB N_A_80_199#_M1004_g 0.0277363f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_29 VPB N_A_80_199#_M1009_g 0.0222235f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_30 VPB N_A_80_199#_c_56_n 0.00504085f $X=-0.19 $Y=1.305 $X2=1.125 $Y2=1.69
cc_31 VPB N_A_80_199#_c_63_n 0.0199736f $X=-0.19 $Y=1.305 $X2=1.632 $Y2=1.92
cc_32 VPB N_A_80_199#_c_59_n 0.00917678f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.235
cc_33 VPB N_B1_M1002_g 0.0234421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB B1 0.00427864f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_35 VPB N_B1_c_127_n 0.00978479f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_36 VPB N_A1_M1000_g 0.0195292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A1 0.0033439f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_38 VPB N_A1_c_161_n 0.00613722f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.56
cc_39 VPB N_A2_M1008_g 0.0279144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB A2 0.0058057f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_41 VPB N_A2_c_201_n 0.0067203f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.995
cc_42 VPB N_VPWR_c_228_n 0.0107835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_229_n 0.0374919f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.56
cc_44 VPB N_VPWR_c_230_n 0.00570708f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_45 VPB N_VPWR_c_231_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.075 $Y2=0.56
cc_46 VPB N_VPWR_c_232_n 0.0148832f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=0.995
cc_47 VPB N_VPWR_c_233_n 0.0277741f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.655
cc_48 VPB N_VPWR_c_234_n 0.0160704f $X=-0.19 $Y=1.305 $X2=1.125 $Y2=0.995
cc_49 VPB N_VPWR_c_227_n 0.0478266f $X=-0.19 $Y=1.305 $X2=1.125 $Y2=1.805
cc_50 VPB N_VPWR_c_236_n 0.00510335f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=0.995
cc_51 VPB N_VPWR_c_237_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.085 $Y2=1.235
cc_52 VPB N_X_c_273_n 0.00401505f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=0.56
cc_53 N_A_80_199#_c_55_n N_B1_c_125_n 0.0240752f $X=1.075 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A_80_199#_c_66_p N_B1_c_125_n 0.0124518f $X=1.675 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_55 N_A_80_199#_c_58_n N_B1_c_125_n 0.00174875f $X=1.125 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_56 N_A_80_199#_c_56_n N_B1_M1002_g 0.00757775f $X=1.125 $Y=1.69 $X2=0 $Y2=0
cc_57 N_A_80_199#_c_63_n N_B1_M1002_g 0.0078995f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_58 N_A_80_199#_M1009_g B1 3.17505e-19 $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_80_199#_c_66_p B1 0.0219068f $X=1.675 $Y=0.74 $X2=0 $Y2=0
cc_60 N_A_80_199#_c_63_n B1 0.0169449f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_61 N_A_80_199#_c_57_n B1 0.0345371f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_80_199#_c_59_n B1 9.95833e-19 $X=1.075 $Y=1.235 $X2=0 $Y2=0
cc_63 N_A_80_199#_c_66_p N_B1_c_127_n 0.0061727f $X=1.675 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A_80_199#_c_63_n N_B1_c_127_n 0.00144331f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_65 N_A_80_199#_c_57_n N_B1_c_127_n 0.00279422f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_80_199#_c_59_n N_B1_c_127_n 0.0182216f $X=1.075 $Y=1.235 $X2=0 $Y2=0
cc_67 N_A_80_199#_c_66_p A1 0.00771051f $X=1.675 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A_80_199#_c_80_p A1 0.0118486f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_69 N_A_80_199#_c_66_p N_A1_c_162_n 0.0016367f $X=1.675 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A_80_199#_c_80_p N_A1_c_162_n 0.00464407f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_71 N_A_80_199#_c_56_n N_VPWR_M1009_s 0.00148542f $X=1.125 $Y=1.69 $X2=0 $Y2=0
cc_72 N_A_80_199#_c_63_n N_VPWR_M1009_s 0.00444135f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_73 N_A_80_199#_M1004_g N_VPWR_c_229_n 0.00544127f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_74 N_A_80_199#_M1004_g N_VPWR_c_230_n 5.30039e-19 $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_75 N_A_80_199#_M1009_g N_VPWR_c_230_n 0.00808779f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_76 N_A_80_199#_c_63_n N_VPWR_c_230_n 0.0320786f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_77 N_A_80_199#_M1004_g N_VPWR_c_232_n 0.00585385f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_78 N_A_80_199#_M1009_g N_VPWR_c_232_n 0.00486043f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_79 N_A_80_199#_c_63_n N_VPWR_c_233_n 0.0197373f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_80 N_A_80_199#_M1002_s N_VPWR_c_227_n 0.00213418f $X=1.515 $Y=1.485 $X2=0
+ $Y2=0
cc_81 N_A_80_199#_M1004_g N_VPWR_c_227_n 0.0114347f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_82 N_A_80_199#_M1009_g N_VPWR_c_227_n 0.00822531f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_83 N_A_80_199#_c_63_n N_VPWR_c_227_n 0.0204043f $X=1.632 $Y=1.92 $X2=0 $Y2=0
cc_84 N_A_80_199#_c_54_n N_X_c_275_n 0.0107114f $X=0.645 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_80_199#_c_59_n N_X_c_275_n 0.00419569f $X=1.075 $Y=1.235 $X2=0 $Y2=0
cc_86 N_A_80_199#_M1004_g N_X_c_273_n 0.0102098f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_80_199#_c_54_n N_X_c_273_n 0.00609067f $X=0.645 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_80_199#_c_55_n N_X_c_273_n 0.00120127f $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_80_199#_c_57_n N_X_c_273_n 0.0448011f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_80_199#_c_58_n N_X_c_273_n 0.00731474f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_80_199#_c_59_n N_X_c_273_n 0.0177218f $X=1.075 $Y=1.235 $X2=0 $Y2=0
cc_92 N_A_80_199#_c_66_p N_VGND_M1007_s 0.00676206f $X=1.675 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_80_199#_c_105_p N_VGND_M1007_s 0.00102707f $X=1.295 $Y=0.74 $X2=0
+ $Y2=0
cc_94 N_A_80_199#_c_58_n N_VGND_M1007_s 6.96297e-19 $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_95 N_A_80_199#_c_54_n N_VGND_c_310_n 0.00752096f $X=0.645 $Y=0.995 $X2=0
+ $Y2=0
cc_96 N_A_80_199#_c_55_n N_VGND_c_310_n 5.0423e-19 $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_80_199#_c_59_n N_VGND_c_310_n 0.00435458f $X=1.075 $Y=1.235 $X2=0
+ $Y2=0
cc_98 N_A_80_199#_c_54_n N_VGND_c_311_n 0.00353537f $X=0.645 $Y=0.995 $X2=0
+ $Y2=0
cc_99 N_A_80_199#_c_55_n N_VGND_c_311_n 0.00486043f $X=1.075 $Y=0.995 $X2=0
+ $Y2=0
cc_100 N_A_80_199#_c_54_n N_VGND_c_312_n 4.98572e-19 $X=0.645 $Y=0.995 $X2=0
+ $Y2=0
cc_101 N_A_80_199#_c_55_n N_VGND_c_312_n 0.00627405f $X=1.075 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_A_80_199#_c_66_p N_VGND_c_312_n 0.00874168f $X=1.675 $Y=0.74 $X2=0
+ $Y2=0
cc_103 N_A_80_199#_c_105_p N_VGND_c_312_n 0.00767611f $X=1.295 $Y=0.74 $X2=0
+ $Y2=0
cc_104 N_A_80_199#_c_59_n N_VGND_c_312_n 2.83666e-19 $X=1.075 $Y=1.235 $X2=0
+ $Y2=0
cc_105 N_A_80_199#_c_66_p N_VGND_c_315_n 0.00298484f $X=1.675 $Y=0.74 $X2=0
+ $Y2=0
cc_106 N_A_80_199#_c_80_p N_VGND_c_315_n 0.0123384f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_107 N_A_80_199#_M1001_d N_VGND_c_317_n 0.0137378f $X=1.64 $Y=0.235 $X2=0
+ $Y2=0
cc_108 N_A_80_199#_c_54_n N_VGND_c_317_n 0.00411309f $X=0.645 $Y=0.995 $X2=0
+ $Y2=0
cc_109 N_A_80_199#_c_55_n N_VGND_c_317_n 0.00822531f $X=1.075 $Y=0.995 $X2=0
+ $Y2=0
cc_110 N_A_80_199#_c_66_p N_VGND_c_317_n 0.00608171f $X=1.675 $Y=0.74 $X2=0
+ $Y2=0
cc_111 N_A_80_199#_c_105_p N_VGND_c_317_n 9.01125e-19 $X=1.295 $Y=0.74 $X2=0
+ $Y2=0
cc_112 N_A_80_199#_c_80_p N_VGND_c_317_n 0.00720706f $X=1.78 $Y=0.42 $X2=0 $Y2=0
cc_113 N_B1_M1002_g N_A1_M1000_g 0.0249266f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_114 B1 N_A1_M1000_g 3.94403e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B1_c_125_n A1 0.00101821f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_116 B1 A1 0.0113526f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_117 N_B1_c_127_n A1 0.00112471f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_118 B1 N_A1_c_161_n 9.77307e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B1_c_127_n N_A1_c_161_n 0.0214253f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_c_125_n N_A1_c_162_n 0.0142151f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_M1002_g N_VPWR_c_230_n 0.00233012f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1002_g N_VPWR_c_231_n 0.00112519f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_VPWR_c_233_n 0.00571722f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_M1002_g N_VPWR_c_227_n 0.0116957f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_125 N_B1_c_125_n N_VGND_c_312_n 0.00415575f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_c_125_n N_VGND_c_315_n 0.00428022f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_c_125_n N_VGND_c_317_n 0.0064108f $X=1.565 $Y=0.995 $X2=0 $Y2=0
cc_128 A1 N_A2_c_199_n 0.00496506f $X=2.45 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_129 N_A1_c_161_n N_A2_c_199_n 0.00863958f $X=2.325 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A1_c_162_n N_A2_c_199_n 0.0253589f $X=2.3 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_131 N_A1_M1000_g N_A2_M1008_g 0.038657f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_132 A1 A2 0.0368368f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_133 N_A1_c_161_n A2 2.52625e-19 $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_134 A1 N_A2_c_201_n 0.00148306f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_135 N_A1_c_161_n N_A2_c_201_n 0.0114029f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A1_M1000_g N_VPWR_c_231_n 0.0078334f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A1_M1000_g N_VPWR_c_233_n 0.00564095f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_M1000_g N_VPWR_c_227_n 0.00506784f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_c_161_n N_A_386_297#_c_292_n 0.00116473f $X=2.325 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A1_M1000_g N_A_386_297#_c_293_n 0.0144238f $X=2.285 $Y=1.985 $X2=0
+ $Y2=0
cc_141 A1 N_A_386_297#_c_293_n 0.0168554f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_142 N_A1_c_161_n N_A_386_297#_c_293_n 4.4906e-19 $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A1_c_162_n N_VGND_c_314_n 0.00160183f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_144 A1 N_VGND_c_315_n 0.0141846f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_145 N_A1_c_162_n N_VGND_c_315_n 0.00518168f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_146 A1 N_VGND_c_317_n 0.0134696f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_147 N_A1_c_162_n N_VGND_c_317_n 0.00982019f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_148 A1 A_458_47# 0.00681103f $X=2.45 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_149 N_A2_M1008_g N_VPWR_c_231_n 0.00887135f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A2_M1008_g N_VPWR_c_234_n 0.00544582f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_M1008_g N_VPWR_c_227_n 0.00581532f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A2_M1008_g N_A_386_297#_c_293_n 0.0171702f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_153 A2 N_A_386_297#_c_293_n 0.00146795f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_154 A2 N_A_386_297#_c_298_n 0.0112544f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A2_c_201_n N_A_386_297#_c_298_n 0.00132222f $X=2.75 $Y=1.155 $X2=0
+ $Y2=0
cc_156 A2 N_VGND_M1005_d 0.00271578f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A2_c_199_n N_VGND_c_314_n 0.010182f $X=2.745 $Y=1.005 $X2=0 $Y2=0
cc_158 A2 N_VGND_c_314_n 0.0205543f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A2_c_201_n N_VGND_c_314_n 9.25957e-19 $X=2.75 $Y=1.155 $X2=0 $Y2=0
cc_160 N_A2_c_199_n N_VGND_c_315_n 0.00525069f $X=2.745 $Y=1.005 $X2=0 $Y2=0
cc_161 N_A2_c_199_n N_VGND_c_317_n 0.00917341f $X=2.745 $Y=1.005 $X2=0 $Y2=0
cc_162 A2 N_VGND_c_317_n 0.00133614f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_163 N_VPWR_c_227_n N_X_M1004_d 0.00396809f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_164 N_VPWR_c_232_n N_X_c_273_n 0.0138731f $X=0.955 $Y=2.72 $X2=0 $Y2=0
cc_165 N_VPWR_c_227_n N_X_c_273_n 0.00878068f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_c_227_n N_A_386_297#_M1002_d 0.00340659f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_167 N_VPWR_c_227_n N_A_386_297#_M1008_d 0.00263722f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_233_n N_A_386_297#_c_302_n 0.0136957f $X=2.355 $Y=2.72 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_227_n N_A_386_297#_c_302_n 0.00858812f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_170 N_VPWR_M1000_d N_A_386_297#_c_293_n 0.00513134f $X=2.36 $Y=1.485 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_231_n N_A_386_297#_c_293_n 0.0158408f $X=2.52 $Y=2.34 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_227_n N_A_386_297#_c_293_n 0.011765f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_173 N_VPWR_c_234_n N_A_386_297#_c_307_n 0.0144241f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_227_n N_A_386_297#_c_307_n 0.00839556f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_175 N_X_c_275_n N_VGND_c_310_n 0.00168574f $X=0.86 $Y=0.73 $X2=0 $Y2=0
cc_176 N_X_c_287_p N_VGND_c_311_n 0.0119756f $X=0.86 $Y=0.42 $X2=0 $Y2=0
cc_177 N_X_c_275_n N_VGND_c_311_n 0.00250975f $X=0.86 $Y=0.73 $X2=0 $Y2=0
cc_178 N_X_M1003_d N_VGND_c_317_n 0.00391594f $X=0.72 $Y=0.235 $X2=0 $Y2=0
cc_179 N_X_c_287_p N_VGND_c_317_n 0.00713507f $X=0.86 $Y=0.42 $X2=0 $Y2=0
cc_180 N_X_c_275_n N_VGND_c_317_n 0.00442355f $X=0.86 $Y=0.73 $X2=0 $Y2=0
cc_181 N_VGND_c_317_n A_458_47# 0.0049739f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

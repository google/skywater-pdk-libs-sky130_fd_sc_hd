# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__and2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.625000 3.155000 0.995000 ;
        RECT 2.900000 0.995000 3.205000 1.325000 ;
        RECT 2.900000 1.325000 3.155000 1.745000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 0.975000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.535000 2.730000 1.745000 ;
        RECT 1.525000 0.495000 1.715000 0.615000 ;
        RECT 1.525000 0.615000 2.730000 0.825000 ;
        RECT 2.440000 0.825000 2.730000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.955000  0.085000 1.285000 0.445000 ;
        RECT 1.885000  0.085000 2.215000 0.445000 ;
        RECT 2.745000  0.085000 3.075000 0.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.090000 2.255000 0.425000 2.635000 ;
        RECT 0.990000 2.275000 1.320000 2.635000 ;
        RECT 1.905000 2.275000 2.235000 2.635000 ;
        RECT 2.745000 2.275000 3.075000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.425000 0.615000 ;
      RECT 0.090000 0.615000 1.355000 0.805000 ;
      RECT 0.165000 0.995000 0.425000 1.325000 ;
      RECT 0.165000 1.325000 0.335000 1.915000 ;
      RECT 0.165000 1.915000 3.505000 2.085000 ;
      RECT 0.515000 1.500000 1.315000 1.745000 ;
      RECT 1.110000 1.435000 1.320000 1.485000 ;
      RECT 1.110000 1.485000 1.315000 1.500000 ;
      RECT 1.145000 0.805000 1.355000 0.995000 ;
      RECT 1.145000 0.995000 2.260000 1.355000 ;
      RECT 1.145000 1.355000 1.320000 1.435000 ;
      RECT 3.330000 0.495000 3.500000 0.675000 ;
      RECT 3.330000 0.675000 3.545000 0.845000 ;
      RECT 3.335000 1.530000 3.545000 1.700000 ;
      RECT 3.335000 1.700000 3.505000 1.915000 ;
      RECT 3.375000 0.845000 3.545000 1.530000 ;
  END
END sky130_fd_sc_hd__and2b_4
END LIBRARY

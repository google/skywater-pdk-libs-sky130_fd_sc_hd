* File: sky130_fd_sc_hd__a311oi_1.pex.spice
* Created: Tue Sep  1 18:54:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A311OI_1%A3 3 6 7 10 12 13
r25 10 13 57.4123 $w=4.4e-07 $l=2.5e-07 $layer=POLY_cond $X=0.325 $Y=1.16
+ $X2=0.325 $Y2=1.41
r26 10 12 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.325 $Y=1.16
+ $X2=0.325 $Y2=0.995
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r28 6 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.41
r29 3 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%A2 3 6 8 9 10 15 16 17
c40 6 0 7.98776e-20 $X=0.895 $Y=1.985
r41 19 28 3.83364 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.697 $Y=0.995
+ $X2=0.697 $Y2=1.16
r42 16 28 6.74005 $w=3.28e-07 $l=1.93e-07 $layer=LI1_cond $X=0.89 $Y=1.16
+ $X2=0.697 $Y2=1.16
r43 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=1.325
r44 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r46 10 19 8.24709 $w=1.93e-07 $l=1.45e-07 $layer=LI1_cond $X=0.697 $Y=0.85
+ $X2=0.697 $Y2=0.995
r47 9 10 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=0.697 $Y=0.51
+ $X2=0.697 $Y2=0.85
r48 8 28 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.697
+ $Y2=1.16
r49 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.895 $Y=1.985
+ $X2=0.895 $Y2=1.325
r50 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.895 $Y=0.56
+ $X2=0.895 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%A1 3 6 9 13 14 16 19 24
c42 24 0 1.1931e-19 $X=1.28 $Y=0.462
r43 16 24 3.20933 $w=3.93e-07 $l=1.1e-07 $layer=LI1_cond $X=1.17 $Y=0.462
+ $X2=1.28 $Y2=0.462
r44 14 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.37 $Y2=1.325
r45 14 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.37 $Y2=0.995
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r47 10 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.28 $Y=1.16 $X2=1.37
+ $Y2=1.16
r48 9 10 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0.995
+ $X2=1.28 $Y2=1.16
r49 8 24 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.28 $Y=0.66 $X2=1.28
+ $Y2=0.462
r50 8 9 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.28 $Y=0.66 $X2=1.28
+ $Y2=0.995
r51 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.325 $Y=1.985
+ $X2=1.325 $Y2=1.325
r52 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.325 $Y=0.56
+ $X2=1.325 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%B1 3 7 10 11 16 18 21
c44 21 0 1.1931e-19 $X=1.85 $Y=0.995
r45 16 18 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=2.09 $Y=2.005
+ $X2=2.09 $Y2=2.21
r46 11 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=1.325
r47 11 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=0.995
r48 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.16 $X2=1.85 $Y2=1.16
r49 8 16 17.4845 $w=1.68e-07 $l=2.68e-07 $layer=LI1_cond $X=1.822 $Y=1.92
+ $X2=2.09 $Y2=1.92
r50 8 10 34.5733 $w=2.23e-07 $l=6.75e-07 $layer=LI1_cond $X=1.822 $Y=1.835
+ $X2=1.822 $Y2=1.16
r51 7 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.56 $X2=1.83
+ $Y2=0.995
r52 3 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.805 $Y=1.985
+ $X2=1.805 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%C1 3 5 7 8 14
c28 3 0 1.18506e-20 $X=2.3 $Y=1.985
r29 12 14 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.325 $Y=1.16
+ $X2=2.53 $Y2=1.16
r30 10 12 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.3 $Y=1.16
+ $X2=2.325 $Y2=1.16
r31 8 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.16 $X2=2.53 $Y2=1.16
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=0.995
+ $X2=2.325 $Y2=1.16
r33 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.325 $Y=0.995
+ $X2=2.325 $Y2=0.56
r34 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.325 $X2=2.3
+ $Y2=1.16
r35 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.3 $Y=1.325 $X2=2.3
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%VPWR 1 2 7 9 15 17 19 26 27 33
r41 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 27 34 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=1.15 $Y2=2.72
r43 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 24 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=2.72 $X2=1.07
+ $Y2=2.72
r45 24 26 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=1.2 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 20 30 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r49 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 19 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.94 $Y=2.72 $X2=1.07
+ $Y2=2.72
r51 19 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.94 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 17 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 13 33 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=2.635
+ $X2=1.07 $Y2=2.72
r55 13 15 24.6002 $w=2.58e-07 $l=5.55e-07 $layer=LI1_cond $X=1.07 $Y=2.635
+ $X2=1.07 $Y2=2.08
r56 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66 $X2=0.26
+ $Y2=2.34
r57 7 30 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r58 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r59 2 15 600 $w=1.7e-07 $l=6.59052e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.485 $X2=1.105 $Y2=2.08
r60 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r61 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%A_109_297# 1 2 9 11 12 14 17
c21 17 0 7.98776e-20 $X=1.535 $Y=2.26
c22 14 0 1.18506e-20 $X=1.455 $Y=2.175
r23 14 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=2.175
+ $X2=1.455 $Y2=2.26
r24 13 14 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.455 $Y=1.745
+ $X2=1.455 $Y2=2.175
r25 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.37 $Y=1.66
+ $X2=1.455 $Y2=1.745
r26 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.37 $Y=1.66 $X2=0.77
+ $Y2=1.66
r27 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.745
+ $X2=0.77 $Y2=1.66
r28 7 9 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.685 $Y=1.745
+ $X2=0.685 $Y2=1.8
r29 2 17 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=1.4
+ $Y=1.485 $X2=1.535 $Y2=2.26
r30 1 9 300 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.685 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%Y 1 2 3 12 14 15 17 20 25 27 28 29 38
r46 28 29 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=2.21
r47 28 38 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=2.53 $Y=1.87 $X2=2.53
+ $Y2=1.74
r48 25 38 3.60138 $w=2.38e-07 $l=7.5e-08 $layer=LI1_cond $X=2.53 $Y=1.665
+ $X2=2.53 $Y2=1.74
r49 22 25 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=1.58
+ $X2=2.53 $Y2=1.58
r50 20 27 6.82058 $w=2.43e-07 $l=1.45e-07 $layer=LI1_cond $X=2.527 $Y=0.655
+ $X2=2.527 $Y2=0.51
r51 18 20 21.9861 $w=1.68e-07 $l=3.37e-07 $layer=LI1_cond $X=2.19 $Y=0.74
+ $X2=2.527 $Y2=0.74
r52 17 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=1.495
+ $X2=2.19 $Y2=1.58
r53 16 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.825
+ $X2=2.19 $Y2=0.74
r54 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.19 $Y=0.825
+ $X2=2.19 $Y2=1.495
r55 14 18 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.74
+ $X2=2.19 $Y2=0.74
r56 14 15 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.105 $Y=0.74
+ $X2=1.705 $Y2=0.74
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=0.655
+ $X2=1.705 $Y2=0.74
r58 10 12 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.62 $Y=0.655
+ $X2=1.62 $Y2=0.42
r59 3 38 300 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_PDIFF $count=2 $X=2.375
+ $Y=1.485 $X2=2.51 $Y2=1.74
r60 2 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.235 $X2=2.535 $Y2=0.56
r61 1 12 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.235 $X2=1.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_1%VGND 1 2 7 9 13 15 17 27 28 34
r43 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r44 28 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r45 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r46 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.07
+ $Y2=0
r47 25 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.99
+ $Y2=0
r48 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r49 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r50 21 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r51 20 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r52 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 18 31 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r54 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r55 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.07
+ $Y2=0
r56 17 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.61
+ $Y2=0
r57 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r58 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r59 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0
r60 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0.4
r61 7 31 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r62 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r63 2 13 182 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.07 $Y2=0.4
r64 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o21ai_4.pex.spice
* Created: Thu Aug 27 14:35:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21AI_4%A1 1 3 6 8 10 13 15 17 20 24 28 31 35 36 38
+ 44 49 52 59
c110 35 0 1.98454e-19 $X=3.53 $Y=1.16
c111 24 0 1.2049e-19 $X=3.51 $Y=1.985
r112 48 59 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=1.35
+ $X2=1.475 $Y2=1.35
r113 47 49 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.31 $Y=1.16 $X2=1.36
+ $Y2=1.16
r114 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.31
+ $Y=1.16 $X2=1.31 $Y2=1.16
r115 45 47 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=1.31 $Y2=1.16
r116 43 45 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=0.63 $Y=1.16 $X2=0.93
+ $Y2=1.16
r117 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.16 $X2=0.63 $Y2=1.16
r118 40 43 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=0.5 $Y=1.16 $X2=0.63
+ $Y2=1.16
r119 38 48 2.85631 $w=6.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.15 $Y=1.35
+ $X2=1.31 $Y2=1.35
r120 38 44 9.283 $w=6.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.15 $Y=1.35 $X2=0.63
+ $Y2=1.35
r121 36 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.16
+ $X2=3.53 $Y2=1.325
r122 36 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.16
+ $X2=3.53 $Y2=0.995
r123 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.53
+ $Y=1.16 $X2=3.53 $Y2=1.16
r124 33 35 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=3.57 $Y=1.515
+ $X2=3.57 $Y2=1.16
r125 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.445 $Y=1.6
+ $X2=3.57 $Y2=1.515
r126 31 59 128.524 $w=1.68e-07 $l=1.97e-06 $layer=LI1_cond $X=3.445 $Y=1.6
+ $X2=1.475 $Y2=1.6
r127 28 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.55 $Y=0.56
+ $X2=3.55 $Y2=0.995
r128 24 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.985
+ $X2=3.51 $Y2=1.325
r129 18 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.16
r130 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.985
r131 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=1.16
r132 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=0.56
r133 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.16
r134 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.985
r135 8 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r136 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=0.56
r137 4 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.325
+ $X2=0.5 $Y2=1.16
r138 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.5 $Y=1.325 $X2=0.5
+ $Y2=1.985
r139 1 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=0.995
+ $X2=0.5 $Y2=1.16
r140 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.5 $Y=0.995 $X2=0.5
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 43 44
c71 43 0 1.2049e-19 $X=2.99 $Y=1.16
c72 22 0 9.53319e-20 $X=3.08 $Y=0.995
r73 42 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.99 $Y=1.16 $X2=3.08
+ $Y2=1.16
r74 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.16 $X2=2.99 $Y2=1.16
r75 40 42 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.65 $Y=1.16
+ $X2=2.99 $Y2=1.16
r76 39 43 16.7628 $w=2.73e-07 $l=4e-07 $layer=LI1_cond $X=2.59 $Y=1.207 $X2=2.99
+ $Y2=1.207
r77 38 40 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.65
+ $Y2=1.16
r78 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.16 $X2=2.59 $Y2=1.16
r79 36 38 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.22 $Y=1.16
+ $X2=2.59 $Y2=1.16
r80 35 39 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=1.207 $X2=2.59
+ $Y2=1.207
r81 34 36 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.16 $Y=1.16 $X2=2.22
+ $Y2=1.16
r82 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.16 $X2=2.16 $Y2=1.16
r83 31 34 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=2.16 $Y2=1.16
r84 29 35 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=1.207 $X2=2.16
+ $Y2=1.207
r85 25 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.325
+ $X2=3.08 $Y2=1.16
r86 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.08 $Y=1.325
+ $X2=3.08 $Y2=1.985
r87 22 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=1.16
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=0.56
r89 18 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.325
+ $X2=2.65 $Y2=1.16
r90 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.65 $Y=1.325
+ $X2=2.65 $Y2=1.985
r91 15 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=0.995
+ $X2=2.65 $Y2=1.16
r92 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.65 $Y=0.995
+ $X2=2.65 $Y2=0.56
r93 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.325
+ $X2=2.22 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.22 $Y=1.325
+ $X2=2.22 $Y2=1.985
r95 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=0.995
+ $X2=2.22 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.22 $Y=0.995
+ $X2=2.22 $Y2=0.56
r97 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.325
+ $X2=1.79 $Y2=1.16
r98 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.79 $Y=1.325 $X2=1.79
+ $Y2=1.985
r99 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=0.995
+ $X2=1.79 $Y2=1.16
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.79 $Y=0.995
+ $X2=1.79 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
c69 1 0 1.03122e-19 $X=3.98 $Y=0.995
r70 39 41 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.09 $Y=1.16 $X2=5.27
+ $Y2=1.16
r71 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.09
+ $Y=1.16 $X2=5.09 $Y2=1.16
r72 37 39 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.84 $Y=1.16
+ $X2=5.09 $Y2=1.16
r73 36 37 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.41 $Y=1.16
+ $X2=4.84 $Y2=1.16
r74 34 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.07 $Y=1.16
+ $X2=4.41 $Y2=1.16
r75 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.07
+ $Y=1.16 $X2=4.07 $Y2=1.16
r76 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.98 $Y=1.16 $X2=4.07
+ $Y2=1.16
r77 29 40 31.9138 $w=2.58e-07 $l=7.2e-07 $layer=LI1_cond $X=4.37 $Y=1.145
+ $X2=5.09 $Y2=1.145
r78 29 35 13.2974 $w=2.58e-07 $l=3e-07 $layer=LI1_cond $X=4.37 $Y=1.145 $X2=4.07
+ $Y2=1.145
r79 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.27 $Y=1.325
+ $X2=5.27 $Y2=1.16
r80 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.27 $Y=1.325
+ $X2=5.27 $Y2=1.985
r81 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=1.16
r82 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.56
r83 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.325
+ $X2=4.84 $Y2=1.16
r84 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.84 $Y=1.325
+ $X2=4.84 $Y2=1.985
r85 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=0.995
+ $X2=4.84 $Y2=1.16
r86 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.84 $Y=0.995
+ $X2=4.84 $Y2=0.56
r87 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.325
+ $X2=4.41 $Y2=1.16
r88 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.41 $Y=1.325
+ $X2=4.41 $Y2=1.985
r89 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=0.995
+ $X2=4.41 $Y2=1.16
r90 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.41 $Y=0.995
+ $X2=4.41 $Y2=0.56
r91 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.325
+ $X2=3.98 $Y2=1.16
r92 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.98 $Y=1.325 $X2=3.98
+ $Y2=1.985
r93 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=1.16
r94 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.98 $Y=0.995 $X2=3.98
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 45 47 66 67 73
r97 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r99 64 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r100 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r101 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r102 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r104 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r105 55 58 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r106 55 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r107 54 57 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r108 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 52 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=2.72
+ $X2=1.145 $Y2=2.72
r110 52 54 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.31 $Y=2.72 $X2=1.61
+ $Y2=2.72
r111 51 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 48 70 4.31589 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r114 48 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 47 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=2.72
+ $X2=1.145 $Y2=2.72
r116 47 50 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.98 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 45 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r119 43 63 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.32 $Y=2.72 $X2=5.29
+ $Y2=2.72
r120 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=2.72
+ $X2=5.485 $Y2=2.72
r121 42 66 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.65 $Y=2.72 $X2=5.75
+ $Y2=2.72
r122 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.65 $Y=2.72
+ $X2=5.485 $Y2=2.72
r123 40 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.46 $Y=2.72 $X2=4.37
+ $Y2=2.72
r124 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=2.72
+ $X2=4.625 $Y2=2.72
r125 39 63 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.79 $Y=2.72 $X2=5.29
+ $Y2=2.72
r126 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=2.72
+ $X2=4.625 $Y2=2.72
r127 37 57 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.63 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 37 38 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.63 $Y=2.72 $X2=3.77
+ $Y2=2.72
r129 36 60 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r130 36 38 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.91 $Y=2.72 $X2=3.77
+ $Y2=2.72
r131 32 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=2.635
+ $X2=5.485 $Y2=2.72
r132 32 34 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.485 $Y=2.635
+ $X2=5.485 $Y2=1.965
r133 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=2.635
+ $X2=4.625 $Y2=2.72
r134 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.625 $Y=2.635
+ $X2=4.625 $Y2=2.34
r135 24 38 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.635
+ $X2=3.77 $Y2=2.72
r136 24 26 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.77 $Y=2.635
+ $X2=3.77 $Y2=2.36
r137 20 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.72
r138 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.34
r139 16 70 3.08278 $w=2.85e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.202 $Y2=2.72
r140 16 18 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.262 $Y2=2
r141 5 34 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=5.345
+ $Y=1.485 $X2=5.485 $Y2=1.965
r142 4 30 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.485 $X2=4.625 $Y2=2.34
r143 3 26 600 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.745 $Y2=2.36
r144 2 22 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.485 $X2=1.145 $Y2=2.34
r145 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=1.485 $X2=0.285 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%A_115_297# 1 2 3 4 15 17 18 20 25
r38 23 25 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=2.435 $Y=2.37
+ $X2=3.295 $Y2=2.37
r39 21 28 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.67 $Y=2.37
+ $X2=1.575 $Y2=2.37
r40 21 23 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=1.67 $Y=2.37
+ $X2=2.435 $Y2=2.37
r41 20 28 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.575 $Y=2.275
+ $X2=1.575 $Y2=2.37
r42 19 20 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=1.575 $Y=2.085
+ $X2=1.575 $Y2=2.275
r43 17 19 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.48 $Y=2
+ $X2=1.575 $Y2=2.085
r44 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.48 $Y=2 $X2=0.81
+ $Y2=2
r45 13 18 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.692 $Y=2.085
+ $X2=0.81 $Y2=2
r46 13 15 10.5436 $w=2.33e-07 $l=2.15e-07 $layer=LI1_cond $X=0.692 $Y=2.085
+ $X2=0.692 $Y2=2.3
r47 4 25 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.485 $X2=3.295 $Y2=2.36
r48 3 23 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.485 $X2=2.435 $Y2=2.36
r49 2 28 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.485 $X2=1.575 $Y2=2.3
r50 1 15 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.485 $X2=0.715 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%Y 1 2 3 4 5 6 19 25 33 35 36 39 41 47 49 52
+ 54
r81 52 54 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=5.63 $Y=0.845
+ $X2=5.63 $Y2=0.85
r82 49 52 2.71052 $w=4.1e-07 $l=1.15e-07 $layer=LI1_cond $X=5.63 $Y=0.73
+ $X2=5.63 $Y2=0.845
r83 49 54 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=5.63 $Y=0.89 $X2=5.63
+ $Y2=0.85
r84 48 49 15.6001 $w=4.08e-07 $l=5.55e-07 $layer=LI1_cond $X=5.63 $Y=1.445
+ $X2=5.63 $Y2=0.89
r85 43 45 0.198374 $w=6.15e-07 $l=1e-08 $layer=LI1_cond $X=4.185 $Y=1.765
+ $X2=4.195 $Y2=1.765
r86 42 47 2.41622 $w=4.47e-07 $l=2.35763e-07 $layer=LI1_cond $X=5.15 $Y=1.572
+ $X2=5.055 $Y2=1.765
r87 41 48 7.30951 $w=2.55e-07 $l=2.60883e-07 $layer=LI1_cond $X=5.425 $Y=1.572
+ $X2=5.63 $Y2=1.445
r88 41 42 12.4283 $w=2.53e-07 $l=2.75e-07 $layer=LI1_cond $X=5.425 $Y=1.572
+ $X2=5.15 $Y2=1.572
r89 37 47 4.54712 $w=1.9e-07 $l=3.2e-07 $layer=LI1_cond $X=5.055 $Y=2.085
+ $X2=5.055 $Y2=1.765
r90 37 39 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=5.055 $Y=2.085
+ $X2=5.055 $Y2=2.3
r91 36 45 1.81094 $w=6.4e-07 $l=9.5e-08 $layer=LI1_cond $X=4.29 $Y=1.765
+ $X2=4.195 $Y2=1.765
r92 35 47 2.41622 $w=4.47e-07 $l=9.5e-08 $layer=LI1_cond $X=4.96 $Y=1.765
+ $X2=5.055 $Y2=1.765
r93 35 36 12.5214 $w=6.38e-07 $l=6.7e-07 $layer=LI1_cond $X=4.96 $Y=1.765
+ $X2=4.29 $Y2=1.765
r94 31 43 7.12972 $w=2.1e-07 $l=3.2e-07 $layer=LI1_cond $X=4.185 $Y=2.085
+ $X2=4.185 $Y2=1.765
r95 31 33 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=4.185 $Y=2.085
+ $X2=4.185 $Y2=2.3
r96 27 30 43.0913 $w=2.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.195 $Y=0.73
+ $X2=5.055 $Y2=0.73
r97 25 49 4.8318 $w=2.3e-07 $l=2.05e-07 $layer=LI1_cond $X=5.425 $Y=0.73
+ $X2=5.63 $Y2=0.73
r98 25 30 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.425 $Y=0.73
+ $X2=5.055 $Y2=0.73
r99 21 24 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.005 $Y=1.94
+ $X2=2.865 $Y2=1.94
r100 19 43 12.1451 $w=6.15e-07 $l=3.2596e-07 $layer=LI1_cond $X=3.935 $Y=1.94
+ $X2=4.185 $Y2=1.765
r101 19 24 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.935 $Y=1.94
+ $X2=2.865 $Y2=1.94
r102 6 47 600 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.485 $X2=5.055 $Y2=1.825
r103 6 39 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.485 $X2=5.055 $Y2=2.3
r104 5 45 600 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.485 $X2=4.195 $Y2=1.825
r105 5 33 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.485 $X2=4.195 $Y2=2.3
r106 4 24 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=1.485 $X2=2.865 $Y2=1.94
r107 3 21 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.485 $X2=2.005 $Y2=1.94
r108 2 30 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.235 $X2=5.055 $Y2=0.7
r109 1 27 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.055
+ $Y=0.235 $X2=4.195 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%A_32_47# 1 2 3 4 5 6 7 22 36 40
r54 38 40 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=4.625 $Y=0.35
+ $X2=5.485 $Y2=0.35
r55 36 38 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=3.86 $Y=0.35
+ $X2=4.625 $Y2=0.35
r56 33 35 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=3.745 $Y=0.615
+ $X2=3.745 $Y2=0.54
r57 32 36 6.89722 $w=1.9e-07 $l=1.55403e-07 $layer=LI1_cond $X=3.745 $Y=0.445
+ $X2=3.86 $Y2=0.35
r58 32 35 4.76009 $w=2.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.745 $Y=0.445
+ $X2=3.745 $Y2=0.54
r59 29 31 46.5277 $w=2.03e-07 $l=8.6e-07 $layer=LI1_cond $X=2.005 $Y=0.717
+ $X2=2.865 $Y2=0.717
r60 27 29 46.5277 $w=2.03e-07 $l=8.6e-07 $layer=LI1_cond $X=1.145 $Y=0.717
+ $X2=2.005 $Y2=0.717
r61 24 27 46.5277 $w=2.03e-07 $l=8.6e-07 $layer=LI1_cond $X=0.285 $Y=0.717
+ $X2=1.145 $Y2=0.717
r62 22 33 6.84582 $w=2.05e-07 $l=1.57972e-07 $layer=LI1_cond $X=3.63 $Y=0.717
+ $X2=3.745 $Y2=0.615
r63 22 31 41.388 $w=2.03e-07 $l=7.65e-07 $layer=LI1_cond $X=3.63 $Y=0.717
+ $X2=2.865 $Y2=0.717
r64 7 40 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.235 $X2=5.485 $Y2=0.36
r65 6 38 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.485
+ $Y=0.235 $X2=4.625 $Y2=0.36
r66 5 35 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.765 $Y2=0.54
r67 4 31 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.235 $X2=2.865 $Y2=0.7
r68 3 29 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.235 $X2=2.005 $Y2=0.7
r69 2 27 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.7
r70 1 24 182 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_4%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 48
+ 54 55 58 61 64
r81 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r82 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r83 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r84 55 65 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=3.45
+ $Y2=0
r85 54 55 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r86 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.295
+ $Y2=0
r87 52 54 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=3.46 $Y=0 $X2=5.75
+ $Y2=0
r88 51 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r89 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r90 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.295
+ $Y2=0
r91 48 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=2.99
+ $Y2=0
r92 47 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r93 47 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r94 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r95 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.575
+ $Y2=0
r96 44 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=2.07
+ $Y2=0
r97 43 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r98 43 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r99 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r100 40 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r101 40 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.15
+ $Y2=0
r102 39 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.575
+ $Y2=0
r103 39 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.15
+ $Y2=0
r104 34 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r105 34 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.23
+ $Y2=0
r106 32 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r107 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r108 30 46 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.07
+ $Y2=0
r109 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.435
+ $Y2=0
r110 29 50 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.99
+ $Y2=0
r111 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.435
+ $Y2=0
r112 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0
r113 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0.36
r114 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0
r115 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0.36
r116 17 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0
r117 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0.36
r118 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r119 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.36
r120 4 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.235 $X2=3.295 $Y2=0.36
r121 3 23 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.235 $X2=2.435 $Y2=0.36
r122 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.575 $Y2=0.36
r123 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.36
.ends


* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s15_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
M1000 VPWR a_282_47# a_394_47# VPB phighvt w=820000u l=150000u
+  ad=1.3732e+12p pd=6.84e+06u as=2.173e+11p ps=2.17e+06u
M1001 a_282_47# a_27_47# VPWR VPB phighvt w=820000u l=150000u
+  ad=2.173e+11p pd=2.17e+06u as=0p ps=0u
M1002 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=8.8045e+11p pd=5.44e+06u as=1.113e+11p ps=1.37e+06u
M1003 X a_394_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1004 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1005 VGND a_282_47# a_394_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1006 X a_394_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1007 a_282_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a31o_1.spice.pex
* Created: Thu Aug 27 14:04:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A31O_1%A_80_21# 1 2 9 12 15 16 17 20 22 30 32 35 37
+ 38 41
r81 37 38 7.14892 $w=4.53e-07 $l=8.5e-08 $layer=LI1_cond $X=2.732 $Y=1.91
+ $X2=2.732 $Y2=1.825
r82 30 42 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.537 $Y=1.16
+ $X2=0.537 $Y2=1.325
r83 30 41 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.537 $Y=1.16
+ $X2=0.537 $Y2=0.995
r84 29 32 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.54 $Y=1.16
+ $X2=0.68 $Y2=1.16
r85 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.16 $X2=0.54 $Y2=1.16
r86 26 38 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.875 $Y=0.825
+ $X2=2.875 $Y2=1.825
r87 23 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.74
+ $X2=2.14 $Y2=0.74
r88 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.79 $Y=0.74
+ $X2=2.875 $Y2=0.825
r89 22 23 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.79 $Y=0.74
+ $X2=2.305 $Y2=0.74
r90 18 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.655
+ $X2=2.14 $Y2=0.74
r91 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.14 $Y=0.655
+ $X2=2.14 $Y2=0.4
r92 16 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.74
+ $X2=2.14 $Y2=0.74
r93 16 17 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=1.975 $Y=0.74
+ $X2=0.765 $Y2=0.74
r94 15 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.995
+ $X2=0.68 $Y2=1.16
r95 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=0.825
+ $X2=0.765 $Y2=0.74
r96 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=0.825
+ $X2=0.68 $Y2=0.995
r97 12 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r98 9 41 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.995
r99 2 37 300 $w=1.7e-07 $l=5.13323e-07 $layer=licon1_PDIFF $count=2 $X=2.475
+ $Y=1.485 $X2=2.67 $Y2=1.91
r100 1 35 182 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.235 $X2=2.14 $Y2=0.74
r101 1 20 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.235 $X2=2.14 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%A3 3 6 8 9 13 14 15
c37 15 0 1.08026e-19 $X=1.02 $Y=0.995
c38 14 0 1.73971e-19 $X=1.02 $Y=1.16
r39 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.02 $Y2=1.325
r40 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.02 $Y2=0.995
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.02
+ $Y=1.16 $X2=1.02 $Y2=1.16
r42 9 25 10.9884 $w=2.13e-07 $l=2.05e-07 $layer=LI1_cond $X=1.132 $Y=1.53
+ $X2=1.132 $Y2=1.325
r43 8 25 6.1189 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=1.087 $Y=1.19
+ $X2=1.087 $Y2=1.325
r44 8 14 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=1.087 $Y=1.19 $X2=1.087
+ $Y2=1.16
r45 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.97 $Y=1.985
+ $X2=0.97 $Y2=1.325
r46 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.97 $Y=0.56 $X2=0.97
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%A2 3 6 8 9 13 14 15
r35 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.16 $X2=1.5
+ $Y2=1.325
r36 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.16 $X2=1.5
+ $Y2=0.995
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.16 $X2=1.5 $Y2=1.16
r38 8 9 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.557 $Y=1.19
+ $X2=1.557 $Y2=1.53
r39 8 14 1.2131 $w=2.83e-07 $l=3e-08 $layer=LI1_cond $X=1.557 $Y=1.19 $X2=1.557
+ $Y2=1.16
r40 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.44 $Y=1.985
+ $X2=1.44 $Y2=1.325
r41 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.44 $Y=0.56 $X2=1.44
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%A1 3 6 8 9 13 14 15
c36 13 0 1.54339e-19 $X=1.98 $Y=1.16
r37 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.16
+ $X2=1.98 $Y2=1.325
r38 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.16
+ $X2=1.98 $Y2=0.995
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.16 $X2=1.98 $Y2=1.16
r40 8 9 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.027 $Y=1.19
+ $X2=2.027 $Y2=1.53
r41 8 14 1.30465 $w=2.63e-07 $l=3e-08 $layer=LI1_cond $X=2.027 $Y=1.19 $X2=2.027
+ $Y2=1.16
r42 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.92 $Y=1.985
+ $X2=1.92 $Y2=1.325
r43 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.92 $Y=0.56 $X2=1.92
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%B1 3 6 8 9 13 15
r28 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.46 $Y2=1.325
r29 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.46 $Y2=0.995
r30 8 9 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.497 $Y=1.16
+ $X2=2.497 $Y2=1.53
r31 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r32 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.4 $Y=1.985 $X2=2.4
+ $Y2=1.325
r33 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.56 $X2=2.4
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%X 1 2 10 13 14 15 16 17 22
c20 14 0 5.37596e-20 $X=0.26 $Y=1.575
c21 10 0 1.08026e-19 $X=0.26 $Y=0.81
r22 17 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.21
+ $X2=0.26 $Y2=2.34
r23 16 17 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.87
+ $X2=0.26 $Y2=2.21
r24 15 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.51
+ $X2=0.26 $Y2=0.385
r25 13 14 5.02519 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=1.575
r26 11 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=1.74
+ $X2=0.26 $Y2=1.87
r27 11 13 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=1.74 $X2=0.26
+ $Y2=1.66
r28 10 14 44.6555 $w=1.88e-07 $l=7.65e-07 $layer=LI1_cond $X=0.19 $Y=0.81
+ $X2=0.19 $Y2=1.575
r29 9 15 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.26 $Y2=0.51
r30 9 10 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.26 $Y2=0.81
r31 2 31 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r32 2 13 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r33 1 22 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%VPWR 1 2 9 15 17 19 24 34 35 38 41
r46 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r47 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r49 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 32 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 31 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.72
+ $X2=1.68 $Y2=2.72
r54 29 31 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.845 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 28 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 28 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 25 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.72 $Y2=2.72
r59 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.68 $Y2=2.72
r61 24 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 19 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.72 $Y2=2.72
r63 19 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 17 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.635
+ $X2=1.68 $Y2=2.72
r67 13 15 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.68 $Y=2.635
+ $X2=1.68 $Y2=2.25
r68 9 12 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.72 $Y=1.66 $X2=0.72
+ $Y2=2.34
r69 7 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.72
r70 7 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=2.635
+ $X2=0.72 $Y2=2.34
r71 2 15 600 $w=1.7e-07 $l=8.43475e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.485 $X2=1.68 $Y2=2.25
r72 1 12 400 $w=1.7e-07 $l=9.36149e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.72 $Y2=2.34
r73 1 9 400 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.72 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%A_209_297# 1 2 7 9 11 13 15
c26 13 0 1.54339e-19 $X=2.2 $Y=1.995
r27 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=1.995 $X2=2.2
+ $Y2=1.91
r28 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.2 $Y=1.995
+ $X2=2.2 $Y2=2.25
r29 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=1.91
+ $X2=1.16 $Y2=1.91
r30 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=1.91
+ $X2=2.2 $Y2=1.91
r31 11 12 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.075 $Y=1.91
+ $X2=1.285 $Y2=1.91
r32 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=1.995 $X2=1.16
+ $Y2=1.91
r33 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.16 $Y=1.995
+ $X2=1.16 $Y2=2.25
r34 2 20 600 $w=1.7e-07 $l=5.00749e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.16 $Y2=1.91
r35 2 15 600 $w=1.7e-07 $l=8.43475e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.16 $Y2=2.25
r36 1 18 600 $w=1.7e-07 $l=4.96488e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.485 $X2=1.2 $Y2=1.91
r37 1 9 600 $w=1.7e-07 $l=8.38928e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.485 $X2=1.2 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r45 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r48 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.64
+ $Y2=0
r50 27 29 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.99
+ $Y2=0
r51 26 37 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r52 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.76
+ $Y2=0
r55 23 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r56 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.64
+ $Y2=0
r57 22 25 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=1.15 $Y2=0
r58 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.76
+ $Y2=0
r59 17 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r60 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0
r63 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0.4
r64 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r65 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.4
r66 2 13 182 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.64 $Y2=0.4
r67 1 9 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.76 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__o2bb2a_1.spice
* Created: Thu Aug 27 14:38:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2bb2a_1.pex.spice"
.subckt sky130_fd_sc_hd__o2bb2a_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_76_199#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.119825 AS=0.169 PD=1.19065 PS=1.82 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1001 A_205_47# N_A1_N_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.0774252 PD=0.735 PS=0.769346 NRD=29.28 NRS=8.568 M=1 R=2.8
+ SA=75000.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_206_369#_M1010_d N_A2_N_M1010_g A_205_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.06615 PD=1.36 PS=0.735 NRD=0 NRS=29.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_489_47#_M1002_d N_A_206_369#_M1002_g N_A_76_199#_M1002_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_B2_M1000_g N_A_489_47#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_489_47#_M1007_d N_B1_M1007_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_76_199#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.205282 AS=0.26 PD=1.88028 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1005 N_A_206_369#_M1005_d N_A1_N_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.129 AS=0.0862183 PD=1.18 PS=0.789718 NRD=118.259 NRS=30.4759 M=1
+ R=2.8 SA=75000.7 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A2_N_M1011_g N_A_206_369#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.20925 AS=0.129 PD=1.345 PS=1.18 NRD=93.7917 NRS=118.259 M=1 R=2.8
+ SA=75001.2 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_76_199#_M1008_d N_A_206_369#_M1008_g N_VPWR_M1011_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0672 AS=0.20925 PD=0.74 PS=1.345 NRD=0 NRS=207.874 M=1
+ R=2.8 SA=75002.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_585_369# N_B2_M1004_g N_A_76_199#_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=21.0987 M=1 R=2.8
+ SA=75002.6 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g A_585_369# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__o2bb2a_1.pxi.spice"
*
.ends
*
*

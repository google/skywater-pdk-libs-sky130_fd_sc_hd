* File: sky130_fd_sc_hd__a21o_4.pex.spice
* Created: Tue Sep  1 18:52:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21O_4%A_84_21# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 38 45 47 48 49 52 56 58 63
c125 58 0 4.87616e-20 $X=4.085 $Y=0.755
r126 71 72 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.355 $Y=1.16
+ $X2=1.785 $Y2=1.16
r127 67 69 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.925 $Y2=1.16
r128 63 65 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.225 $Y=0.57
+ $X2=4.225 $Y2=0.755
r129 59 61 3.05 $w=1.7e-07 $l=9.80051e-08 $layer=LI1_cond $X=3.045 $Y=0.755
+ $X2=2.96 $Y2=0.727
r130 58 65 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.085 $Y=0.755
+ $X2=4.225 $Y2=0.755
r131 58 59 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.085 $Y=0.755
+ $X2=3.045 $Y2=0.755
r132 54 61 3.05 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=2.96 $Y=0.84 $X2=2.96
+ $Y2=0.727
r133 54 56 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.96 $Y=0.84
+ $X2=2.96 $Y2=1.62
r134 50 61 3.05 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=2.96 $Y=0.615 $X2=2.96
+ $Y2=0.727
r135 50 52 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.96 $Y=0.615
+ $X2=2.96 $Y2=0.42
r136 48 61 3.05 $w=1.7e-07 $l=9.75705e-08 $layer=LI1_cond $X=2.875 $Y=0.7
+ $X2=2.96 $Y2=0.727
r137 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.875 $Y=0.7
+ $X2=2.205 $Y2=0.7
r138 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=0.785
+ $X2=2.205 $Y2=0.7
r139 46 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.12 $Y=0.785
+ $X2=2.12 $Y2=0.995
r140 45 72 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=1.785 $Y2=1.16
r141 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.84
+ $Y=1.16 $X2=1.84 $Y2=1.16
r142 41 71 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=1.355 $Y2=1.16
r143 41 69 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=0.925 $Y2=1.16
r144 40 44 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.16 $Y=1.16
+ $X2=1.84 $Y2=1.16
r145 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.16 $X2=1.16 $Y2=1.16
r146 38 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.035 $Y=1.16
+ $X2=2.12 $Y2=0.995
r147 38 44 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.035 $Y=1.16
+ $X2=1.84 $Y2=1.16
r148 34 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.16
r149 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.985
r150 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=0.995
+ $X2=1.785 $Y2=1.16
r151 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.785 $Y=0.995
+ $X2=1.785 $Y2=0.56
r152 27 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.325
+ $X2=1.355 $Y2=1.16
r153 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.355 $Y=1.325
+ $X2=1.355 $Y2=1.985
r154 24 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=0.995
+ $X2=1.355 $Y2=1.16
r155 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.355 $Y=0.995
+ $X2=1.355 $Y2=0.56
r156 20 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.325
+ $X2=0.925 $Y2=1.16
r157 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.325
+ $X2=0.925 $Y2=1.985
r158 17 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=0.995
+ $X2=0.925 $Y2=1.16
r159 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.925 $Y=0.995
+ $X2=0.925 $Y2=0.56
r160 13 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r161 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.985
r162 10 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=1.16
r163 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=0.56
r164 3 56 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.62
r165 2 63 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.085
+ $Y=0.235 $X2=4.22 $Y2=0.57
r166 1 61 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.76
r167 1 52 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%B1 1 3 6 8 10 13 15 22
r49 21 22 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=3.17 $Y2=1.16
r50 18 21 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.62 $Y=1.16 $X2=2.75
+ $Y2=1.16
r51 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.16 $X2=2.62 $Y2=1.16
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.325
+ $X2=3.17 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.17 $Y=1.325
+ $X2=3.17 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=0.995
+ $X2=3.17 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.17 $Y=0.995
+ $X2=3.17 $Y2=0.56
r56 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.325
+ $X2=2.75 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.325 $X2=2.75
+ $Y2=1.985
r58 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=0.995
+ $X2=2.75 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.995 $X2=2.75
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%A2 3 7 10 13 16 17 18 21 23 29 30 32 36 38 40
c85 21 0 1.32673e-19 $X=3.59 $Y=1.16
r86 32 40 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=1.595
+ $X2=4.81 $Y2=1.51
r87 32 40 1.52122 $w=2.48e-07 $l=3.3e-08 $layer=LI1_cond $X=4.81 $Y=1.477
+ $X2=4.81 $Y2=1.51
r88 30 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.91 $Y=1.16
+ $X2=4.91 $Y2=1.325
r89 30 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.91 $Y=1.16
+ $X2=4.91 $Y2=0.995
r90 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.91
+ $Y=1.16 $X2=4.91 $Y2=1.16
r91 26 32 8.62027 $w=2.48e-07 $l=1.87e-07 $layer=LI1_cond $X=4.81 $Y=1.29
+ $X2=4.81 $Y2=1.477
r92 25 29 4.90401 $w=2.33e-07 $l=1e-07 $layer=LI1_cond $X=4.81 $Y=1.172 $X2=4.91
+ $Y2=1.172
r93 25 26 0.335614 $w=2.5e-07 $l=1.18e-07 $layer=LI1_cond $X=4.81 $Y=1.172
+ $X2=4.81 $Y2=1.29
r94 21 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.16
+ $X2=3.59 $Y2=0.995
r95 20 23 6.17535 $w=2.63e-07 $l=1.42e-07 $layer=LI1_cond $X=3.59 $Y=1.142
+ $X2=3.732 $Y2=1.142
r96 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.16 $X2=3.59 $Y2=1.16
r97 17 32 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=1.595
+ $X2=4.81 $Y2=1.595
r98 17 18 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.685 $Y=1.595
+ $X2=3.82 $Y2=1.595
r99 16 18 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=3.732 $Y=1.51
+ $X2=3.82 $Y2=1.595
r100 15 23 3.18883 $w=1.75e-07 $l=1.33e-07 $layer=LI1_cond $X=3.732 $Y=1.275
+ $X2=3.732 $Y2=1.142
r101 15 16 14.8935 $w=1.73e-07 $l=2.35e-07 $layer=LI1_cond $X=3.732 $Y=1.275
+ $X2=3.732 $Y2=1.51
r102 13 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.85 $Y=1.985
+ $X2=4.85 $Y2=1.325
r103 10 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.85 $Y=0.56
+ $X2=4.85 $Y2=0.995
r104 7 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.63 $Y=0.56
+ $X2=3.63 $Y2=0.995
r105 1 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.325
+ $X2=3.59 $Y2=1.16
r106 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.59 $Y=1.325
+ $X2=3.59 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%A1 1 3 6 8 10 13 15 22
c45 8 0 4.87616e-20 $X=4.43 $Y=0.995
r46 20 22 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.19 $Y=1.16
+ $X2=4.43 $Y2=1.16
r47 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=1.16 $X2=4.19 $Y2=1.16
r48 17 20 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.01 $Y=1.16 $X2=4.19
+ $Y2=1.16
r49 15 21 8.69768 $w=2.63e-07 $l=2e-07 $layer=LI1_cond $X=4.39 $Y=1.142 $X2=4.19
+ $Y2=1.142
r50 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.43 $Y=1.325
+ $X2=4.43 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.43 $Y=1.325
+ $X2=4.43 $Y2=1.985
r52 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=0.56
r54 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.325
+ $X2=4.01 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.01 $Y=1.325 $X2=4.01
+ $Y2=1.985
r56 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=0.995
+ $X2=4.01 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.01 $Y=0.995 $X2=4.01
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%VPWR 1 2 3 4 5 16 18 22 26 32 36 39 40 42 43
+ 44 46 51 67 68 74 77
r97 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r98 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r99 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r100 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r101 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r102 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r104 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r105 59 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r106 58 61 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r108 56 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.04 $Y2=2.72
r109 56 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.53 $Y2=2.72
r110 55 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r111 55 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.14 $Y2=2.72
r114 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.61 $Y2=2.72
r115 51 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.04 $Y2=2.72
r116 51 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r117 50 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 47 71 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.222 $Y2=2.72
r120 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 46 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.14 $Y2=2.72
r122 46 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 44 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r125 42 64 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=2.72
+ $X2=4.37 $Y2=2.72
r126 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=2.72
+ $X2=4.64 $Y2=2.72
r127 41 67 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.805 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=2.72
+ $X2=4.64 $Y2=2.72
r129 39 61 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.45 $Y2=2.72
r130 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.8 $Y2=2.72
r131 38 64 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.965 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=2.72
+ $X2=3.8 $Y2=2.72
r133 34 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=2.635
+ $X2=4.64 $Y2=2.72
r134 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.64 $Y=2.635
+ $X2=4.64 $Y2=2.36
r135 30 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=2.635 $X2=3.8
+ $Y2=2.72
r136 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.8 $Y=2.635
+ $X2=3.8 $Y2=2.36
r137 26 29 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.04 $Y=1.68
+ $X2=2.04 $Y2=2.36
r138 24 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r139 24 29 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.36
r140 20 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.72
r141 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.02
r142 16 71 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.222 $Y2=2.72
r143 16 18 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.28 $Y2=2.02
r144 5 36 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.485 $X2=4.64 $Y2=2.36
r145 4 32 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=1.485 $X2=3.8 $Y2=2.36
r146 3 29 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.485 $X2=2 $Y2=2.36
r147 3 26 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.485 $X2=2 $Y2=1.68
r148 2 22 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.485 $X2=1.14 $Y2=2.02
r149 1 18 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%X 1 2 3 4 15 17 21 23 25 27 32 38
r45 35 38 1.35638 $w=4.83e-07 $l=5.5e-08 $layer=LI1_cond $X=0.387 $Y=1.585
+ $X2=0.387 $Y2=1.53
r46 32 35 2.90768 $w=3.27e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.47 $Y=1.67
+ $X2=0.387 $Y2=1.585
r47 32 38 0.369921 $w=4.83e-07 $l=1.5e-08 $layer=LI1_cond $X=0.387 $Y=1.515
+ $X2=0.387 $Y2=1.53
r48 29 32 18.0028 $w=4.83e-07 $l=7.3e-07 $layer=LI1_cond $X=0.387 $Y=0.785
+ $X2=0.387 $Y2=1.515
r49 25 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.755
+ $X2=1.61 $Y2=1.67
r50 25 27 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.61 $Y=1.755
+ $X2=1.61 $Y2=2.02
r51 24 32 3.78066 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=0.795 $Y=1.67
+ $X2=0.47 $Y2=1.67
r52 23 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.485 $Y=1.67
+ $X2=1.61 $Y2=1.67
r53 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.485 $Y=1.67
+ $X2=0.795 $Y2=1.67
r54 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.71 $Y=0.7 $X2=1.57
+ $Y2=0.7
r55 17 29 9.10402 $w=1.7e-07 $l=2.82319e-07 $layer=LI1_cond $X=0.63 $Y=0.7
+ $X2=0.387 $Y2=0.785
r56 17 19 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.63 $Y=0.7 $X2=0.71
+ $Y2=0.7
r57 13 32 2.90768 $w=3.27e-07 $l=2.79285e-07 $layer=LI1_cond $X=0.71 $Y=1.755
+ $X2=0.47 $Y2=1.67
r58 13 15 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.71 $Y=1.755
+ $X2=0.71 $Y2=2.02
r59 4 31 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.485 $X2=1.57 $Y2=1.67
r60 4 27 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.485 $X2=1.57 $Y2=2.02
r61 3 32 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.485 $X2=0.71 $Y2=1.67
r62 3 15 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.485 $X2=0.71 $Y2=2.02
r63 2 21 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.7
r64 1 19 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%A_483_297# 1 2 3 4 15 17 18 21 27 31 33 39 43
+ 45
c61 27 0 1.32673e-19 $X=4.135 $Y=1.935
r62 37 45 3.22182 $w=2.92e-07 $l=1.01833e-07 $layer=LI1_cond $X=5.232 $Y=1.85
+ $X2=5.195 $Y2=1.935
r63 37 39 9.94265 $w=2.53e-07 $l=2.2e-07 $layer=LI1_cond $X=5.232 $Y=1.85
+ $X2=5.232 $Y2=1.63
r64 34 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=1.935
+ $X2=4.22 $Y2=1.935
r65 33 45 3.35233 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.03 $Y=1.935
+ $X2=5.195 $Y2=1.935
r66 33 34 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.03 $Y=1.935
+ $X2=4.305 $Y2=1.935
r67 29 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.22 $Y=2.02 $X2=4.22
+ $Y2=1.935
r68 29 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.22 $Y=2.02
+ $X2=4.22 $Y2=2.3
r69 28 41 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.465 $Y=1.935
+ $X2=3.375 $Y2=1.935
r70 27 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=1.935
+ $X2=4.22 $Y2=1.935
r71 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.135 $Y=1.935
+ $X2=3.465 $Y2=1.935
r72 24 26 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=3.375 $Y=2.295
+ $X2=3.375 $Y2=2.055
r73 23 41 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=2.02
+ $X2=3.375 $Y2=1.935
r74 23 26 2.15657 $w=1.78e-07 $l=3.5e-08 $layer=LI1_cond $X=3.375 $Y=2.02
+ $X2=3.375 $Y2=2.055
r75 19 41 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=1.85
+ $X2=3.375 $Y2=1.935
r76 19 21 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=3.375 $Y=1.85
+ $X2=3.375 $Y2=1.61
r77 17 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.285 $Y=2.38
+ $X2=3.375 $Y2=2.295
r78 17 18 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.285 $Y=2.38
+ $X2=2.625 $Y2=2.38
r79 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.54 $Y=2.295
+ $X2=2.625 $Y2=2.38
r80 13 15 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.54 $Y=2.295
+ $X2=2.54 $Y2=1.86
r81 4 45 300 $w=1.7e-07 $l=6.05124e-07 $layer=licon1_PDIFF $count=2 $X=4.925
+ $Y=1.485 $X2=5.195 $Y2=1.97
r82 4 39 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.485 $X2=5.195 $Y2=1.63
r83 3 43 600 $w=1.7e-07 $l=5.13079e-07 $layer=licon1_PDIFF $count=1 $X=4.085
+ $Y=1.485 $X2=4.22 $Y2=1.935
r84 3 31 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.085
+ $Y=1.485 $X2=4.22 $Y2=2.3
r85 2 26 600 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.485 $X2=3.38 $Y2=2.055
r86 2 21 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.485 $X2=3.38 $Y2=1.61
r87 1 15 300 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=2 $X=2.415
+ $Y=1.485 $X2=2.54 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_4%VGND 1 2 3 4 5 16 18 22 26 30 33 34 35 37 47
+ 60 61 67 72 78 80
r87 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r88 76 78 9.47869 $w=5.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.685 $Y2=0.18
r89 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r90 74 76 0.225675 $w=5.28e-07 $l=1e-08 $layer=LI1_cond $X=2.52 $Y=0.18 $X2=2.53
+ $Y2=0.18
r91 71 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r92 70 74 10.1554 $w=5.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.07 $Y=0.18
+ $X2=2.52 $Y2=0.18
r93 70 72 9.59153 $w=5.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.07 $Y=0.18
+ $X2=1.91 $Y2=0.18
r94 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r95 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r96 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r97 58 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r98 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r99 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r100 55 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r101 54 57 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r102 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r103 52 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r104 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.585 $Y=0
+ $X2=3.91 $Y2=0
r105 51 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r106 51 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r107 50 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.99 $Y=0
+ $X2=2.685 $Y2=0
r108 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r109 47 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r110 47 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0
+ $X2=2.99 $Y2=0
r111 46 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r112 46 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r113 45 72 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.91
+ $Y2=0
r114 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r115 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r116 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.61 $Y2=0
r117 41 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r118 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r119 38 64 4.84988 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r120 38 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.69
+ $Y2=0
r121 37 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r122 37 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.69 $Y2=0
r123 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r124 35 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r125 33 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.945 $Y=0
+ $X2=4.83 $Y2=0
r126 33 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.085
+ $Y2=0
r127 32 60 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.29
+ $Y2=0
r128 32 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.085
+ $Y2=0
r129 28 34 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=0.085
+ $X2=5.085 $Y2=0
r130 28 30 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.085 $Y=0.085
+ $X2=5.085 $Y2=0.38
r131 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r132 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.36
r133 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r134 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.36
r135 16 64 3.00127 $w=3.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.222 $Y2=0
r136 16 18 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.36
r137 5 30 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.925
+ $Y=0.235 $X2=5.06 $Y2=0.38
r138 4 26 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.42 $Y2=0.36
r139 3 74 91 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.235 $X2=2.52 $Y2=0.36
r140 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.36
r141 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__bufbuf_16.pex.spice
* Created: Thu Aug 27 14:10:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%A 1 3 6 8 14
r25 11 14 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r26 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r27 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r29 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%A_109_47# 1 2 9 13 17 21 25 29 33 35 37 42
+ 47 50 51 52 57
c94 47 0 1.44067e-19 $X=1.96 $Y=1.16
c95 29 0 1.25206e-19 $X=2.25 $Y=1.985
c96 25 0 1.25206e-19 $X=2.25 $Y=0.56
r97 53 55 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.41 $Y=1.16 $X2=1.83
+ $Y2=1.16
r98 48 57 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=1.96 $Y=1.16
+ $X2=2.25 $Y2=1.16
r99 48 55 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=1.96 $Y=1.16
+ $X2=1.83 $Y2=1.16
r100 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.96
+ $Y=1.16 $X2=1.96 $Y2=1.16
r101 45 52 1.92922 $w=2e-07 $l=1.18e-07 $layer=LI1_cond $X=0.845 $Y=1.175
+ $X2=0.727 $Y2=1.175
r102 45 47 61.8318 $w=1.98e-07 $l=1.115e-06 $layer=LI1_cond $X=0.845 $Y=1.175
+ $X2=1.96 $Y2=1.175
r103 43 52 4.50812 $w=2.35e-07 $l=1e-07 $layer=LI1_cond $X=0.727 $Y=1.275
+ $X2=0.727 $Y2=1.175
r104 43 51 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.727 $Y=1.275
+ $X2=0.727 $Y2=1.445
r105 42 52 4.50812 $w=2.35e-07 $l=1e-07 $layer=LI1_cond $X=0.727 $Y=1.075
+ $X2=0.727 $Y2=1.175
r106 42 50 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.727 $Y=1.075
+ $X2=0.727 $Y2=0.905
r107 37 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.63
+ $X2=0.68 $Y2=2.31
r108 35 51 6.73378 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.61
+ $X2=0.68 $Y2=1.445
r109 35 37 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=0.68 $Y=1.61 $X2=0.68
+ $Y2=1.63
r110 31 50 6.73378 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.68 $Y2=0.905
r111 31 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.68 $Y2=0.4
r112 27 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.16
r113 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.985
r114 23 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=1.16
r115 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r116 19 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.16
r117 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.985
r118 15 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=1.16
r119 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=0.56
r120 11 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.16
r121 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.985
r122 7 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.16
r123 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r124 2 39 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.31
r125 2 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.63
r126 1 33 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%A_215_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 72 73 74 77 81 86 88 94 98 101 103 112
c204 112 0 1.44067e-19 $X=4.77 $Y=1.16
c205 94 0 1.39258e-19 $X=4.5 $Y=1.16
c206 59 0 1.25206e-19 $X=4.77 $Y=1.985
c207 55 0 1.25206e-19 $X=4.77 $Y=0.56
r208 109 110 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.35 $Y2=1.16
r209 108 109 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.51 $Y=1.16
+ $X2=3.93 $Y2=1.16
r210 107 108 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.09 $Y=1.16
+ $X2=3.51 $Y2=1.16
r211 95 112 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=4.5 $Y=1.16
+ $X2=4.77 $Y2=1.16
r212 95 110 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=4.5 $Y=1.16
+ $X2=4.35 $Y2=1.16
r213 94 95 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.5
+ $Y=1.16 $X2=4.5 $Y2=1.16
r214 92 107 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.8 $Y=1.16
+ $X2=3.09 $Y2=1.16
r215 92 104 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=2.8 $Y=1.16
+ $X2=2.67 $Y2=1.16
r216 91 94 94.2727 $w=1.98e-07 $l=1.7e-06 $layer=LI1_cond $X=2.8 $Y=1.175
+ $X2=4.5 $Y2=1.175
r217 91 92 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.8
+ $Y=1.16 $X2=2.8 $Y2=1.16
r218 89 103 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.175
+ $X2=2.46 $Y2=1.175
r219 89 91 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.545 $Y=1.175
+ $X2=2.8 $Y2=1.175
r220 88 101 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.445
+ $X2=2.46 $Y2=1.53
r221 87 103 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.46 $Y=1.275
+ $X2=2.46 $Y2=1.175
r222 87 88 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.46 $Y=1.275
+ $X2=2.46 $Y2=1.445
r223 86 103 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.46 $Y=1.075
+ $X2=2.46 $Y2=1.175
r224 85 98 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.46 $Y2=0.82
r225 85 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.46 $Y2=1.075
r226 81 83 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.04 $Y=1.63
+ $X2=2.04 $Y2=2.31
r227 79 101 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.04 $Y=1.53
+ $X2=2.46 $Y2=1.53
r228 79 81 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.04 $Y=1.615
+ $X2=2.04 $Y2=1.63
r229 75 98 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.04 $Y=0.82
+ $X2=2.46 $Y2=0.82
r230 75 77 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=0.735
+ $X2=2.04 $Y2=0.4
r231 73 79 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.53
+ $X2=2.04 $Y2=1.53
r232 73 74 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.875 $Y=1.53
+ $X2=1.365 $Y2=1.53
r233 71 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.82
+ $X2=2.04 $Y2=0.82
r234 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.875 $Y=0.82
+ $X2=1.365 $Y2=0.82
r235 67 69 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.63 $X2=1.2
+ $Y2=2.31
r236 65 74 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.365 $Y2=1.53
r237 65 67 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.2 $Y2=1.63
r238 61 72 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.365 $Y2=0.82
r239 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.4
r240 57 112 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.16
r241 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.985
r242 53 112 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=1.16
r243 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=0.56
r244 49 110 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.16
r245 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.985
r246 45 110 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r247 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
r248 41 109 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.16
r249 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.985
r250 37 109 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=1.16
r251 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=0.56
r252 33 108 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.16
r253 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.985
r254 29 108 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=1.16
r255 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=0.56
r256 25 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.16
r257 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r258 21 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=1.16
r259 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=0.56
r260 17 104 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.16
r261 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r262 13 104 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=1.16
r263 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=0.56
r264 4 83 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2.31
r265 4 81 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.63
r266 3 69 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.31
r267 3 67 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.63
r268 2 77 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.4
r269 1 63 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%A_549_47# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 153 157 158 159 160 163 167 171 173 177 181 186 188 194 197 198
+ 200 203 205 224
c464 224 0 1.39258e-19 $X=11.49 $Y=1.16
c465 160 0 1.25206e-19 $X=3.045 $Y=1.53
c466 158 0 1.25206e-19 $X=3.045 $Y=0.82
r467 221 222 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=10.65 $Y=1.16
+ $X2=11.07 $Y2=1.16
r468 220 221 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=10.23 $Y=1.16
+ $X2=10.65 $Y2=1.16
r469 219 220 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.81 $Y=1.16
+ $X2=10.23 $Y2=1.16
r470 218 219 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.39 $Y=1.16
+ $X2=9.81 $Y2=1.16
r471 217 218 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.97 $Y=1.16
+ $X2=9.39 $Y2=1.16
r472 216 217 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.55 $Y=1.16
+ $X2=8.97 $Y2=1.16
r473 215 216 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.13 $Y=1.16
+ $X2=8.55 $Y2=1.16
r474 214 215 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.71 $Y=1.16
+ $X2=8.13 $Y2=1.16
r475 213 214 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.29 $Y=1.16
+ $X2=7.71 $Y2=1.16
r476 212 213 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.87 $Y=1.16
+ $X2=7.29 $Y2=1.16
r477 211 212 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.87 $Y2=1.16
r478 210 211 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.03 $Y=1.16
+ $X2=6.45 $Y2=1.16
r479 209 210 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=6.03 $Y2=1.16
r480 195 224 91.0912 $w=2.7e-07 $l=4.1e-07 $layer=POLY_cond $X=11.08 $Y=1.16
+ $X2=11.49 $Y2=1.16
r481 195 222 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=11.08 $Y=1.16
+ $X2=11.07 $Y2=1.16
r482 194 195 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=11.08
+ $Y=1.16 $X2=11.08 $Y2=1.16
r483 192 209 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=5.3 $Y=1.16
+ $X2=5.61 $Y2=1.16
r484 192 206 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=5.3 $Y=1.16
+ $X2=5.19 $Y2=1.16
r485 191 194 320.527 $w=1.98e-07 $l=5.78e-06 $layer=LI1_cond $X=5.3 $Y=1.175
+ $X2=11.08 $Y2=1.175
r486 191 192 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=5.3
+ $Y=1.16 $X2=5.3 $Y2=1.16
r487 189 205 0.866423 $w=2e-07 $l=8.8e-08 $layer=LI1_cond $X=5.065 $Y=1.175
+ $X2=4.977 $Y2=1.175
r488 189 191 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.065 $Y=1.175
+ $X2=5.3 $Y2=1.175
r489 188 203 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.977 $Y=1.445
+ $X2=4.977 $Y2=1.53
r490 187 205 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=4.977 $Y=1.275
+ $X2=4.977 $Y2=1.175
r491 187 188 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.977 $Y=1.275
+ $X2=4.977 $Y2=1.445
r492 186 205 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=4.977 $Y=1.075
+ $X2=4.977 $Y2=1.175
r493 185 200 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.977 $Y=0.905
+ $X2=4.977 $Y2=0.82
r494 185 186 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.977 $Y=0.905
+ $X2=4.977 $Y2=1.075
r495 181 183 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.56 $Y=1.63
+ $X2=4.56 $Y2=2.31
r496 179 203 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=4.56 $Y=1.53
+ $X2=4.977 $Y2=1.53
r497 179 181 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.56 $Y2=1.63
r498 175 200 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=4.56 $Y=0.82
+ $X2=4.977 $Y2=0.82
r499 175 177 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.735
+ $X2=4.56 $Y2=0.4
r500 174 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=1.53
+ $X2=3.72 $Y2=1.53
r501 173 179 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.53
+ $X2=4.56 $Y2=1.53
r502 173 174 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.395 $Y=1.53
+ $X2=3.885 $Y2=1.53
r503 172 197 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0.82
+ $X2=3.72 $Y2=0.82
r504 171 175 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0.82
+ $X2=4.56 $Y2=0.82
r505 171 172 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.395 $Y=0.82
+ $X2=3.885 $Y2=0.82
r506 167 169 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.72 $Y=1.63
+ $X2=3.72 $Y2=2.31
r507 165 198 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.615
+ $X2=3.72 $Y2=1.53
r508 165 167 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.72 $Y=1.615
+ $X2=3.72 $Y2=1.63
r509 161 197 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.735
+ $X2=3.72 $Y2=0.82
r510 161 163 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.72 $Y=0.735
+ $X2=3.72 $Y2=0.4
r511 159 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=1.53
+ $X2=3.72 $Y2=1.53
r512 159 160 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.555 $Y=1.53
+ $X2=3.045 $Y2=1.53
r513 157 197 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0.82
+ $X2=3.72 $Y2=0.82
r514 157 158 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.555 $Y=0.82
+ $X2=3.045 $Y2=0.82
r515 153 155 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.88 $Y=1.63
+ $X2=2.88 $Y2=2.31
r516 151 160 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.88 $Y=1.615
+ $X2=3.045 $Y2=1.53
r517 151 153 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.88 $Y=1.615
+ $X2=2.88 $Y2=1.63
r518 147 158 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.88 $Y=0.735
+ $X2=3.045 $Y2=0.82
r519 147 149 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.88 $Y=0.735
+ $X2=2.88 $Y2=0.4
r520 143 224 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.49 $Y=1.295
+ $X2=11.49 $Y2=1.16
r521 143 145 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=11.49 $Y=1.295
+ $X2=11.49 $Y2=1.985
r522 139 224 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.49 $Y=1.025
+ $X2=11.49 $Y2=1.16
r523 139 141 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.49 $Y=1.025
+ $X2=11.49 $Y2=0.56
r524 135 222 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.07 $Y=1.295
+ $X2=11.07 $Y2=1.16
r525 135 137 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=11.07 $Y=1.295
+ $X2=11.07 $Y2=1.985
r526 131 222 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.07 $Y=1.025
+ $X2=11.07 $Y2=1.16
r527 131 133 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.07 $Y=1.025
+ $X2=11.07 $Y2=0.56
r528 127 221 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.65 $Y=1.295
+ $X2=10.65 $Y2=1.16
r529 127 129 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.65 $Y=1.295
+ $X2=10.65 $Y2=1.985
r530 123 221 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.65 $Y=1.025
+ $X2=10.65 $Y2=1.16
r531 123 125 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.65 $Y=1.025
+ $X2=10.65 $Y2=0.56
r532 119 220 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.23 $Y=1.295
+ $X2=10.23 $Y2=1.16
r533 119 121 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.23 $Y=1.295
+ $X2=10.23 $Y2=1.985
r534 115 220 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.23 $Y=1.025
+ $X2=10.23 $Y2=1.16
r535 115 117 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.23 $Y=1.025
+ $X2=10.23 $Y2=0.56
r536 111 219 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.81 $Y=1.295
+ $X2=9.81 $Y2=1.16
r537 111 113 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.81 $Y=1.295
+ $X2=9.81 $Y2=1.985
r538 107 219 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.81 $Y=1.025
+ $X2=9.81 $Y2=1.16
r539 107 109 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.81 $Y=1.025
+ $X2=9.81 $Y2=0.56
r540 103 218 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.39 $Y=1.295
+ $X2=9.39 $Y2=1.16
r541 103 105 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.39 $Y=1.295
+ $X2=9.39 $Y2=1.985
r542 99 218 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.39 $Y=1.025
+ $X2=9.39 $Y2=1.16
r543 99 101 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.39 $Y=1.025
+ $X2=9.39 $Y2=0.56
r544 95 217 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.97 $Y=1.295
+ $X2=8.97 $Y2=1.16
r545 95 97 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.97 $Y=1.295
+ $X2=8.97 $Y2=1.985
r546 91 217 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.97 $Y=1.025
+ $X2=8.97 $Y2=1.16
r547 91 93 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.97 $Y=1.025
+ $X2=8.97 $Y2=0.56
r548 87 216 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.55 $Y=1.295
+ $X2=8.55 $Y2=1.16
r549 87 89 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.55 $Y=1.295
+ $X2=8.55 $Y2=1.985
r550 83 216 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.55 $Y=1.025
+ $X2=8.55 $Y2=1.16
r551 83 85 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.55 $Y=1.025
+ $X2=8.55 $Y2=0.56
r552 79 215 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.13 $Y=1.295
+ $X2=8.13 $Y2=1.16
r553 79 81 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.13 $Y=1.295
+ $X2=8.13 $Y2=1.985
r554 75 215 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.13 $Y=1.025
+ $X2=8.13 $Y2=1.16
r555 75 77 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.13 $Y=1.025
+ $X2=8.13 $Y2=0.56
r556 71 214 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.71 $Y=1.295
+ $X2=7.71 $Y2=1.16
r557 71 73 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.71 $Y=1.295
+ $X2=7.71 $Y2=1.985
r558 67 214 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.71 $Y=1.025
+ $X2=7.71 $Y2=1.16
r559 67 69 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.71 $Y=1.025
+ $X2=7.71 $Y2=0.56
r560 63 213 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.29 $Y=1.295
+ $X2=7.29 $Y2=1.16
r561 63 65 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.29 $Y=1.295
+ $X2=7.29 $Y2=1.985
r562 59 213 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.29 $Y=1.025
+ $X2=7.29 $Y2=1.16
r563 59 61 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.29 $Y=1.025
+ $X2=7.29 $Y2=0.56
r564 55 212 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.87 $Y=1.295
+ $X2=6.87 $Y2=1.16
r565 55 57 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.87 $Y=1.295
+ $X2=6.87 $Y2=1.985
r566 51 212 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.87 $Y=1.025
+ $X2=6.87 $Y2=1.16
r567 51 53 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.87 $Y=1.025
+ $X2=6.87 $Y2=0.56
r568 47 211 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.45 $Y=1.295
+ $X2=6.45 $Y2=1.16
r569 47 49 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.45 $Y=1.295
+ $X2=6.45 $Y2=1.985
r570 43 211 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.45 $Y=1.025
+ $X2=6.45 $Y2=1.16
r571 43 45 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.45 $Y=1.025
+ $X2=6.45 $Y2=0.56
r572 39 210 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.03 $Y=1.295
+ $X2=6.03 $Y2=1.16
r573 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.03 $Y=1.295
+ $X2=6.03 $Y2=1.985
r574 35 210 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.03 $Y=1.025
+ $X2=6.03 $Y2=1.16
r575 35 37 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.03 $Y=1.025
+ $X2=6.03 $Y2=0.56
r576 31 209 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.16
r577 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.985
r578 27 209 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=1.16
r579 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=0.56
r580 23 206 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.16
r581 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.985
r582 19 206 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=1.16
r583 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=0.56
r584 6 183 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.31
r585 6 181 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.63
r586 5 169 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2.31
r587 5 167 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=1.63
r588 4 155 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2.31
r589 4 153 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.63
r590 3 177 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.4
r591 2 163 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.4
r592 1 149 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 43
+ 45 51 55 59 63 67 69 73 77 81 85 89 93 95 99 101 103 106 107 109 110 112 113
+ 114 115 117 118 120 121 123 124 126 127 128 129 130 132 166 175 178 181 185
+ 188
r192 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r193 181 182 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r194 178 179 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r195 175 176 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r196 172 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r197 170 185 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r198 170 182 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=10.81 $Y2=2.72
r199 169 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r200 167 181 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.945 $Y=2.72
+ $X2=10.86 $Y2=2.72
r201 167 169 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.945 $Y=2.72
+ $X2=11.27 $Y2=2.72
r202 166 184 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=11.615 $Y=2.72
+ $X2=11.787 $Y2=2.72
r203 166 169 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.615 $Y=2.72
+ $X2=11.27 $Y2=2.72
r204 165 182 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r205 164 165 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r206 162 165 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r207 161 162 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r208 159 162 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r209 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r210 156 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r211 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r212 153 156 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r213 153 179 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r214 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r215 150 178 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.82 $Y2=2.72
r216 150 152 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=6.21 $Y2=2.72
r217 149 179 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r218 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r219 146 149 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r220 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r221 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r222 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r223 140 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r224 140 176 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r225 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r226 137 175 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.62 $Y2=2.72
r227 137 139 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=2.07 $Y2=2.72
r228 136 176 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r229 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r230 133 172 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r231 133 135 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r232 132 175 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=1.62 $Y2=2.72
r233 132 135 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=0.69 $Y2=2.72
r234 130 136 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r235 130 188 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r236 128 164 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=9.935 $Y=2.72
+ $X2=9.89 $Y2=2.72
r237 128 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.935 $Y=2.72
+ $X2=10.02 $Y2=2.72
r238 126 161 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.095 $Y=2.72
+ $X2=8.97 $Y2=2.72
r239 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.095 $Y=2.72
+ $X2=9.18 $Y2=2.72
r240 125 164 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=9.265 $Y=2.72
+ $X2=9.89 $Y2=2.72
r241 125 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=2.72
+ $X2=9.18 $Y2=2.72
r242 123 158 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.255 $Y=2.72
+ $X2=8.05 $Y2=2.72
r243 123 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.255 $Y=2.72
+ $X2=8.34 $Y2=2.72
r244 122 161 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.425 $Y=2.72
+ $X2=8.97 $Y2=2.72
r245 122 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=2.72
+ $X2=8.34 $Y2=2.72
r246 120 155 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.415 $Y=2.72
+ $X2=7.13 $Y2=2.72
r247 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=2.72
+ $X2=7.5 $Y2=2.72
r248 119 158 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.585 $Y=2.72
+ $X2=8.05 $Y2=2.72
r249 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=2.72
+ $X2=7.5 $Y2=2.72
r250 117 152 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.21 $Y2=2.72
r251 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.66 $Y2=2.72
r252 116 155 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.745 $Y=2.72
+ $X2=7.13 $Y2=2.72
r253 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=2.72
+ $X2=6.66 $Y2=2.72
r254 114 148 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.83 $Y2=2.72
r255 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.98 $Y2=2.72
r256 112 145 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=2.72
+ $X2=3.91 $Y2=2.72
r257 112 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2.72
+ $X2=4.14 $Y2=2.72
r258 111 148 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.83 $Y2=2.72
r259 111 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.14 $Y2=2.72
r260 109 142 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=2.99 $Y2=2.72
r261 109 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.3 $Y2=2.72
r262 108 145 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.91 $Y2=2.72
r263 108 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.3 $Y2=2.72
r264 106 139 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.07 $Y2=2.72
r265 106 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.46 $Y2=2.72
r266 105 142 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.99 $Y2=2.72
r267 105 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.46 $Y2=2.72
r268 101 184 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=11.7 $Y=2.635
+ $X2=11.787 $Y2=2.72
r269 101 103 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.7 $Y=2.635
+ $X2=11.7 $Y2=2
r270 97 181 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.86 $Y=2.635
+ $X2=10.86 $Y2=2.72
r271 97 99 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.86 $Y=2.635
+ $X2=10.86 $Y2=2
r272 96 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.105 $Y=2.72
+ $X2=10.02 $Y2=2.72
r273 95 181 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.775 $Y=2.72
+ $X2=10.86 $Y2=2.72
r274 95 96 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.775 $Y=2.72
+ $X2=10.105 $Y2=2.72
r275 91 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.02 $Y=2.635
+ $X2=10.02 $Y2=2.72
r276 91 93 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.02 $Y=2.635
+ $X2=10.02 $Y2=2
r277 87 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.18 $Y=2.635
+ $X2=9.18 $Y2=2.72
r278 87 89 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.18 $Y=2.635
+ $X2=9.18 $Y2=2
r279 83 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.34 $Y=2.635
+ $X2=8.34 $Y2=2.72
r280 83 85 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.34 $Y=2.635
+ $X2=8.34 $Y2=2
r281 79 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=2.635
+ $X2=7.5 $Y2=2.72
r282 79 81 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.5 $Y=2.635
+ $X2=7.5 $Y2=2
r283 75 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2.72
r284 75 77 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2
r285 71 178 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r286 71 73 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2
r287 70 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.98 $Y2=2.72
r288 69 178 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.82 $Y2=2.72
r289 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.065 $Y2=2.72
r290 65 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r291 65 67 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2
r292 61 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.72
r293 61 63 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2
r294 57 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2.72
r295 57 59 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2
r296 53 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.72
r297 53 55 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2
r298 49 175 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r299 49 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2
r300 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r301 43 172 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r302 43 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r303 14 103 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=11.565
+ $Y=1.485 $X2=11.7 $Y2=2
r304 13 99 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=10.725
+ $Y=1.485 $X2=10.86 $Y2=2
r305 12 93 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.885
+ $Y=1.485 $X2=10.02 $Y2=2
r306 11 89 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.045
+ $Y=1.485 $X2=9.18 $Y2=2
r307 10 85 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.205
+ $Y=1.485 $X2=8.34 $Y2=2
r308 9 81 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=2
r309 8 77 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=2
r310 7 73 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2
r311 6 67 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2
r312 5 63 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2
r313 4 59 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2
r314 3 55 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2
r315 2 51 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2
r316 1 48 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r317 1 45 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 50 53 57 58 59 60 61 62 65 69 71 73 74 77 81 83 87 91 95 97 101 105 109 111
+ 115 119 123 125 129 133 137 139 143 147 151 153 159 160 163 164 165 166 167
+ 168 169 170 171 172 173 174 176 177
c337 60 0 1.25206e-19 $X=5.565 $Y=1.53
c338 58 0 1.25206e-19 $X=5.565 $Y=0.82
r339 176 177 8.74426 $w=4.23e-07 $l=2.55e-07 $layer=LI1_cond $X=11.747 $Y=1.19
+ $X2=11.747 $Y2=1.445
r340 175 176 12.8802 $w=2.53e-07 $l=2.85e-07 $layer=LI1_cond $X=11.747 $Y=0.905
+ $X2=11.747 $Y2=1.19
r341 154 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.445 $Y=1.53
+ $X2=11.28 $Y2=1.53
r342 153 177 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.62 $Y=1.53
+ $X2=11.747 $Y2=1.53
r343 153 154 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=11.62 $Y=1.53
+ $X2=11.445 $Y2=1.53
r344 152 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.445 $Y=0.82
+ $X2=11.28 $Y2=0.82
r345 151 175 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=11.62 $Y=0.82
+ $X2=11.747 $Y2=0.905
r346 151 152 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=11.62 $Y=0.82
+ $X2=11.445 $Y2=0.82
r347 147 149 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.28 $Y=1.63
+ $X2=11.28 $Y2=2.31
r348 145 174 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.28 $Y=1.615
+ $X2=11.28 $Y2=1.53
r349 145 147 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.28 $Y=1.615
+ $X2=11.28 $Y2=1.63
r350 141 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.28 $Y=0.735
+ $X2=11.28 $Y2=0.82
r351 141 143 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.28 $Y=0.735
+ $X2=11.28 $Y2=0.4
r352 140 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.605 $Y=1.53
+ $X2=10.44 $Y2=1.53
r353 139 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.115 $Y=1.53
+ $X2=11.28 $Y2=1.53
r354 139 140 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.115 $Y=1.53
+ $X2=10.605 $Y2=1.53
r355 138 171 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.605 $Y=0.82
+ $X2=10.44 $Y2=0.82
r356 137 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.115 $Y=0.82
+ $X2=11.28 $Y2=0.82
r357 137 138 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.115 $Y=0.82
+ $X2=10.605 $Y2=0.82
r358 133 135 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.44 $Y=1.63
+ $X2=10.44 $Y2=2.31
r359 131 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.44 $Y=1.615
+ $X2=10.44 $Y2=1.53
r360 131 133 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=10.44 $Y=1.615
+ $X2=10.44 $Y2=1.63
r361 127 171 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.44 $Y=0.735
+ $X2=10.44 $Y2=0.82
r362 127 129 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.44 $Y=0.735
+ $X2=10.44 $Y2=0.4
r363 126 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.765 $Y=1.53
+ $X2=9.6 $Y2=1.53
r364 125 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.275 $Y=1.53
+ $X2=10.44 $Y2=1.53
r365 125 126 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.275 $Y=1.53
+ $X2=9.765 $Y2=1.53
r366 124 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.765 $Y=0.82
+ $X2=9.6 $Y2=0.82
r367 123 171 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.275 $Y=0.82
+ $X2=10.44 $Y2=0.82
r368 123 124 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.275 $Y=0.82
+ $X2=9.765 $Y2=0.82
r369 119 121 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.6 $Y=1.63
+ $X2=9.6 $Y2=2.31
r370 117 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.6 $Y=1.615
+ $X2=9.6 $Y2=1.53
r371 117 119 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=9.6 $Y=1.615
+ $X2=9.6 $Y2=1.63
r372 113 169 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.6 $Y=0.735
+ $X2=9.6 $Y2=0.82
r373 113 115 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.6 $Y=0.735
+ $X2=9.6 $Y2=0.4
r374 112 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=1.53
+ $X2=8.76 $Y2=1.53
r375 111 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=1.53
+ $X2=9.6 $Y2=1.53
r376 111 112 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.435 $Y=1.53
+ $X2=8.925 $Y2=1.53
r377 110 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=0.82
+ $X2=8.76 $Y2=0.82
r378 109 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=0.82
+ $X2=9.6 $Y2=0.82
r379 109 110 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.435 $Y=0.82
+ $X2=8.925 $Y2=0.82
r380 105 107 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.76 $Y=1.63
+ $X2=8.76 $Y2=2.31
r381 103 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=1.615
+ $X2=8.76 $Y2=1.53
r382 103 105 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.76 $Y=1.615
+ $X2=8.76 $Y2=1.63
r383 99 167 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=0.735
+ $X2=8.76 $Y2=0.82
r384 99 101 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.76 $Y=0.735
+ $X2=8.76 $Y2=0.4
r385 98 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=1.53
+ $X2=7.92 $Y2=1.53
r386 97 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=1.53
+ $X2=8.76 $Y2=1.53
r387 97 98 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.595 $Y=1.53
+ $X2=8.085 $Y2=1.53
r388 96 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=0.82
+ $X2=7.92 $Y2=0.82
r389 95 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=0.82
+ $X2=8.76 $Y2=0.82
r390 95 96 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.595 $Y=0.82
+ $X2=8.085 $Y2=0.82
r391 91 93 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.92 $Y=1.63
+ $X2=7.92 $Y2=2.31
r392 89 166 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=1.615
+ $X2=7.92 $Y2=1.53
r393 89 91 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.92 $Y=1.615
+ $X2=7.92 $Y2=1.63
r394 85 165 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=0.735
+ $X2=7.92 $Y2=0.82
r395 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=0.735
+ $X2=7.92 $Y2=0.4
r396 84 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=1.53
+ $X2=7.08 $Y2=1.53
r397 83 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=1.53
+ $X2=7.92 $Y2=1.53
r398 83 84 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.755 $Y=1.53
+ $X2=7.245 $Y2=1.53
r399 82 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=0.82
+ $X2=7.08 $Y2=0.82
r400 81 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=0.82
+ $X2=7.92 $Y2=0.82
r401 81 82 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.755 $Y=0.82
+ $X2=7.245 $Y2=0.82
r402 77 79 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.08 $Y=1.63
+ $X2=7.08 $Y2=2.31
r403 75 164 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=1.615
+ $X2=7.08 $Y2=1.53
r404 75 77 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.08 $Y=1.615
+ $X2=7.08 $Y2=1.63
r405 74 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=0.735
+ $X2=7.08 $Y2=0.82
r406 73 162 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=7.08 $Y=0.425
+ $X2=7.08 $Y2=0.4
r407 73 74 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=7.08 $Y=0.425
+ $X2=7.08 $Y2=0.735
r408 72 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=1.53
+ $X2=6.24 $Y2=1.53
r409 71 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=1.53
+ $X2=7.08 $Y2=1.53
r410 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.915 $Y=1.53
+ $X2=6.405 $Y2=1.53
r411 70 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0.82
+ $X2=6.24 $Y2=0.82
r412 69 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0.82
+ $X2=7.08 $Y2=0.82
r413 69 70 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.915 $Y=0.82
+ $X2=6.405 $Y2=0.82
r414 65 67 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.24 $Y=1.63
+ $X2=6.24 $Y2=2.31
r415 63 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=1.615
+ $X2=6.24 $Y2=1.53
r416 63 65 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.24 $Y=1.615
+ $X2=6.24 $Y2=1.63
r417 62 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=0.735
+ $X2=6.24 $Y2=0.82
r418 61 158 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=6.24 $Y=0.425
+ $X2=6.24 $Y2=0.4
r419 61 62 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.24 $Y=0.425
+ $X2=6.24 $Y2=0.735
r420 59 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=1.53
+ $X2=6.24 $Y2=1.53
r421 59 60 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.075 $Y=1.53
+ $X2=5.565 $Y2=1.53
r422 57 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0.82
+ $X2=6.24 $Y2=0.82
r423 57 58 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.075 $Y=0.82
+ $X2=5.565 $Y2=0.82
r424 53 55 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.4 $Y=1.63 $X2=5.4
+ $Y2=2.31
r425 51 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.4 $Y=1.615
+ $X2=5.565 $Y2=1.53
r426 51 53 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.4 $Y=1.615
+ $X2=5.4 $Y2=1.63
r427 50 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.4 $Y=0.735
+ $X2=5.565 $Y2=0.82
r428 49 156 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=5.4 $Y=0.425
+ $X2=5.4 $Y2=0.4
r429 49 50 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=5.4 $Y=0.425 $X2=5.4
+ $Y2=0.735
r430 16 149 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=11.145
+ $Y=1.485 $X2=11.28 $Y2=2.31
r431 16 147 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.145
+ $Y=1.485 $X2=11.28 $Y2=1.63
r432 15 135 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=10.305
+ $Y=1.485 $X2=10.44 $Y2=2.31
r433 15 133 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.305
+ $Y=1.485 $X2=10.44 $Y2=1.63
r434 14 121 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.465
+ $Y=1.485 $X2=9.6 $Y2=2.31
r435 14 119 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.465
+ $Y=1.485 $X2=9.6 $Y2=1.63
r436 13 107 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.485 $X2=8.76 $Y2=2.31
r437 13 105 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.485 $X2=8.76 $Y2=1.63
r438 12 93 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=7.785
+ $Y=1.485 $X2=7.92 $Y2=2.31
r439 12 91 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.785
+ $Y=1.485 $X2=7.92 $Y2=1.63
r440 11 79 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=2.31
r441 11 77 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=1.63
r442 10 67 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=2.31
r443 10 65 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.63
r444 9 55 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=2.31
r445 9 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.63
r446 8 143 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=11.145
+ $Y=0.235 $X2=11.28 $Y2=0.4
r447 7 129 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=10.305
+ $Y=0.235 $X2=10.44 $Y2=0.4
r448 6 115 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=9.465
+ $Y=0.235 $X2=9.6 $Y2=0.4
r449 5 101 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.625
+ $Y=0.235 $X2=8.76 $Y2=0.4
r450 4 87 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=7.785
+ $Y=0.235 $X2=7.92 $Y2=0.4
r451 3 162 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.4
r452 2 158 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.4
r453 1 156 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 43
+ 45 49 53 57 61 65 67 71 75 79 83 87 91 93 97 99 101 104 105 107 108 110 111
+ 112 113 115 116 118 119 121 122 124 125 126 127 128 130 164 173 176 179 183
+ 186
r226 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r227 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r228 176 177 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r229 173 174 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r230 170 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r231 168 183 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r232 168 180 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=10.81 $Y2=0
r233 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r234 165 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.945 $Y=0
+ $X2=10.86 $Y2=0
r235 165 167 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.945 $Y=0
+ $X2=11.27 $Y2=0
r236 164 182 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=11.615 $Y=0
+ $X2=11.787 $Y2=0
r237 164 167 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.615 $Y=0
+ $X2=11.27 $Y2=0
r238 163 180 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r239 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r240 160 163 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r241 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r242 157 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r243 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r244 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r245 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r246 151 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r247 151 177 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r248 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r249 148 176 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=5.82 $Y2=0
r250 148 150 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.21 $Y2=0
r251 147 177 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r252 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r253 144 147 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r254 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r255 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r256 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r257 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r258 138 174 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r259 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r260 135 173 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=1.62 $Y2=0
r261 135 137 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r262 134 174 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r263 133 134 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r264 131 170 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r265 131 133 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.69 $Y2=0
r266 130 173 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=1.62 $Y2=0
r267 130 133 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=0.69 $Y2=0
r268 128 134 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r269 128 186 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r270 126 162 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=9.935 $Y=0
+ $X2=9.89 $Y2=0
r271 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.935 $Y=0
+ $X2=10.02 $Y2=0
r272 124 159 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=8.97 $Y2=0
r273 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=9.18 $Y2=0
r274 123 162 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=9.265 $Y=0
+ $X2=9.89 $Y2=0
r275 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=0
+ $X2=9.18 $Y2=0
r276 121 156 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.255 $Y=0
+ $X2=8.05 $Y2=0
r277 121 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.255 $Y=0
+ $X2=8.34 $Y2=0
r278 120 159 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.425 $Y=0
+ $X2=8.97 $Y2=0
r279 120 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=0
+ $X2=8.34 $Y2=0
r280 118 153 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.415 $Y=0
+ $X2=7.13 $Y2=0
r281 118 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=0 $X2=7.5
+ $Y2=0
r282 117 156 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.585 $Y=0
+ $X2=8.05 $Y2=0
r283 117 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.5
+ $Y2=0
r284 115 150 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.21 $Y2=0
r285 115 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.66 $Y2=0
r286 114 153 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.13 $Y2=0
r287 114 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.66 $Y2=0
r288 112 146 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.83 $Y2=0
r289 112 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.98 $Y2=0
r290 110 143 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=0
+ $X2=3.91 $Y2=0
r291 110 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0
+ $X2=4.14 $Y2=0
r292 109 146 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.83 $Y2=0
r293 109 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.14 $Y2=0
r294 107 140 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=0
+ $X2=2.99 $Y2=0
r295 107 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.3
+ $Y2=0
r296 106 143 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=3.91 $Y2=0
r297 106 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.3
+ $Y2=0
r298 104 137 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.07 $Y2=0
r299 104 105 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.46 $Y2=0
r300 103 140 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=0
+ $X2=2.99 $Y2=0
r301 103 105 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0
+ $X2=2.46 $Y2=0
r302 99 182 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=11.7 $Y=0.085
+ $X2=11.787 $Y2=0
r303 99 101 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.7 $Y=0.085
+ $X2=11.7 $Y2=0.4
r304 95 179 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.86 $Y=0.085
+ $X2=10.86 $Y2=0
r305 95 97 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.86 $Y=0.085
+ $X2=10.86 $Y2=0.4
r306 94 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.105 $Y=0
+ $X2=10.02 $Y2=0
r307 93 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.775 $Y=0
+ $X2=10.86 $Y2=0
r308 93 94 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.775 $Y=0
+ $X2=10.105 $Y2=0
r309 89 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.02 $Y=0.085
+ $X2=10.02 $Y2=0
r310 89 91 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.02 $Y=0.085
+ $X2=10.02 $Y2=0.4
r311 85 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.18 $Y=0.085
+ $X2=9.18 $Y2=0
r312 85 87 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.18 $Y=0.085
+ $X2=9.18 $Y2=0.4
r313 81 122 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.34 $Y=0.085
+ $X2=8.34 $Y2=0
r314 81 83 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.34 $Y=0.085
+ $X2=8.34 $Y2=0.4
r315 77 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0
r316 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.4
r317 73 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0
r318 73 75 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0.4
r319 69 176 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r320 69 71 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.4
r321 68 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r322 67 176 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.82
+ $Y2=0
r323 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.065 $Y2=0
r324 63 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r325 63 65 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.4
r326 59 111 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r327 59 61 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.4
r328 55 108 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0
r329 55 57 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.4
r330 51 105 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r331 51 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.4
r332 47 173 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r333 47 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.4
r334 43 170 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r335 43 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r336 14 101 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=11.565
+ $Y=0.235 $X2=11.7 $Y2=0.4
r337 13 97 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=10.725
+ $Y=0.235 $X2=10.86 $Y2=0.4
r338 12 91 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.885
+ $Y=0.235 $X2=10.02 $Y2=0.4
r339 11 87 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.045
+ $Y=0.235 $X2=9.18 $Y2=0.4
r340 10 83 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.205
+ $Y=0.235 $X2=8.34 $Y2=0.4
r341 9 79 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.4
r342 8 75 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.4
r343 7 71 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.4
r344 6 65 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.4
r345 5 61 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.4
r346 4 57 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.4
r347 3 53 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.4
r348 2 49 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.4
r349 1 45 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__nor4b_2.pex.spice
* Created: Thu Aug 27 14:33:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4B_2%A 1 3 6 8 10 13 15 16 17 26
c44 26 0 1.30704e-19 $X=0.89 $Y=1.16
r45 24 26 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.625 $Y=1.16
+ $X2=0.89 $Y2=1.16
r46 21 24 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.625 $Y2=1.16
r47 16 17 26.9351 $w=2.08e-07 $l=5.1e-07 $layer=LI1_cond $X=0.625 $Y=1.18
+ $X2=1.135 $Y2=1.18
r48 16 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.16 $X2=0.625 $Y2=1.16
r49 15 16 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.215 $Y=1.18
+ $X2=0.625 $Y2=1.18
r50 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r52 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r54 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r56 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%B 1 3 6 8 10 13 15 16 17 26
c43 17 0 1.30704e-19 $X=2.445 $Y=1.105
r44 24 26 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.73 $Y2=1.16
r45 21 24 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.585 $Y2=1.16
r46 16 17 25.0866 $w=2.08e-07 $l=4.75e-07 $layer=LI1_cond $X=2.055 $Y=1.18
+ $X2=2.53 $Y2=1.18
r47 15 16 24.8225 $w=2.08e-07 $l=4.7e-07 $layer=LI1_cond $X=1.585 $Y=1.18
+ $X2=2.055 $Y2=1.18
r48 15 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.16 $X2=1.585 $Y2=1.16
r49 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r50 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r51 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r52 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r53 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r54 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r55 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%C 1 3 6 8 10 13 15 16 24
c45 24 0 3.0059e-19 $X=3.125 $Y=1.16
r46 22 24 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=2.98 $Y=1.16
+ $X2=3.125 $Y2=1.16
r47 19 22 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.705 $Y=1.16
+ $X2=2.98 $Y2=1.16
r48 15 16 24.8225 $w=2.08e-07 $l=4.7e-07 $layer=LI1_cond $X=2.98 $Y=1.18
+ $X2=3.45 $Y2=1.18
r49 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r50 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.325
+ $X2=3.125 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.125 $Y=1.325
+ $X2=3.125 $Y2=1.985
r52 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=0.995
+ $X2=3.125 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.125 $Y=0.995
+ $X2=3.125 $Y2=0.56
r54 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.325
+ $X2=2.705 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.705 $Y=1.325
+ $X2=2.705 $Y2=1.985
r56 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%A_694_21# 1 2 7 9 12 14 16 19 21 26 30 31 35
+ 39 40
c71 21 0 3.09582e-19 $X=4.04 $Y=1.16
r72 39 40 11.2584 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=4.642 $Y=2.285
+ $X2=4.642 $Y2=2.035
r73 35 37 11.0961 $w=3.53e-07 $l=2.45e-07 $layer=LI1_cond $X=4.642 $Y=0.66
+ $X2=4.642 $Y2=0.905
r74 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.485
+ $Y=1.16 $X2=4.485 $Y2=1.16
r75 27 30 0.716491 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.55 $Y=1.245
+ $X2=4.485 $Y2=1.16
r76 27 40 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.55 $Y=1.245
+ $X2=4.55 $Y2=2.035
r77 26 30 0.716491 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.55 $Y=1.075
+ $X2=4.485 $Y2=1.16
r78 26 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.55 $Y=1.075
+ $X2=4.55 $Y2=0.905
r79 22 24 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.545 $Y=1.16
+ $X2=3.965 $Y2=1.16
r80 21 31 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.04 $Y=1.16
+ $X2=4.485 $Y2=1.16
r81 21 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=1.16
+ $X2=3.965 $Y2=1.16
r82 17 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.325
+ $X2=3.965 $Y2=1.16
r83 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.965 $Y=1.325
+ $X2=3.965 $Y2=1.985
r84 14 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=0.995
+ $X2=3.965 $Y2=1.16
r85 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.965 $Y=0.995
+ $X2=3.965 $Y2=0.56
r86 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=1.325
+ $X2=3.545 $Y2=1.16
r87 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.545 $Y=1.325
+ $X2=3.545 $Y2=1.985
r88 7 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=0.995
+ $X2=3.545 $Y2=1.16
r89 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.545 $Y=0.995
+ $X2=3.545 $Y2=0.56
r90 2 39 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=4.57
+ $Y=2.065 $X2=4.695 $Y2=2.285
r91 1 35 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.465 $X2=4.695 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%D_N 3 6 8 11 13 14 15 20 22
r31 14 15 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.31 $Y=1.53
+ $X2=5.31 $Y2=1.87
r32 14 22 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=5.31 $Y=1.53
+ $X2=5.31 $Y2=1.285
r33 13 22 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.31 $Y=1.18
+ $X2=5.31 $Y2=1.285
r34 11 21 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.967 $Y=1.16
+ $X2=4.967 $Y2=1.325
r35 11 20 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.967 $Y=1.16
+ $X2=4.967 $Y2=0.995
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.97
+ $Y=1.16 $X2=4.97 $Y2=1.16
r37 8 13 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=1.18
+ $X2=5.31 $Y2=1.18
r38 8 10 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=5.185 $Y=1.18
+ $X2=4.97 $Y2=1.18
r39 6 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.905 $Y=2.275
+ $X2=4.905 $Y2=1.325
r40 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.905 $Y=0.675
+ $X2=4.905 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%A_27_297# 1 2 3 12 16 17 20 22 26 29
r42 24 26 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.94 $Y=1.625
+ $X2=1.94 $Y2=1.63
r43 23 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=1.54
+ $X2=1.1 $Y2=1.54
r44 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.775 $Y=1.54
+ $X2=1.94 $Y2=1.625
r45 22 23 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.775 $Y=1.54
+ $X2=1.225 $Y2=1.54
r46 18 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.625
+ $X2=1.1 $Y2=1.54
r47 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.1 $Y=1.625 $X2=1.1
+ $Y2=2.3
r48 16 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=1.54
+ $X2=1.1 $Y2=1.54
r49 16 17 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=1.54
+ $X2=0.425 $Y2=1.54
r50 12 14 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.63
+ $X2=0.255 $Y2=2.31
r51 10 17 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.425 $Y2=1.54
r52 10 12 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.255 $Y2=1.63
r53 3 26 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.63
r54 2 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.62
r55 2 20 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.3
r56 1 14 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r57 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%VPWR 1 2 9 13 15 16 17 18 20 34 36
r58 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r60 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r61 30 31 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r62 28 31 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r63 28 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 27 30 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r65 27 28 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 25 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=0.7 $Y2=2.72
r67 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 20 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.7 $Y2=2.72
r69 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 16 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r73 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.99 $Y=2.72
+ $X2=5.115 $Y2=2.72
r74 15 33 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=5.24 $Y=2.72 $X2=5.29
+ $Y2=2.72
r75 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.24 $Y=2.72
+ $X2=5.115 $Y2=2.72
r76 11 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=2.635
+ $X2=5.115 $Y2=2.72
r77 11 13 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.115 $Y=2.635
+ $X2=5.115 $Y2=2.3
r78 7 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r79 7 9 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r80 2 13 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=2.065 $X2=5.115 $Y2=2.3
r81 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%A_277_297# 1 2 9 11 12 15
r19 13 15 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.935 $Y=2.295
+ $X2=2.935 $Y2=1.96
r20 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.83 $Y=2.38
+ $X2=2.935 $Y2=2.295
r21 11 12 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=2.83 $Y=2.38
+ $X2=1.605 $Y2=2.38
r22 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.5 $Y=2.295
+ $X2=1.605 $Y2=2.38
r23 7 9 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=1.5 $Y=2.295 $X2=1.5
+ $Y2=1.96
r24 2 15 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=1.485 $X2=2.915 $Y2=1.96
r25 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%A_474_297# 1 2 3 12 14 15 16 17 18 22
r41 20 22 15.7579 $w=2.43e-07 $l=3.35e-07 $layer=LI1_cond $X=4.172 $Y=2.295
+ $X2=4.172 $Y2=1.96
r42 19 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.46 $Y=2.38
+ $X2=3.335 $Y2=2.38
r43 18 20 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=4.05 $Y=2.38
+ $X2=4.172 $Y2=2.295
r44 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.05 $Y=2.38 $X2=3.46
+ $Y2=2.38
r45 17 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=2.295
+ $X2=3.335 $Y2=2.38
r46 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.625
+ $X2=3.335 $Y2=1.54
r47 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.335 $Y=1.625
+ $X2=3.335 $Y2=2.295
r48 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.21 $Y=1.54
+ $X2=3.335 $Y2=1.54
r49 14 15 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.21 $Y=1.54
+ $X2=2.66 $Y2=1.54
r50 10 15 8.24022 $w=1.7e-07 $l=2.31633e-07 $layer=LI1_cond $X=2.467 $Y=1.625
+ $X2=2.66 $Y2=1.54
r51 10 12 0.149668 $w=3.83e-07 $l=5e-09 $layer=LI1_cond $X=2.467 $Y=1.625
+ $X2=2.467 $Y2=1.63
r52 3 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.04
+ $Y=1.485 $X2=4.175 $Y2=1.96
r53 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.485 $X2=3.335 $Y2=2.3
r54 2 25 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.485 $X2=3.335 $Y2=1.62
r55 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.37
+ $Y=1.485 $X2=2.495 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%Y 1 2 3 4 5 18 20 21 24 26 30 32 36 42 43 44
+ 45 46 56 58 62
c99 58 0 1.50811e-19 $X=3.91 $Y=1.53
c100 45 0 3.0059e-19 $X=3.825 $Y=1.105
c101 44 0 1.58772e-19 $X=3.755 $Y=0.815
r102 58 59 2.67406 $w=4.03e-07 $l=7.5e-08 $layer=LI1_cond $X=3.832 $Y=1.53
+ $X2=3.832 $Y2=1.455
r103 46 62 2.41871 $w=4.03e-07 $l=8.5e-08 $layer=LI1_cond $X=3.832 $Y=1.535
+ $X2=3.832 $Y2=1.62
r104 46 58 0.142277 $w=4.03e-07 $l=5e-09 $layer=LI1_cond $X=3.832 $Y=1.535
+ $X2=3.832 $Y2=1.53
r105 46 59 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=3.875 $Y=1.45
+ $X2=3.875 $Y2=1.455
r106 45 51 2.3409 $w=3.18e-07 $l=6.5e-08 $layer=LI1_cond $X=3.875 $Y=1.17
+ $X2=3.875 $Y2=1.235
r107 45 56 4.90503 $w=3.18e-07 $l=9.5e-08 $layer=LI1_cond $X=3.875 $Y=1.17
+ $X2=3.875 $Y2=1.075
r108 45 46 7.0227 $w=3.18e-07 $l=1.95e-07 $layer=LI1_cond $X=3.875 $Y=1.255
+ $X2=3.875 $Y2=1.45
r109 45 51 0.720277 $w=3.18e-07 $l=2e-08 $layer=LI1_cond $X=3.875 $Y=1.255
+ $X2=3.875 $Y2=1.235
r110 40 44 3.67302 $w=2.67e-07 $l=1.16962e-07 $layer=LI1_cond $X=3.817 $Y=0.905
+ $X2=3.755 $Y2=0.815
r111 40 56 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=3.817 $Y=0.905
+ $X2=3.817 $Y2=1.075
r112 34 44 3.67302 $w=2.67e-07 $l=9e-08 $layer=LI1_cond $X=3.755 $Y=0.725
+ $X2=3.755 $Y2=0.815
r113 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.755 $Y=0.725
+ $X2=3.755 $Y2=0.39
r114 33 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0.815
+ $X2=2.915 $Y2=0.815
r115 32 44 2.80098 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=0.815
+ $X2=3.755 $Y2=0.815
r116 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.59 $Y=0.815
+ $X2=3.08 $Y2=0.815
r117 28 43 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.915 $Y=0.725
+ $X2=2.915 $Y2=0.815
r118 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.915 $Y=0.725
+ $X2=2.915 $Y2=0.39
r119 27 42 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0.815
+ $X2=1.52 $Y2=0.815
r120 26 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0.815
+ $X2=2.915 $Y2=0.815
r121 26 27 65.6212 $w=1.78e-07 $l=1.065e-06 $layer=LI1_cond $X=2.75 $Y=0.815
+ $X2=1.685 $Y2=0.815
r122 22 42 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.52 $Y=0.725
+ $X2=1.52 $Y2=0.815
r123 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=0.725
+ $X2=1.52 $Y2=0.39
r124 20 42 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=1.52 $Y2=0.815
r125 20 21 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=0.845 $Y2=0.815
r126 16 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.845 $Y2=0.815
r127 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.68 $Y2=0.39
r128 5 62 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.62
+ $Y=1.485 $X2=3.755 $Y2=1.62
r129 4 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.62
+ $Y=0.235 $X2=3.755 $Y2=0.39
r130 3 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.78
+ $Y=0.235 $X2=2.915 $Y2=0.39
r131 2 24 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r132 1 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_2%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 43 44
+ 46 47 49 50 51 52 53 54 76 82 88
r86 87 88 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.235
+ $X2=2.58 $Y2=0.235
r87 84 87 7.94271 $w=6.38e-07 $l=4.25e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.495 $Y2=0.235
r88 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r89 81 84 2.42953 $w=6.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.94 $Y=0.235
+ $X2=2.07 $Y2=0.235
r90 81 82 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.235
+ $X2=1.855 $Y2=0.235
r91 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r92 73 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r93 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r94 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r95 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r96 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r97 67 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r98 66 88 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.58
+ $Y2=0
r99 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r100 63 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r101 62 82 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.855
+ $Y2=0
r102 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r103 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r104 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r105 56 78 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r106 56 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r107 54 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r108 54 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r109 52 72 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.99 $Y=0 $X2=4.83
+ $Y2=0
r110 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.99 $Y=0 $X2=5.115
+ $Y2=0
r111 51 75 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=5.24 $Y=0 $X2=5.29
+ $Y2=0
r112 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.24 $Y=0 $X2=5.115
+ $Y2=0
r113 49 69 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.91
+ $Y2=0
r114 49 50 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.192
+ $Y2=0
r115 48 72 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.83 $Y2=0
r116 48 50 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.192 $Y2=0
r117 46 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=2.99
+ $Y2=0
r118 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.335
+ $Y2=0
r119 45 69 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.91
+ $Y2=0
r120 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.335
+ $Y2=0
r121 43 58 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r122 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r123 42 62 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r124 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r125 38 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0
r126 38 40 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0.66
r127 34 50 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.192 $Y=0.085
+ $X2=4.192 $Y2=0
r128 34 36 16.5011 $w=2.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.192 $Y=0.085
+ $X2=4.192 $Y2=0.39
r129 30 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0
r130 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0.39
r131 26 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r132 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.39
r133 22 78 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r134 22 24 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.39
r135 7 40 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=4.98
+ $Y=0.465 $X2=5.115 $Y2=0.66
r136 6 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.04
+ $Y=0.235 $X2=4.175 $Y2=0.39
r137 5 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.235 $X2=3.335 $Y2=0.39
r138 4 87 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.37
+ $Y=0.235 $X2=2.495 $Y2=0.39
r139 3 81 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r140 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r141 1 24 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__nor3b_4.spice.pex
* Created: Thu Aug 27 14:32:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR3B_4%C_N 1 3 6 8 14 17
c26 1 0 1.59348e-19 $X=0.49 $Y=0.995
r27 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.49 $Y2=1.16
r28 8 17 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.18 $X2=0.23
+ $Y2=1.18
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r30 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r31 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r32 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r33 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 45
r73 43 45 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=2.17 $Y2=1.16
r74 41 43 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.75 $Y=1.16
+ $X2=2.02 $Y2=1.16
r75 39 41 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.34 $Y=1.16
+ $X2=1.75 $Y2=1.16
r76 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.16 $X2=1.34 $Y2=1.16
r77 37 39 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.33 $Y=1.16 $X2=1.34
+ $Y2=1.16
r78 35 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r79 30 31 27.1991 $w=2.08e-07 $l=5.15e-07 $layer=LI1_cond $X=2.02 $Y=1.18
+ $X2=2.535 $Y2=1.18
r80 30 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.02
+ $Y=1.16 $X2=2.02 $Y2=1.16
r81 29 30 21.3896 $w=2.08e-07 $l=4.05e-07 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=2.02 $Y2=1.18
r82 29 40 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=1.34 $Y2=1.18
r83 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r85 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
r87 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r89 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r91 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r93 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r95 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325 $X2=0.91
+ $Y2=1.985
r97 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995 $X2=0.91
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 39 41
c75 39 0 1.61212e-19 $X=3.88 $Y=1.16
r76 40 41 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.95 $Y=1.16
+ $X2=4.37 $Y2=1.16
r77 38 40 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.88 $Y=1.16 $X2=3.95
+ $Y2=1.16
r78 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r79 36 38 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.53 $Y=1.16
+ $X2=3.88 $Y2=1.16
r80 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.2 $Y=1.16 $X2=3.53
+ $Y2=1.16
r81 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.16 $X2=3.2 $Y2=1.16
r82 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.11 $Y=1.16 $X2=3.2
+ $Y2=1.16
r83 29 39 21.3896 $w=2.08e-07 $l=4.05e-07 $layer=LI1_cond $X=3.475 $Y=1.18
+ $X2=3.88 $Y2=1.18
r84 29 35 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.475 $Y=1.18
+ $X2=3.2 $Y2=1.18
r85 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.16
r86 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.985
r87 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=1.16
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=0.56
r89 18 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.325
+ $X2=3.95 $Y2=1.16
r90 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.95 $Y=1.325
+ $X2=3.95 $Y2=1.985
r91 15 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=1.16
r92 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=0.56
r93 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.985
r95 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=0.56
r97 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r98 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325 $X2=3.11
+ $Y2=1.985
r99 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=1.16
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 39 41 43 46 47 50 51 56 61 65 72
c157 72 0 1.61212e-19 $X=6.05 $Y=1.16
r158 69 70 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.21 $Y=1.16
+ $X2=5.63 $Y2=1.16
r159 57 72 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.9 $Y=1.16
+ $X2=6.05 $Y2=1.16
r160 57 70 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.9 $Y=1.16
+ $X2=5.63 $Y2=1.16
r161 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.9
+ $Y=1.16 $X2=5.9 $Y2=1.16
r162 54 69 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.88 $Y=1.16
+ $X2=5.21 $Y2=1.16
r163 54 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.88 $Y=1.16 $X2=4.79
+ $Y2=1.16
r164 53 56 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=4.88 $Y=1.18
+ $X2=5.9 $Y2=1.18
r165 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.88
+ $Y=1.16 $X2=4.88 $Y2=1.16
r166 51 53 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=4.705 $Y=1.18
+ $X2=4.88 $Y2=1.18
r167 49 51 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.62 $Y=1.285
+ $X2=4.705 $Y2=1.18
r168 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.62 $Y=1.285
+ $X2=4.62 $Y2=1.455
r169 48 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=1.54
+ $X2=0.7 $Y2=1.54
r170 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.535 $Y=1.54
+ $X2=4.62 $Y2=1.455
r171 47 48 244.652 $w=1.68e-07 $l=3.75e-06 $layer=LI1_cond $X=4.535 $Y=1.54
+ $X2=0.785 $Y2=1.54
r172 46 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.455 $X2=0.7
+ $Y2=1.54
r173 45 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.905
+ $X2=0.7 $Y2=0.82
r174 45 46 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.7 $Y=0.905
+ $X2=0.7 $Y2=1.455
r175 44 64 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.257 $Y2=1.54
r176 43 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.615 $Y=1.54
+ $X2=0.7 $Y2=1.54
r177 43 44 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.615 $Y=1.54
+ $X2=0.405 $Y2=1.54
r178 39 64 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=1.625
+ $X2=0.257 $Y2=1.54
r179 39 41 26.3695 $w=2.93e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=1.625
+ $X2=0.257 $Y2=2.3
r180 35 61 27.5968 $w=1.68e-07 $l=4.23e-07 $layer=LI1_cond $X=0.277 $Y=0.82
+ $X2=0.7 $Y2=0.82
r181 35 37 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=0.277 $Y=0.735
+ $X2=0.277 $Y2=0.39
r182 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=1.325
+ $X2=6.05 $Y2=1.16
r183 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.05 $Y=1.325
+ $X2=6.05 $Y2=1.985
r184 28 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=0.995
+ $X2=6.05 $Y2=1.16
r185 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.05 $Y=0.995
+ $X2=6.05 $Y2=0.56
r186 24 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.16
r187 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.985
r188 21 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=1.16
r189 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=0.56
r190 17 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.16
r191 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.985
r192 14 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=1.16
r193 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=0.56
r194 10 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.16
r195 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.985
r196 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=1.16
r197 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=0.56
r198 2 64 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r199 2 41 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r200 1 37 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r96 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r97 46 47 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r98 44 47 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=2.53 $Y=2.72 $X2=6.67
+ $Y2=2.72
r99 43 46 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=6.67 $Y2=2.72
r100 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r101 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r102 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r103 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r104 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 35 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r107 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r108 30 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r109 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r110 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r112 26 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.07 $Y2=2.72
r113 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.38 $Y2=2.72
r114 25 43 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.53 $Y2=2.72
r115 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.38 $Y2=2.72
r116 23 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.54 $Y2=2.72
r118 22 40 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.54 $Y2=2.72
r120 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2.72
r121 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2.3
r122 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.72
r123 14 16 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.3
r124 10 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r125 10 12 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=1.96
r126 3 20 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=2.3
r127 2 16 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2.3
r128 1 12 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%A_197_297# 1 2 3 4 15 19 21 24 26 27 32
r48 32 35 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.16 $Y=1.88 $X2=4.16
+ $Y2=1.96
r49 27 30 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.32 $Y=1.88 $X2=3.32
+ $Y2=1.96
r50 22 27 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=1.88
+ $X2=3.32 $Y2=1.88
r51 21 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=1.88
+ $X2=4.16 $Y2=1.88
r52 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.035 $Y=1.88
+ $X2=3.445 $Y2=1.88
r53 20 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=1.88
+ $X2=1.96 $Y2=1.88
r54 19 27 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.195 $Y=1.88
+ $X2=3.32 $Y2=1.88
r55 19 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.195 $Y=1.88
+ $X2=2.085 $Y2=1.88
r56 16 24 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.88
+ $X2=1.12 $Y2=1.88
r57 15 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.88
+ $X2=1.96 $Y2=1.88
r58 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.88
+ $X2=1.245 $Y2=1.88
r59 4 35 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.485 $X2=4.16 $Y2=1.96
r60 3 30 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=1.96
r61 2 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.96
r62 1 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%A_555_297# 1 2 3 4 5 16 18 22 24 28 30 34 37
+ 42 46 47
r60 42 44 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.74 $Y=2.3 $X2=3.74
+ $Y2=2.38
r61 37 39 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.9 $Y=2.3 $X2=2.9
+ $Y2=2.38
r62 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.26 $Y=2.295
+ $X2=6.26 $Y2=1.96
r63 31 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=2.38
+ $X2=5.42 $Y2=2.38
r64 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.135 $Y=2.38
+ $X2=6.26 $Y2=2.295
r65 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.135 $Y=2.38
+ $X2=5.545 $Y2=2.38
r66 26 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=2.295
+ $X2=5.42 $Y2=2.38
r67 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.42 $Y=2.295
+ $X2=5.42 $Y2=1.96
r68 25 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.705 $Y=2.38
+ $X2=4.58 $Y2=2.38
r69 24 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=2.38
+ $X2=5.42 $Y2=2.38
r70 24 25 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.295 $Y=2.38
+ $X2=4.705 $Y2=2.38
r71 20 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=2.295
+ $X2=4.58 $Y2=2.38
r72 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.58 $Y=2.295
+ $X2=4.58 $Y2=1.96
r73 19 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.865 $Y=2.38
+ $X2=3.74 $Y2=2.38
r74 18 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.455 $Y=2.38
+ $X2=4.58 $Y2=2.38
r75 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.455 $Y=2.38
+ $X2=3.865 $Y2=2.38
r76 17 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.025 $Y=2.38
+ $X2=2.9 $Y2=2.38
r77 16 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.615 $Y=2.38
+ $X2=3.74 $Y2=2.38
r78 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.615 $Y=2.38
+ $X2=3.025 $Y2=2.38
r79 5 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.125
+ $Y=1.485 $X2=6.26 $Y2=1.96
r80 4 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.485 $X2=5.42 $Y2=1.96
r81 3 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=1.485 $X2=4.58 $Y2=1.96
r82 2 42 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.485 $X2=3.74 $Y2=2.3
r83 1 37 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.485 $X2=2.9 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 41 45 47
+ 51 55 57 61 65 67 70 73 74 75 76 78 79 81 82 84 85
c180 30 0 1.59348e-19 $X=1.285 $Y=0.815
r181 83 85 14.5805 $w=2.05e-07 $l=2.45e-07 $layer=LI1_cond $X=6.657 $Y=1.625
+ $X2=6.657 $Y2=1.87
r182 83 84 3.43356 $w=2.72e-07 $l=1.13666e-07 $layer=LI1_cond $X=6.657 $Y=1.625
+ $X2=6.59 $Y2=1.54
r183 70 84 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=1.455
+ $X2=6.59 $Y2=1.54
r184 69 82 3.39178 $w=2.92e-07 $l=9e-08 $layer=LI1_cond $X=6.59 $Y=0.905
+ $X2=6.59 $Y2=0.815
r185 69 70 18.6425 $w=3.38e-07 $l=5.5e-07 $layer=LI1_cond $X=6.59 $Y=0.905
+ $X2=6.59 $Y2=1.455
r186 68 79 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.005 $Y=0.815
+ $X2=5.84 $Y2=0.815
r187 67 82 3.13665 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=6.42 $Y=0.815
+ $X2=6.59 $Y2=0.815
r188 67 68 25.5707 $w=1.78e-07 $l=4.15e-07 $layer=LI1_cond $X=6.42 $Y=0.815
+ $X2=6.005 $Y2=0.815
r189 66 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.965 $Y=1.54
+ $X2=5.84 $Y2=1.54
r190 65 84 3.08518 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.42 $Y=1.54
+ $X2=6.59 $Y2=1.54
r191 65 66 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.42 $Y=1.54
+ $X2=5.965 $Y2=1.54
r192 59 79 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.84 $Y=0.725
+ $X2=5.84 $Y2=0.815
r193 59 61 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.84 $Y=0.725
+ $X2=5.84 $Y2=0.39
r194 58 76 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0.815
+ $X2=5 $Y2=0.815
r195 57 79 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=0.815
+ $X2=5.84 $Y2=0.815
r196 57 58 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.675 $Y=0.815
+ $X2=5.165 $Y2=0.815
r197 56 78 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.125 $Y=1.54 $X2=5
+ $Y2=1.54
r198 55 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.715 $Y=1.54
+ $X2=5.84 $Y2=1.54
r199 55 56 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.715 $Y=1.54
+ $X2=5.125 $Y2=1.54
r200 49 76 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5 $Y=0.725 $X2=5
+ $Y2=0.815
r201 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5 $Y=0.725 $X2=5
+ $Y2=0.39
r202 48 75 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0.815
+ $X2=4.16 $Y2=0.815
r203 47 76 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.815
+ $X2=5 $Y2=0.815
r204 47 48 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.835 $Y=0.815
+ $X2=4.325 $Y2=0.815
r205 43 75 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.16 $Y=0.725
+ $X2=4.16 $Y2=0.815
r206 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.16 $Y=0.725
+ $X2=4.16 $Y2=0.39
r207 42 74 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=0.815
+ $X2=3.32 $Y2=0.815
r208 41 75 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0.815
+ $X2=4.16 $Y2=0.815
r209 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.995 $Y=0.815
+ $X2=3.485 $Y2=0.815
r210 37 74 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.32 $Y=0.725
+ $X2=3.32 $Y2=0.815
r211 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.32 $Y=0.725
+ $X2=3.32 $Y2=0.39
r212 36 73 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0.815
+ $X2=1.96 $Y2=0.815
r213 35 74 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0.815
+ $X2=3.32 $Y2=0.815
r214 35 36 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=3.155 $Y=0.815
+ $X2=2.125 $Y2=0.815
r215 31 73 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.96 $Y=0.725
+ $X2=1.96 $Y2=0.815
r216 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.96 $Y=0.725
+ $X2=1.96 $Y2=0.39
r217 29 73 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0.815
+ $X2=1.96 $Y2=0.815
r218 29 30 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.795 $Y=0.815
+ $X2=1.285 $Y2=0.815
r219 25 30 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.12 $Y=0.725
+ $X2=1.285 $Y2=0.815
r220 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.12 $Y=0.725
+ $X2=1.12 $Y2=0.39
r221 8 81 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.705
+ $Y=1.485 $X2=5.84 $Y2=1.62
r222 7 78 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5 $Y2=1.62
r223 6 61 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.705
+ $Y=0.235 $X2=5.84 $Y2=0.39
r224 5 51 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.39
r225 4 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.39
r226 3 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.185
+ $Y=0.235 $X2=3.32 $Y2=0.39
r227 2 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r228 1 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_4%VGND 1 2 3 4 5 6 7 26 30 34 38 42 44 48 51
+ 52 54 55 57 58 59 60 61 83 84 87 92 95 97 100
r118 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r119 94 95 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.235
+ $X2=2.985 $Y2=0.235
r120 90 94 6.91483 $w=6.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.9 $Y2=0.235
r121 90 92 11.7251 $w=6.38e-07 $l=2.35e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.295 $Y2=0.235
r122 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r123 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r124 84 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r125 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r126 81 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.345 $Y=0 $X2=6.26
+ $Y2=0
r127 81 83 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.345 $Y=0
+ $X2=6.67 $Y2=0
r128 80 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r129 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r130 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r131 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r132 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r133 74 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r134 73 95 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=2.985 $Y2=0
r135 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r136 70 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r137 69 92 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.07 $Y=0
+ $X2=2.295 $Y2=0
r138 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r139 66 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r140 66 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r141 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r142 63 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r143 63 65 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=0
+ $X2=1.15 $Y2=0
r144 61 88 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r145 61 100 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r146 59 79 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.29
+ $Y2=0
r147 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.42
+ $Y2=0
r148 57 76 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=0
+ $X2=4.37 $Y2=0
r149 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=0 $X2=4.58
+ $Y2=0
r150 56 79 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=5.29 $Y2=0
r151 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.58
+ $Y2=0
r152 54 73 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.655 $Y=0
+ $X2=3.45 $Y2=0
r153 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.74
+ $Y2=0
r154 53 76 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.825 $Y=0
+ $X2=4.37 $Y2=0
r155 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.74
+ $Y2=0
r156 51 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r157 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.54
+ $Y2=0
r158 50 69 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.625 $Y=0
+ $X2=2.07 $Y2=0
r159 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.54
+ $Y2=0
r160 46 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=0.085
+ $X2=6.26 $Y2=0
r161 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.26 $Y=0.085
+ $X2=6.26 $Y2=0.39
r162 45 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=0 $X2=5.42
+ $Y2=0
r163 44 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0 $X2=6.26
+ $Y2=0
r164 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.175 $Y=0
+ $X2=5.505 $Y2=0
r165 40 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=0.085
+ $X2=5.42 $Y2=0
r166 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.42 $Y=0.085
+ $X2=5.42 $Y2=0.39
r167 36 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r168 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.39
r169 32 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0.085
+ $X2=3.74 $Y2=0
r170 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.74 $Y=0.085
+ $X2=3.74 $Y2=0.39
r171 28 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0
r172 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0.39
r173 24 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r174 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.39
r175 7 48 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.125
+ $Y=0.235 $X2=6.26 $Y2=0.39
r176 6 42 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.235 $X2=5.42 $Y2=0.39
r177 5 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.39
r178 4 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.235 $X2=3.74 $Y2=0.39
r179 3 94 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.235 $X2=2.9 $Y2=0.39
r180 2 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r181 1 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends


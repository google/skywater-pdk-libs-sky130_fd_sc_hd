# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlrtn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595000 0.255000 5.925000 0.485000 ;
        RECT 5.655000 1.875000 5.925000 2.465000 ;
        RECT 5.755000 0.485000 5.925000 0.765000 ;
        RECT 5.755000 0.765000 6.355000 0.865000 ;
        RECT 5.755000 1.425000 6.355000 1.500000 ;
        RECT 5.755000 1.500000 5.925000 1.875000 ;
        RECT 5.760000 1.415000 6.355000 1.425000 ;
        RECT 5.765000 1.410000 6.355000 1.415000 ;
        RECT 5.770000 0.865000 6.355000 0.890000 ;
        RECT 5.775000 1.385000 6.355000 1.410000 ;
        RECT 5.785000 0.890000 6.355000 1.385000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.480000 0.995000 5.170000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.875000  0.085000 2.205000 0.445000 ;
        RECT 3.735000  0.085000 4.070000 0.530000 ;
        RECT 5.095000  0.085000 5.425000 0.485000 ;
        RECT 6.095000  0.085000 6.355000 0.595000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.955000 1.835000 2.270000 2.635000 ;
        RECT 3.800000 2.135000 4.110000 2.635000 ;
        RECT 4.280000 2.135000 4.560000 2.635000 ;
        RECT 5.090000 1.875000 5.460000 2.635000 ;
        RECT 6.095000 1.670000 6.355000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.780000 0.805000 ;
      RECT 0.175000 1.795000 0.780000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.780000 1.070000 ;
      RECT 0.610000 1.070000 0.840000 1.400000 ;
      RECT 0.610000 1.400000 0.780000 1.795000 ;
      RECT 1.015000 0.345000 1.185000 1.685000 ;
      RECT 1.015000 1.685000 1.240000 2.465000 ;
      RECT 1.455000 1.495000 2.140000 1.665000 ;
      RECT 1.455000 1.665000 1.785000 2.415000 ;
      RECT 1.535000 0.345000 1.705000 0.615000 ;
      RECT 1.535000 0.615000 2.140000 0.765000 ;
      RECT 1.535000 0.765000 2.340000 0.785000 ;
      RECT 1.960000 0.785000 2.340000 1.095000 ;
      RECT 1.960000 1.095000 2.140000 1.495000 ;
      RECT 2.470000 1.355000 2.755000 2.005000 ;
      RECT 2.675000 0.705000 3.095000 1.145000 ;
      RECT 2.775000 2.255000 3.605000 2.425000 ;
      RECT 2.810000 0.365000 3.500000 0.535000 ;
      RECT 2.925000 1.145000 3.095000 1.415000 ;
      RECT 2.925000 1.415000 3.265000 1.995000 ;
      RECT 3.330000 0.535000 3.500000 1.025000 ;
      RECT 3.330000 1.025000 4.310000 1.245000 ;
      RECT 3.435000 1.245000 4.310000 1.325000 ;
      RECT 3.435000 1.325000 3.605000 2.255000 ;
      RECT 3.820000 1.535000 5.585000 1.705000 ;
      RECT 3.820000 1.705000 4.920000 1.865000 ;
      RECT 4.240000 0.255000 4.590000 0.655000 ;
      RECT 4.240000 0.655000 5.585000 0.825000 ;
      RECT 4.730000 1.865000 4.920000 2.465000 ;
      RECT 5.350000 0.995000 5.615000 1.325000 ;
      RECT 5.415000 0.825000 5.585000 0.995000 ;
      RECT 5.415000 1.325000 5.585000 1.535000 ;
    LAYER mcon ;
      RECT 0.610000 1.445000 0.780000 1.615000 ;
      RECT 1.070000 1.785000 1.240000 1.955000 ;
      RECT 2.470000 1.785000 2.640000 1.955000 ;
      RECT 2.930000 1.445000 3.100000 1.615000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_2

* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_2.pex.spice
* Created: Tue Sep  1 19:11:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%A 3 7 11 13 15 19 21 22 23
r56 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1
+ $Y=1.16 $X2=1 $Y2=1.16
r57 32 34 10.3656 $w=2.79e-07 $l=6e-08 $layer=POLY_cond $X=0.94 $Y=1.16 $X2=1
+ $Y2=1.16
r58 28 30 30.233 $w=2.79e-07 $l=1.75e-07 $layer=POLY_cond $X=0.32 $Y=1.16
+ $X2=0.495 $Y2=1.16
r59 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.16 $X2=0.32 $Y2=1.16
r60 23 35 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=1.177 $X2=1
+ $Y2=1.177
r61 22 35 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=0.69 $Y=1.177 $X2=1
+ $Y2=1.177
r62 22 29 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=1.177
+ $X2=0.32 $Y2=1.177
r63 21 29 4.60977 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=0.23 $Y=1.177 $X2=0.32
+ $Y2=1.177
r64 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.37 $Y=1.025
+ $X2=1.37 $Y2=0.445
r65 13 17 2.5914 $w=2.79e-07 $l=1.5e-08 $layer=POLY_cond $X=1.355 $Y=1.16
+ $X2=1.37 $Y2=1.16
r66 13 34 61.3298 $w=2.79e-07 $l=3.55e-07 $layer=POLY_cond $X=1.355 $Y=1.16
+ $X2=1 $Y2=1.16
r67 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.355 $Y=1.295
+ $X2=1.355 $Y2=1.985
r68 9 32 17.2686 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.94 $Y=1.015
+ $X2=0.94 $Y2=1.16
r69 9 11 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.94 $Y=1.015
+ $X2=0.94 $Y2=0.445
r70 5 32 2.5914 $w=2.79e-07 $l=1.5e-08 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.94 $Y2=1.16
r71 5 30 74.2867 $w=2.79e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.495 $Y2=1.16
r72 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.925 $Y=1.295
+ $X2=0.925 $Y2=1.985
r73 1 30 17.2686 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.495 $Y=1.305
+ $X2=0.495 $Y2=1.16
r74 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.495 $Y=1.305
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%Y 1 2 3 12 14 15 18 22 24 26 27
+ 28 29 30 31 37 38
c68 37 0 8.53357e-20 $X=1.615 $Y=0.895
r69 31 38 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=1.545
+ $X2=1.615 $Y2=1.46
r70 31 38 0.329269 $w=2.78e-07 $l=8e-09 $layer=LI1_cond $X=1.615 $Y=1.452
+ $X2=1.615 $Y2=1.46
r71 30 31 10.7836 $w=2.78e-07 $l=2.62e-07 $layer=LI1_cond $X=1.615 $Y=1.19
+ $X2=1.615 $Y2=1.452
r72 29 37 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.81
+ $X2=1.615 $Y2=0.895
r73 29 30 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=0.915
+ $X2=1.615 $Y2=1.19
r74 29 37 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=1.615 $Y=0.915
+ $X2=1.615 $Y2=0.895
r75 26 29 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=1.615 $Y2=0.81
r76 26 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=1.25 $Y2=0.81
r77 25 28 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.235 $Y=1.545
+ $X2=1.14 $Y2=1.545
r78 24 31 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.475 $Y=1.545
+ $X2=1.615 $Y2=1.545
r79 24 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.475 $Y=1.545
+ $X2=1.235 $Y2=1.545
r80 20 28 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.63
+ $X2=1.14 $Y2=1.545
r81 20 22 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=1.14 $Y=1.63 $X2=1.14
+ $Y2=1.83
r82 16 27 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.137 $Y=0.725
+ $X2=1.25 $Y2=0.81
r83 16 18 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=1.137 $Y=0.725
+ $X2=1.137 $Y2=0.445
r84 14 28 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.045 $Y=1.545
+ $X2=1.14 $Y2=1.545
r85 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.045 $Y=1.545
+ $X2=0.375 $Y2=1.545
r86 10 15 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.265 $Y=1.63
+ $X2=0.375 $Y2=1.545
r87 10 12 10.4768 $w=2.18e-07 $l=2e-07 $layer=LI1_cond $X=0.265 $Y=1.63
+ $X2=0.265 $Y2=1.83
r88 3 22 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.485 $X2=1.14 $Y2=1.83
r89 2 12 300 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=1.83
r90 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.155 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%KAPWR 1 2 7 13 14 18 21 26
r39 17 26 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.57 $Y=2.21
+ $X2=1.57 $Y2=1.965
r40 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.585 $Y=2.21
+ $X2=1.585 $Y2=2.21
r41 13 18 0.230264 $w=2e-07 $l=3e-07 $layer=MET1_cond $X=0.54 $Y=2.24 $X2=0.24
+ $Y2=2.24
r42 12 21 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.71 $Y=2.21
+ $X2=0.71 $Y2=1.965
r43 11 14 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.685 $Y=2.21
+ $X2=0.83 $Y2=2.21
r44 11 13 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.685 $Y=2.21
+ $X2=0.54 $Y2=2.21
r45 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.685 $Y=2.21
+ $X2=0.685 $Y2=2.21
r46 7 16 0.077601 $w=2.52e-07 $l=1.59295e-07 $layer=MET1_cond $X=1.44 $Y=2.24
+ $X2=1.585 $Y2=2.21
r47 7 14 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=1.44 $Y=2.24 $X2=0.83
+ $Y2=2.24
r48 2 26 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=1.485 $X2=1.57 $Y2=1.965
r49 1 21 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.485 $X2=0.71 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%VGND 1 2 9 11 13 15 17 22 28 32
c24 11 0 8.53357e-20 $X=1.585 $Y=0.085
r25 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r26 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r27 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r28 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r29 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r30 23 28 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.707
+ $Y2=0
r31 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.15
+ $Y2=0
r32 22 31 4.79676 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.63
+ $Y2=0
r33 22 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.15
+ $Y2=0
r34 17 28 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.707
+ $Y2=0
r35 17 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.23
+ $Y2=0
r36 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r37 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r38 11 31 2.96942 $w=3.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.63 $Y2=0
r39 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.585 $Y2=0.39
r40 7 28 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0
r41 7 9 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0.445
r42 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.39
r43 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.725 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%VPWR 1 8 9
r25 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72 $X2=1.61
+ $Y2=2.72
r26 4 8 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=1.61
+ $Y2=2.72
r27 1 9 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 1 4 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends


* File: sky130_fd_sc_hd__ha_1.pxi.spice
* Created: Thu Aug 27 14:21:59 2020
* 
x_PM_SKY130_FD_SC_HD__HA_1%A_79_21# N_A_79_21#_M1003_s N_A_79_21#_M1005_d
+ N_A_79_21#_c_92_n N_A_79_21#_M1012_g N_A_79_21#_M1011_g N_A_79_21#_c_93_n
+ N_A_79_21#_c_94_n N_A_79_21#_c_95_n N_A_79_21#_c_96_n N_A_79_21#_c_102_n
+ N_A_79_21#_c_103_n N_A_79_21#_c_97_n N_A_79_21#_c_98_n N_A_79_21#_c_104_n
+ PM_SKY130_FD_SC_HD__HA_1%A_79_21#
x_PM_SKY130_FD_SC_HD__HA_1%A_250_199# N_A_250_199#_M1004_s N_A_250_199#_M1009_d
+ N_A_250_199#_M1005_g N_A_250_199#_M1003_g N_A_250_199#_M1010_g
+ N_A_250_199#_M1013_g N_A_250_199#_c_161_n N_A_250_199#_c_162_n
+ N_A_250_199#_c_163_n N_A_250_199#_c_172_n N_A_250_199#_c_173_n
+ N_A_250_199#_c_174_n N_A_250_199#_c_164_n N_A_250_199#_c_176_n
+ N_A_250_199#_c_165_n N_A_250_199#_c_166_n N_A_250_199#_c_167_n
+ N_A_250_199#_c_168_n N_A_250_199#_c_169_n PM_SKY130_FD_SC_HD__HA_1%A_250_199#
x_PM_SKY130_FD_SC_HD__HA_1%B N_B_M1001_g N_B_M1002_g N_B_c_292_n N_B_M1009_g
+ N_B_c_293_n N_B_M1004_g N_B_c_294_n B B B N_B_c_300_n N_B_c_301_n N_B_c_302_n
+ B PM_SKY130_FD_SC_HD__HA_1%B
x_PM_SKY130_FD_SC_HD__HA_1%A N_A_M1008_g N_A_c_376_n N_A_M1007_g N_A_M1006_g
+ N_A_M1000_g A A N_A_c_379_n PM_SKY130_FD_SC_HD__HA_1%A
x_PM_SKY130_FD_SC_HD__HA_1%SUM N_SUM_M1012_s N_SUM_M1011_s SUM SUM SUM SUM SUM
+ SUM N_SUM_c_457_n SUM SUM PM_SKY130_FD_SC_HD__HA_1%SUM
x_PM_SKY130_FD_SC_HD__HA_1%VPWR N_VPWR_M1011_d N_VPWR_M1007_d N_VPWR_M1000_d
+ N_VPWR_c_488_n N_VPWR_c_477_n VPWR N_VPWR_c_478_n N_VPWR_c_479_n
+ N_VPWR_c_476_n N_VPWR_c_481_n N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n
+ N_VPWR_c_485_n PM_SKY130_FD_SC_HD__HA_1%VPWR
x_PM_SKY130_FD_SC_HD__HA_1%COUT N_COUT_M1010_d N_COUT_M1013_d N_COUT_c_544_n
+ N_COUT_c_542_n COUT COUT COUT N_COUT_c_543_n PM_SKY130_FD_SC_HD__HA_1%COUT
x_PM_SKY130_FD_SC_HD__HA_1%VGND N_VGND_M1012_d N_VGND_M1002_d N_VGND_M1006_d
+ N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n VGND N_VGND_c_567_n
+ N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n
+ N_VGND_c_573_n N_VGND_c_574_n PM_SKY130_FD_SC_HD__HA_1%VGND
x_PM_SKY130_FD_SC_HD__HA_1%A_297_47# N_A_297_47#_M1003_d N_A_297_47#_M1008_d
+ N_A_297_47#_c_649_n N_A_297_47#_c_634_n N_A_297_47#_c_635_n
+ N_A_297_47#_c_642_n PM_SKY130_FD_SC_HD__HA_1%A_297_47#
cc_1 VNB N_A_79_21#_c_92_n 0.0229166f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_93_n 0.0116115f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.16
cc_3 VNB N_A_79_21#_c_94_n 0.03421f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_4 VNB N_A_79_21#_c_95_n 0.00956187f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.075
cc_5 VNB N_A_79_21#_c_96_n 0.00125104f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.935
cc_6 VNB N_A_79_21#_c_97_n 0.0103009f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.51
cc_7 VNB N_A_79_21#_c_98_n 0.00195951f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.16
cc_8 VNB N_A_250_199#_M1003_g 0.0327009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_250_199#_c_161_n 0.0383161f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.935
cc_10 VNB N_A_250_199#_c_162_n 0.00118612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_250_199#_c_163_n 0.00840268f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.51
cc_12 VNB N_A_250_199#_c_164_n 0.00579852f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_13 VNB N_A_250_199#_c_165_n 0.00146092f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_14 VNB N_A_250_199#_c_166_n 0.0248692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_250_199#_c_167_n 0.00288254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_250_199#_c_168_n 0.0225749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_250_199#_c_169_n 0.0199171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_M1002_g 0.0409724f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_19 VNB N_B_c_292_n 0.0249467f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_20 VNB N_B_c_293_n 0.017225f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_21 VNB N_B_c_294_n 0.0258978f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.075
cc_22 VNB N_A_M1008_g 0.0406098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_c_376_n 0.0247949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_M1006_g 0.0359067f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_25 VNB A 0.00269502f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_26 VNB N_A_c_379_n 0.0175665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB SUM 0.0065071f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_28 VNB N_SUM_c_457_n 0.0136819f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=2.02
cc_29 VNB SUM 0.0237503f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.16
cc_30 VNB N_VPWR_c_476_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_31 VNB N_COUT_c_542_n 0.02217f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_32 VNB N_COUT_c_543_n 0.0203973f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.51
cc_33 VNB N_VGND_c_564_n 0.0060017f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_34 VNB N_VGND_c_565_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_35 VNB N_VGND_c_566_n 0.00513775f $X=-0.19 $Y=-0.24 $X2=1.045 $Y2=1.075
cc_36 VNB N_VGND_c_567_n 0.0182914f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=2.02
cc_37 VNB N_VGND_c_568_n 0.0287637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_569_n 0.0425743f $X=-0.19 $Y=-0.24 $X2=1.595 $Y2=2.19
cc_39 VNB N_VGND_c_570_n 0.0182496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_571_n 0.260866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_572_n 0.00375078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_573_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_574_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_297_47#_c_634_n 0.0059863f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_45 VNB N_A_297_47#_c_635_n 0.00293934f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_46 VPB N_A_79_21#_M1011_g 0.0261089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_47 VPB N_A_79_21#_c_94_n 0.00913593f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_48 VPB N_A_79_21#_c_96_n 0.0150233f $X=-0.19 $Y=1.305 $X2=1.045 $Y2=1.935
cc_49 VPB N_A_79_21#_c_102_n 0.00586191f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=2.02
cc_50 VPB N_A_79_21#_c_103_n 0.00171804f $X=-0.19 $Y=1.305 $X2=1.13 $Y2=2.02
cc_51 VPB N_A_79_21#_c_104_n 0.00738039f $X=-0.19 $Y=1.305 $X2=1.595 $Y2=2.02
cc_52 VPB N_A_250_199#_M1005_g 0.0556072f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_53 VPB N_A_250_199#_M1013_g 0.0228008f $X=-0.19 $Y=1.305 $X2=1.045 $Y2=1.075
cc_54 VPB N_A_250_199#_c_172_n 0.00221691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_250_199#_c_173_n 0.00474958f $X=-0.19 $Y=1.305 $X2=1.595 $Y2=2.19
cc_56 VPB N_A_250_199#_c_174_n 0.00306113f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_250_199#_c_164_n 0.00199884f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_58 VPB N_A_250_199#_c_176_n 0.00218475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_250_199#_c_165_n 2.9289e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_60 VPB N_A_250_199#_c_166_n 0.00530782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_250_199#_c_168_n 0.00462376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_B_M1001_g 0.0236854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B_M1002_g 0.0100915f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_64 VPB N_B_c_292_n 0.0132711f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_65 VPB N_B_M1009_g 0.0216213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB B 0.00502263f $X=-0.19 $Y=1.305 $X2=1.045 $Y2=1.935
cc_67 VPB N_B_c_300_n 0.0324837f $X=-0.19 $Y=1.305 $X2=1.595 $Y2=2.02
cc_68 VPB N_B_c_301_n 0.0174043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_B_c_302_n 0.0425861f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_70 VPB B 0.0026068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_c_376_n 0.0247562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_M1007_g 0.0417572f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_73 VPB N_A_M1000_g 0.0422213f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_74 VPB A 0.00339211f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_75 VPB A 0.0113595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_c_379_n 0.0197435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB SUM 0.0065071f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_78 VPB SUM 0.0269238f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_79 VPB SUM 0.0124231f $X=-0.19 $Y=1.305 $X2=1.045 $Y2=1.16
cc_80 VPB N_VPWR_c_477_n 0.00456988f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_81 VPB N_VPWR_c_478_n 0.018869f $X=-0.19 $Y=1.305 $X2=1.045 $Y2=1.16
cc_82 VPB N_VPWR_c_479_n 0.0181937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_476_n 0.043974f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_84 VPB N_VPWR_c_481_n 0.0182363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_482_n 0.0202593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_483_n 0.0319616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_484_n 0.0198334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_485_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_COUT_c_544_n 0.00666696f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_90 VPB N_COUT_c_542_n 0.0117188f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_91 VPB COUT 0.0270182f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_92 N_A_79_21#_c_96_n N_A_250_199#_M1005_g 0.0206262f $X=1.045 $Y=1.935 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_102_n N_A_250_199#_M1005_g 0.0138745f $X=1.51 $Y=2.02 $X2=0
+ $Y2=0
cc_94 N_A_79_21#_c_104_n N_A_250_199#_M1005_g 2.60173e-19 $X=1.595 $Y=2.02 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_95_n N_A_250_199#_M1003_g 0.0084221f $X=1.045 $Y=1.075 $X2=0
+ $Y2=0
cc_96 N_A_79_21#_c_97_n N_A_250_199#_M1003_g 4.49111e-19 $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_c_95_n N_A_250_199#_c_165_n 0.00718969f $X=1.045 $Y=1.075 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_96_n N_A_250_199#_c_165_n 0.00568393f $X=1.045 $Y=1.935 $X2=0
+ $Y2=0
cc_99 N_A_79_21#_c_102_n N_A_250_199#_c_165_n 0.00425848f $X=1.51 $Y=2.02 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_98_n N_A_250_199#_c_165_n 0.0136441f $X=1.045 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_c_94_n N_A_250_199#_c_166_n 0.00652051f $X=0.655 $Y=1.16 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_95_n N_A_250_199#_c_166_n 7.0804e-19 $X=1.045 $Y=1.075 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_c_96_n N_A_250_199#_c_166_n 7.0804e-19 $X=1.045 $Y=1.935 $X2=0
+ $Y2=0
cc_104 N_A_79_21#_c_102_n N_A_250_199#_c_166_n 0.00232016f $X=1.51 $Y=2.02 $X2=0
+ $Y2=0
cc_105 N_A_79_21#_c_97_n N_A_250_199#_c_166_n 0.00120572f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_c_98_n N_A_250_199#_c_166_n 0.00165735f $X=1.045 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_79_21#_c_104_n N_A_250_199#_c_166_n 2.37457e-19 $X=1.595 $Y=2.02
+ $X2=0 $Y2=0
cc_108 N_A_79_21#_c_104_n N_B_M1001_g 8.97627e-19 $X=1.595 $Y=2.02 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_104_n B 0.0204239f $X=1.595 $Y=2.02 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_92_n SUM 0.00323429f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_79_21#_M1011_g SUM 0.00328979f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_79_21#_M1011_g SUM 0.00778907f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_92_n N_SUM_c_457_n 0.00407486f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_92_n SUM 0.0173447f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_93_n SUM 0.0136576f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_95_n SUM 0.00571705f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_96_n SUM 0.00809204f $X=1.045 $Y=1.935 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_102_n N_VPWR_M1011_d 0.00124571f $X=1.51 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_79_21#_c_103_n N_VPWR_M1011_d 0.0025543f $X=1.13 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_79_21#_c_93_n N_VPWR_c_488_n 0.0104923f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_94_n N_VPWR_c_488_n 0.00466049f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_96_n N_VPWR_c_488_n 0.0313449f $X=1.045 $Y=1.935 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_103_n N_VPWR_c_488_n 0.0139466f $X=1.13 $Y=2.02 $X2=0 $Y2=0
cc_124 N_A_79_21#_M1005_d N_VPWR_c_476_n 0.00417627f $X=1.46 $Y=2.065 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_M1011_g N_VPWR_c_476_n 0.0117832f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_102_n N_VPWR_c_476_n 0.00767696f $X=1.51 $Y=2.02 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_103_n N_VPWR_c_476_n 8.91481e-19 $X=1.13 $Y=2.02 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_104_n N_VPWR_c_476_n 0.00599338f $X=1.595 $Y=2.02 $X2=0
+ $Y2=0
cc_129 N_A_79_21#_M1011_g N_VPWR_c_481_n 0.00543342f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_79_21#_M1011_g N_VPWR_c_482_n 0.00480473f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_79_21#_c_102_n N_VPWR_c_482_n 0.00924191f $X=1.51 $Y=2.02 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_103_n N_VPWR_c_482_n 0.0141558f $X=1.13 $Y=2.02 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_102_n N_VPWR_c_483_n 0.00308156f $X=1.51 $Y=2.02 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_104_n N_VPWR_c_483_n 0.00644334f $X=1.595 $Y=2.02 $X2=0
+ $Y2=0
cc_135 N_A_79_21#_c_92_n N_VGND_c_564_n 0.00442456f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_93_n N_VGND_c_564_n 0.0137319f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_94_n N_VGND_c_564_n 0.00488398f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_95_n N_VGND_c_564_n 0.0156913f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_97_n N_VGND_c_564_n 0.0259068f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_92_n N_VGND_c_567_n 0.00543728f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_97_n N_VGND_c_568_n 0.013655f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_142 N_A_79_21#_M1003_s N_VGND_c_571_n 0.00390713f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_79_21#_c_92_n N_VGND_c_571_n 0.011787f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_97_n N_VGND_c_571_n 0.0116462f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_95_n N_A_297_47#_c_635_n 0.00598365f $X=1.045 $Y=1.075 $X2=0
+ $Y2=0
cc_146 N_A_79_21#_c_97_n N_A_297_47#_c_635_n 0.00121593f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_147 N_A_250_199#_M1005_g N_B_M1002_g 0.00677382f $X=1.385 $Y=2.275 $X2=0
+ $Y2=0
cc_148 N_A_250_199#_M1003_g N_B_M1002_g 0.0262193f $X=1.41 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_250_199#_c_161_n N_B_M1002_g 0.0130752f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_150 N_A_250_199#_c_165_n N_B_M1002_g 0.00115517f $X=1.385 $Y=1.06 $X2=0 $Y2=0
cc_151 N_A_250_199#_c_166_n N_B_M1002_g 0.0186141f $X=1.385 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_250_199#_c_161_n N_B_c_292_n 0.00492578f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_153 N_A_250_199#_c_167_n N_B_c_292_n 0.00924318f $X=3.085 $Y=0.8 $X2=0 $Y2=0
cc_154 N_A_250_199#_c_172_n N_B_M1009_g 0.00701263f $X=3.435 $Y=2.19 $X2=0 $Y2=0
cc_155 N_A_250_199#_c_162_n N_B_c_293_n 0.00234105f $X=3.085 $Y=0.51 $X2=0 $Y2=0
cc_156 N_A_250_199#_c_163_n N_B_c_293_n 0.00444942f $X=3.835 $Y=0.8 $X2=0 $Y2=0
cc_157 N_A_250_199#_c_163_n N_B_c_294_n 0.0079839f $X=3.835 $Y=0.8 $X2=0 $Y2=0
cc_158 N_A_250_199#_c_167_n N_B_c_294_n 0.00933316f $X=3.085 $Y=0.8 $X2=0 $Y2=0
cc_159 N_A_250_199#_M1005_g B 0.00155561f $X=1.385 $Y=2.275 $X2=0 $Y2=0
cc_160 N_A_250_199#_c_161_n B 0.0223589f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_161 N_A_250_199#_M1005_g B 8.3268e-19 $X=1.385 $Y=2.275 $X2=0 $Y2=0
cc_162 N_A_250_199#_M1005_g N_B_c_300_n 0.0373968f $X=1.385 $Y=2.275 $X2=0 $Y2=0
cc_163 N_A_250_199#_c_161_n N_B_c_300_n 0.00165507f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_164 N_A_250_199#_c_161_n N_B_c_301_n 0.00548196f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_165 N_A_250_199#_c_174_n N_B_c_301_n 0.00325047f $X=3.52 $Y=1.87 $X2=0 $Y2=0
cc_166 N_A_250_199#_c_176_n N_B_c_301_n 0.00388358f $X=3.92 $Y=1.785 $X2=0 $Y2=0
cc_167 N_A_250_199#_c_174_n N_B_c_302_n 0.00453475f $X=3.52 $Y=1.87 $X2=0 $Y2=0
cc_168 N_A_250_199#_M1005_g B 5.44018e-19 $X=1.385 $Y=2.275 $X2=0 $Y2=0
cc_169 N_A_250_199#_c_161_n N_A_M1008_g 0.00925764f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_170 N_A_250_199#_c_162_n N_A_M1008_g 3.5555e-19 $X=3.085 $Y=0.51 $X2=0 $Y2=0
cc_171 N_A_250_199#_c_167_n N_A_M1008_g 9.46444e-19 $X=3.085 $Y=0.8 $X2=0 $Y2=0
cc_172 N_A_250_199#_c_161_n N_A_c_376_n 0.0120469f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_173 N_A_250_199#_c_163_n N_A_M1006_g 0.0159476f $X=3.835 $Y=0.8 $X2=0 $Y2=0
cc_174 N_A_250_199#_c_164_n N_A_M1006_g 0.00411404f $X=3.92 $Y=1.325 $X2=0 $Y2=0
cc_175 N_A_250_199#_c_167_n N_A_M1006_g 0.00159259f $X=3.085 $Y=0.8 $X2=0 $Y2=0
cc_176 N_A_250_199#_c_168_n N_A_M1006_g 0.0199937f $X=4.075 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_250_199#_c_169_n N_A_M1006_g 0.0196549f $X=4.075 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_250_199#_c_172_n N_A_M1000_g 0.00277205f $X=3.435 $Y=2.19 $X2=0 $Y2=0
cc_179 N_A_250_199#_c_173_n N_A_M1000_g 0.0154589f $X=3.835 $Y=1.87 $X2=0 $Y2=0
cc_180 N_A_250_199#_c_163_n A 0.0184671f $X=3.835 $Y=0.8 $X2=0 $Y2=0
cc_181 N_A_250_199#_c_173_n A 0.00524875f $X=3.835 $Y=1.87 $X2=0 $Y2=0
cc_182 N_A_250_199#_c_174_n A 0.0144887f $X=3.52 $Y=1.87 $X2=0 $Y2=0
cc_183 N_A_250_199#_c_164_n A 0.0156083f $X=3.92 $Y=1.325 $X2=0 $Y2=0
cc_184 N_A_250_199#_c_176_n A 0.0156352f $X=3.92 $Y=1.785 $X2=0 $Y2=0
cc_185 N_A_250_199#_c_167_n A 0.00640198f $X=3.085 $Y=0.8 $X2=0 $Y2=0
cc_186 N_A_250_199#_c_168_n A 2.32088e-19 $X=4.075 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_250_199#_c_161_n A 0.0484719f $X=3 $Y=1.06 $X2=0 $Y2=0
cc_188 N_A_250_199#_c_163_n A 0.00674865f $X=3.835 $Y=0.8 $X2=0 $Y2=0
cc_189 N_A_250_199#_c_174_n A 5.22199e-19 $X=3.52 $Y=1.87 $X2=0 $Y2=0
cc_190 N_A_250_199#_c_167_n A 0.0130791f $X=3.085 $Y=0.8 $X2=0 $Y2=0
cc_191 N_A_250_199#_M1013_g N_A_c_379_n 0.0292551f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_250_199#_c_163_n N_A_c_379_n 0.00122233f $X=3.835 $Y=0.8 $X2=0 $Y2=0
cc_193 N_A_250_199#_c_173_n N_A_c_379_n 3.03728e-19 $X=3.835 $Y=1.87 $X2=0 $Y2=0
cc_194 N_A_250_199#_c_174_n N_A_c_379_n 0.00114807f $X=3.52 $Y=1.87 $X2=0 $Y2=0
cc_195 N_A_250_199#_c_176_n N_A_c_379_n 0.00496915f $X=3.92 $Y=1.785 $X2=0 $Y2=0
cc_196 N_A_250_199#_c_173_n N_VPWR_M1000_d 0.00397523f $X=3.835 $Y=1.87 $X2=0
+ $Y2=0
cc_197 N_A_250_199#_c_176_n N_VPWR_M1000_d 0.00529043f $X=3.92 $Y=1.785 $X2=0
+ $Y2=0
cc_198 N_A_250_199#_M1005_g N_VPWR_c_488_n 0.00520245f $X=1.385 $Y=2.275 $X2=0
+ $Y2=0
cc_199 N_A_250_199#_M1013_g N_VPWR_c_477_n 0.00287759f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_250_199#_c_173_n N_VPWR_c_477_n 0.0190723f $X=3.835 $Y=1.87 $X2=0
+ $Y2=0
cc_201 N_A_250_199#_c_172_n N_VPWR_c_478_n 0.00679825f $X=3.435 $Y=2.19 $X2=0
+ $Y2=0
cc_202 N_A_250_199#_M1013_g N_VPWR_c_479_n 0.00543342f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_250_199#_M1009_d N_VPWR_c_476_n 0.00485007f $X=3.29 $Y=2.065 $X2=0
+ $Y2=0
cc_204 N_A_250_199#_M1005_g N_VPWR_c_476_n 0.00710884f $X=1.385 $Y=2.275 $X2=0
+ $Y2=0
cc_205 N_A_250_199#_M1013_g N_VPWR_c_476_n 0.0106163f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_250_199#_c_172_n N_VPWR_c_476_n 0.00605484f $X=3.435 $Y=2.19 $X2=0
+ $Y2=0
cc_207 N_A_250_199#_c_173_n N_VPWR_c_476_n 0.00843536f $X=3.835 $Y=1.87 $X2=0
+ $Y2=0
cc_208 N_A_250_199#_M1005_g N_VPWR_c_482_n 0.00882152f $X=1.385 $Y=2.275 $X2=0
+ $Y2=0
cc_209 N_A_250_199#_M1005_g N_VPWR_c_483_n 0.00422112f $X=1.385 $Y=2.275 $X2=0
+ $Y2=0
cc_210 N_A_250_199#_M1013_g N_COUT_c_544_n 0.00324226f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_250_199#_M1013_g N_COUT_c_542_n 0.003653f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_250_199#_c_164_n N_COUT_c_542_n 0.0305823f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_213 N_A_250_199#_c_176_n N_COUT_c_542_n 0.00835575f $X=3.92 $Y=1.785 $X2=0
+ $Y2=0
cc_214 N_A_250_199#_c_168_n N_COUT_c_542_n 0.00754383f $X=4.075 $Y=1.16 $X2=0
+ $Y2=0
cc_215 N_A_250_199#_c_169_n N_COUT_c_542_n 0.00245797f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_216 N_A_250_199#_M1013_g COUT 0.00902992f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_250_199#_c_172_n COUT 0.00442841f $X=3.435 $Y=2.19 $X2=0 $Y2=0
cc_218 N_A_250_199#_c_169_n N_COUT_c_543_n 0.00857862f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_250_199#_c_163_n N_VGND_M1006_d 0.00140691f $X=3.835 $Y=0.8 $X2=0
+ $Y2=0
cc_220 N_A_250_199#_c_164_n N_VGND_M1006_d 0.00223361f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_221 N_A_250_199#_M1003_g N_VGND_c_564_n 0.00468029f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A_250_199#_M1003_g N_VGND_c_565_n 0.00155517f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_250_199#_c_163_n N_VGND_c_566_n 0.00481848f $X=3.835 $Y=0.8 $X2=0
+ $Y2=0
cc_224 N_A_250_199#_c_164_n N_VGND_c_566_n 0.0140595f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_225 N_A_250_199#_c_168_n N_VGND_c_566_n 2.60901e-19 $X=4.075 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_250_199#_c_169_n N_VGND_c_566_n 0.00287759f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_250_199#_M1003_g N_VGND_c_568_n 0.00585385f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_228 N_A_250_199#_c_162_n N_VGND_c_569_n 0.00732874f $X=3.085 $Y=0.51 $X2=0
+ $Y2=0
cc_229 N_A_250_199#_c_163_n N_VGND_c_569_n 0.00852444f $X=3.835 $Y=0.8 $X2=0
+ $Y2=0
cc_230 N_A_250_199#_c_169_n N_VGND_c_570_n 0.00543728f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_250_199#_M1004_s N_VGND_c_571_n 0.00344181f $X=2.96 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_250_199#_M1003_g N_VGND_c_571_n 0.0122169f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_233 N_A_250_199#_c_162_n N_VGND_c_571_n 0.00616598f $X=3.085 $Y=0.51 $X2=0
+ $Y2=0
cc_234 N_A_250_199#_c_163_n N_VGND_c_571_n 0.0143447f $X=3.835 $Y=0.8 $X2=0
+ $Y2=0
cc_235 N_A_250_199#_c_164_n N_VGND_c_571_n 7.42202e-19 $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_236 N_A_250_199#_c_169_n N_VGND_c_571_n 0.0106176f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_250_199#_c_161_n N_A_297_47#_c_634_n 0.0620304f $X=3 $Y=1.06 $X2=0
+ $Y2=0
cc_238 N_A_250_199#_c_162_n N_A_297_47#_c_634_n 0.00689583f $X=3.085 $Y=0.51
+ $X2=0 $Y2=0
cc_239 N_A_250_199#_M1003_g N_A_297_47#_c_635_n 0.00183499f $X=1.41 $Y=0.445
+ $X2=0 $Y2=0
cc_240 N_A_250_199#_c_161_n N_A_297_47#_c_635_n 0.0139109f $X=3 $Y=1.06 $X2=0
+ $Y2=0
cc_241 N_A_250_199#_c_162_n N_A_297_47#_c_642_n 0.0101661f $X=3.085 $Y=0.51
+ $X2=0 $Y2=0
cc_242 N_B_M1002_g N_A_M1008_g 0.033214f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_243 N_B_c_294_n N_A_M1008_g 0.00587607f $X=3.295 $Y=0.81 $X2=0 $Y2=0
cc_244 N_B_M1002_g N_A_c_376_n 0.015002f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_245 N_B_c_292_n N_A_c_376_n 0.0156246f $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_246 B N_A_c_376_n 0.00529165f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_247 N_B_c_300_n N_A_c_376_n 0.0206333f $X=1.935 $Y=1.66 $X2=0 $Y2=0
cc_248 N_B_c_301_n N_A_c_376_n 0.00761419f $X=3 $Y=1.74 $X2=0 $Y2=0
cc_249 N_B_M1001_g N_A_M1007_g 0.0212295f $X=1.805 $Y=2.275 $X2=0 $Y2=0
cc_250 N_B_c_292_n N_A_M1007_g 2.44403e-19 $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_251 N_B_M1009_g N_A_M1007_g 0.00701339f $X=3.215 $Y=2.275 $X2=0 $Y2=0
cc_252 N_B_c_301_n N_A_M1007_g 0.0159047f $X=3 $Y=1.74 $X2=0 $Y2=0
cc_253 N_B_c_302_n N_A_M1007_g 0.0105516f $X=3.06 $Y=1.75 $X2=0 $Y2=0
cc_254 B N_A_M1007_g 0.0125548f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_255 N_B_c_292_n N_A_M1006_g 0.00608316f $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_256 N_B_c_293_n N_A_M1006_g 0.0489147f $X=3.295 $Y=0.735 $X2=0 $Y2=0
cc_257 N_B_c_292_n N_A_M1000_g 0.00684541f $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_258 N_B_c_301_n N_A_M1000_g 0.0012153f $X=3 $Y=1.74 $X2=0 $Y2=0
cc_259 N_B_c_302_n N_A_M1000_g 0.0212445f $X=3.06 $Y=1.75 $X2=0 $Y2=0
cc_260 N_B_c_292_n A 0.00455059f $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_261 N_B_M1002_g A 2.66956e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_262 N_B_c_292_n A 0.0103042f $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_263 N_B_c_294_n A 0.00369869f $X=3.295 $Y=0.81 $X2=0 $Y2=0
cc_264 B A 0.0111024f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_265 N_B_c_301_n A 0.0594272f $X=3 $Y=1.74 $X2=0 $Y2=0
cc_266 N_B_c_302_n A 0.00767616f $X=3.06 $Y=1.75 $X2=0 $Y2=0
cc_267 N_B_c_292_n N_A_c_379_n 0.0214366f $X=3.06 $Y=1.575 $X2=0 $Y2=0
cc_268 N_B_c_294_n N_A_c_379_n 0.00122993f $X=3.295 $Y=0.81 $X2=0 $Y2=0
cc_269 N_B_M1009_g N_VPWR_c_478_n 0.00585385f $X=3.215 $Y=2.275 $X2=0 $Y2=0
cc_270 N_B_M1001_g N_VPWR_c_476_n 0.0101036f $X=1.805 $Y=2.275 $X2=0 $Y2=0
cc_271 N_B_M1009_g N_VPWR_c_476_n 0.01139f $X=3.215 $Y=2.275 $X2=0 $Y2=0
cc_272 N_B_c_302_n N_VPWR_c_476_n 4.7105e-19 $X=3.06 $Y=1.75 $X2=0 $Y2=0
cc_273 B N_VPWR_c_476_n 0.0109814f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_274 N_B_M1001_g N_VPWR_c_483_n 0.00544863f $X=1.805 $Y=2.275 $X2=0 $Y2=0
cc_275 B N_VPWR_c_483_n 0.0121947f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_276 N_B_M1009_g N_VPWR_c_484_n 0.00233344f $X=3.215 $Y=2.275 $X2=0 $Y2=0
cc_277 N_B_c_301_n N_VPWR_c_484_n 0.0244055f $X=3 $Y=1.74 $X2=0 $Y2=0
cc_278 N_B_c_302_n N_VPWR_c_484_n 0.00569434f $X=3.06 $Y=1.75 $X2=0 $Y2=0
cc_279 B A_376_413# 0.00776224f $X=2.07 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_280 N_B_M1002_g N_VGND_c_565_n 0.00853463f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_281 N_B_M1002_g N_VGND_c_568_n 0.00339367f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_282 N_B_c_293_n N_VGND_c_569_n 0.00436487f $X=3.295 $Y=0.735 $X2=0 $Y2=0
cc_283 N_B_c_294_n N_VGND_c_569_n 9.28424e-19 $X=3.295 $Y=0.81 $X2=0 $Y2=0
cc_284 N_B_M1002_g N_VGND_c_571_n 0.00401529f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_285 N_B_c_293_n N_VGND_c_571_n 0.007316f $X=3.295 $Y=0.735 $X2=0 $Y2=0
cc_286 N_B_c_294_n N_VGND_c_571_n 4.54057e-19 $X=3.295 $Y=0.81 $X2=0 $Y2=0
cc_287 N_B_M1002_g N_A_297_47#_c_634_n 0.0107229f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_288 N_B_c_294_n N_A_297_47#_c_634_n 6.87069e-19 $X=3.295 $Y=0.81 $X2=0 $Y2=0
cc_289 N_A_M1000_g N_VPWR_c_477_n 0.00165904f $X=3.655 $Y=2.275 $X2=0 $Y2=0
cc_290 N_A_M1000_g N_VPWR_c_478_n 0.00585385f $X=3.655 $Y=2.275 $X2=0 $Y2=0
cc_291 N_A_M1007_g N_VPWR_c_476_n 0.011637f $X=2.355 $Y=2.275 $X2=0 $Y2=0
cc_292 N_A_M1000_g N_VPWR_c_476_n 0.00620294f $X=3.655 $Y=2.275 $X2=0 $Y2=0
cc_293 N_A_M1007_g N_VPWR_c_483_n 0.00468308f $X=2.355 $Y=2.275 $X2=0 $Y2=0
cc_294 N_A_M1007_g N_VPWR_c_484_n 0.00388256f $X=2.355 $Y=2.275 $X2=0 $Y2=0
cc_295 N_A_M1000_g COUT 6.63503e-19 $X=3.655 $Y=2.275 $X2=0 $Y2=0
cc_296 N_A_M1006_g N_COUT_c_543_n 8.90179e-19 $X=3.655 $Y=0.445 $X2=0 $Y2=0
cc_297 N_A_M1008_g N_VGND_c_565_n 0.0112612f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_M1006_g N_VGND_c_566_n 0.00302106f $X=3.655 $Y=0.445 $X2=0 $Y2=0
cc_299 N_A_M1008_g N_VGND_c_569_n 0.00339367f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_300 N_A_M1006_g N_VGND_c_569_n 0.00436487f $X=3.655 $Y=0.445 $X2=0 $Y2=0
cc_301 N_A_M1008_g N_VGND_c_571_n 0.00536411f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_302 N_A_M1006_g N_VGND_c_571_n 0.00586581f $X=3.655 $Y=0.445 $X2=0 $Y2=0
cc_303 N_A_M1008_g N_A_297_47#_c_634_n 0.0119639f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_304 N_A_c_376_n N_A_297_47#_c_634_n 5.41705e-19 $X=2.355 $Y=1.565 $X2=0 $Y2=0
cc_305 N_SUM_M1011_s N_VPWR_c_476_n 0.00212516f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_306 SUM N_VPWR_c_476_n 0.0122965f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_307 SUM N_VPWR_c_481_n 0.016214f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_308 N_SUM_c_457_n N_VGND_c_567_n 0.0154152f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_309 N_SUM_M1012_s N_VGND_c_571_n 0.0021362f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_310 N_SUM_c_457_n N_VGND_c_571_n 0.012194f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_311 N_VPWR_c_476_n A_376_413# 0.00767593f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_312 N_VPWR_c_476_n N_COUT_M1013_d 0.00212516f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_313 N_VPWR_c_479_n COUT 0.0164862f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_476_n COUT 0.0124843f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_315 N_COUT_c_543_n N_VGND_c_570_n 0.015624f $X=4.34 $Y=0.4 $X2=0 $Y2=0
cc_316 N_COUT_M1010_d N_VGND_c_571_n 0.0021362f $X=4.205 $Y=0.235 $X2=0 $Y2=0
cc_317 N_COUT_c_543_n N_VGND_c_571_n 0.0123641f $X=4.34 $Y=0.4 $X2=0 $Y2=0
cc_318 N_VGND_c_571_n N_A_297_47#_M1003_d 0.00416801f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_319 N_VGND_c_571_n N_A_297_47#_M1008_d 0.003754f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_568_n N_A_297_47#_c_649_n 0.00701792f $X=1.875 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_571_n N_A_297_47#_c_649_n 0.00608739f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_M1002_d N_A_297_47#_c_634_n 0.00159539f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_VGND_c_565_n N_A_297_47#_c_634_n 0.0159625f $X=2.04 $Y=0.38 $X2=0 $Y2=0
cc_324 N_VGND_c_568_n N_A_297_47#_c_634_n 0.00243651f $X=1.875 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_569_n N_A_297_47#_c_634_n 0.00243651f $X=3.755 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_571_n N_A_297_47#_c_634_n 0.00990569f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_569_n N_A_297_47#_c_642_n 0.00713694f $X=3.755 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_571_n N_A_297_47#_c_642_n 0.00608739f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_571_n A_674_47# 0.00269901f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24

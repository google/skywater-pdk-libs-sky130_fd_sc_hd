* File: sky130_fd_sc_hd__einvn_1.pxi.spice
* Created: Thu Aug 27 14:20:08 2020
* 
x_PM_SKY130_FD_SC_HD__EINVN_1%TE_B N_TE_B_M1005_g N_TE_B_c_42_n N_TE_B_M1002_g
+ N_TE_B_c_43_n N_TE_B_c_48_n N_TE_B_M1000_g TE_B TE_B N_TE_B_c_44_n
+ PM_SKY130_FD_SC_HD__EINVN_1%TE_B
x_PM_SKY130_FD_SC_HD__EINVN_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1002_s
+ N_A_27_47#_M1003_g N_A_27_47#_c_80_n N_A_27_47#_c_86_n N_A_27_47#_c_81_n
+ N_A_27_47#_c_82_n N_A_27_47#_c_95_n N_A_27_47#_c_87_n N_A_27_47#_c_83_n
+ N_A_27_47#_c_84_n N_A_27_47#_c_115_p N_A_27_47#_c_89_n N_A_27_47#_c_85_n
+ PM_SKY130_FD_SC_HD__EINVN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVN_1%A N_A_c_139_n N_A_M1001_g N_A_M1004_g A A A
+ N_A_c_141_n PM_SKY130_FD_SC_HD__EINVN_1%A
x_PM_SKY130_FD_SC_HD__EINVN_1%VPWR N_VPWR_M1002_d N_VPWR_c_168_n VPWR
+ N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_167_n N_VPWR_c_172_n
+ PM_SKY130_FD_SC_HD__EINVN_1%VPWR
x_PM_SKY130_FD_SC_HD__EINVN_1%Z N_Z_M1001_d N_Z_M1004_d Z Z Z Z
+ PM_SKY130_FD_SC_HD__EINVN_1%Z
x_PM_SKY130_FD_SC_HD__EINVN_1%VGND N_VGND_M1005_d VGND N_VGND_c_232_n
+ N_VGND_c_233_n N_VGND_c_234_n N_VGND_c_235_n PM_SKY130_FD_SC_HD__EINVN_1%VGND
cc_1 VNB N_TE_B_M1005_g 0.0416983f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_TE_B_c_42_n 0.0294103f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.41
cc_3 VNB N_TE_B_c_43_n 0.0165134f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.335
cc_4 VNB N_TE_B_c_44_n 0.0164024f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_5 VNB N_A_27_47#_c_80_n 0.0141471f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.985
cc_6 VNB N_A_27_47#_c_81_n 0.0010873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_82_n 0.00995565f $X=-0.19 $Y=-0.24 $X2=0.407 $Y2=1.16
cc_8 VNB N_A_27_47#_c_83_n 0.00569771f $X=-0.19 $Y=-0.24 $X2=0.297 $Y2=1.19
cc_9 VNB N_A_27_47#_c_84_n 0.029031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_85_n 0.0184211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_139_n 0.0192724f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_12 VNB A 0.0205666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_c_141_n 0.0344588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_167_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0.407 $Y2=1.335
cc_15 VNB Z 0.00247112f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.335
cc_16 VNB Z 0.0149239f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.41
cc_17 VNB N_VGND_c_232_n 0.0227443f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.985
cc_18 VNB N_VGND_c_233_n 0.14235f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_VGND_c_234_n 0.014818f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_20 VNB N_VGND_c_235_n 0.0184163f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_TE_B_c_42_n 0.00850781f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.41
cc_22 VPB N_TE_B_M1002_g 0.0430975f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_23 VPB N_TE_B_c_43_n 0.0119894f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.335
cc_24 VPB N_TE_B_c_48_n 0.0178796f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.41
cc_25 VPB N_TE_B_c_44_n 0.0201207f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_26 VPB N_A_27_47#_c_86_n 0.0156843f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_27 VPB N_A_27_47#_c_87_n 0.0076959f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_28 VPB N_A_27_47#_c_84_n 0.0103109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_27_47#_c_89_n 0.0015164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_M1004_g 0.0263993f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_31 VPB A 0.0127322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_c_141_n 0.00992195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_168_n 0.00294119f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_34 VPB N_VPWR_c_169_n 0.0148836f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.335
cc_35 VPB N_VPWR_c_170_n 0.0364623f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_36 VPB N_VPWR_c_167_n 0.0438487f $X=-0.19 $Y=1.305 $X2=0.407 $Y2=1.335
cc_37 VPB N_VPWR_c_172_n 0.00522083f $X=-0.19 $Y=1.305 $X2=0.297 $Y2=1.19
cc_38 VPB Z 0.00131752f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.335
cc_39 VPB Z 0.0296293f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.985
cc_40 N_TE_B_M1005_g N_A_27_47#_c_81_n 0.0157631f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_41 N_TE_B_c_43_n N_A_27_47#_c_81_n 0.00392316f $X=0.87 $Y=1.335 $X2=0 $Y2=0
cc_42 N_TE_B_c_44_n N_A_27_47#_c_81_n 0.0107574f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_43 N_TE_B_c_42_n N_A_27_47#_c_82_n 6.91349e-19 $X=0.47 $Y=1.41 $X2=0 $Y2=0
cc_44 N_TE_B_c_44_n N_A_27_47#_c_82_n 0.0261211f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_45 N_TE_B_M1002_g N_A_27_47#_c_95_n 0.0126027f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_46 N_TE_B_c_43_n N_A_27_47#_c_95_n 0.00121726f $X=0.87 $Y=1.335 $X2=0 $Y2=0
cc_47 N_TE_B_c_48_n N_A_27_47#_c_95_n 0.00165029f $X=0.945 $Y=1.41 $X2=0 $Y2=0
cc_48 N_TE_B_c_44_n N_A_27_47#_c_95_n 0.0098503f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_49 N_TE_B_c_42_n N_A_27_47#_c_87_n 2.97054e-19 $X=0.47 $Y=1.41 $X2=0 $Y2=0
cc_50 N_TE_B_c_44_n N_A_27_47#_c_87_n 0.0244556f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_51 N_TE_B_M1005_g N_A_27_47#_c_83_n 0.00557175f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_52 N_TE_B_c_44_n N_A_27_47#_c_83_n 0.0622599f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_53 N_TE_B_c_42_n N_A_27_47#_c_84_n 0.002621f $X=0.47 $Y=1.41 $X2=0 $Y2=0
cc_54 N_TE_B_c_43_n N_A_27_47#_c_84_n 0.0042336f $X=0.87 $Y=1.335 $X2=0 $Y2=0
cc_55 N_TE_B_c_42_n N_A_27_47#_c_89_n 0.00557175f $X=0.47 $Y=1.41 $X2=0 $Y2=0
cc_56 N_TE_B_M1002_g N_A_27_47#_c_89_n 0.00599241f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_57 N_TE_B_c_43_n N_A_27_47#_c_89_n 0.0194212f $X=0.87 $Y=1.335 $X2=0 $Y2=0
cc_58 N_TE_B_c_48_n N_A_27_47#_c_89_n 0.0170018f $X=0.945 $Y=1.41 $X2=0 $Y2=0
cc_59 N_TE_B_M1002_g N_VPWR_c_168_n 0.00697722f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_60 N_TE_B_c_48_n N_VPWR_c_168_n 0.00322148f $X=0.945 $Y=1.41 $X2=0 $Y2=0
cc_61 N_TE_B_M1002_g N_VPWR_c_169_n 0.00413026f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_62 N_TE_B_c_48_n N_VPWR_c_170_n 0.00583607f $X=0.945 $Y=1.41 $X2=0 $Y2=0
cc_63 N_TE_B_M1002_g N_VPWR_c_167_n 0.00573844f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_64 N_TE_B_c_48_n N_VPWR_c_167_n 0.0119966f $X=0.945 $Y=1.41 $X2=0 $Y2=0
cc_65 N_TE_B_c_43_n Z 8.72145e-19 $X=0.87 $Y=1.335 $X2=0 $Y2=0
cc_66 N_TE_B_c_48_n Z 0.00374975f $X=0.945 $Y=1.41 $X2=0 $Y2=0
cc_67 N_TE_B_M1005_g N_VGND_c_233_n 0.00562917f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_68 N_TE_B_M1005_g N_VGND_c_234_n 0.00407353f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_69 N_TE_B_M1005_g N_VGND_c_235_n 0.00835269f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_27_47#_c_83_n N_A_c_139_n 4.01394e-19 $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_71 N_A_27_47#_c_85_n N_A_c_139_n 0.0326628f $X=1.387 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_27_47#_c_89_n N_A_M1004_g 0.00167204f $X=1.067 $Y=1.615 $X2=0 $Y2=0
cc_73 N_A_27_47#_c_83_n N_A_c_141_n 2.71115e-19 $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_84_n N_A_c_141_n 0.0203629f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_95_n N_VPWR_M1002_d 0.00503058f $X=0.685 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_27_47#_c_115_p N_VPWR_M1002_d 0.0033419f $X=0.777 $Y=1.895 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_27_47#_c_89_n N_VPWR_M1002_d 0.00113704f $X=1.067 $Y=1.615 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_27_47#_c_95_n N_VPWR_c_168_n 0.0173986f $X=0.685 $Y=1.98 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_86_n N_VPWR_c_169_n 0.0186589f $X=0.227 $Y=2.065 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_95_n N_VPWR_c_169_n 0.00248249f $X=0.685 $Y=1.98 $X2=0 $Y2=0
cc_81 N_A_27_47#_M1002_s N_VPWR_c_167_n 0.00219164f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_82 N_A_27_47#_c_86_n N_VPWR_c_167_n 0.0108489f $X=0.227 $Y=2.065 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_95_n N_VPWR_c_167_n 0.00554215f $X=0.685 $Y=1.98 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_89_n A_204_297# 0.00683858f $X=1.067 $Y=1.615 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_27_47#_c_83_n Z 0.0633001f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_84_n Z 0.00210987f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_85_n Z 0.00162044f $X=1.387 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_85_n Z 0.00469892f $X=1.387 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_84_n Z 0.00402899f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_89_n Z 0.0333849f $X=1.067 $Y=1.615 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_81_n N_VGND_M1005_d 0.0110485f $X=0.685 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_27_47#_c_83_n N_VGND_M1005_d 0.00319369f $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_27_47#_M1005_s N_VGND_c_233_n 0.00217724f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_80_n N_VGND_c_233_n 0.0108288f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_81_n N_VGND_c_233_n 0.00899476f $X=0.685 $Y=0.7 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_80_n N_VGND_c_234_n 0.0185662f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_81_n N_VGND_c_234_n 0.00272761f $X=0.685 $Y=0.7 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_81_n N_VGND_c_235_n 0.0630544f $X=0.685 $Y=0.7 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_85_n N_VGND_c_235_n 0.0192481f $X=1.387 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_M1004_g N_VPWR_c_170_n 0.00357877f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_M1004_g N_VPWR_c_167_n 0.00755644f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_102 A N_Z_M1001_d 0.00356078f $X=1.98 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_103 A N_Z_M1004_d 0.00430356f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A_c_139_n Z 0.0134264f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_M1004_g Z 0.01863f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_106 A Z 0.0611504f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_107 N_A_c_141_n Z 0.00763089f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_c_139_n Z 0.0139163f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_109 A Z 0.0201989f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_110 N_A_c_141_n Z 0.00215351f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_M1004_g Z 0.0325596f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_112 A Z 0.0219813f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_113 N_A_c_141_n Z 0.00206064f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_139_n N_VGND_c_232_n 0.00357877f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_139_n N_VGND_c_233_n 0.00634206f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_c_139_n N_VGND_c_235_n 0.00200069f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_117 N_VPWR_c_167_n A_204_297# 0.00666001f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_118 N_VPWR_c_167_n N_Z_M1004_d 0.00209344f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_119 N_VPWR_c_170_n Z 0.07654f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_120 N_VPWR_c_167_n Z 0.0444626f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_121 A_204_297# Z 0.00436656f $X=1.02 $Y=1.485 $X2=1.355 $Y2=0.56
cc_122 A_204_297# Z 0.0338836f $X=1.02 $Y=1.485 $X2=0.26 $Y2=0.445
cc_123 Z N_VGND_c_232_n 0.0357203f $X=1.98 $Y=0.425 $X2=0 $Y2=0
cc_124 N_Z_M1001_d N_VGND_c_233_n 0.00209344f $X=1.905 $Y=0.235 $X2=0 $Y2=0
cc_125 Z N_VGND_c_233_n 0.0217513f $X=1.98 $Y=0.425 $X2=0 $Y2=0
cc_126 Z A_286_47# 0.00273439f $X=1.52 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_127 Z A_286_47# 0.00470202f $X=1.98 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_128 N_VGND_c_233_n A_286_47# 0.00844528f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24

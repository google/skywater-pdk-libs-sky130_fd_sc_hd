* File: sky130_fd_sc_hd__a32oi_4.spice
* Created: Thu Aug 27 14:05:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a32oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a32oi_4  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1014 N_A_27_47#_M1014_d N_B2_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1021 N_A_27_47#_M1021_d N_B2_M1021_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1025 N_A_27_47#_M1021_d N_B2_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1038 N_A_27_47#_M1038_d N_B2_M1038_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1022 N_Y_M1022_d N_B1_M1022_g N_A_27_47#_M1038_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1028 N_Y_M1022_d N_B1_M1028_g N_A_27_47#_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1032 N_Y_M1032_d N_B1_M1032_g N_A_27_47#_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1033 N_Y_M1032_d N_B1_M1033_g N_A_27_47#_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_803_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1013_d N_A1_M1015_g N_A_803_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1023_d N_A1_M1023_g N_A_803_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1029 N_Y_M1023_d N_A1_M1029_g N_A_803_47#_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.13325 PD=0.92 PS=1.06 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1016 N_A_803_47#_M1029_s N_A2_M1016_g N_A_1249_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13325 AS=0.08775 PD=1.06 PS=0.92 NRD=24.912 NRS=0 M=1 R=4.33333
+ SA=75002 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1018 N_A_803_47#_M1018_d N_A2_M1018_g N_A_1249_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.4 SB=75001 A=0.0975 P=1.6 MULT=1
MM1026 N_A_803_47#_M1018_d N_A2_M1026_g N_A_1249_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.8 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1030 N_A_803_47#_M1030_d N_A2_M1030_g N_A_1249_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A3_M1009_g N_A_1249_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A3_M1011_g N_A_1249_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1011_d N_A3_M1017_g N_A_1249_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A3_M1019_g N_A_1249_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75009.3 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1002_d N_B2_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75008.9 A=0.15 P=2.3 MULT=1
MM1027 N_Y_M1027_d N_B2_M1027_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75008.5 A=0.15 P=2.3 MULT=1
MM1034 N_Y_M1027_d N_B2_M1034_g N_A_27_297#_M1034_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75008.1 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_A_27_297#_M1034_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75007.7 A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1000_d N_B1_M1006_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75007.2 A=0.15 P=2.3 MULT=1
MM1031 N_Y_M1031_d N_B1_M1031_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75006.8 A=0.15 P=2.3 MULT=1
MM1035 N_Y_M1031_d N_B1_M1035_g N_A_27_297#_M1035_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75006.4 A=0.15 P=2.3 MULT=1
MM1004 N_A_27_297#_M1035_s N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.135 PD=1.29 PS=1.27 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75006 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_297#_M1008_d N_A1_M1008_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75005.5 A=0.15 P=2.3 MULT=1
MM1012 N_A_27_297#_M1008_d N_A1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.3375 PD=1.27 PS=1.675 NRD=0 NRS=5.8903 M=1 R=6.66667 SA=75004.4
+ SB=75005.1 A=0.15 P=2.3 MULT=1
MM1039 N_A_27_297#_M1039_d N_A1_M1039_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2525 AS=0.3375 PD=1.505 PS=1.675 NRD=0 NRS=4.9053 M=1 R=6.66667
+ SA=75005.2 SB=75004.3 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_27_297#_M1039_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.2525 PD=1.27 PS=1.505 NRD=0 NRS=45.2903 M=1 R=6.66667 SA=75005.9
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1003_d N_A2_M1024_g N_A_27_297#_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.3
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1036 N_VPWR_M1036_d N_A2_M1036_g N_A_27_297#_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.7
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1037 N_VPWR_M1036_d N_A2_M1037_g N_A_27_297#_M1037_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.395 PD=1.27 PS=1.79 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.1
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1001 N_A_27_297#_M1037_s N_A3_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.395 AS=0.135 PD=1.79 PS=1.27 NRD=101.435 NRS=0 M=1 R=6.66667 SA=75008.1
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_297#_M1007_d N_A3_M1007_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1010 N_A_27_297#_M1007_d N_A3_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_A_27_297#_M1020_d N_A3_M1020_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.8525 P=24.21
*
.include "sky130_fd_sc_hd__a32oi_4.pxi.spice"
*
.ends
*
*

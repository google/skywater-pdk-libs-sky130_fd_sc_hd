* File: sky130_fd_sc_hd__o2111a_1.spice
* Created: Thu Aug 27 14:33:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2111a_1.pex.spice"
.subckt sky130_fd_sc_hd__o2111a_1  VNB VPB D1 C1 B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_79_21#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 A_306_47# N_D1_M1004_g N_A_79_21#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.19825 PD=1.015 PS=1.91 NRD=23.532 NRS=7.38 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1005 A_409_47# N_C1_M1005_g A_306_47# VNB NSHORT L=0.15 W=0.65 AD=0.118625
+ AS=0.118625 PD=1.015 PS=1.015 NRD=23.532 NRS=23.532 M=1 R=4.33333 SA=75000.7
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_A_512_47#_M1001_d N_B1_M1001_g A_409_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.118625 PD=1.26 PS=1.015 NRD=61.836 NRS=23.532 M=1 R=4.33333
+ SA=75001.3 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_512_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.19825 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_512_47#_M1009_d N_A1_M1009_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.08775 PD=1.83 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_A_79_21#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3825 AS=0.26 PD=1.765 PS=2.52 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1008 N_A_79_21#_M1008_d N_D1_M1008_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.2175 AS=0.3825 PD=1.435 PS=1.765 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75001.1 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_C1_M1002_g N_A_79_21#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.305 AS=0.2175 PD=1.61 PS=1.435 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75001.7
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_A_79_21#_M1006_d N_B1_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.2125 AS=0.305 PD=1.425 PS=1.61 NRD=29.55 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 A_676_297# N_A2_M1000_g N_A_79_21#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.2125 PD=1.21 PS=1.425 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75003
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_676_297# VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75003.4 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_64 VPB 0 1.11775e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__o2111a_1.pxi.spice"
*
.ends
*
*

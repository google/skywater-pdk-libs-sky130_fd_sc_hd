* File: sky130_fd_sc_hd__einvn_4.spice.pex
* Created: Thu Aug 27 14:20:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVN_4%TE_B 1 3 6 8 10 12 13 15 17 18 20 22 23 25
+ 27 28 31 32 33 40
c79 32 0 7.37964e-20 $X=1.785 $Y=1.395
c80 31 0 7.37964e-20 $X=1.365 $Y=1.395
c81 28 0 2.52753e-20 $X=0.945 $Y=1.25
c82 23 0 2.02538e-19 $X=2.13 $Y=1.395
c83 18 0 1.51809e-19 $X=1.71 $Y=1.395
c84 6 0 1.13048e-19 $X=0.47 $Y=1.985
r85 39 40 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.545 $Y2=1.16
r86 36 39 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r87 33 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r88 28 30 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.945 $Y=1.25
+ $X2=0.945 $Y2=1.395
r89 25 27 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.205 $Y=1.47
+ $X2=2.205 $Y2=2.015
r90 24 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.86 $Y=1.395
+ $X2=1.785 $Y2=1.395
r91 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.13 $Y=1.395
+ $X2=2.205 $Y2=1.47
r92 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.13 $Y=1.395
+ $X2=1.86 $Y2=1.395
r93 20 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.785 $Y=1.47
+ $X2=1.785 $Y2=1.395
r94 20 22 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.785 $Y=1.47
+ $X2=1.785 $Y2=2.015
r95 19 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.44 $Y=1.395
+ $X2=1.365 $Y2=1.395
r96 18 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=1.395
+ $X2=1.785 $Y2=1.395
r97 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.71 $Y=1.395
+ $X2=1.44 $Y2=1.395
r98 15 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.365 $Y=1.47
+ $X2=1.365 $Y2=1.395
r99 15 17 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.365 $Y=1.47
+ $X2=1.365 $Y2=2.015
r100 14 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.395
+ $X2=0.945 $Y2=1.395
r101 13 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.395
+ $X2=1.365 $Y2=1.395
r102 13 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.29 $Y=1.395
+ $X2=1.02 $Y2=1.395
r103 10 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=1.47
+ $X2=0.945 $Y2=1.395
r104 10 12 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.945 $Y=1.47
+ $X2=0.945 $Y2=2.015
r105 8 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.25
+ $X2=0.945 $Y2=1.25
r106 8 40 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.87 $Y=1.25
+ $X2=0.545 $Y2=1.25
r107 4 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r108 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r109 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r110 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 26 27 32 34 35 37 40 51 52
c102 25 0 8.8865e-20 $X=1.83 $Y=1.035
c103 15 0 1.87534e-19 $X=2.175 $Y=1.035
c104 10 0 9.82445e-20 $X=1.755 $Y=1.035
r105 41 52 22.4813 $w=2.68e-07 $l=1.25e-07 $layer=POLY_cond $X=2.625 $Y=1.16
+ $X2=2.625 $Y2=1.035
r106 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.16 $X2=2.625 $Y2=1.16
r107 38 51 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=0.68 $Y2=1.16
r108 38 40 62.1621 $w=3.28e-07 $l=1.78e-06 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=2.625 $Y2=1.16
r109 36 51 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=1.16
r110 36 37 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=1.495
r111 35 51 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.995
+ $X2=0.68 $Y2=1.16
r112 34 35 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=0.825
+ $X2=0.68 $Y2=0.995
r113 30 37 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.215 $Y=1.58
+ $X2=0.68 $Y2=1.58
r114 30 32 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.215 $Y=1.665
+ $X2=0.215 $Y2=1.815
r115 27 34 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.215 $Y=0.74
+ $X2=0.68 $Y2=0.74
r116 27 29 4.45769 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.56
r117 22 52 22.7584 $w=2.68e-07 $l=9.48683e-08 $layer=POLY_cond $X=2.67 $Y=0.96
+ $X2=2.625 $Y2=1.035
r118 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.67 $Y=0.96 $X2=2.67
+ $Y2=0.56
r119 21 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.325 $Y=1.035
+ $X2=2.25 $Y2=1.035
r120 20 52 16.3317 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.49 $Y=1.035
+ $X2=2.625 $Y2=1.035
r121 20 21 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.035
+ $X2=2.325 $Y2=1.035
r122 17 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=0.96
+ $X2=2.25 $Y2=1.035
r123 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.25 $Y=0.96 $X2=2.25
+ $Y2=0.56
r124 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.035
+ $X2=1.83 $Y2=1.035
r125 15 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.175 $Y=1.035
+ $X2=2.25 $Y2=1.035
r126 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.175 $Y=1.035
+ $X2=1.905 $Y2=1.035
r127 12 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=0.96
+ $X2=1.83 $Y2=1.035
r128 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.83 $Y=0.96 $X2=1.83
+ $Y2=0.56
r129 10 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.035
+ $X2=1.83 $Y2=1.035
r130 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.755 $Y=1.035
+ $X2=1.485 $Y2=1.035
r131 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=0.96
+ $X2=1.485 $Y2=1.035
r132 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.41 $Y=0.96 $X2=1.41
+ $Y2=0.56
r133 2 32 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.815
r134 1 29 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 35 36
+ 40
r69 36 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=1.16 $X2=4.82 $Y2=1.16
r70 35 36 8.02825 $w=4.43e-07 $l=3.1e-07 $layer=LI1_cond $X=4.752 $Y=0.85
+ $X2=4.752 $Y2=1.16
r71 33 34 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.985 $Y=1.16
+ $X2=4.405 $Y2=1.16
r72 32 33 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.565 $Y=1.16
+ $X2=3.985 $Y2=1.16
r73 30 32 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.145 $Y=1.16
+ $X2=3.565 $Y2=1.16
r74 29 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.48 $Y=1.16
+ $X2=4.82 $Y2=1.16
r75 29 34 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.48 $Y=1.16
+ $X2=4.405 $Y2=1.16
r76 25 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.325
+ $X2=4.405 $Y2=1.16
r77 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.405 $Y=1.325
+ $X2=4.405 $Y2=1.985
r78 22 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=0.995
+ $X2=4.405 $Y2=1.16
r79 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.405 $Y=0.995
+ $X2=4.405 $Y2=0.56
r80 18 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.325
+ $X2=3.985 $Y2=1.16
r81 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.985 $Y=1.325
+ $X2=3.985 $Y2=1.985
r82 15 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=0.995
+ $X2=3.985 $Y2=1.16
r83 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.985 $Y=0.995
+ $X2=3.985 $Y2=0.56
r84 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.16
r85 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.985
r86 8 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=1.16
r87 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=0.56
r88 4 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=1.16
r89 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=1.985
r90 1 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=1.16
r91 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%VPWR 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r69 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r71 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r73 42 45 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r74 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 41 44 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 39 54 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.64 $Y=2.72
+ $X2=2.445 $Y2=2.72
r78 39 41 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.64 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r82 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=1.575 $Y2=2.72
r83 35 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=2.07 $Y2=2.72
r84 34 54 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.445 $Y2=2.72
r85 34 37 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.07 $Y2=2.72
r86 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r87 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r90 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.575 $Y2=2.72
r92 29 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r93 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r94 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 18 54 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=2.635
+ $X2=2.445 $Y2=2.72
r98 18 20 18.7641 $w=3.88e-07 $l=6.35e-07 $layer=LI1_cond $X=2.445 $Y=2.635
+ $X2=2.445 $Y2=2
r99 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.72
r100 14 16 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.02
r101 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r102 10 12 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.02
r103 3 20 300 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=2 $X=2.28
+ $Y=1.545 $X2=2.415 $Y2=2
r104 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.44
+ $Y=1.545 $X2=1.575 $Y2=2.02
r105 1 12 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%A_204_309# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 42 44 45
c61 26 0 1.87534e-19 $X=2.81 $Y=1.58
c62 21 0 1.13048e-19 $X=1.24 $Y=1.58
c63 20 0 1.8711e-19 $X=1.91 $Y=1.58
r64 40 42 12.4308 $w=4.43e-07 $l=4.8e-07 $layer=LI1_cond $X=4.752 $Y=2.295
+ $X2=4.752 $Y2=1.815
r65 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=2.38
+ $X2=3.775 $Y2=2.38
r66 38 40 8.76165 $w=1.7e-07 $l=2.61063e-07 $layer=LI1_cond $X=4.53 $Y=2.38
+ $X2=4.752 $Y2=2.295
r67 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.53 $Y=2.38
+ $X2=3.86 $Y2=2.38
r68 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=2.295
+ $X2=3.775 $Y2=2.38
r69 34 36 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.775 $Y=2.295
+ $X2=3.775 $Y2=1.815
r70 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.38
+ $X2=3.775 $Y2=2.38
r71 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.69 $Y=2.38
+ $X2=3.02 $Y2=2.38
r72 29 33 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.915 $Y=2.295
+ $X2=3.02 $Y2=2.38
r73 29 31 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=2.915 $Y=2.295
+ $X2=2.915 $Y2=1.815
r74 28 31 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.915 $Y=1.665
+ $X2=2.915 $Y2=1.815
r75 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.58
+ $X2=1.995 $Y2=1.58
r76 26 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.81 $Y=1.58
+ $X2=2.915 $Y2=1.665
r77 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.81 $Y=1.58
+ $X2=2.08 $Y2=1.58
r78 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=1.665
+ $X2=1.995 $Y2=1.58
r79 22 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.995 $Y=1.665
+ $X2=1.995 $Y2=1.815
r80 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=1.58
+ $X2=1.995 $Y2=1.58
r81 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.91 $Y=1.58
+ $X2=1.24 $Y2=1.58
r82 16 21 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.127 $Y=1.665
+ $X2=1.24 $Y2=1.58
r83 16 18 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.127 $Y=1.665
+ $X2=1.127 $Y2=1.815
r84 5 42 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=1.485 $X2=4.615 $Y2=1.815
r85 4 36 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=3.64
+ $Y=1.485 $X2=3.775 $Y2=1.815
r86 3 31 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.485 $X2=2.935 $Y2=1.815
r87 2 24 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.545 $X2=1.995 $Y2=1.815
r88 1 18 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.545 $X2=1.155 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%Z 1 2 3 4 15 19 21 23 39
r39 23 39 3.97209 $w=8.58e-07 $l=2.8e-07 $layer=LI1_cond $X=3.915 $Y=1.05
+ $X2=4.195 $Y2=1.05
r40 21 23 6.52558 $w=8.58e-07 $l=4.6e-07 $layer=LI1_cond $X=3.455 $Y=1.05
+ $X2=3.915 $Y2=1.05
r41 21 30 1.4186 $w=8.58e-07 $l=1e-07 $layer=LI1_cond $X=3.455 $Y=1.05 $X2=3.355
+ $Y2=1.05
r42 17 39 6.40395 $w=3.3e-07 $l=4.3e-07 $layer=LI1_cond $X=4.195 $Y=1.48
+ $X2=4.195 $Y2=1.05
r43 17 19 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.195 $Y=1.48
+ $X2=4.195 $Y2=1.61
r44 13 30 6.40395 $w=3.3e-07 $l=4.3e-07 $layer=LI1_cond $X=3.355 $Y=1.48
+ $X2=3.355 $Y2=1.05
r45 13 15 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.355 $Y=1.48
+ $X2=3.355 $Y2=1.61
r46 4 19 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=4.06
+ $Y=1.485 $X2=4.195 $Y2=1.61
r47 3 15 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.485 $X2=3.355 $Y2=1.61
r48 2 39 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.195 $Y2=0.74
r49 1 30 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.235 $X2=3.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r74 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r75 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r76 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r77 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r78 42 45 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=4.83
+ $Y2=0
r79 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r80 41 44 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.83
+ $Y2=0
r81 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r82 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.46
+ $Y2=0
r83 39 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.99
+ $Y2=0
r84 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r85 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r86 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r87 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r88 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.07
+ $Y2=0
r89 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.46
+ $Y2=0
r90 34 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.07
+ $Y2=0
r91 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r92 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r93 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r94 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r95 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r96 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r97 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.15
+ $Y2=0
r98 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r99 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r100 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r101 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r102 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r103 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.36
r104 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r105 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.36
r106 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r107 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r108 3 20 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.36
r109 2 16 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.36
r110 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_4%A_215_47# 1 2 3 4 5 16 19 20 21 24 29 30 34
+ 36
c61 36 0 1.50694e-19 $X=2.04 $Y=0.74
c62 24 0 5.18434e-20 $X=2.825 $Y=0.74
c63 20 0 2.52753e-20 $X=1.285 $Y=0.74
c64 19 0 2.99402e-19 $X=1.955 $Y=0.74
r65 32 34 47.7762 $w=1.93e-07 $l=8.4e-07 $layer=LI1_cond $X=3.775 $Y=0.352
+ $X2=4.615 $Y2=0.352
r66 30 32 44.3636 $w=1.93e-07 $l=7.8e-07 $layer=LI1_cond $X=2.995 $Y=0.352
+ $X2=3.775 $Y2=0.352
r67 27 29 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.91 $Y=0.655
+ $X2=2.91 $Y2=0.56
r68 26 30 6.85817 $w=1.95e-07 $l=1.33918e-07 $layer=LI1_cond $X=2.91 $Y=0.45
+ $X2=2.995 $Y2=0.352
r69 26 29 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.91 $Y=0.45
+ $X2=2.91 $Y2=0.56
r70 25 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=0.74
+ $X2=2.04 $Y2=0.74
r71 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.825 $Y=0.74
+ $X2=2.91 $Y2=0.655
r72 24 25 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.825 $Y=0.74
+ $X2=2.125 $Y2=0.74
r73 21 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.655
+ $X2=2.04 $Y2=0.74
r74 21 23 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.04 $Y=0.655
+ $X2=2.04 $Y2=0.56
r75 19 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=2.04 $Y2=0.74
r76 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=1.285 $Y2=0.74
r77 16 20 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.15 $Y=0.655
+ $X2=1.285 $Y2=0.74
r78 16 18 4.29259 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=0.655
+ $X2=1.15 $Y2=0.56
r79 5 34 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.235 $X2=4.615 $Y2=0.365
r80 4 32 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.775 $Y2=0.365
r81 3 29 182 $w=1.7e-07 $l=3.99061e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.91 $Y2=0.56
r82 2 23 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.56
r83 1 18 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.56
.ends


* File: sky130_fd_sc_hd__and4bb_2.pxi.spice
* Created: Thu Aug 27 14:09:09 2020
* 
x_PM_SKY130_FD_SC_HD__AND4BB_2%A_N N_A_N_M1013_g N_A_N_M1005_g A_N A_N
+ N_A_N_c_92_n PM_SKY130_FD_SC_HD__AND4BB_2%A_N
x_PM_SKY130_FD_SC_HD__AND4BB_2%A_174_21# N_A_174_21#_M1010_s N_A_174_21#_M1002_d
+ N_A_174_21#_M1006_d N_A_174_21#_c_117_n N_A_174_21#_M1003_g
+ N_A_174_21#_M1000_g N_A_174_21#_c_118_n N_A_174_21#_M1015_g
+ N_A_174_21#_M1001_g N_A_174_21#_c_119_n N_A_174_21#_c_120_n
+ N_A_174_21#_c_121_n N_A_174_21#_c_204_p N_A_174_21#_c_138_p
+ N_A_174_21#_c_122_n N_A_174_21#_c_143_p N_A_174_21#_c_129_n
+ N_A_174_21#_c_130_n N_A_174_21#_c_181_p N_A_174_21#_c_123_n
+ PM_SKY130_FD_SC_HD__AND4BB_2%A_174_21#
x_PM_SKY130_FD_SC_HD__AND4BB_2%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1005_s
+ N_A_27_47#_c_222_n N_A_27_47#_M1002_g N_A_27_47#_c_223_n N_A_27_47#_M1010_g
+ N_A_27_47#_c_305_p N_A_27_47#_c_229_n N_A_27_47#_c_224_n N_A_27_47#_c_258_n
+ N_A_27_47#_c_231_n N_A_27_47#_c_232_n N_A_27_47#_c_225_n N_A_27_47#_c_226_n
+ PM_SKY130_FD_SC_HD__AND4BB_2%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4BB_2%A_505_280# N_A_505_280#_M1008_d
+ N_A_505_280#_M1007_d N_A_505_280#_M1011_g N_A_505_280#_M1012_g
+ N_A_505_280#_c_318_n N_A_505_280#_c_319_n N_A_505_280#_c_320_n
+ N_A_505_280#_c_331_n N_A_505_280#_c_321_n N_A_505_280#_c_314_n
+ N_A_505_280#_c_323_n N_A_505_280#_c_324_n N_A_505_280#_c_315_n
+ N_A_505_280#_c_325_n PM_SKY130_FD_SC_HD__AND4BB_2%A_505_280#
x_PM_SKY130_FD_SC_HD__AND4BB_2%C N_C_M1009_g N_C_M1006_g C C C N_C_c_387_n
+ N_C_c_388_n PM_SKY130_FD_SC_HD__AND4BB_2%C
x_PM_SKY130_FD_SC_HD__AND4BB_2%D N_D_M1004_g N_D_M1014_g D D D N_D_c_427_n
+ PM_SKY130_FD_SC_HD__AND4BB_2%D
x_PM_SKY130_FD_SC_HD__AND4BB_2%B_N N_B_N_M1008_g N_B_N_M1007_g B_N B_N
+ N_B_N_c_471_n N_B_N_c_472_n PM_SKY130_FD_SC_HD__AND4BB_2%B_N
x_PM_SKY130_FD_SC_HD__AND4BB_2%VPWR N_VPWR_M1005_d N_VPWR_M1001_d N_VPWR_M1012_d
+ N_VPWR_M1014_d N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n VPWR
+ N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_505_n
+ N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ PM_SKY130_FD_SC_HD__AND4BB_2%VPWR
x_PM_SKY130_FD_SC_HD__AND4BB_2%X N_X_M1003_s N_X_M1000_s X X X N_X_c_584_n X
+ PM_SKY130_FD_SC_HD__AND4BB_2%X
x_PM_SKY130_FD_SC_HD__AND4BB_2%VGND N_VGND_M1013_d N_VGND_M1015_d N_VGND_M1004_d
+ N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n VGND N_VGND_c_609_n
+ N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n N_VGND_c_614_n
+ N_VGND_c_615_n N_VGND_c_616_n PM_SKY130_FD_SC_HD__AND4BB_2%VGND
cc_1 VNB N_A_N_M1013_g 0.0369733f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.0024619f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_92_n 0.0444604f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_174_21#_c_117_n 0.0162441f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_174_21#_c_118_n 0.0180659f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_6 VNB N_A_174_21#_c_119_n 0.00107364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_174_21#_c_120_n 0.0449654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_174_21#_c_121_n 0.00679851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_174_21#_c_122_n 0.00455999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_174_21#_c_123_n 0.00143078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_222_n 0.0570294f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_12 VNB N_A_27_47#_c_223_n 0.0169709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_224_n 0.00346791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_225_n 0.00787965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_226_n 0.00270383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_505_280#_M1011_g 0.04429f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_17 VNB N_A_505_280#_c_314_n 0.0330596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_505_280#_c_315_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_C_M1006_g 0.00965768f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_20 VNB C 0.00711595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_C_c_387_n 0.02576f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_22 VNB N_C_c_388_n 0.0166213f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_23 VNB N_D_M1004_g 0.0299741f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_24 VNB D 0.00743717f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_25 VNB N_D_c_427_n 0.0186932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B_N_M1007_g 0.0112547f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_27 VNB B_N 0.00547409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_B_N_c_471_n 0.0295815f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_29 VNB N_B_N_c_472_n 0.0205749f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_30 VNB N_VPWR_c_505_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_584_n 6.38923e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_606_n 0.00210688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_607_n 0.00547513f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_608_n 0.00237268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_609_n 0.0151362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_610_n 0.01464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_611_n 0.0589856f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_612_n 0.0150402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_613_n 0.241773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_614_n 0.00506835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_615_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_616_n 0.00353967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_A_N_M1005_g 0.0597241f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_44 VPB A_N 0.0159685f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_45 VPB N_A_N_c_92_n 0.0118271f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_46 VPB N_A_174_21#_M1000_g 0.0187091f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_47 VPB N_A_174_21#_M1001_g 0.0221938f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.53
cc_48 VPB N_A_174_21#_c_119_n 0.00227696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_174_21#_c_120_n 0.0106905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_174_21#_c_122_n 0.00492861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_174_21#_c_129_n 0.00586258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_174_21#_c_130_n 0.00485593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_222_n 0.0156104f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_54 VPB N_A_27_47#_M1002_g 0.055785f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_55 VPB N_A_27_47#_c_229_n 9.19263e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_224_n 0.00160467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_231_n 0.0112733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_232_n 0.00301495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_226_n 3.66935e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_505_280#_M1011_g 0.00519402f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_61 VPB N_A_505_280#_M1012_g 0.0272104f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_62 VPB N_A_505_280#_c_318_n 0.0215189f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_63 VPB N_A_505_280#_c_319_n 0.00151961f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_505_280#_c_320_n 0.00819307f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_65 VPB N_A_505_280#_c_321_n 0.0147617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_505_280#_c_314_n 0.0297444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_505_280#_c_323_n 9.82358e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_505_280#_c_324_n 0.0291413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_505_280#_c_325_n 0.0112142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_C_M1006_g 0.0471038f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_71 VPB N_D_M1014_g 0.0465585f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_72 VPB D 0.00245404f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_73 VPB N_D_c_427_n 0.00943794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B_N_M1007_g 0.0608713f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_75 VPB B_N 0.00376338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_506_n 0.00224652f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_77 VPB N_VPWR_c_507_n 4.06791e-19 $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_78 VPB N_VPWR_c_508_n 0.00281836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_509_n 0.01518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_510_n 0.0130834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_511_n 0.017432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_512_n 0.014294f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_505_n 0.0453327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_514_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_515_n 0.0177703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_516_n 0.0158558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_517_n 0.00449449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_518_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_X_c_584_n 0.00137385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 N_A_N_M1013_g N_A_174_21#_c_117_n 0.0217878f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_N_M1005_g N_A_174_21#_M1000_g 0.0217878f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_92 N_A_N_c_92_n N_A_174_21#_c_120_n 0.0217878f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_N_M1005_g N_A_27_47#_c_229_n 0.00114093f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_94 N_A_N_M1013_g N_A_27_47#_c_224_n 0.00954277f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_N_M1005_g N_A_27_47#_c_224_n 0.0187175f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_96 A_N N_A_27_47#_c_224_n 0.0447039f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A_N_c_92_n N_A_27_47#_c_224_n 0.00844587f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_N_M1005_g N_A_27_47#_c_231_n 0.0158393f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_99 A_N N_A_27_47#_c_231_n 0.00987856f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_N_c_92_n N_A_27_47#_c_231_n 0.00220498f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_N_M1013_g N_A_27_47#_c_225_n 0.0147979f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_102 A_N N_A_27_47#_c_225_n 0.0112557f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A_N_c_92_n N_A_27_47#_c_225_n 0.00348632f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_N_M1005_g N_VPWR_c_506_n 0.00836134f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_105 N_A_N_M1005_g N_VPWR_c_509_n 0.00342834f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_106 N_A_N_M1005_g N_VPWR_c_505_n 0.00495667f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_107 N_A_N_M1013_g N_X_c_584_n 0.00108796f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_N_M1013_g N_VGND_c_606_n 0.00832549f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_N_M1013_g N_VGND_c_609_n 0.00339367f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_N_M1013_g N_VGND_c_613_n 0.00489827f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_174_21#_c_118_n N_A_27_47#_c_222_n 0.00542216f $X=1.365 $Y=0.995
+ $X2=0 $Y2=0
cc_112 N_A_174_21#_c_119_n N_A_27_47#_c_222_n 0.00224166f $X=1.5 $Y=1.16 $X2=0
+ $Y2=0
cc_113 N_A_174_21#_c_120_n N_A_27_47#_c_222_n 0.0217715f $X=1.5 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_A_174_21#_c_121_n N_A_27_47#_c_222_n 0.00622732f $X=2.01 $Y=0.72 $X2=0
+ $Y2=0
cc_115 N_A_174_21#_c_138_p N_A_27_47#_c_222_n 0.00111522f $X=2.095 $Y=0.42 $X2=0
+ $Y2=0
cc_116 N_A_174_21#_c_122_n N_A_27_47#_c_222_n 0.0181905f $X=2.32 $Y=1.915 $X2=0
+ $Y2=0
cc_117 N_A_174_21#_c_123_n N_A_27_47#_c_222_n 0.0148805f $X=2.32 $Y=0.72 $X2=0
+ $Y2=0
cc_118 N_A_174_21#_M1001_g N_A_27_47#_M1002_g 0.0122305f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_174_21#_c_122_n N_A_27_47#_M1002_g 0.0135713f $X=2.32 $Y=1.915 $X2=0
+ $Y2=0
cc_120 N_A_174_21#_c_143_p N_A_27_47#_M1002_g 0.00399216f $X=2.48 $Y=2.3 $X2=0
+ $Y2=0
cc_121 N_A_174_21#_c_130_n N_A_27_47#_M1002_g 0.00750077f $X=2.565 $Y=2 $X2=0
+ $Y2=0
cc_122 N_A_174_21#_c_123_n N_A_27_47#_c_223_n 0.00716984f $X=2.32 $Y=0.72 $X2=0
+ $Y2=0
cc_123 N_A_174_21#_c_117_n N_A_27_47#_c_224_n 0.0107584f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_174_21#_M1000_g N_A_27_47#_c_258_n 0.0156881f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_174_21#_M1001_g N_A_27_47#_c_258_n 0.0164169f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_174_21#_c_119_n N_A_27_47#_c_258_n 0.00426092f $X=1.5 $Y=1.16 $X2=0
+ $Y2=0
cc_127 N_A_174_21#_c_120_n N_A_27_47#_c_258_n 0.00212863f $X=1.5 $Y=1.16 $X2=0
+ $Y2=0
cc_128 N_A_174_21#_c_122_n N_A_27_47#_c_258_n 0.00149407f $X=2.32 $Y=1.915 $X2=0
+ $Y2=0
cc_129 N_A_174_21#_c_130_n N_A_27_47#_c_258_n 0.00763398f $X=2.565 $Y=2 $X2=0
+ $Y2=0
cc_130 N_A_174_21#_M1001_g N_A_27_47#_c_232_n 0.00725878f $X=1.365 $Y=1.985
+ $X2=0 $Y2=0
cc_131 N_A_174_21#_c_122_n N_A_27_47#_c_232_n 0.0249959f $X=2.32 $Y=1.915 $X2=0
+ $Y2=0
cc_132 N_A_174_21#_c_117_n N_A_27_47#_c_225_n 0.00144547f $X=0.945 $Y=0.995
+ $X2=0 $Y2=0
cc_133 N_A_174_21#_c_119_n N_A_27_47#_c_226_n 0.0247586f $X=1.5 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_174_21#_c_120_n N_A_27_47#_c_226_n 0.00224902f $X=1.5 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_174_21#_c_121_n N_A_27_47#_c_226_n 0.0212431f $X=2.01 $Y=0.72 $X2=0
+ $Y2=0
cc_136 N_A_174_21#_c_122_n N_A_27_47#_c_226_n 0.0234288f $X=2.32 $Y=1.915 $X2=0
+ $Y2=0
cc_137 N_A_174_21#_c_122_n N_A_505_280#_M1011_g 0.0066264f $X=2.32 $Y=1.915
+ $X2=0 $Y2=0
cc_138 N_A_174_21#_c_123_n N_A_505_280#_M1011_g 0.0015643f $X=2.32 $Y=0.72 $X2=0
+ $Y2=0
cc_139 N_A_174_21#_c_122_n N_A_505_280#_M1012_g 0.00345887f $X=2.32 $Y=1.915
+ $X2=0 $Y2=0
cc_140 N_A_174_21#_c_129_n N_A_505_280#_M1012_g 0.011676f $X=3.245 $Y=2 $X2=0
+ $Y2=0
cc_141 N_A_174_21#_c_129_n N_A_505_280#_c_318_n 0.0504461f $X=3.245 $Y=2 $X2=0
+ $Y2=0
cc_142 N_A_174_21#_c_129_n N_A_505_280#_c_331_n 0.014171f $X=3.245 $Y=2 $X2=0
+ $Y2=0
cc_143 N_A_174_21#_c_122_n N_A_505_280#_c_323_n 0.0247306f $X=2.32 $Y=1.915
+ $X2=0 $Y2=0
cc_144 N_A_174_21#_c_129_n N_A_505_280#_c_323_n 0.0124104f $X=3.245 $Y=2 $X2=0
+ $Y2=0
cc_145 N_A_174_21#_c_122_n N_A_505_280#_c_324_n 0.00196674f $X=2.32 $Y=1.915
+ $X2=0 $Y2=0
cc_146 N_A_174_21#_c_129_n N_A_505_280#_c_324_n 4.63768e-19 $X=3.245 $Y=2 $X2=0
+ $Y2=0
cc_147 N_A_174_21#_c_130_n N_A_505_280#_c_324_n 0.00186806f $X=2.565 $Y=2 $X2=0
+ $Y2=0
cc_148 N_A_174_21#_c_129_n N_C_M1006_g 0.0109911f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_149 N_A_174_21#_c_122_n C 0.017111f $X=2.32 $Y=1.915 $X2=0 $Y2=0
cc_150 N_A_174_21#_c_123_n C 0.00635323f $X=2.32 $Y=0.72 $X2=0 $Y2=0
cc_151 N_A_174_21#_c_129_n N_D_M1014_g 0.00127967f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_152 N_A_174_21#_c_129_n N_VPWR_M1012_d 0.00169766f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_153 N_A_174_21#_M1000_g N_VPWR_c_506_n 0.00170957f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_174_21#_c_129_n N_VPWR_c_507_n 0.0166541f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_155 N_A_174_21#_c_143_p N_VPWR_c_510_n 0.0111381f $X=2.48 $Y=2.3 $X2=0 $Y2=0
cc_156 N_A_174_21#_c_130_n N_VPWR_c_510_n 0.004756f $X=2.565 $Y=2 $X2=0 $Y2=0
cc_157 N_A_174_21#_c_129_n N_VPWR_c_511_n 0.00244309f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_158 N_A_174_21#_c_181_p N_VPWR_c_511_n 0.0112274f $X=3.33 $Y=2.3 $X2=0 $Y2=0
cc_159 N_A_174_21#_M1002_d N_VPWR_c_505_n 0.00310074f $X=2.295 $Y=2.065 $X2=0
+ $Y2=0
cc_160 N_A_174_21#_M1006_d N_VPWR_c_505_n 0.00405853f $X=3.195 $Y=2.065 $X2=0
+ $Y2=0
cc_161 N_A_174_21#_M1000_g N_VPWR_c_505_n 0.00587767f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_174_21#_M1001_g N_VPWR_c_505_n 0.00662463f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_174_21#_c_143_p N_VPWR_c_505_n 0.00637602f $X=2.48 $Y=2.3 $X2=0 $Y2=0
cc_164 N_A_174_21#_c_129_n N_VPWR_c_505_n 0.00568161f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_165 N_A_174_21#_c_130_n N_VPWR_c_505_n 0.00844957f $X=2.565 $Y=2 $X2=0 $Y2=0
cc_166 N_A_174_21#_c_181_p N_VPWR_c_505_n 0.00643448f $X=3.33 $Y=2.3 $X2=0 $Y2=0
cc_167 N_A_174_21#_M1000_g N_VPWR_c_515_n 0.00429465f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_174_21#_M1001_g N_VPWR_c_515_n 0.00429465f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_174_21#_M1001_g N_VPWR_c_516_n 0.00422273f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_174_21#_c_143_p N_VPWR_c_516_n 0.0127668f $X=2.48 $Y=2.3 $X2=0 $Y2=0
cc_171 N_A_174_21#_M1000_g X 0.00376127f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_174_21#_M1001_g X 0.00462904f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_174_21#_c_117_n N_X_c_584_n 0.0128832f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_174_21#_M1000_g N_X_c_584_n 0.00417667f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_174_21#_c_118_n N_X_c_584_n 0.00189608f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_174_21#_M1001_g N_X_c_584_n 0.0018922f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_174_21#_c_119_n N_X_c_584_n 0.0327519f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_174_21#_c_120_n N_X_c_584_n 0.0196534f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_174_21#_c_119_n N_VGND_M1015_d 0.0011856f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_174_21#_c_121_n N_VGND_M1015_d 0.00496608f $X=2.01 $Y=0.72 $X2=0
+ $Y2=0
cc_181 N_A_174_21#_c_204_p N_VGND_M1015_d 9.26568e-19 $X=1.585 $Y=0.72 $X2=0
+ $Y2=0
cc_182 N_A_174_21#_c_117_n N_VGND_c_606_n 0.0016047f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_174_21#_c_117_n N_VGND_c_607_n 4.69742e-19 $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_174_21#_c_118_n N_VGND_c_607_n 0.00781637f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_174_21#_c_120_n N_VGND_c_607_n 5.29514e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_174_21#_c_121_n N_VGND_c_607_n 0.0118298f $X=2.01 $Y=0.72 $X2=0 $Y2=0
cc_187 N_A_174_21#_c_204_p N_VGND_c_607_n 0.00936203f $X=1.585 $Y=0.72 $X2=0
+ $Y2=0
cc_188 N_A_174_21#_c_138_p N_VGND_c_607_n 0.0117639f $X=2.095 $Y=0.42 $X2=0
+ $Y2=0
cc_189 N_A_174_21#_c_117_n N_VGND_c_610_n 0.00579312f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_174_21#_c_118_n N_VGND_c_610_n 0.0046653f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_174_21#_c_121_n N_VGND_c_611_n 0.00810179f $X=2.01 $Y=0.72 $X2=0
+ $Y2=0
cc_192 N_A_174_21#_c_138_p N_VGND_c_611_n 0.0111381f $X=2.095 $Y=0.42 $X2=0
+ $Y2=0
cc_193 N_A_174_21#_M1010_s N_VGND_c_613_n 0.00242518f $X=1.97 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_A_174_21#_c_117_n N_VGND_c_613_n 0.0104929f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_174_21#_c_118_n N_VGND_c_613_n 0.00789179f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_174_21#_c_121_n N_VGND_c_613_n 0.0140091f $X=2.01 $Y=0.72 $X2=0 $Y2=0
cc_197 N_A_174_21#_c_204_p N_VGND_c_613_n 8.47748e-19 $X=1.585 $Y=0.72 $X2=0
+ $Y2=0
cc_198 N_A_174_21#_c_138_p N_VGND_c_613_n 0.00637602f $X=2.095 $Y=0.42 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_222_n N_A_505_280#_M1011_g 0.0171282f $X=2.22 $Y=1.325 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_223_n N_A_505_280#_M1011_g 0.0519442f $X=2.305 $Y=0.73 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_M1002_g N_A_505_280#_M1012_g 0.0190229f $X=2.22 $Y=2.275 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_M1002_g N_A_505_280#_c_323_n 3.55433e-19 $X=2.22 $Y=2.275
+ $X2=0 $Y2=0
cc_203 N_A_27_47#_M1002_g N_A_505_280#_c_324_n 0.0178959f $X=2.22 $Y=2.275 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_224_n N_VPWR_M1005_d 0.00470101f $X=0.585 $Y=1.885 $X2=-0.19
+ $Y2=-0.24
cc_205 N_A_27_47#_c_258_n N_VPWR_M1005_d 0.00697892f $X=1.755 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A_27_47#_c_231_n N_VPWR_M1005_d 6.83486e-19 $X=0.67 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_207 N_A_27_47#_c_258_n N_VPWR_M1001_d 0.0163189f $X=1.755 $Y=1.97 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_232_n N_VPWR_M1001_d 0.0131812f $X=1.84 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_231_n N_VPWR_c_506_n 0.0174546f $X=0.67 $Y=1.97 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1002_g N_VPWR_c_507_n 5.01338e-19 $X=2.22 $Y=2.275 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_229_n N_VPWR_c_509_n 0.0111968f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_231_n N_VPWR_c_509_n 0.00271686f $X=0.67 $Y=1.97 $X2=0 $Y2=0
cc_213 N_A_27_47#_M1002_g N_VPWR_c_510_n 0.00460953f $X=2.22 $Y=2.275 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1005_s N_VPWR_c_505_n 0.00367799f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1002_g N_VPWR_c_505_n 0.00695597f $X=2.22 $Y=2.275 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_229_n N_VPWR_c_505_n 0.00638769f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_258_n N_VPWR_c_505_n 0.0183628f $X=1.755 $Y=1.97 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_231_n N_VPWR_c_505_n 0.00561995f $X=0.67 $Y=1.97 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_258_n N_VPWR_c_515_n 0.00883322f $X=1.755 $Y=1.97 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1002_g N_VPWR_c_516_n 0.0079638f $X=2.22 $Y=2.275 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_258_n N_VPWR_c_516_n 0.0294416f $X=1.755 $Y=1.97 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_258_n N_X_M1000_s 0.00438154f $X=1.755 $Y=1.97 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_224_n X 0.00772116f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_258_n X 0.0166092f $X=1.755 $Y=1.97 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_232_n X 0.00606944f $X=1.84 $Y=1.885 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_224_n N_X_c_584_n 0.031619f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_232_n N_X_c_584_n 0.00661005f $X=1.84 $Y=1.885 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_225_n N_X_c_584_n 0.00764158f $X=0.585 $Y=0.72 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_224_n N_VGND_M1013_d 0.00104998f $X=0.585 $Y=1.885 $X2=-0.19
+ $Y2=-0.24
cc_230 N_A_27_47#_c_225_n N_VGND_M1013_d 0.00280791f $X=0.585 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_231 N_A_27_47#_c_225_n N_VGND_c_606_n 0.00721829f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_223_n N_VGND_c_607_n 0.00280581f $X=2.305 $Y=0.73 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_305_p N_VGND_c_609_n 0.0111381f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_225_n N_VGND_c_609_n 0.00247038f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_222_n N_VGND_c_611_n 5.49187e-19 $X=2.22 $Y=1.325 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_223_n N_VGND_c_611_n 0.00425094f $X=2.305 $Y=0.73 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1013_s N_VGND_c_613_n 0.0036562f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_223_n N_VGND_c_613_n 0.0070255f $X=2.305 $Y=0.73 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_305_p N_VGND_c_613_n 0.00637602f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_225_n N_VGND_c_613_n 0.0049411f $X=0.585 $Y=0.72 $X2=0 $Y2=0
cc_241 N_A_505_280#_M1011_g N_C_M1006_g 0.0110838f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_505_280#_M1012_g N_C_M1006_g 0.0247753f $X=2.69 $Y=2.275 $X2=0 $Y2=0
cc_243 N_A_505_280#_c_318_n N_C_M1006_g 0.0114425f $X=3.585 $Y=1.66 $X2=0 $Y2=0
cc_244 N_A_505_280#_c_319_n N_C_M1006_g 8.42713e-19 $X=3.67 $Y=1.915 $X2=0 $Y2=0
cc_245 N_A_505_280#_c_323_n N_C_M1006_g 0.0011047f $X=2.66 $Y=1.565 $X2=0 $Y2=0
cc_246 N_A_505_280#_c_324_n N_C_M1006_g 0.0173401f $X=2.66 $Y=1.565 $X2=0 $Y2=0
cc_247 N_A_505_280#_M1011_g C 0.0109549f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_248 N_A_505_280#_c_318_n C 0.0138456f $X=3.585 $Y=1.66 $X2=0 $Y2=0
cc_249 N_A_505_280#_M1011_g N_C_c_387_n 0.0189174f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A_505_280#_c_318_n N_C_c_387_n 0.00122881f $X=3.585 $Y=1.66 $X2=0 $Y2=0
cc_251 N_A_505_280#_M1011_g N_C_c_388_n 0.0274655f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_252 N_A_505_280#_c_318_n N_D_M1014_g 0.0133391f $X=3.585 $Y=1.66 $X2=0 $Y2=0
cc_253 N_A_505_280#_c_319_n N_D_M1014_g 0.00466067f $X=3.67 $Y=1.915 $X2=0 $Y2=0
cc_254 N_A_505_280#_c_331_n N_D_M1014_g 0.0052306f $X=3.755 $Y=2 $X2=0 $Y2=0
cc_255 N_A_505_280#_c_318_n D 0.024484f $X=3.585 $Y=1.66 $X2=0 $Y2=0
cc_256 N_A_505_280#_c_318_n N_D_c_427_n 0.00268438f $X=3.585 $Y=1.66 $X2=0 $Y2=0
cc_257 N_A_505_280#_c_318_n N_B_N_M1007_g 0.00187263f $X=3.585 $Y=1.66 $X2=0
+ $Y2=0
cc_258 N_A_505_280#_c_319_n N_B_N_M1007_g 0.00151892f $X=3.67 $Y=1.915 $X2=0
+ $Y2=0
cc_259 N_A_505_280#_c_320_n N_B_N_M1007_g 0.0162963f $X=4.255 $Y=2 $X2=0 $Y2=0
cc_260 N_A_505_280#_c_314_n N_B_N_M1007_g 0.0219335f $X=4.43 $Y=1.915 $X2=0
+ $Y2=0
cc_261 N_A_505_280#_c_320_n B_N 0.0108555f $X=4.255 $Y=2 $X2=0 $Y2=0
cc_262 N_A_505_280#_c_314_n B_N 0.0407278f $X=4.43 $Y=1.915 $X2=0 $Y2=0
cc_263 N_A_505_280#_c_314_n N_B_N_c_471_n 0.00753248f $X=4.43 $Y=1.915 $X2=0
+ $Y2=0
cc_264 N_A_505_280#_c_314_n N_B_N_c_472_n 0.00582504f $X=4.43 $Y=1.915 $X2=0
+ $Y2=0
cc_265 N_A_505_280#_c_320_n N_VPWR_M1014_d 0.00255903f $X=4.255 $Y=2 $X2=0 $Y2=0
cc_266 N_A_505_280#_c_331_n N_VPWR_M1014_d 0.00150236f $X=3.755 $Y=2 $X2=0 $Y2=0
cc_267 N_A_505_280#_M1012_g N_VPWR_c_507_n 0.00673272f $X=2.69 $Y=2.275 $X2=0
+ $Y2=0
cc_268 N_A_505_280#_c_320_n N_VPWR_c_508_n 0.020494f $X=4.255 $Y=2 $X2=0 $Y2=0
cc_269 N_A_505_280#_M1012_g N_VPWR_c_510_n 0.00339367f $X=2.69 $Y=2.275 $X2=0
+ $Y2=0
cc_270 N_A_505_280#_c_331_n N_VPWR_c_511_n 0.00264874f $X=3.755 $Y=2 $X2=0 $Y2=0
cc_271 N_A_505_280#_c_320_n N_VPWR_c_512_n 0.00244309f $X=4.255 $Y=2 $X2=0 $Y2=0
cc_272 N_A_505_280#_c_321_n N_VPWR_c_512_n 0.0179115f $X=4.34 $Y=2.3 $X2=0 $Y2=0
cc_273 N_A_505_280#_M1007_d N_VPWR_c_505_n 0.00226392f $X=4.205 $Y=2.065 $X2=0
+ $Y2=0
cc_274 N_A_505_280#_M1012_g N_VPWR_c_505_n 0.00408948f $X=2.69 $Y=2.275 $X2=0
+ $Y2=0
cc_275 N_A_505_280#_c_320_n N_VPWR_c_505_n 0.00564956f $X=4.255 $Y=2 $X2=0 $Y2=0
cc_276 N_A_505_280#_c_331_n N_VPWR_c_505_n 0.0048944f $X=3.755 $Y=2 $X2=0 $Y2=0
cc_277 N_A_505_280#_c_321_n N_VPWR_c_505_n 0.00991723f $X=4.34 $Y=2.3 $X2=0
+ $Y2=0
cc_278 N_A_505_280#_M1012_g N_VPWR_c_516_n 5.15836e-19 $X=2.69 $Y=2.275 $X2=0
+ $Y2=0
cc_279 N_A_505_280#_M1011_g N_VGND_c_611_n 0.00585385f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_280 N_A_505_280#_c_315_n N_VGND_c_612_n 0.0170867f $X=4.43 $Y=0.42 $X2=0
+ $Y2=0
cc_281 N_A_505_280#_M1008_d N_VGND_c_613_n 0.00335808f $X=4.205 $Y=0.235 $X2=0
+ $Y2=0
cc_282 N_A_505_280#_M1011_g N_VGND_c_613_n 0.0107924f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_283 N_A_505_280#_c_315_n N_VGND_c_613_n 0.00982816f $X=4.43 $Y=0.42 $X2=0
+ $Y2=0
cc_284 C N_D_M1004_g 6.64279e-19 $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_285 N_C_c_387_n N_D_M1004_g 0.0153811f $X=3.09 $Y=0.94 $X2=0 $Y2=0
cc_286 N_C_c_388_n N_D_M1004_g 0.0310338f $X=3.09 $Y=0.775 $X2=0 $Y2=0
cc_287 N_C_M1006_g N_D_M1014_g 0.0396448f $X=3.12 $Y=2.275 $X2=0 $Y2=0
cc_288 N_C_M1006_g D 0.00390559f $X=3.12 $Y=2.275 $X2=0 $Y2=0
cc_289 C D 0.063959f $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_290 N_C_c_387_n D 0.00211845f $X=3.09 $Y=0.94 $X2=0 $Y2=0
cc_291 N_C_c_388_n D 0.00209165f $X=3.09 $Y=0.775 $X2=0 $Y2=0
cc_292 N_C_M1006_g N_D_c_427_n 0.0148835f $X=3.12 $Y=2.275 $X2=0 $Y2=0
cc_293 C N_D_c_427_n 2.07553e-19 $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_294 N_C_c_387_n N_D_c_427_n 0.00183531f $X=3.09 $Y=0.94 $X2=0 $Y2=0
cc_295 N_C_M1006_g N_VPWR_c_507_n 0.00786314f $X=3.12 $Y=2.275 $X2=0 $Y2=0
cc_296 N_C_M1006_g N_VPWR_c_511_n 0.00339367f $X=3.12 $Y=2.275 $X2=0 $Y2=0
cc_297 N_C_M1006_g N_VPWR_c_505_n 0.00397127f $X=3.12 $Y=2.275 $X2=0 $Y2=0
cc_298 C N_VGND_c_611_n 0.00777064f $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_299 N_C_c_387_n N_VGND_c_611_n 7.49045e-19 $X=3.09 $Y=0.94 $X2=0 $Y2=0
cc_300 N_C_c_388_n N_VGND_c_611_n 0.00417173f $X=3.09 $Y=0.775 $X2=0 $Y2=0
cc_301 C N_VGND_c_613_n 0.00857114f $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_302 N_C_c_387_n N_VGND_c_613_n 7.02243e-19 $X=3.09 $Y=0.94 $X2=0 $Y2=0
cc_303 N_C_c_388_n N_VGND_c_613_n 0.00631876f $X=3.09 $Y=0.775 $X2=0 $Y2=0
cc_304 C A_548_47# 0.00393403f $X=2.91 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_305 N_D_M1014_g N_B_N_M1007_g 0.0256765f $X=3.54 $Y=2.275 $X2=0 $Y2=0
cc_306 D N_B_N_M1007_g 7.19391e-19 $X=3.37 $Y=0.425 $X2=0 $Y2=0
cc_307 N_D_c_427_n N_B_N_M1007_g 0.00977166f $X=3.57 $Y=1.24 $X2=0 $Y2=0
cc_308 N_D_M1004_g B_N 0.00104867f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_309 D B_N 0.0439528f $X=3.37 $Y=0.425 $X2=0 $Y2=0
cc_310 N_D_c_427_n B_N 0.00181173f $X=3.57 $Y=1.24 $X2=0 $Y2=0
cc_311 N_D_M1004_g N_B_N_c_471_n 0.0108356f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_312 D N_B_N_c_471_n 8.47201e-19 $X=3.37 $Y=0.425 $X2=0 $Y2=0
cc_313 N_D_c_427_n N_B_N_c_471_n 9.76608e-19 $X=3.57 $Y=1.24 $X2=0 $Y2=0
cc_314 N_D_M1004_g N_B_N_c_472_n 0.0109584f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_315 D N_B_N_c_472_n 0.00218067f $X=3.37 $Y=0.425 $X2=0 $Y2=0
cc_316 N_D_M1014_g N_VPWR_c_507_n 0.00116396f $X=3.54 $Y=2.275 $X2=0 $Y2=0
cc_317 N_D_M1014_g N_VPWR_c_508_n 0.005234f $X=3.54 $Y=2.275 $X2=0 $Y2=0
cc_318 N_D_M1014_g N_VPWR_c_511_n 0.00553297f $X=3.54 $Y=2.275 $X2=0 $Y2=0
cc_319 N_D_M1014_g N_VPWR_c_505_n 0.0101794f $X=3.54 $Y=2.275 $X2=0 $Y2=0
cc_320 N_D_M1004_g N_VGND_c_608_n 0.00689445f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_321 N_D_M1004_g N_VGND_c_611_n 0.00390689f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_322 D N_VGND_c_611_n 0.00833675f $X=3.37 $Y=0.425 $X2=0 $Y2=0
cc_323 N_D_M1004_g N_VGND_c_613_n 0.00586074f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_324 D N_VGND_c_613_n 0.00983187f $X=3.37 $Y=0.425 $X2=0 $Y2=0
cc_325 D A_639_47# 0.00274529f $X=3.37 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_326 N_B_N_M1007_g N_VPWR_c_508_n 0.00860639f $X=4.13 $Y=2.275 $X2=0 $Y2=0
cc_327 N_B_N_M1007_g N_VPWR_c_512_n 0.00339367f $X=4.13 $Y=2.275 $X2=0 $Y2=0
cc_328 N_B_N_M1007_g N_VPWR_c_505_n 0.00489827f $X=4.13 $Y=2.275 $X2=0 $Y2=0
cc_329 B_N N_VGND_c_608_n 0.0175645f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_330 N_B_N_c_471_n N_VGND_c_608_n 6.04781e-19 $X=4.09 $Y=0.93 $X2=0 $Y2=0
cc_331 N_B_N_c_472_n N_VGND_c_608_n 0.00974832f $X=4.09 $Y=0.765 $X2=0 $Y2=0
cc_332 N_B_N_c_471_n N_VGND_c_612_n 3.50417e-19 $X=4.09 $Y=0.93 $X2=0 $Y2=0
cc_333 N_B_N_c_472_n N_VGND_c_612_n 0.0046653f $X=4.09 $Y=0.765 $X2=0 $Y2=0
cc_334 B_N N_VGND_c_613_n 0.00435768f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_335 N_B_N_c_471_n N_VGND_c_613_n 4.58436e-19 $X=4.09 $Y=0.93 $X2=0 $Y2=0
cc_336 N_B_N_c_472_n N_VGND_c_613_n 0.00607644f $X=4.09 $Y=0.765 $X2=0 $Y2=0
cc_337 N_VPWR_c_505_n N_X_M1000_s 0.00327078f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_338 N_X_c_584_n N_VGND_c_610_n 0.0134454f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_339 N_X_M1003_s N_VGND_c_613_n 0.0038878f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_340 N_X_c_584_n N_VGND_c_613_n 0.00849738f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_341 N_VGND_c_613_n A_476_47# 0.00818821f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_342 N_VGND_c_613_n A_548_47# 0.00851002f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_343 N_VGND_c_613_n A_639_47# 0.00700839f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__fa_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.240000 1.275000 ;
        RECT 0.910000 1.275000 1.080000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.230000 1.030000 2.620000 1.360000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.250000 0.955000 4.625000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.885000 1.035000 6.325000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.010000 1.075000 1.300000 1.120000 ;
        RECT 1.010000 1.120000 6.380000 1.260000 ;
        RECT 1.010000 1.260000 1.300000 1.305000 ;
        RECT 2.390000 1.075000 2.680000 1.120000 ;
        RECT 2.390000 1.260000 2.680000 1.305000 ;
        RECT 4.250000 1.075000 4.540000 1.120000 ;
        RECT 4.250000 1.260000 4.540000 1.305000 ;
        RECT 6.090000 1.075000 6.380000 1.120000 ;
        RECT 6.090000 1.260000 6.380000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 1.445000 1.700000 1.880000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.200000 1.435000 3.560000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.635000 1.445000 6.055000 1.765000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.470000 1.415000 1.760000 1.460000 ;
        RECT 1.470000 1.460000 5.920000 1.600000 ;
        RECT 1.470000 1.600000 1.760000 1.645000 ;
        RECT 3.330000 1.415000 3.620000 1.460000 ;
        RECT 3.330000 1.600000 3.620000 1.645000 ;
        RECT 5.630000 1.415000 5.920000 1.460000 ;
        RECT 5.630000 1.600000 5.920000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.670000 1.105000 2.040000 1.275000 ;
        RECT 1.870000 1.275000 2.040000 1.595000 ;
        RECT 1.870000 1.595000 2.960000 1.765000 ;
        RECT 2.790000 0.965000 3.955000 1.250000 ;
        RECT 2.790000 1.250000 2.960000 1.595000 ;
        RECT 3.785000 1.250000 3.955000 1.515000 ;
        RECT 3.785000 1.515000 5.405000 1.685000 ;
        RECT 5.155000 1.685000 5.405000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.830000 ;
        RECT 0.085000 0.830000 0.260000 1.485000 ;
        RECT 0.085000 1.485000 0.345000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.840000 0.255000 7.240000 0.810000 ;
        RECT 6.840000 1.485000 7.240000 2.465000 ;
        RECT 6.910000 0.810000 7.240000 1.485000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.360000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 2.300000  0.085000 2.630000 0.445000 ;
        RECT 3.240000  0.085000 3.570000 0.490000 ;
        RECT 4.080000  0.085000 4.410000 0.445000 ;
        RECT 6.265000  0.085000 6.595000 0.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.515000 2.150000 0.765000 2.635000 ;
        RECT 2.300000 2.275000 2.630000 2.635000 ;
        RECT 3.240000 2.255000 3.570000 2.635000 ;
        RECT 4.080000 2.275000 4.410000 2.635000 ;
        RECT 6.340000 2.275000 6.670000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.430000 0.995000 0.685000 1.325000 ;
      RECT 0.515000 0.635000 1.710000 0.805000 ;
      RECT 0.515000 0.805000 0.685000 0.995000 ;
      RECT 0.515000 1.325000 0.685000 1.625000 ;
      RECT 0.515000 1.625000 1.105000 1.945000 ;
      RECT 0.935000 1.945000 1.105000 2.065000 ;
      RECT 0.935000 2.065000 1.710000 2.465000 ;
      RECT 1.110000 0.255000 1.710000 0.635000 ;
      RECT 1.470000 0.805000 1.710000 0.935000 ;
      RECT 1.960000 0.255000 2.130000 0.615000 ;
      RECT 1.960000 0.615000 2.970000 0.785000 ;
      RECT 1.960000 1.935000 3.035000 2.105000 ;
      RECT 1.960000 2.105000 2.130000 2.465000 ;
      RECT 2.800000 0.255000 2.970000 0.615000 ;
      RECT 2.800000 2.105000 3.035000 2.465000 ;
      RECT 3.740000 0.255000 3.910000 0.615000 ;
      RECT 3.740000 0.615000 4.750000 0.785000 ;
      RECT 3.740000 1.935000 4.750000 2.105000 ;
      RECT 3.740000 2.105000 3.910000 2.465000 ;
      RECT 4.580000 0.255000 4.750000 0.615000 ;
      RECT 4.580000 2.105000 4.750000 2.465000 ;
      RECT 4.795000 0.955000 5.460000 1.125000 ;
      RECT 4.965000 0.765000 5.460000 0.955000 ;
      RECT 5.085000 0.255000 6.095000 0.505000 ;
      RECT 5.085000 0.505000 5.255000 0.595000 ;
      RECT 5.085000 2.125000 6.170000 2.465000 ;
      RECT 5.925000 0.505000 6.095000 0.615000 ;
      RECT 5.925000 0.615000 6.665000 0.785000 ;
      RECT 6.000000 1.935000 6.665000 2.105000 ;
      RECT 6.000000 2.105000 6.170000 2.125000 ;
      RECT 6.495000 0.785000 6.665000 0.995000 ;
      RECT 6.495000 0.995000 6.740000 1.325000 ;
      RECT 6.495000 1.325000 6.665000 1.935000 ;
    LAYER mcon ;
      RECT 1.530000 0.765000 1.700000 0.935000 ;
      RECT 5.230000 0.765000 5.400000 0.935000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 5.460000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 5.170000 0.735000 5.460000 0.780000 ;
      RECT 5.170000 0.920000 5.460000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_1

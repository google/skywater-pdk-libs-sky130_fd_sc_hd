* File: sky130_fd_sc_hd__clkdlybuf4s50_1.pex.spice
* Created: Thu Aug 27 14:12:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A 3 7 9 12 13
r29 12 15 43.9584 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.38 $Y=1.16
+ $X2=0.38 $Y2=1.31
r30 12 14 43.1341 $w=3.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.38 $Y=1.16
+ $X2=0.38 $Y2=1.015
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.16 $X2=0.37 $Y2=1.16
r32 9 13 7.23627 $w=2.13e-07 $l=1.35e-07 $layer=LI1_cond $X=0.235 $Y=1.182
+ $X2=0.37 $Y2=1.182
r33 7 15 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.48 $Y=1.985
+ $X2=0.48 $Y2=1.31
r34 3 14 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.48 $Y=0.445
+ $X2=0.48 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_27_47# 1 2 9 13 17 21 23 24 25 26
+ 29 30
r69 30 34 13.7388 $w=6.1e-07 $l=1.35e-07 $layer=POLY_cond $X=1.11 $Y=1.16
+ $X2=1.11 $Y2=1.295
r70 30 33 13.7388 $w=6.1e-07 $l=1.35e-07 $layer=POLY_cond $X=1.11 $Y=1.16
+ $X2=1.11 $Y2=1.025
r71 29 31 12.5253 $w=3.75e-07 $l=3.85e-07 $layer=LI1_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=1.545
r72 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.16 $X2=0.97 $Y2=1.16
r73 27 29 11.0613 $w=3.75e-07 $l=3.4e-07 $layer=LI1_cond $X=0.92 $Y=0.82
+ $X2=0.92 $Y2=1.16
r74 25 31 5.38787 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.705 $Y=1.545
+ $X2=0.92 $Y2=1.545
r75 25 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.705 $Y=1.545
+ $X2=0.43 $Y2=1.545
r76 23 27 5.38787 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.705 $Y=0.82
+ $X2=0.92 $Y2=0.82
r77 23 24 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.705 $Y=0.82
+ $X2=0.415 $Y2=0.82
r78 19 26 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.257 $Y=1.63
+ $X2=0.43 $Y2=1.545
r79 19 21 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=1.63
+ $X2=0.257 $Y2=1.965
r80 15 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.25 $Y=0.735
+ $X2=0.415 $Y2=0.82
r81 15 17 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.25 $Y=0.735 $X2=0.25
+ $Y2=0.435
r82 13 34 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.165 $Y=2.075
+ $X2=1.165 $Y2=1.295
r83 9 33 49.7577 $w=5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.165 $Y=0.56
+ $X2=1.165 $Y2=1.025
r84 2 21 300 $w=1.7e-07 $l=5.4111e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=1.965
r85 1 17 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_283_47# 1 2 9 13 15 16 19 23 27 30
c54 30 0 7.48979e-20 $X=1.555 $Y=1.195
c55 27 0 7.91693e-20 $X=2.075 $Y=1.16
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.16 $X2=2.075 $Y2=1.16
r57 25 30 2.57785 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=1.73 $Y=1.195
+ $X2=1.555 $Y2=1.195
r58 25 27 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=1.73 $Y=1.195
+ $X2=2.075 $Y2=1.195
r59 21 30 3.87184 $w=3.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.32
+ $X2=1.555 $Y2=1.195
r60 21 23 21.2379 $w=3.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.555 $Y=1.32
+ $X2=1.555 $Y2=1.965
r61 17 30 3.87184 $w=3.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.07
+ $X2=1.555 $Y2=1.195
r62 17 19 20.9086 $w=3.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.555 $Y=1.07
+ $X2=1.555 $Y2=0.435
r63 15 28 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.075 $Y2=1.16
r64 15 16 14.3442 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.465 $Y2=1.16
r65 11 16 11.9087 $w=5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.465 $Y=1.295
+ $X2=2.465 $Y2=1.16
r66 11 13 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.465 $Y=1.295
+ $X2=2.465 $Y2=2.075
r67 7 16 11.9087 $w=5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.465 $Y=1.025
+ $X2=2.465 $Y2=1.16
r68 7 9 49.7577 $w=5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.465 $Y=1.025
+ $X2=2.465 $Y2=0.56
r69 2 23 300 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.665 $X2=1.555 $Y2=1.965
r70 1 19 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.55 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%A_390_47# 1 2 9 13 17 21 23 24 27 28
+ 33
c58 28 0 7.91693e-20 $X=3.075 $Y=1.16
r59 28 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.16
+ $X2=3.075 $Y2=1.325
r60 28 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.16
+ $X2=3.075 $Y2=0.995
r61 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.075
+ $Y=1.16 $X2=3.075 $Y2=1.16
r62 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.58 $Y=1.16
+ $X2=3.075 $Y2=1.16
r63 24 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=1.495
+ $X2=2.495 $Y2=1.58
r64 23 25 9.01297 $w=2.9e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.495 $Y=1.325
+ $X2=2.41 $Y2=1.16
r65 23 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.495 $Y=1.325
+ $X2=2.495 $Y2=1.495
r66 19 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.115 $Y=1.58
+ $X2=2.495 $Y2=1.58
r67 19 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.115 $Y=1.665
+ $X2=2.115 $Y2=1.96
r68 15 25 18.3554 $w=2.9e-07 $l=5.58346e-07 $layer=LI1_cond $X=2.115 $Y=0.73
+ $X2=2.41 $Y2=1.16
r69 15 17 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.115 $Y=0.73
+ $X2=2.115 $Y2=0.435
r70 13 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.115 $Y=1.985
+ $X2=3.115 $Y2=1.325
r71 9 36 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.115 $Y=0.445
+ $X2=3.115 $Y2=0.995
r72 2 21 300 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=2 $X=1.95
+ $Y=1.665 $X2=2.075 $Y2=1.96
r73 1 17 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.235 $X2=2.075 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.765 $Y2=2.72
r51 25 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.765 $Y2=2.72
r53 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r54 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 16 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.855 $Y2=2.72
r58 15 33 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=2.855 $Y2=2.72
r60 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=2.635
+ $X2=2.855 $Y2=2.72
r61 11 13 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.855 $Y=2.635
+ $X2=2.855 $Y2=1.965
r62 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.72
r63 7 9 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=1.965
r64 2 13 300 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=1.665 $X2=2.855 $Y2=1.965
r65 1 9 300 $w=1.7e-07 $l=5.755e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.765 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%X 1 2 7 8 9 10 11 12 36 44
r14 28 44 0.626018 $w=4.03e-07 $l=2.2e-08 $layer=LI1_cond $X=3.392 $Y=1.892
+ $X2=3.392 $Y2=1.87
r15 12 31 7.11385 $w=4.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.392 $Y=2.21
+ $X2=3.392 $Y2=1.96
r16 11 44 0.910572 $w=4.03e-07 $l=3.2e-08 $layer=LI1_cond $X=3.392 $Y=1.838
+ $X2=3.392 $Y2=1.87
r17 11 42 5.88868 $w=4.03e-07 $l=1.48e-07 $layer=LI1_cond $X=3.392 $Y=1.838
+ $X2=3.392 $Y2=1.69
r18 11 31 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=3.392 $Y=1.923
+ $X2=3.392 $Y2=1.96
r19 11 28 0.882117 $w=4.03e-07 $l=3.1e-08 $layer=LI1_cond $X=3.392 $Y=1.923
+ $X2=3.392 $Y2=1.892
r20 10 42 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=3.47 $Y=1.53
+ $X2=3.47 $Y2=1.69
r21 9 10 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=3.47 $Y=1.19 $X2=3.47
+ $Y2=1.53
r22 8 9 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=3.47 $Y=0.85 $X2=3.47
+ $Y2=1.19
r23 8 40 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=3.47 $Y=0.85 $X2=3.47
+ $Y2=0.64
r24 7 40 5.37648 $w=4.03e-07 $l=1.3e-07 $layer=LI1_cond $X=3.392 $Y=0.51
+ $X2=3.392 $Y2=0.64
r25 7 36 2.13415 $w=4.03e-07 $l=7.5e-08 $layer=LI1_cond $X=3.392 $Y=0.51
+ $X2=3.392 $Y2=0.435
r26 2 31 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=3.19
+ $Y=1.485 $X2=3.345 $Y2=1.96
r27 1 36 182 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.235 $X2=3.345 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r47 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r50 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r51 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r52 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r53 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r54 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r55 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r56 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.15
+ $Y2=0
r57 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r58 20 22 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.23
+ $Y2=0
r59 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r60 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r61 16 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.53
+ $Y2=0
r62 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r63 15 33 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.45
+ $Y2=0
r64 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r65 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r66 11 13 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.435
r67 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r68 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.435
r69 2 13 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.435
r70 1 9 182 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.75 $Y2=0.435
.ends


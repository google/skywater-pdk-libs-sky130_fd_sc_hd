* File: sky130_fd_sc_hd__dlxbn_2.pxi.spice
* Created: Thu Aug 27 14:17:56 2020
* 
x_PM_SKY130_FD_SC_HD__DLXBN_2%GATE_N N_GATE_N_c_174_n N_GATE_N_c_169_n
+ N_GATE_N_M1022_g N_GATE_N_c_175_n N_GATE_N_M1008_g N_GATE_N_c_170_n
+ N_GATE_N_c_176_n GATE_N GATE_N N_GATE_N_c_172_n N_GATE_N_c_173_n
+ PM_SKY130_FD_SC_HD__DLXBN_2%GATE_N
x_PM_SKY130_FD_SC_HD__DLXBN_2%A_27_47# N_A_27_47#_M1022_s N_A_27_47#_M1008_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_M1006_g N_A_27_47#_M1015_g
+ N_A_27_47#_c_366_p N_A_27_47#_c_213_n N_A_27_47#_c_214_n N_A_27_47#_c_224_n
+ N_A_27_47#_c_225_n N_A_27_47#_c_226_n N_A_27_47#_c_215_n N_A_27_47#_c_216_n
+ N_A_27_47#_c_217_n N_A_27_47#_c_218_n N_A_27_47#_c_228_n N_A_27_47#_c_229_n
+ N_A_27_47#_c_230_n N_A_27_47#_c_231_n N_A_27_47#_c_232_n N_A_27_47#_c_219_n
+ N_A_27_47#_c_220_n N_A_27_47#_c_234_n N_A_27_47#_c_221_n
+ PM_SKY130_FD_SC_HD__DLXBN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DLXBN_2%D N_D_M1024_g N_D_M1005_g D N_D_c_381_n
+ N_D_c_382_n PM_SKY130_FD_SC_HD__DLXBN_2%D
x_PM_SKY130_FD_SC_HD__DLXBN_2%A_303_47# N_A_303_47#_M1024_s N_A_303_47#_M1005_s
+ N_A_303_47#_M1003_g N_A_303_47#_M1004_g N_A_303_47#_c_427_n
+ N_A_303_47#_c_420_n N_A_303_47#_c_428_n N_A_303_47#_c_429_n
+ N_A_303_47#_c_421_n N_A_303_47#_c_422_n N_A_303_47#_c_423_n
+ N_A_303_47#_c_424_n N_A_303_47#_c_425_n PM_SKY130_FD_SC_HD__DLXBN_2%A_303_47#
x_PM_SKY130_FD_SC_HD__DLXBN_2%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1013_g N_A_193_47#_c_502_n N_A_193_47#_c_503_n
+ N_A_193_47#_M1016_g N_A_193_47#_c_509_n N_A_193_47#_c_505_n
+ N_A_193_47#_c_511_n N_A_193_47#_c_512_n N_A_193_47#_c_513_n
+ N_A_193_47#_c_514_n N_A_193_47#_c_515_n N_A_193_47#_c_516_n
+ N_A_193_47#_c_517_n PM_SKY130_FD_SC_HD__DLXBN_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DLXBN_2%A_728_21# N_A_728_21#_M1002_s N_A_728_21#_M1014_s
+ N_A_728_21#_M1007_g N_A_728_21#_M1020_g N_A_728_21#_c_615_n
+ N_A_728_21#_M1019_g N_A_728_21#_M1001_g N_A_728_21#_c_616_n
+ N_A_728_21#_M1023_g N_A_728_21#_M1011_g N_A_728_21#_c_617_n
+ N_A_728_21#_c_618_n N_A_728_21#_c_619_n N_A_728_21#_c_630_n
+ N_A_728_21#_c_620_n N_A_728_21#_M1009_g N_A_728_21#_c_631_n
+ N_A_728_21#_M1025_g N_A_728_21#_c_632_n N_A_728_21#_c_633_n
+ N_A_728_21#_c_634_n N_A_728_21#_c_725_p N_A_728_21#_c_688_p
+ N_A_728_21#_c_621_n N_A_728_21#_c_635_n N_A_728_21#_c_622_n
+ N_A_728_21#_c_652_p N_A_728_21#_c_648_p N_A_728_21#_c_654_p
+ PM_SKY130_FD_SC_HD__DLXBN_2%A_728_21#
x_PM_SKY130_FD_SC_HD__DLXBN_2%A_565_413# N_A_565_413#_M1006_d
+ N_A_565_413#_M1013_d N_A_565_413#_c_746_n N_A_565_413#_M1002_g
+ N_A_565_413#_M1014_g N_A_565_413#_c_747_n N_A_565_413#_c_748_n
+ N_A_565_413#_c_757_n N_A_565_413#_c_760_n N_A_565_413#_c_749_n
+ N_A_565_413#_c_750_n N_A_565_413#_c_755_n N_A_565_413#_c_751_n
+ PM_SKY130_FD_SC_HD__DLXBN_2%A_565_413#
x_PM_SKY130_FD_SC_HD__DLXBN_2%A_1223_47# N_A_1223_47#_M1009_s
+ N_A_1223_47#_M1025_s N_A_1223_47#_c_829_n N_A_1223_47#_M1017_g
+ N_A_1223_47#_M1012_g N_A_1223_47#_c_830_n N_A_1223_47#_c_831_n
+ N_A_1223_47#_M1021_g N_A_1223_47#_M1018_g N_A_1223_47#_c_834_n
+ N_A_1223_47#_c_835_n N_A_1223_47#_c_840_n N_A_1223_47#_c_836_n
+ N_A_1223_47#_c_856_n PM_SKY130_FD_SC_HD__DLXBN_2%A_1223_47#
x_PM_SKY130_FD_SC_HD__DLXBN_2%VPWR N_VPWR_M1008_d N_VPWR_M1005_d N_VPWR_M1020_d
+ N_VPWR_M1014_d N_VPWR_M1011_s N_VPWR_M1025_d N_VPWR_M1018_d N_VPWR_c_909_n
+ N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n N_VPWR_c_914_n
+ N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_917_n VPWR N_VPWR_c_918_n
+ N_VPWR_c_919_n N_VPWR_c_920_n N_VPWR_c_921_n N_VPWR_c_922_n N_VPWR_c_923_n
+ N_VPWR_c_924_n N_VPWR_c_925_n N_VPWR_c_926_n N_VPWR_c_927_n N_VPWR_c_928_n
+ N_VPWR_c_929_n N_VPWR_c_908_n PM_SKY130_FD_SC_HD__DLXBN_2%VPWR
x_PM_SKY130_FD_SC_HD__DLXBN_2%Q N_Q_M1019_s N_Q_M1001_d N_Q_c_1040_n
+ N_Q_c_1038_n N_Q_c_1039_n N_Q_c_1048_n Q Q Q Q PM_SKY130_FD_SC_HD__DLXBN_2%Q
x_PM_SKY130_FD_SC_HD__DLXBN_2%Q_N N_Q_N_M1017_s N_Q_N_M1012_s N_Q_N_c_1067_n
+ N_Q_N_c_1076_n N_Q_N_c_1069_n Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_HD__DLXBN_2%Q_N
x_PM_SKY130_FD_SC_HD__DLXBN_2%VGND N_VGND_M1022_d N_VGND_M1024_d N_VGND_M1007_d
+ N_VGND_M1002_d N_VGND_M1023_d N_VGND_M1009_d N_VGND_M1021_d N_VGND_c_1096_n
+ N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n N_VGND_c_1100_n
+ N_VGND_c_1101_n N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n VGND
+ N_VGND_c_1105_n N_VGND_c_1106_n N_VGND_c_1107_n N_VGND_c_1108_n
+ N_VGND_c_1109_n N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n
+ N_VGND_c_1117_n PM_SKY130_FD_SC_HD__DLXBN_2%VGND
cc_1 VNB N_GATE_N_c_169_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_170_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_172_n 0.0210048f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_173_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0398906f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_213_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_8 VNB N_A_27_47#_c_214_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_215_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_216_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_217_n 0.0271287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_218_n 0.00378508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_219_n 0.0231162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_220_n 0.0176114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_221_n 0.00469707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1024_g 0.0259397f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_M1005_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_381_n 0.00419114f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_382_n 0.0423288f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_20 VNB N_A_303_47#_M1004_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_303_47#_c_420_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_303_47#_c_421_n 0.00496114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_303_47#_c_422_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_24 VNB N_A_303_47#_c_423_n 0.00269182f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_25 VNB N_A_303_47#_c_424_n 0.0274388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_303_47#_c_425_n 0.01709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_502_n 0.0133385f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_28 VNB N_A_193_47#_c_503_n 0.00520223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_M1016_g 0.0464035f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_30 VNB N_A_193_47#_c_505_n 0.0142766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_728_21#_M1007_g 0.0478162f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_728_21#_c_615_n 0.0160878f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_33 VNB N_A_728_21#_c_616_n 0.0195704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_728_21#_c_617_n 0.0394189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_728_21#_c_618_n 0.0283804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_728_21#_c_619_n 0.0342221f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_37 VNB N_A_728_21#_c_620_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_728_21#_c_621_n 0.00252501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_728_21#_c_622_n 0.00281539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_565_413#_c_746_n 0.0195151f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_41 VNB N_A_565_413#_c_747_n 0.0442039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_565_413#_c_748_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_43 VNB N_A_565_413#_c_749_n 0.00691811f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_44 VNB N_A_565_413#_c_750_n 0.0118438f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_45 VNB N_A_565_413#_c_751_n 0.00194757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1223_47#_c_829_n 0.0169457f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_47 VNB N_A_1223_47#_c_830_n 0.01318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1223_47#_c_831_n 0.0191396f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_49 VNB N_A_1223_47#_M1021_g 0.0238416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1223_47#_M1018_g 5.18715e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1223_47#_c_834_n 0.0128325f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_52 VNB N_A_1223_47#_c_835_n 0.00948496f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_53 VNB N_A_1223_47#_c_836_n 0.0051319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_908_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_Q_c_1038_n 0.00105223f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_56 VNB N_Q_N_c_1067_n 0.00121852f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_57 VNB Q_N 0.0155028f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_58 VNB N_VGND_c_1096_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_59 VNB N_VGND_c_1097_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_60 VNB N_VGND_c_1098_n 0.0115286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1099_n 0.0197453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1100_n 0.00194728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1101_n 0.00828166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1102_n 0.00254474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1103_n 0.00991007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1104_n 0.0315363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1105_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1106_n 0.0278111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1107_n 0.0412073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1108_n 0.0157972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1109_n 0.0183601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1110_n 0.0153174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1111_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1112_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1113_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1114_n 0.00423916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1115_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1116_n 0.00440331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1117_n 0.400895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VPB N_GATE_N_c_174_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_81 VPB N_GATE_N_c_175_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_82 VPB N_GATE_N_c_176_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_83 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_84 VPB N_GATE_N_c_172_n 0.0106763f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_85 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_86 VPB N_A_27_47#_M1015_g 0.0212472f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_87 VPB N_A_27_47#_c_224_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_225_n 0.00556025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_47#_c_226_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_27_47#_c_215_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_27_47#_c_228_n 0.0289584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_47#_c_229_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_27_47#_c_230_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_47#_c_231_n 0.0035222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_c_232_n 0.0037442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_27_47#_c_219_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_47#_c_234_n 0.0330434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_27_47#_c_221_n 2.971e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_D_M1005_g 0.0463366f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_100 VPB N_D_c_381_n 0.00235652f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_101 VPB N_A_303_47#_M1004_g 0.0366887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_303_47#_c_427_n 0.00736238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_303_47#_c_428_n 0.00415091f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_104 VPB N_A_303_47#_c_429_n 0.00297469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_303_47#_c_422_n 0.00361895f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_106 VPB N_A_193_47#_M1013_g 0.0316829f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_107 VPB N_A_193_47#_c_502_n 0.0172364f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_108 VPB N_A_193_47#_c_503_n 0.00687211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_193_47#_c_509_n 0.0117991f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_110 VPB N_A_193_47#_c_505_n 0.00814268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_193_47#_c_511_n 0.00297592f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_112 VPB N_A_193_47#_c_512_n 0.00564475f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_113 VPB N_A_193_47#_c_513_n 0.00239973f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_114 VPB N_A_193_47#_c_514_n 0.00732901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_193_47#_c_515_n 0.00114133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_193_47#_c_516_n 0.0104341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_193_47#_c_517_n 0.0126899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_728_21#_M1007_g 0.0155525f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_119 VPB N_A_728_21#_M1020_g 0.0240498f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_120 VPB N_A_728_21#_M1001_g 0.0186895f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_121 VPB N_A_728_21#_M1011_g 0.0224764f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_122 VPB N_A_728_21#_c_617_n 0.0194636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_728_21#_c_618_n 0.00558514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_728_21#_c_619_n 6.08077e-19 $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_125 VPB N_A_728_21#_c_630_n 0.0170715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_728_21#_c_631_n 0.0183859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_728_21#_c_632_n 0.0184988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_728_21#_c_633_n 0.00678594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_728_21#_c_634_n 0.0413724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_728_21#_c_635_n 0.00368741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_728_21#_c_622_n 0.00281539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_565_413#_M1014_g 0.0223351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_565_413#_c_747_n 0.015753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_565_413#_c_748_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_135 VPB N_A_565_413#_c_755_n 0.00517422f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_136 VPB N_A_565_413#_c_751_n 0.00167692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_1223_47#_M1012_g 0.0198362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_1223_47#_c_831_n 0.00570712f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_139 VPB N_A_1223_47#_M1018_g 0.0265634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_1223_47#_c_840_n 0.0150603f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_141 VPB N_A_1223_47#_c_836_n 0.0054092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_909_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_143 VPB N_VPWR_c_910_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_144 VPB N_VPWR_c_911_n 0.00966208f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_912_n 0.0177191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_913_n 0.00189136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_914_n 0.0114544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_915_n 0.00281522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_916_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_917_n 0.0425526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_918_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_919_n 0.0301497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_920_n 0.0406078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_921_n 0.0153766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_922_n 0.0183604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_923_n 0.0153174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_924_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_925_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_926_n 0.00574408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_927_n 0.00421326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_928_n 0.00516749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_929_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_908_n 0.0655254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_Q_c_1039_n 0.00153052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_Q_N_c_1069_n 0.00222189f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_166 VPB Q_N 0.00509848f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_167 N_GATE_N_c_169_n N_A_27_47#_M1010_g 0.0187834f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_168 N_GATE_N_c_173_n N_A_27_47#_M1010_g 0.00419721f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_169 N_GATE_N_c_176_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_170 N_GATE_N_c_172_n N_A_27_47#_M1000_g 0.00527139f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_171 N_GATE_N_c_169_n N_A_27_47#_c_213_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_172 N_GATE_N_c_170_n N_A_27_47#_c_213_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_173 N_GATE_N_c_170_n N_A_27_47#_c_214_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_174 GATE_N N_A_27_47#_c_214_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_175 N_GATE_N_c_172_n N_A_27_47#_c_214_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_176 N_GATE_N_c_175_n N_A_27_47#_c_224_n 0.0135489f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_177 N_GATE_N_c_176_n N_A_27_47#_c_224_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_178 N_GATE_N_c_175_n N_A_27_47#_c_226_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_179 N_GATE_N_c_176_n N_A_27_47#_c_226_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_180 GATE_N N_A_27_47#_c_226_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_181 N_GATE_N_c_172_n N_A_27_47#_c_226_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_182 N_GATE_N_c_172_n N_A_27_47#_c_215_n 0.00319349f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_183 N_GATE_N_c_170_n N_A_27_47#_c_216_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_184 GATE_N N_A_27_47#_c_216_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_185 N_GATE_N_c_173_n N_A_27_47#_c_216_n 0.00151818f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_186 N_GATE_N_c_174_n N_A_27_47#_c_229_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_187 N_GATE_N_c_176_n N_A_27_47#_c_229_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_188 GATE_N N_A_27_47#_c_229_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_189 N_GATE_N_c_174_n N_A_27_47#_c_230_n 7.602e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_176_n N_A_27_47#_c_230_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_191 GATE_N N_A_27_47#_c_219_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_192 N_GATE_N_c_172_n N_A_27_47#_c_219_n 0.0165768f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_193 N_GATE_N_c_175_n N_VPWR_c_909_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_194 N_GATE_N_c_175_n N_VPWR_c_918_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_195 N_GATE_N_c_175_n N_VPWR_c_908_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_196 N_GATE_N_c_169_n N_VGND_c_1096_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_197 N_GATE_N_c_169_n N_VGND_c_1105_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_198 N_GATE_N_c_170_n N_VGND_c_1105_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_199 N_GATE_N_c_169_n N_VGND_c_1117_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_228_n N_D_M1005_g 0.00583826f $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_228_n N_D_c_381_n 0.0087134f $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1010_g N_D_c_382_n 0.00488997f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_228_n N_A_303_47#_M1004_g 0.00493352f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_221_n N_A_303_47#_M1004_g 0.00369716f $X=3.115 $Y=1.415
+ $X2=0 $Y2=0
cc_205 N_A_27_47#_c_228_n N_A_303_47#_c_428_n 0.0116478f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_228_n N_A_303_47#_c_429_n 0.0115915f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_217_n N_A_303_47#_c_421_n 9.56555e-19 $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_218_n N_A_303_47#_c_421_n 0.0129081f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_228_n N_A_303_47#_c_421_n 0.00675641f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_221_n N_A_303_47#_c_421_n 0.00178567f $X=3.115 $Y=1.415
+ $X2=0 $Y2=0
cc_211 N_A_27_47#_c_228_n N_A_303_47#_c_422_n 0.0108506f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_217_n N_A_303_47#_c_424_n 0.0117556f $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_218_n N_A_303_47#_c_424_n 9.50608e-19 $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_228_n N_A_303_47#_c_424_n 0.00107604f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_221_n N_A_303_47#_c_424_n 9.9633e-19 $X=3.115 $Y=1.415 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_217_n N_A_303_47#_c_425_n 0.00200147f $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_218_n N_A_303_47#_c_425_n 2.04855e-19 $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_220_n N_A_303_47#_c_425_n 0.0197936f $X=2.82 $Y=0.705 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_M1015_g N_A_193_47#_M1013_g 0.014011f $X=3.355 $Y=2.275 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_225_n N_A_193_47#_M1013_g 0.00220245f $X=3.2 $Y=1.74 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_218_n N_A_193_47#_c_502_n 7.03475e-19 $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_228_n N_A_193_47#_c_502_n 0.00144279f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_231_n N_A_193_47#_c_502_n 0.00140497f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_232_n N_A_193_47#_c_502_n 0.0049391f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_234_n N_A_193_47#_c_502_n 0.0184089f $X=3.355 $Y=1.74 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_221_n N_A_193_47#_c_502_n 0.01293f $X=3.115 $Y=1.415 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_217_n N_A_193_47#_c_503_n 0.0186665f $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_218_n N_A_193_47#_c_503_n 0.00136525f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_217_n N_A_193_47#_M1016_g 0.0192792f $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_218_n N_A_193_47#_M1016_g 0.00256371f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_220_n N_A_193_47#_M1016_g 0.0126141f $X=2.82 $Y=0.705 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_221_n N_A_193_47#_M1016_g 0.0049729f $X=3.115 $Y=1.415 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_228_n N_A_193_47#_c_509_n 0.00274258f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_231_n N_A_193_47#_c_509_n 7.88621e-19 $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_232_n N_A_193_47#_c_509_n 0.00220245f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_234_n N_A_193_47#_c_509_n 0.0160512f $X=3.355 $Y=1.74 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1010_g N_A_193_47#_c_505_n 0.00782494f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_213_n N_A_193_47#_c_505_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_215_n N_A_193_47#_c_505_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_216_n N_A_193_47#_c_505_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_228_n N_A_193_47#_c_505_n 0.0185373f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_229_n N_A_193_47#_c_505_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_230_n N_A_193_47#_c_505_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_224_n N_A_193_47#_c_511_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_228_n N_A_193_47#_c_511_n 0.00195186f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_219_n N_A_193_47#_c_511_n 0.00782494f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_228_n N_A_193_47#_c_512_n 0.0887801f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1000_g N_A_193_47#_c_513_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_224_n N_A_193_47#_c_513_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_228_n N_A_193_47#_c_513_n 0.0259095f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_230_n N_A_193_47#_c_513_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1000_g N_A_193_47#_c_514_n 0.00782494f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_225_n N_A_193_47#_c_515_n 0.00155445f $X=3.2 $Y=1.74 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_228_n N_A_193_47#_c_515_n 0.0255946f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_228_n N_A_193_47#_c_516_n 0.00169866f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_231_n N_A_193_47#_c_516_n 0.00124306f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_221_n N_A_193_47#_c_516_n 0.00220245f $X=3.115 $Y=1.415
+ $X2=0 $Y2=0
cc_258 N_A_27_47#_c_217_n N_A_193_47#_c_517_n 4.0812e-19 $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_218_n N_A_193_47#_c_517_n 0.00161882f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_228_n N_A_193_47#_c_517_n 0.0240266f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_231_n N_A_193_47#_c_517_n 0.00272314f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_234_n N_A_193_47#_c_517_n 2.5966e-19 $X=3.355 $Y=1.74 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_221_n N_A_193_47#_c_517_n 0.0454941f $X=3.115 $Y=1.415 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_232_n N_A_728_21#_M1007_g 4.9921e-19 $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_221_n N_A_728_21#_M1007_g 2.17095e-19 $X=3.115 $Y=1.415
+ $X2=0 $Y2=0
cc_266 N_A_27_47#_M1015_g N_A_728_21#_M1020_g 0.0313447f $X=3.355 $Y=2.275 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_225_n N_A_728_21#_c_634_n 8.09252e-19 $X=3.2 $Y=1.74 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_234_n N_A_728_21#_c_634_n 0.0313447f $X=3.355 $Y=1.74 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_217_n N_A_565_413#_c_757_n 0.00144439f $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_218_n N_A_565_413#_c_757_n 0.0162478f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_220_n N_A_565_413#_c_757_n 0.00412044f $X=2.82 $Y=0.705
+ $X2=0 $Y2=0
cc_272 N_A_27_47#_M1015_g N_A_565_413#_c_760_n 0.0116262f $X=3.355 $Y=2.275
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_c_225_n N_A_565_413#_c_760_n 0.016081f $X=3.2 $Y=1.74 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_231_n N_A_565_413#_c_760_n 0.00173361f $X=3.035 $Y=1.53
+ $X2=0 $Y2=0
cc_275 N_A_27_47#_c_234_n N_A_565_413#_c_760_n 0.00111122f $X=3.355 $Y=1.74
+ $X2=0 $Y2=0
cc_276 N_A_27_47#_c_218_n N_A_565_413#_c_749_n 0.0184898f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_218_n N_A_565_413#_c_750_n 0.0027819f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_234_n N_A_565_413#_c_750_n 0.00291146f $X=3.355 $Y=1.74
+ $X2=0 $Y2=0
cc_279 N_A_27_47#_c_221_n N_A_565_413#_c_750_n 0.016104f $X=3.115 $Y=1.415 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_231_n N_A_565_413#_c_755_n 0.00130345f $X=3.035 $Y=1.53
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_232_n N_A_565_413#_c_755_n 0.0359174f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_234_n N_A_565_413#_c_755_n 0.00856317f $X=3.355 $Y=1.74
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_221_n N_A_565_413#_c_755_n 0.00353544f $X=3.115 $Y=1.415
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_c_224_n N_VPWR_M1008_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_285 N_A_27_47#_M1000_g N_VPWR_c_909_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_224_n N_VPWR_c_909_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_226_n N_VPWR_c_909_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_229_n N_VPWR_c_909_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_228_n N_VPWR_c_910_n 0.0019389f $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_224_n N_VPWR_c_918_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_226_n N_VPWR_c_918_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_292 N_A_27_47#_M1000_g N_VPWR_c_919_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1015_g N_VPWR_c_920_n 0.00366111f $X=3.355 $Y=2.275 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1000_g N_VPWR_c_908_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1015_g N_VPWR_c_908_n 0.00549379f $X=3.355 $Y=2.275 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_224_n N_VPWR_c_908_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_226_n N_VPWR_c_908_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_213_n N_VGND_M1022_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_27_47#_M1010_g N_VGND_c_1096_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_213_n N_VGND_c_1096_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_215_n N_VGND_c_1096_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_219_n N_VGND_c_1096_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_220_n N_VGND_c_1097_n 0.00174223f $X=2.82 $Y=0.705 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_366_p N_VGND_c_1105_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_213_n N_VGND_c_1105_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1010_g N_VGND_c_1106_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_217_n N_VGND_c_1107_n 9.43262e-19 $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_218_n N_VGND_c_1107_n 0.00182549f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_220_n N_VGND_c_1107_n 0.00425892f $X=2.82 $Y=0.705 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1022_s N_VGND_c_1117_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_M1010_g N_VGND_c_1117_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_366_p N_VGND_c_1117_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_213_n N_VGND_c_1117_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_217_n N_VGND_c_1117_n 0.00121904f $X=2.82 $Y=0.87 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_218_n N_VGND_c_1117_n 0.00328555f $X=3.03 $Y=0.87 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_220_n N_VGND_c_1117_n 0.00628992f $X=2.82 $Y=0.705 $X2=0
+ $Y2=0
cc_317 N_D_c_382_n N_A_303_47#_M1004_g 0.0382098f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_318 N_D_M1005_g N_A_303_47#_c_427_n 0.012851f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_319 N_D_M1024_g N_A_303_47#_c_420_n 0.0144498f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_320 N_D_c_381_n N_A_303_47#_c_420_n 0.00627239f $X=1.645 $Y=1.04 $X2=0 $Y2=0
cc_321 N_D_c_382_n N_A_303_47#_c_420_n 0.00123166f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_322 N_D_M1005_g N_A_303_47#_c_428_n 0.00794545f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_323 N_D_M1005_g N_A_303_47#_c_429_n 0.00412429f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_324 N_D_c_381_n N_A_303_47#_c_429_n 0.0229667f $X=1.645 $Y=1.04 $X2=0 $Y2=0
cc_325 N_D_c_382_n N_A_303_47#_c_429_n 0.00131849f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_326 N_D_M1024_g N_A_303_47#_c_421_n 0.00563568f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_327 N_D_c_381_n N_A_303_47#_c_421_n 0.0107593f $X=1.645 $Y=1.04 $X2=0 $Y2=0
cc_328 N_D_c_381_n N_A_303_47#_c_422_n 0.0164827f $X=1.645 $Y=1.04 $X2=0 $Y2=0
cc_329 N_D_c_382_n N_A_303_47#_c_422_n 0.00552652f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_330 N_D_M1024_g N_A_303_47#_c_423_n 0.00120855f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_331 N_D_c_381_n N_A_303_47#_c_423_n 0.0138491f $X=1.645 $Y=1.04 $X2=0 $Y2=0
cc_332 N_D_c_382_n N_A_303_47#_c_423_n 0.0042466f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_333 N_D_M1024_g N_A_303_47#_c_424_n 0.0197208f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_334 N_D_M1024_g N_A_303_47#_c_425_n 0.015283f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_335 N_D_M1024_g N_A_193_47#_c_505_n 0.00199368f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_336 N_D_M1005_g N_A_193_47#_c_505_n 0.00451505f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_337 N_D_c_381_n N_A_193_47#_c_505_n 0.0200106f $X=1.645 $Y=1.04 $X2=0 $Y2=0
cc_338 N_D_c_382_n N_A_193_47#_c_505_n 0.00254748f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_339 N_D_M1005_g N_A_193_47#_c_511_n 0.00137923f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_340 N_D_M1005_g N_A_193_47#_c_512_n 0.00294239f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_341 N_D_M1005_g N_VPWR_c_910_n 0.00304701f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_342 N_D_M1005_g N_VPWR_c_919_n 0.00543342f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_343 N_D_M1005_g N_VPWR_c_908_n 0.00734866f $X=1.85 $Y=2.165 $X2=0 $Y2=0
cc_344 N_D_M1024_g N_VGND_c_1097_n 0.0110406f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_345 N_D_M1024_g N_VGND_c_1106_n 0.00337001f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_346 N_D_M1024_g N_VGND_c_1117_n 0.0053254f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_347 N_D_c_382_n N_VGND_c_1117_n 0.00103829f $X=1.85 $Y=1.04 $X2=0 $Y2=0
cc_348 N_A_303_47#_M1004_g N_A_193_47#_M1013_g 0.0342299f $X=2.27 $Y=2.165 $X2=0
+ $Y2=0
cc_349 N_A_303_47#_M1004_g N_A_193_47#_c_503_n 0.0248238f $X=2.27 $Y=2.165 $X2=0
+ $Y2=0
cc_350 N_A_303_47#_c_427_n N_A_193_47#_c_505_n 0.00103987f $X=1.64 $Y=1.99 $X2=0
+ $Y2=0
cc_351 N_A_303_47#_c_429_n N_A_193_47#_c_505_n 0.0082816f $X=1.805 $Y=1.58 $X2=0
+ $Y2=0
cc_352 N_A_303_47#_c_423_n N_A_193_47#_c_505_n 0.0184284f $X=1.64 $Y=0.51 $X2=0
+ $Y2=0
cc_353 N_A_303_47#_c_427_n N_A_193_47#_c_511_n 0.0439827f $X=1.64 $Y=1.99 $X2=0
+ $Y2=0
cc_354 N_A_303_47#_M1004_g N_A_193_47#_c_512_n 0.00365242f $X=2.27 $Y=2.165
+ $X2=0 $Y2=0
cc_355 N_A_303_47#_c_427_n N_A_193_47#_c_512_n 0.0228727f $X=1.64 $Y=1.99 $X2=0
+ $Y2=0
cc_356 N_A_303_47#_c_428_n N_A_193_47#_c_512_n 0.00551435f $X=1.99 $Y=1.58 $X2=0
+ $Y2=0
cc_357 N_A_303_47#_c_427_n N_A_193_47#_c_513_n 0.00270021f $X=1.64 $Y=1.99 $X2=0
+ $Y2=0
cc_358 N_A_303_47#_M1004_g N_A_193_47#_c_515_n 0.00149195f $X=2.27 $Y=2.165
+ $X2=0 $Y2=0
cc_359 N_A_303_47#_M1004_g N_A_193_47#_c_517_n 0.00673436f $X=2.27 $Y=2.165
+ $X2=0 $Y2=0
cc_360 N_A_303_47#_c_428_n N_A_193_47#_c_517_n 0.00754519f $X=1.99 $Y=1.58 $X2=0
+ $Y2=0
cc_361 N_A_303_47#_c_422_n N_A_193_47#_c_517_n 0.00645446f $X=2.075 $Y=1.495
+ $X2=0 $Y2=0
cc_362 N_A_303_47#_c_425_n N_A_565_413#_c_757_n 6.54613e-19 $X=2.275 $Y=0.765
+ $X2=0 $Y2=0
cc_363 N_A_303_47#_M1004_g N_VPWR_c_910_n 0.0223997f $X=2.27 $Y=2.165 $X2=0
+ $Y2=0
cc_364 N_A_303_47#_c_427_n N_VPWR_c_910_n 0.0232987f $X=1.64 $Y=1.99 $X2=0 $Y2=0
cc_365 N_A_303_47#_c_428_n N_VPWR_c_910_n 0.013562f $X=1.99 $Y=1.58 $X2=0 $Y2=0
cc_366 N_A_303_47#_c_427_n N_VPWR_c_919_n 0.0159418f $X=1.64 $Y=1.99 $X2=0 $Y2=0
cc_367 N_A_303_47#_M1004_g N_VPWR_c_920_n 0.00212864f $X=2.27 $Y=2.165 $X2=0
+ $Y2=0
cc_368 N_A_303_47#_M1005_s N_VPWR_c_908_n 0.00174533f $X=1.515 $Y=1.845 $X2=0
+ $Y2=0
cc_369 N_A_303_47#_M1004_g N_VPWR_c_908_n 0.00262666f $X=2.27 $Y=2.165 $X2=0
+ $Y2=0
cc_370 N_A_303_47#_c_427_n N_VPWR_c_908_n 0.00576627f $X=1.64 $Y=1.99 $X2=0
+ $Y2=0
cc_371 N_A_303_47#_c_421_n N_VGND_M1024_d 0.00156939f $X=2.075 $Y=1.095 $X2=0
+ $Y2=0
cc_372 N_A_303_47#_c_420_n N_VGND_c_1097_n 0.00259081f $X=1.99 $Y=0.7 $X2=0
+ $Y2=0
cc_373 N_A_303_47#_c_421_n N_VGND_c_1097_n 0.0141976f $X=2.075 $Y=1.095 $X2=0
+ $Y2=0
cc_374 N_A_303_47#_c_425_n N_VGND_c_1097_n 0.00964732f $X=2.275 $Y=0.765 $X2=0
+ $Y2=0
cc_375 N_A_303_47#_c_420_n N_VGND_c_1106_n 0.00255672f $X=1.99 $Y=0.7 $X2=0
+ $Y2=0
cc_376 N_A_303_47#_c_423_n N_VGND_c_1106_n 0.00711582f $X=1.64 $Y=0.51 $X2=0
+ $Y2=0
cc_377 N_A_303_47#_c_424_n N_VGND_c_1107_n 9.84895e-19 $X=2.275 $Y=0.93 $X2=0
+ $Y2=0
cc_378 N_A_303_47#_c_425_n N_VGND_c_1107_n 0.0046653f $X=2.275 $Y=0.765 $X2=0
+ $Y2=0
cc_379 N_A_303_47#_M1024_s N_VGND_c_1117_n 0.00283248f $X=1.515 $Y=0.235 $X2=0
+ $Y2=0
cc_380 N_A_303_47#_c_420_n N_VGND_c_1117_n 0.00473142f $X=1.99 $Y=0.7 $X2=0
+ $Y2=0
cc_381 N_A_303_47#_c_421_n N_VGND_c_1117_n 0.00552372f $X=2.075 $Y=1.095 $X2=0
+ $Y2=0
cc_382 N_A_303_47#_c_423_n N_VGND_c_1117_n 0.00607883f $X=1.64 $Y=0.51 $X2=0
+ $Y2=0
cc_383 N_A_303_47#_c_424_n N_VGND_c_1117_n 0.00117722f $X=2.275 $Y=0.93 $X2=0
+ $Y2=0
cc_384 N_A_303_47#_c_425_n N_VGND_c_1117_n 0.00454932f $X=2.275 $Y=0.765 $X2=0
+ $Y2=0
cc_385 N_A_193_47#_M1016_g N_A_728_21#_M1007_g 0.0429763f $X=3.24 $Y=0.415 $X2=0
+ $Y2=0
cc_386 N_A_193_47#_M1016_g N_A_565_413#_c_757_n 0.0125662f $X=3.24 $Y=0.415
+ $X2=0 $Y2=0
cc_387 N_A_193_47#_M1013_g N_A_565_413#_c_760_n 0.00281839f $X=2.75 $Y=2.275
+ $X2=0 $Y2=0
cc_388 N_A_193_47#_M1016_g N_A_565_413#_c_749_n 0.00562201f $X=3.24 $Y=0.415
+ $X2=0 $Y2=0
cc_389 N_A_193_47#_M1016_g N_A_565_413#_c_750_n 0.00348305f $X=3.24 $Y=0.415
+ $X2=0 $Y2=0
cc_390 N_A_193_47#_M1013_g N_A_565_413#_c_755_n 8.05921e-19 $X=2.75 $Y=2.275
+ $X2=0 $Y2=0
cc_391 N_A_193_47#_c_502_n N_A_565_413#_c_755_n 6.71539e-19 $X=3.165 $Y=1.32
+ $X2=0 $Y2=0
cc_392 N_A_193_47#_c_512_n N_VPWR_M1005_d 6.81311e-19 $X=2.43 $Y=1.87 $X2=0
+ $Y2=0
cc_393 N_A_193_47#_c_514_n N_VPWR_c_909_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_394 N_A_193_47#_M1013_g N_VPWR_c_910_n 0.00357414f $X=2.75 $Y=2.275 $X2=0
+ $Y2=0
cc_395 N_A_193_47#_c_512_n N_VPWR_c_910_n 0.0171797f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_396 N_A_193_47#_c_515_n N_VPWR_c_910_n 0.0013481f $X=2.575 $Y=1.87 $X2=0
+ $Y2=0
cc_397 N_A_193_47#_c_517_n N_VPWR_c_910_n 0.00972665f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_398 N_A_193_47#_c_514_n N_VPWR_c_919_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_399 N_A_193_47#_M1013_g N_VPWR_c_920_n 0.00487021f $X=2.75 $Y=2.275 $X2=0
+ $Y2=0
cc_400 N_A_193_47#_c_517_n N_VPWR_c_920_n 0.00456724f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_401 N_A_193_47#_M1013_g N_VPWR_c_908_n 0.00815857f $X=2.75 $Y=2.275 $X2=0
+ $Y2=0
cc_402 N_A_193_47#_c_512_n N_VPWR_c_908_n 0.0527463f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_403 N_A_193_47#_c_513_n N_VPWR_c_908_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_404 N_A_193_47#_c_514_n N_VPWR_c_908_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_405 N_A_193_47#_c_515_n N_VPWR_c_908_n 0.0151013f $X=2.575 $Y=1.87 $X2=0
+ $Y2=0
cc_406 N_A_193_47#_c_517_n N_VPWR_c_908_n 0.00403974f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_407 N_A_193_47#_c_512_n A_469_369# 0.00119229f $X=2.43 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_408 N_A_193_47#_c_515_n A_469_369# 0.00120144f $X=2.575 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_409 N_A_193_47#_c_517_n A_469_369# 0.0030615f $X=2.69 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_410 N_A_193_47#_M1016_g N_VGND_c_1098_n 0.0018373f $X=3.24 $Y=0.415 $X2=0
+ $Y2=0
cc_411 N_A_193_47#_c_505_n N_VGND_c_1106_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_412 N_A_193_47#_M1016_g N_VGND_c_1107_n 0.0037981f $X=3.24 $Y=0.415 $X2=0
+ $Y2=0
cc_413 N_A_193_47#_M1010_d N_VGND_c_1117_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_414 N_A_193_47#_M1016_g N_VGND_c_1117_n 0.00555936f $X=3.24 $Y=0.415 $X2=0
+ $Y2=0
cc_415 N_A_193_47#_c_505_n N_VGND_c_1117_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_416 N_A_728_21#_c_615_n N_A_565_413#_c_746_n 0.0209154f $X=5.09 $Y=0.995
+ $X2=0 $Y2=0
cc_417 N_A_728_21#_c_621_n N_A_565_413#_c_746_n 0.00671379f $X=4.495 $Y=0.995
+ $X2=0 $Y2=0
cc_418 N_A_728_21#_M1001_g N_A_565_413#_M1014_g 0.0230216f $X=5.09 $Y=1.985
+ $X2=0 $Y2=0
cc_419 N_A_728_21#_c_634_n N_A_565_413#_M1014_g 0.00346217f $X=3.945 $Y=1.7
+ $X2=0 $Y2=0
cc_420 N_A_728_21#_c_635_n N_A_565_413#_M1014_g 0.00755466f $X=4.495 $Y=1.535
+ $X2=0 $Y2=0
cc_421 N_A_728_21#_c_648_p N_A_565_413#_M1014_g 3.06193e-19 $X=4.445 $Y=1.755
+ $X2=0 $Y2=0
cc_422 N_A_728_21#_M1007_g N_A_565_413#_c_747_n 0.0214321f $X=3.715 $Y=0.445
+ $X2=0 $Y2=0
cc_423 N_A_728_21#_c_633_n N_A_565_413#_c_747_n 0.00879412f $X=4.36 $Y=1.7 $X2=0
+ $Y2=0
cc_424 N_A_728_21#_c_634_n N_A_565_413#_c_747_n 0.00487525f $X=3.945 $Y=1.7
+ $X2=0 $Y2=0
cc_425 N_A_728_21#_c_652_p N_A_565_413#_c_747_n 0.00203472f $X=4.47 $Y=0.825
+ $X2=0 $Y2=0
cc_426 N_A_728_21#_c_648_p N_A_565_413#_c_747_n 0.00212837f $X=4.445 $Y=1.755
+ $X2=0 $Y2=0
cc_427 N_A_728_21#_c_654_p N_A_565_413#_c_747_n 0.0181635f $X=4.495 $Y=1.16
+ $X2=0 $Y2=0
cc_428 N_A_728_21#_c_618_n N_A_565_413#_c_748_n 0.0216214f $X=5.585 $Y=1.16
+ $X2=0 $Y2=0
cc_429 N_A_728_21#_c_622_n N_A_565_413#_c_748_n 0.0218433f $X=5.075 $Y=1.16
+ $X2=0 $Y2=0
cc_430 N_A_728_21#_M1007_g N_A_565_413#_c_757_n 0.00148607f $X=3.715 $Y=0.445
+ $X2=0 $Y2=0
cc_431 N_A_728_21#_M1020_g N_A_565_413#_c_760_n 0.00369776f $X=3.715 $Y=2.275
+ $X2=0 $Y2=0
cc_432 N_A_728_21#_M1007_g N_A_565_413#_c_749_n 0.00598699f $X=3.715 $Y=0.445
+ $X2=0 $Y2=0
cc_433 N_A_728_21#_M1007_g N_A_565_413#_c_750_n 0.00570022f $X=3.715 $Y=0.445
+ $X2=0 $Y2=0
cc_434 N_A_728_21#_M1007_g N_A_565_413#_c_755_n 0.0114233f $X=3.715 $Y=0.445
+ $X2=0 $Y2=0
cc_435 N_A_728_21#_M1020_g N_A_565_413#_c_755_n 0.0143765f $X=3.715 $Y=2.275
+ $X2=0 $Y2=0
cc_436 N_A_728_21#_c_633_n N_A_565_413#_c_755_n 0.022954f $X=4.36 $Y=1.7 $X2=0
+ $Y2=0
cc_437 N_A_728_21#_c_634_n N_A_565_413#_c_755_n 0.00824307f $X=3.945 $Y=1.7
+ $X2=0 $Y2=0
cc_438 N_A_728_21#_M1007_g N_A_565_413#_c_751_n 0.0170014f $X=3.715 $Y=0.445
+ $X2=0 $Y2=0
cc_439 N_A_728_21#_c_633_n N_A_565_413#_c_751_n 0.02399f $X=4.36 $Y=1.7 $X2=0
+ $Y2=0
cc_440 N_A_728_21#_c_634_n N_A_565_413#_c_751_n 0.006103f $X=3.945 $Y=1.7 $X2=0
+ $Y2=0
cc_441 N_A_728_21#_c_654_p N_A_565_413#_c_751_n 0.0254258f $X=4.495 $Y=1.16
+ $X2=0 $Y2=0
cc_442 N_A_728_21#_c_619_n N_A_1223_47#_c_829_n 0.00249753f $X=6.32 $Y=1.325
+ $X2=0 $Y2=0
cc_443 N_A_728_21#_c_620_n N_A_1223_47#_c_829_n 0.0159717f $X=6.45 $Y=0.73 $X2=0
+ $Y2=0
cc_444 N_A_728_21#_c_630_n N_A_1223_47#_M1012_g 0.00638756f $X=6.32 $Y=1.62
+ $X2=0 $Y2=0
cc_445 N_A_728_21#_c_632_n N_A_1223_47#_M1012_g 0.0124781f $X=6.45 $Y=1.695
+ $X2=0 $Y2=0
cc_446 N_A_728_21#_c_619_n N_A_1223_47#_c_831_n 0.0132452f $X=6.32 $Y=1.325
+ $X2=0 $Y2=0
cc_447 N_A_728_21#_c_616_n N_A_1223_47#_c_835_n 0.00524028f $X=5.51 $Y=0.995
+ $X2=0 $Y2=0
cc_448 N_A_728_21#_c_619_n N_A_1223_47#_c_835_n 0.0139898f $X=6.32 $Y=1.325
+ $X2=0 $Y2=0
cc_449 N_A_728_21#_c_620_n N_A_1223_47#_c_835_n 0.00969929f $X=6.45 $Y=0.73
+ $X2=0 $Y2=0
cc_450 N_A_728_21#_M1011_g N_A_1223_47#_c_840_n 0.00523864f $X=5.51 $Y=1.985
+ $X2=0 $Y2=0
cc_451 N_A_728_21#_c_630_n N_A_1223_47#_c_840_n 0.0101898f $X=6.32 $Y=1.62 $X2=0
+ $Y2=0
cc_452 N_A_728_21#_c_631_n N_A_1223_47#_c_840_n 0.00975787f $X=6.45 $Y=1.77
+ $X2=0 $Y2=0
cc_453 N_A_728_21#_c_632_n N_A_1223_47#_c_840_n 0.0102457f $X=6.45 $Y=1.695
+ $X2=0 $Y2=0
cc_454 N_A_728_21#_c_619_n N_A_1223_47#_c_836_n 0.00562989f $X=6.32 $Y=1.325
+ $X2=0 $Y2=0
cc_455 N_A_728_21#_c_632_n N_A_1223_47#_c_836_n 0.0046403f $X=6.45 $Y=1.695
+ $X2=0 $Y2=0
cc_456 N_A_728_21#_c_617_n N_A_1223_47#_c_856_n 0.0139296f $X=6.245 $Y=1.16
+ $X2=0 $Y2=0
cc_457 N_A_728_21#_c_619_n N_A_1223_47#_c_856_n 0.00895211f $X=6.32 $Y=1.325
+ $X2=0 $Y2=0
cc_458 N_A_728_21#_M1020_g N_VPWR_c_911_n 0.00454869f $X=3.715 $Y=2.275 $X2=0
+ $Y2=0
cc_459 N_A_728_21#_c_633_n N_VPWR_c_911_n 0.0154822f $X=4.36 $Y=1.7 $X2=0 $Y2=0
cc_460 N_A_728_21#_c_634_n N_VPWR_c_911_n 0.00545641f $X=3.945 $Y=1.7 $X2=0
+ $Y2=0
cc_461 N_A_728_21#_c_688_p N_VPWR_c_911_n 0.0196384f $X=4.445 $Y=2.27 $X2=0
+ $Y2=0
cc_462 N_A_728_21#_c_688_p N_VPWR_c_912_n 0.0112378f $X=4.445 $Y=2.27 $X2=0
+ $Y2=0
cc_463 N_A_728_21#_M1001_g N_VPWR_c_913_n 0.0171275f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_464 N_A_728_21#_M1011_g N_VPWR_c_913_n 8.65231e-19 $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_465 N_A_728_21#_c_618_n N_VPWR_c_913_n 0.00157349f $X=5.585 $Y=1.16 $X2=0
+ $Y2=0
cc_466 N_A_728_21#_c_622_n N_VPWR_c_913_n 0.020301f $X=5.075 $Y=1.16 $X2=0 $Y2=0
cc_467 N_A_728_21#_M1011_g N_VPWR_c_914_n 0.00312709f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_468 N_A_728_21#_c_617_n N_VPWR_c_914_n 0.0042583f $X=6.245 $Y=1.16 $X2=0
+ $Y2=0
cc_469 N_A_728_21#_c_631_n N_VPWR_c_914_n 0.00329695f $X=6.45 $Y=1.77 $X2=0
+ $Y2=0
cc_470 N_A_728_21#_c_631_n N_VPWR_c_915_n 0.00537515f $X=6.45 $Y=1.77 $X2=0
+ $Y2=0
cc_471 N_A_728_21#_M1020_g N_VPWR_c_920_n 0.00541489f $X=3.715 $Y=2.275 $X2=0
+ $Y2=0
cc_472 N_A_728_21#_M1001_g N_VPWR_c_921_n 0.0046653f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_728_21#_M1011_g N_VPWR_c_921_n 0.00541763f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_474 N_A_728_21#_c_631_n N_VPWR_c_922_n 0.00541359f $X=6.45 $Y=1.77 $X2=0
+ $Y2=0
cc_475 N_A_728_21#_M1014_s N_VPWR_c_908_n 0.0023739f $X=4.32 $Y=1.485 $X2=0
+ $Y2=0
cc_476 N_A_728_21#_M1020_g N_VPWR_c_908_n 0.0106979f $X=3.715 $Y=2.275 $X2=0
+ $Y2=0
cc_477 N_A_728_21#_M1001_g N_VPWR_c_908_n 0.00789179f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_478 N_A_728_21#_M1011_g N_VPWR_c_908_n 0.010828f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_479 N_A_728_21#_c_631_n N_VPWR_c_908_n 0.0110094f $X=6.45 $Y=1.77 $X2=0 $Y2=0
cc_480 N_A_728_21#_c_633_n N_VPWR_c_908_n 0.00898578f $X=4.36 $Y=1.7 $X2=0 $Y2=0
cc_481 N_A_728_21#_c_634_n N_VPWR_c_908_n 0.00110429f $X=3.945 $Y=1.7 $X2=0
+ $Y2=0
cc_482 N_A_728_21#_c_688_p N_VPWR_c_908_n 0.00827281f $X=4.445 $Y=2.27 $X2=0
+ $Y2=0
cc_483 N_A_728_21#_c_616_n N_Q_c_1040_n 0.009438f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_484 N_A_728_21#_c_618_n N_Q_c_1040_n 0.00217272f $X=5.585 $Y=1.16 $X2=0 $Y2=0
cc_485 N_A_728_21#_c_615_n N_Q_c_1038_n 0.00349798f $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_486 N_A_728_21#_c_616_n N_Q_c_1038_n 0.00491792f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_487 N_A_728_21#_c_618_n N_Q_c_1038_n 8.95338e-19 $X=5.585 $Y=1.16 $X2=0 $Y2=0
cc_488 N_A_728_21#_M1001_g N_Q_c_1039_n 0.00349798f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_489 N_A_728_21#_M1011_g N_Q_c_1039_n 0.00491792f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_490 N_A_728_21#_c_618_n N_Q_c_1039_n 9.16513e-19 $X=5.585 $Y=1.16 $X2=0 $Y2=0
cc_491 N_A_728_21#_M1011_g N_Q_c_1048_n 0.0079195f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_492 N_A_728_21#_c_618_n N_Q_c_1048_n 0.00226238f $X=5.585 $Y=1.16 $X2=0 $Y2=0
cc_493 N_A_728_21#_M1011_g Q 0.0103096f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_494 N_A_728_21#_c_617_n Q 0.0270569f $X=6.245 $Y=1.16 $X2=0 $Y2=0
cc_495 N_A_728_21#_c_618_n Q 0.0217813f $X=5.585 $Y=1.16 $X2=0 $Y2=0
cc_496 N_A_728_21#_c_622_n Q 0.0274156f $X=5.075 $Y=1.16 $X2=0 $Y2=0
cc_497 N_A_728_21#_M1007_g N_VGND_c_1098_n 0.018542f $X=3.715 $Y=0.445 $X2=0
+ $Y2=0
cc_498 N_A_728_21#_c_725_p N_VGND_c_1098_n 0.023358f $X=4.445 $Y=0.58 $X2=0
+ $Y2=0
cc_499 N_A_728_21#_c_725_p N_VGND_c_1099_n 0.00652583f $X=4.445 $Y=0.58 $X2=0
+ $Y2=0
cc_500 N_A_728_21#_c_615_n N_VGND_c_1100_n 0.0136528f $X=5.09 $Y=0.995 $X2=0
+ $Y2=0
cc_501 N_A_728_21#_c_616_n N_VGND_c_1100_n 0.00108124f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_728_21#_c_618_n N_VGND_c_1100_n 0.00157349f $X=5.585 $Y=1.16 $X2=0
+ $Y2=0
cc_503 N_A_728_21#_c_622_n N_VGND_c_1100_n 0.020301f $X=5.075 $Y=1.16 $X2=0
+ $Y2=0
cc_504 N_A_728_21#_c_616_n N_VGND_c_1101_n 0.00312709f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_728_21#_c_617_n N_VGND_c_1101_n 0.0044252f $X=6.245 $Y=1.16 $X2=0
+ $Y2=0
cc_506 N_A_728_21#_c_620_n N_VGND_c_1101_n 0.00316893f $X=6.45 $Y=0.73 $X2=0
+ $Y2=0
cc_507 N_A_728_21#_c_620_n N_VGND_c_1102_n 0.00420958f $X=6.45 $Y=0.73 $X2=0
+ $Y2=0
cc_508 N_A_728_21#_M1007_g N_VGND_c_1107_n 0.0046653f $X=3.715 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_728_21#_c_615_n N_VGND_c_1108_n 0.0046653f $X=5.09 $Y=0.995 $X2=0
+ $Y2=0
cc_510 N_A_728_21#_c_616_n N_VGND_c_1108_n 0.00509502f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_511 N_A_728_21#_c_619_n N_VGND_c_1109_n 2.96334e-19 $X=6.32 $Y=1.325 $X2=0
+ $Y2=0
cc_512 N_A_728_21#_c_620_n N_VGND_c_1109_n 0.00541359f $X=6.45 $Y=0.73 $X2=0
+ $Y2=0
cc_513 N_A_728_21#_M1002_s N_VGND_c_1117_n 0.00370868f $X=4.32 $Y=0.235 $X2=0
+ $Y2=0
cc_514 N_A_728_21#_M1007_g N_VGND_c_1117_n 0.00813035f $X=3.715 $Y=0.445 $X2=0
+ $Y2=0
cc_515 N_A_728_21#_c_615_n N_VGND_c_1117_n 0.00796766f $X=5.09 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_A_728_21#_c_616_n N_VGND_c_1117_n 0.00972138f $X=5.51 $Y=0.995 $X2=0
+ $Y2=0
cc_517 N_A_728_21#_c_620_n N_VGND_c_1117_n 0.0110992f $X=6.45 $Y=0.73 $X2=0
+ $Y2=0
cc_518 N_A_728_21#_c_725_p N_VGND_c_1117_n 0.00762661f $X=4.445 $Y=0.58 $X2=0
+ $Y2=0
cc_519 N_A_565_413#_c_760_n N_VPWR_c_910_n 0.00489615f $X=3.5 $Y=2.34 $X2=0
+ $Y2=0
cc_520 N_A_565_413#_M1014_g N_VPWR_c_911_n 0.00250378f $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_521 N_A_565_413#_M1014_g N_VPWR_c_912_n 0.00585385f $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_522 N_A_565_413#_M1014_g N_VPWR_c_913_n 0.00272345f $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_523 N_A_565_413#_c_760_n N_VPWR_c_920_n 0.0343719f $X=3.5 $Y=2.34 $X2=0 $Y2=0
cc_524 N_A_565_413#_M1013_d N_VPWR_c_908_n 0.00699187f $X=2.825 $Y=2.065 $X2=0
+ $Y2=0
cc_525 N_A_565_413#_M1014_g N_VPWR_c_908_n 0.0120037f $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_526 N_A_565_413#_c_760_n N_VPWR_c_908_n 0.0265731f $X=3.5 $Y=2.34 $X2=0 $Y2=0
cc_527 N_A_565_413#_c_760_n A_686_413# 0.00145479f $X=3.5 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_528 N_A_565_413#_c_755_n A_686_413# 0.00208506f $X=3.585 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_529 N_A_565_413#_c_757_n N_VGND_c_1097_n 0.00209539f $X=3.35 $Y=0.45 $X2=0
+ $Y2=0
cc_530 N_A_565_413#_c_746_n N_VGND_c_1098_n 0.00488932f $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_565_413#_c_747_n N_VGND_c_1098_n 0.00207331f $X=4.58 $Y=1.16 $X2=0
+ $Y2=0
cc_532 N_A_565_413#_c_757_n N_VGND_c_1098_n 0.01074f $X=3.35 $Y=0.45 $X2=0 $Y2=0
cc_533 N_A_565_413#_c_749_n N_VGND_c_1098_n 0.0166369f $X=3.435 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_A_565_413#_c_751_n N_VGND_c_1098_n 0.0283975f $X=4.135 $Y=1.16 $X2=0
+ $Y2=0
cc_535 N_A_565_413#_c_746_n N_VGND_c_1099_n 0.00585385f $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_A_565_413#_c_746_n N_VGND_c_1100_n 0.00253505f $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_537 N_A_565_413#_c_757_n N_VGND_c_1107_n 0.0221606f $X=3.35 $Y=0.45 $X2=0
+ $Y2=0
cc_538 N_A_565_413#_M1006_d N_VGND_c_1117_n 0.00237979f $X=2.885 $Y=0.235 $X2=0
+ $Y2=0
cc_539 N_A_565_413#_c_746_n N_VGND_c_1117_n 0.0120818f $X=4.655 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_A_565_413#_c_757_n N_VGND_c_1117_n 0.0222941f $X=3.35 $Y=0.45 $X2=0
+ $Y2=0
cc_541 N_A_565_413#_c_757_n A_663_47# 0.00369541f $X=3.35 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_542 N_A_565_413#_c_749_n A_663_47# 0.00128174f $X=3.435 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_543 N_A_1223_47#_c_840_n N_VPWR_c_914_n 0.0516742f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_544 N_A_1223_47#_M1012_g N_VPWR_c_915_n 0.0114729f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_545 N_A_1223_47#_c_831_n N_VPWR_c_915_n 0.00244466f $X=7 $Y=1.16 $X2=0 $Y2=0
cc_546 N_A_1223_47#_M1018_g N_VPWR_c_915_n 7.50282e-19 $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_547 N_A_1223_47#_c_840_n N_VPWR_c_915_n 0.0464059f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_548 N_A_1223_47#_c_836_n N_VPWR_c_915_n 0.00959603f $X=6.84 $Y=1.16 $X2=0
+ $Y2=0
cc_549 N_A_1223_47#_M1018_g N_VPWR_c_917_n 0.00312874f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_550 N_A_1223_47#_c_840_n N_VPWR_c_922_n 0.0210382f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_551 N_A_1223_47#_M1012_g N_VPWR_c_923_n 0.0046653f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_552 N_A_1223_47#_M1018_g N_VPWR_c_923_n 0.00541359f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_553 N_A_1223_47#_M1025_s N_VPWR_c_908_n 0.00209319f $X=6.115 $Y=1.845 $X2=0
+ $Y2=0
cc_554 N_A_1223_47#_M1012_g N_VPWR_c_908_n 0.00798142f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_555 N_A_1223_47#_M1018_g N_VPWR_c_908_n 0.0105084f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_556 N_A_1223_47#_c_840_n N_VPWR_c_908_n 0.0124268f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_557 N_A_1223_47#_c_835_n N_Q_c_1040_n 0.00857632f $X=6.24 $Y=0.51 $X2=0 $Y2=0
cc_558 N_A_1223_47#_c_835_n N_Q_c_1038_n 0.00510033f $X=6.24 $Y=0.51 $X2=0 $Y2=0
cc_559 N_A_1223_47#_c_840_n N_Q_c_1039_n 0.0118252f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_560 N_A_1223_47#_c_840_n Q 0.00368257f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_561 N_A_1223_47#_c_856_n Q 0.0274156f $X=6.24 $Y=1.16 $X2=0 $Y2=0
cc_562 N_A_1223_47#_c_829_n N_Q_N_c_1067_n 0.00421369f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_563 N_A_1223_47#_c_830_n N_Q_N_c_1067_n 0.00306399f $X=7.275 $Y=1.16 $X2=0
+ $Y2=0
cc_564 N_A_1223_47#_M1021_g N_Q_N_c_1067_n 0.00803505f $X=7.35 $Y=0.56 $X2=0
+ $Y2=0
cc_565 N_A_1223_47#_c_834_n N_Q_N_c_1067_n 0.00120998f $X=7.35 $Y=1.16 $X2=0
+ $Y2=0
cc_566 N_A_1223_47#_c_836_n N_Q_N_c_1067_n 0.00463694f $X=6.84 $Y=1.16 $X2=0
+ $Y2=0
cc_567 N_A_1223_47#_M1021_g N_Q_N_c_1076_n 0.00202845f $X=7.35 $Y=0.56 $X2=0
+ $Y2=0
cc_568 N_A_1223_47#_M1012_g N_Q_N_c_1069_n 9.04394e-19 $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_569 N_A_1223_47#_c_830_n N_Q_N_c_1069_n 0.0097645f $X=7.275 $Y=1.16 $X2=0
+ $Y2=0
cc_570 N_A_1223_47#_c_831_n N_Q_N_c_1069_n 0.00309279f $X=7 $Y=1.16 $X2=0 $Y2=0
cc_571 N_A_1223_47#_M1018_g N_Q_N_c_1069_n 0.0104283f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_572 N_A_1223_47#_c_834_n N_Q_N_c_1069_n 6.77984e-19 $X=7.35 $Y=1.16 $X2=0
+ $Y2=0
cc_573 N_A_1223_47#_c_840_n N_Q_N_c_1069_n 0.00268711f $X=6.24 $Y=2 $X2=0 $Y2=0
cc_574 N_A_1223_47#_c_836_n N_Q_N_c_1069_n 0.0227962f $X=6.84 $Y=1.16 $X2=0
+ $Y2=0
cc_575 N_A_1223_47#_M1021_g Q_N 0.0061015f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_576 N_A_1223_47#_M1018_g Q_N 0.0115188f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_577 N_A_1223_47#_M1018_g Q_N 0.00643425f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_578 N_A_1223_47#_c_834_n Q_N 0.0130776f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_579 N_A_1223_47#_c_835_n N_VGND_c_1101_n 0.0237866f $X=6.24 $Y=0.51 $X2=0
+ $Y2=0
cc_580 N_A_1223_47#_c_829_n N_VGND_c_1102_n 0.00787161f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_581 N_A_1223_47#_c_831_n N_VGND_c_1102_n 0.00255976f $X=7 $Y=1.16 $X2=0 $Y2=0
cc_582 N_A_1223_47#_M1021_g N_VGND_c_1102_n 6.5116e-19 $X=7.35 $Y=0.56 $X2=0
+ $Y2=0
cc_583 N_A_1223_47#_c_835_n N_VGND_c_1102_n 0.0213546f $X=6.24 $Y=0.51 $X2=0
+ $Y2=0
cc_584 N_A_1223_47#_c_836_n N_VGND_c_1102_n 0.0104995f $X=6.84 $Y=1.16 $X2=0
+ $Y2=0
cc_585 N_A_1223_47#_M1021_g N_VGND_c_1104_n 0.00312874f $X=7.35 $Y=0.56 $X2=0
+ $Y2=0
cc_586 N_A_1223_47#_c_835_n N_VGND_c_1109_n 0.0210709f $X=6.24 $Y=0.51 $X2=0
+ $Y2=0
cc_587 N_A_1223_47#_c_829_n N_VGND_c_1110_n 0.0046653f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_588 N_A_1223_47#_M1021_g N_VGND_c_1110_n 0.00541359f $X=7.35 $Y=0.56 $X2=0
+ $Y2=0
cc_589 N_A_1223_47#_M1009_s N_VGND_c_1117_n 0.00210122f $X=6.115 $Y=0.235 $X2=0
+ $Y2=0
cc_590 N_A_1223_47#_c_829_n N_VGND_c_1117_n 0.00798142f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_591 N_A_1223_47#_M1021_g N_VGND_c_1117_n 0.0105084f $X=7.35 $Y=0.56 $X2=0
+ $Y2=0
cc_592 N_A_1223_47#_c_835_n N_VGND_c_1117_n 0.0124992f $X=6.24 $Y=0.51 $X2=0
+ $Y2=0
cc_593 N_VPWR_c_908_n A_469_369# 0.00373974f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_594 N_VPWR_c_908_n A_686_413# 0.00170472f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_595 N_VPWR_c_908_n N_Q_M1001_d 0.00389051f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_596 N_VPWR_c_921_n Q 0.0142437f $X=5.635 $Y=2.72 $X2=0 $Y2=0
cc_597 N_VPWR_c_908_n Q 0.00930022f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_598 N_VPWR_c_914_n Q 0.00941311f $X=5.72 $Y=2 $X2=0 $Y2=0
cc_599 N_VPWR_c_908_n N_Q_N_M1012_s 0.00397872f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_600 N_VPWR_c_923_n Q_N 0.0155342f $X=7.475 $Y=2.72 $X2=0 $Y2=0
cc_601 N_VPWR_c_908_n Q_N 0.00961085f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_602 N_VPWR_c_917_n Q_N 0.021861f $X=7.56 $Y=1.66 $X2=0 $Y2=0
cc_603 Q N_VGND_c_1101_n 0.0103416f $X=5.73 $Y=1.105 $X2=0 $Y2=0
cc_604 N_Q_c_1040_n N_VGND_c_1108_n 0.00790409f $X=5.415 $Y=0.825 $X2=0 $Y2=0
cc_605 N_Q_M1019_s N_VGND_c_1117_n 0.00409776f $X=5.165 $Y=0.235 $X2=0 $Y2=0
cc_606 N_Q_c_1040_n N_VGND_c_1117_n 0.00934436f $X=5.415 $Y=0.825 $X2=0 $Y2=0
cc_607 Q_N N_VGND_c_1104_n 0.021861f $X=7.555 $Y=1.105 $X2=0 $Y2=0
cc_608 Q_N N_VGND_c_1110_n 0.0155f $X=7.095 $Y=0.425 $X2=0 $Y2=0
cc_609 N_Q_N_M1017_s N_VGND_c_1117_n 0.00397872f $X=7 $Y=0.235 $X2=0 $Y2=0
cc_610 Q_N N_VGND_c_1117_n 0.0096031f $X=7.095 $Y=0.425 $X2=0 $Y2=0
cc_611 N_VGND_c_1117_n A_469_47# 0.0139156f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_612 N_VGND_c_1117_n A_663_47# 0.00687059f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__inv_6.spice
* Created: Tue Sep  1 19:10:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__inv_6.pex.spice"
.subckt sky130_fd_sc_hd__inv_6  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.247 PD=0.92 PS=2.06 NRD=0 NRS=21.228 M=1 R=4.33333 SA=75000.3
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1010_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1755 PD=0.92 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.43
+ AS=0.135 PD=2.86 PS=1.27 NRD=32.4853 NRS=0 M=1 R=6.66667 SA=75000.4 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1001_d N_A_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.2 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1006 N_VPWR_M1003_d N_A_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.27
+ AS=0.135 PD=2.54 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__inv_6.pxi.spice"
*
.ends
*
*

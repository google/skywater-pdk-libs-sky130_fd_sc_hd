* File: sky130_fd_sc_hd__sdlclkp_2.spice.SKY130_FD_SC_HD__SDLCLKP_2.pxi
* Created: Thu Aug 27 14:47:46 2020
* 
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%SCE N_SCE_M1023_g N_SCE_M1011_g SCE SCE
+ N_SCE_c_142_n PM_SKY130_FD_SC_HD__SDLCLKP_2%SCE
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%GATE N_GATE_M1003_g N_GATE_M1010_g GATE GATE
+ N_GATE_c_168_n N_GATE_c_169_n PM_SKY130_FD_SC_HD__SDLCLKP_2%GATE
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%A_257_147# N_A_257_147#_M1020_d
+ N_A_257_147#_M1007_d N_A_257_147#_M1005_g N_A_257_147#_M1009_g
+ N_A_257_147#_M1016_g N_A_257_147#_M1001_g N_A_257_147#_c_211_n
+ N_A_257_147#_c_212_n N_A_257_147#_c_213_n N_A_257_147#_c_214_n
+ N_A_257_147#_c_215_n N_A_257_147#_c_222_n N_A_257_147#_c_216_n
+ N_A_257_147#_c_217_n N_A_257_147#_c_218_n N_A_257_147#_c_219_n
+ N_A_257_147#_c_224_n N_A_257_147#_c_236_n N_A_257_147#_c_225_n
+ N_A_257_147#_c_226_n N_A_257_147#_c_227_n N_A_257_147#_c_228_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%A_257_147#
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%A_257_243# N_A_257_243#_M1016_s
+ N_A_257_243#_M1001_s N_A_257_243#_M1021_g N_A_257_243#_c_389_n
+ N_A_257_243#_c_390_n N_A_257_243#_M1017_g N_A_257_243#_c_391_n
+ N_A_257_243#_c_392_n N_A_257_243#_c_393_n N_A_257_243#_c_405_n
+ N_A_257_243#_c_432_n N_A_257_243#_c_394_n N_A_257_243#_c_395_n
+ N_A_257_243#_c_396_n N_A_257_243#_c_397_n N_A_257_243#_c_398_n
+ N_A_257_243#_c_399_n N_A_257_243#_c_400_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%A_257_243#
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%A_465_315# N_A_465_315#_M1006_d
+ N_A_465_315#_M1000_d N_A_465_315#_M1018_g N_A_465_315#_M1012_g
+ N_A_465_315#_M1014_g N_A_465_315#_M1008_g N_A_465_315#_c_516_n
+ N_A_465_315#_c_511_n N_A_465_315#_c_530_n N_A_465_315#_c_518_n
+ N_A_465_315#_c_519_n N_A_465_315#_c_520_n N_A_465_315#_c_541_n
+ N_A_465_315#_c_542_n N_A_465_315#_c_521_n N_A_465_315#_c_522_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%A_465_315#
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%A_287_413# N_A_287_413#_M1005_d
+ N_A_287_413#_M1021_d N_A_287_413#_c_637_n N_A_287_413#_M1006_g
+ N_A_287_413#_M1000_g N_A_287_413#_c_648_n N_A_287_413#_c_652_n
+ N_A_287_413#_c_643_n N_A_287_413#_c_638_n N_A_287_413#_c_639_n
+ N_A_287_413#_c_640_n N_A_287_413#_c_641_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%A_287_413#
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%CLK N_CLK_M1020_g N_CLK_c_736_n N_CLK_M1007_g
+ N_CLK_M1015_g N_CLK_M1022_g N_CLK_c_739_n N_CLK_c_740_n N_CLK_c_741_n CLK
+ N_CLK_c_742_n N_CLK_c_747_n N_CLK_c_743_n N_CLK_c_744_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%CLK
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%A_1020_47# N_A_1020_47#_M1014_s
+ N_A_1020_47#_M1008_d N_A_1020_47#_c_816_n N_A_1020_47#_M1002_g
+ N_A_1020_47#_M1013_g N_A_1020_47#_c_817_n N_A_1020_47#_M1004_g
+ N_A_1020_47#_M1019_g N_A_1020_47#_c_827_n N_A_1020_47#_c_818_n
+ N_A_1020_47#_c_819_n N_A_1020_47#_c_820_n N_A_1020_47#_c_821_n
+ N_A_1020_47#_c_822_n PM_SKY130_FD_SC_HD__SDLCLKP_2%A_1020_47#
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%VPWR N_VPWR_M1011_s N_VPWR_M1018_d
+ N_VPWR_M1001_d N_VPWR_M1008_s N_VPWR_M1022_d N_VPWR_M1019_d N_VPWR_c_899_n
+ N_VPWR_c_900_n N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n
+ N_VPWR_c_905_n VPWR N_VPWR_c_906_n N_VPWR_c_907_n N_VPWR_c_908_n
+ N_VPWR_c_909_n N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_898_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%VPWR
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%A_27_47# N_A_27_47#_M1023_s N_A_27_47#_M1010_d
+ N_A_27_47#_M1003_d N_A_27_47#_c_1000_n N_A_27_47#_c_1001_n N_A_27_47#_c_1002_n
+ N_A_27_47#_c_1003_n N_A_27_47#_c_1012_n N_A_27_47#_c_1020_n
+ N_A_27_47#_c_1025_n PM_SKY130_FD_SC_HD__SDLCLKP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%GCLK N_GCLK_M1002_s N_GCLK_M1013_s
+ N_GCLK_c_1052_n N_GCLK_c_1061_n N_GCLK_c_1063_n N_GCLK_c_1054_n
+ N_GCLK_c_1069_n GCLK GCLK GCLK GCLK N_GCLK_c_1073_n GCLK
+ PM_SKY130_FD_SC_HD__SDLCLKP_2%GCLK
x_PM_SKY130_FD_SC_HD__SDLCLKP_2%VGND N_VGND_M1023_d N_VGND_M1012_d
+ N_VGND_M1016_d N_VGND_M1015_d N_VGND_M1004_d N_VGND_c_1082_n N_VGND_c_1083_n
+ N_VGND_c_1084_n N_VGND_c_1085_n N_VGND_c_1086_n VGND N_VGND_c_1087_n
+ N_VGND_c_1088_n N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n
+ N_VGND_c_1092_n N_VGND_c_1093_n N_VGND_c_1094_n N_VGND_c_1095_n
+ N_VGND_c_1096_n PM_SKY130_FD_SC_HD__SDLCLKP_2%VGND
cc_1 VNB N_SCE_M1023_g 0.0353283f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB SCE 0.0152509f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_SCE_c_142_n 0.0345609f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_GATE_M1010_g 0.0276674f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_5 VNB N_GATE_c_168_n 0.0274229f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_6 VNB N_GATE_c_169_n 0.00458727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_257_147#_M1005_g 0.0195404f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_257_147#_M1016_g 0.0380294f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_9 VNB N_A_257_147#_c_211_n 0.00683453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_257_147#_c_212_n 0.026946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_257_147#_c_213_n 0.00464205f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_257_147#_c_214_n 0.00396482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_257_147#_c_215_n 8.01096e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_257_147#_c_216_n 0.00256965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_257_147#_c_217_n 0.00348885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_257_147#_c_218_n 0.00214693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_257_147#_c_219_n 0.0237398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_257_243#_c_389_n 0.0152184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_257_243#_c_390_n 0.00503808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_257_243#_c_391_n 0.0111999f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_21 VNB N_A_257_243#_c_392_n 0.00809335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_257_243#_c_393_n 0.00729754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_257_243#_c_394_n 0.00830168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_257_243#_c_395_n 0.00127255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_257_243#_c_396_n 0.00222987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_257_243#_c_397_n 0.00452491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_257_243#_c_398_n 0.0269987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_257_243#_c_399_n 0.00250527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_257_243#_c_400_n 0.0189173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_465_315#_M1012_g 0.044686f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_31 VNB N_A_465_315#_M1014_g 0.045986f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_32 VNB N_A_465_315#_c_511_n 0.00906762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_287_413#_c_637_n 0.0210888f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_34 VNB N_A_287_413#_c_638_n 0.0018369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_287_413#_c_639_n 0.00624625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_287_413#_c_640_n 0.00187427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_287_413#_c_641_n 0.0292321f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_CLK_c_736_n 0.0202615f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_39 VNB N_CLK_M1015_g 0.0239752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_CLK_M1022_g 0.00619163f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_41 VNB N_CLK_c_739_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_42 VNB N_CLK_c_740_n 0.0291162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_CLK_c_741_n 0.0222729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_CLK_c_742_n 0.0155137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_CLK_c_743_n 0.0285934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_CLK_c_744_n 4.99148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1020_47#_c_816_n 0.0168764f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_48 VNB N_A_1020_47#_c_817_n 0.021509f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_49 VNB N_A_1020_47#_c_818_n 0.00485525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1020_47#_c_819_n 0.00372843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1020_47#_c_820_n 0.00205783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1020_47#_c_821_n 9.59822e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1020_47#_c_822_n 0.0418221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_898_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_27_47#_c_1000_n 0.0141546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_27_47#_c_1001_n 0.00400734f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_57 VNB N_A_27_47#_c_1002_n 0.00595497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_27_47#_c_1003_n 0.0102175f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_59 VNB N_GCLK_c_1052_n 7.54805e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB GCLK 0.0152892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1082_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1083_n 0.00566378f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.53
cc_63 VNB N_VGND_c_1084_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1085_n 0.0100062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1086_n 0.0316357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1087_n 0.0142589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1088_n 0.0434128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1089_n 0.0279198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1090_n 0.0156497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1091_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1092_n 0.00663229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1093_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1094_n 0.0259865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1095_n 0.0143885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1096_n 0.363701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VPB N_SCE_M1011_g 0.0419446f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_77 VPB SCE 0.0188506f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_78 VPB N_SCE_c_142_n 0.0111553f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_79 VPB N_GATE_M1003_g 0.036273f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_80 VPB GATE 0.00670128f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_81 VPB N_GATE_c_168_n 0.00607012f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_82 VPB N_GATE_c_169_n 8.45903e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_257_147#_M1009_g 0.0211245f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_84 VPB N_A_257_147#_c_215_n 0.00360704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_257_147#_c_222_n 0.00578607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_257_147#_c_219_n 0.00647809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_257_147#_c_224_n 0.0169863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_257_147#_c_225_n 0.00400932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_257_147#_c_226_n 0.00220035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_257_147#_c_227_n 0.0266048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_257_147#_c_228_n 0.0457093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_257_243#_M1021_g 0.0505653f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_93 VPB N_A_257_243#_c_389_n 0.0163673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_257_243#_c_390_n 0.00221973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_257_243#_c_393_n 0.00526869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_257_243#_c_405_n 0.00370903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_465_315#_M1018_g 0.022326f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_98 VPB N_A_465_315#_M1012_g 0.0170562f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_99 VPB N_A_465_315#_M1014_g 0.00538896f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_100 VPB N_A_465_315#_M1008_g 0.0229485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_465_315#_c_516_n 0.0033307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_465_315#_c_511_n 0.0039663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_465_315#_c_518_n 0.0151849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_465_315#_c_519_n 0.0052362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_465_315#_c_520_n 0.0310341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_465_315#_c_521_n 0.00438062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_465_315#_c_522_n 0.0296818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_287_413#_M1000_g 0.0243607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_287_413#_c_643_n 0.0134653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_287_413#_c_639_n 0.00269176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_287_413#_c_640_n 0.00386605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_287_413#_c_641_n 0.00831864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_CLK_M1022_g 0.0363646f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_114 VPB N_CLK_c_742_n 0.00856676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_CLK_c_747_n 0.0479145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_CLK_c_744_n 2.37095e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_1020_47#_M1013_g 0.018228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_1020_47#_M1019_g 0.0253024f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_119 VPB N_A_1020_47#_c_820_n 0.00858661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_1020_47#_c_822_n 0.00819567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_899_n 0.0098838f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_122 VPB N_VPWR_c_900_n 0.0318765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_901_n 0.00217586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_902_n 0.00998035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_903_n 0.0449692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_904_n 0.0141605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_905_n 0.0139062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_906_n 0.0340438f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_907_n 0.0135884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_908_n 0.0156552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_909_n 0.0487185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_910_n 0.0137909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_911_n 0.00455555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_912_n 0.00521963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_898_n 0.0446009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_1001_n 0.00313483f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_137 VPB N_GCLK_c_1054_n 0.00109645f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_138 VPB GCLK 0.00449873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 N_SCE_M1011_g N_GATE_M1003_g 0.0495309f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_140 N_SCE_M1023_g N_GATE_M1010_g 0.0256093f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_141 N_SCE_c_142_n GATE 4.13522e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_142 N_SCE_c_142_n N_GATE_c_168_n 0.0495309f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_143 N_SCE_M1023_g N_GATE_c_169_n 4.13522e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_144 N_SCE_M1011_g N_VPWR_c_900_n 0.00472725f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_145 SCE N_VPWR_c_900_n 0.0237825f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_146 N_SCE_c_142_n N_VPWR_c_900_n 0.00105941f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_147 N_SCE_M1011_g N_VPWR_c_909_n 0.00539841f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_148 N_SCE_M1011_g N_VPWR_c_898_n 0.0103231f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_149 N_SCE_M1023_g N_A_27_47#_c_1001_n 0.00890447f $X=0.47 $Y=0.445 $X2=0
+ $Y2=0
cc_150 N_SCE_M1011_g N_A_27_47#_c_1001_n 0.0182361f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_151 SCE N_A_27_47#_c_1001_n 0.0499681f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_152 N_SCE_c_142_n N_A_27_47#_c_1001_n 0.00726295f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_153 N_SCE_M1023_g N_A_27_47#_c_1003_n 0.0159826f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_154 SCE N_A_27_47#_c_1003_n 0.0214425f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_155 N_SCE_c_142_n N_A_27_47#_c_1003_n 0.00349016f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_156 N_SCE_M1011_g N_A_27_47#_c_1012_n 0.0070608f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_157 N_SCE_M1023_g N_VGND_c_1082_n 0.00809304f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_158 N_SCE_M1023_g N_VGND_c_1087_n 0.00337001f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_159 N_SCE_M1023_g N_VGND_c_1096_n 0.00485988f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_160 N_GATE_M1010_g N_A_257_147#_M1005_g 0.0143632f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_161 N_GATE_M1010_g N_A_257_147#_c_211_n 9.82505e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_162 N_GATE_c_168_n N_A_257_147#_c_211_n 0.00116699f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_GATE_c_169_n N_A_257_147#_c_211_n 0.0305181f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_GATE_M1010_g N_A_257_147#_c_212_n 0.0095729f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_165 N_GATE_c_168_n N_A_257_147#_c_212_n 6.18885e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_GATE_c_169_n N_A_257_147#_c_212_n 3.98477e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_167 GATE N_A_257_147#_c_236_n 0.00134565f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_168 N_GATE_c_169_n N_A_257_147#_c_236_n 2.00479e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_GATE_M1003_g N_A_257_147#_c_225_n 4.36779e-19 $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_170 GATE N_A_257_147#_c_225_n 0.0404082f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_171 N_GATE_c_169_n N_A_257_147#_c_225_n 0.00784692f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_172 GATE N_A_257_243#_M1021_g 0.00459698f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_173 N_GATE_M1003_g N_A_257_243#_c_390_n 0.0258836f $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_174 N_GATE_c_168_n N_A_257_243#_c_390_n 0.00719003f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_175 N_GATE_c_169_n N_A_257_243#_c_390_n 0.00194283f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_GATE_M1003_g N_VPWR_c_909_n 0.00357877f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_177 N_GATE_M1003_g N_VPWR_c_898_n 0.00536442f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_178 GATE N_A_27_47#_M1003_d 0.00345627f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_179 N_GATE_M1010_g N_A_27_47#_c_1001_n 0.00390472f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_GATE_c_168_n N_A_27_47#_c_1001_n 0.00960649f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_GATE_c_169_n N_A_27_47#_c_1001_n 0.0754313f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_182 N_GATE_M1010_g N_A_27_47#_c_1002_n 0.0123694f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_183 N_GATE_c_168_n N_A_27_47#_c_1002_n 0.00311345f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_GATE_c_169_n N_A_27_47#_c_1002_n 0.028952f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_185 N_GATE_M1003_g N_A_27_47#_c_1020_n 0.0145681f $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_186 GATE N_A_27_47#_c_1020_n 0.0261201f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_187 N_GATE_M1010_g N_VGND_c_1082_n 0.00763365f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_188 N_GATE_M1010_g N_VGND_c_1088_n 0.00337001f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_189 N_GATE_M1010_g N_VGND_c_1096_n 0.00408452f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_257_147#_M1009_g N_A_257_243#_M1021_g 0.0138034f $X=1.84 $Y=2.275
+ $X2=0 $Y2=0
cc_191 N_A_257_147#_c_225_n N_A_257_243#_M1021_g 0.0149237f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_192 N_A_257_147#_c_227_n N_A_257_243#_M1021_g 0.021304f $X=1.78 $Y=1.74 $X2=0
+ $Y2=0
cc_193 N_A_257_147#_c_218_n N_A_257_243#_c_389_n 0.0105586f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_194 N_A_257_147#_c_224_n N_A_257_243#_c_389_n 0.00213361f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_195 N_A_257_147#_c_225_n N_A_257_243#_c_389_n 0.00868281f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_196 N_A_257_147#_c_227_n N_A_257_243#_c_389_n 0.0180583f $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_197 N_A_257_147#_c_212_n N_A_257_243#_c_390_n 0.0227923f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_198 N_A_257_147#_c_218_n N_A_257_243#_c_390_n 0.0043361f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_199 N_A_257_147#_c_225_n N_A_257_243#_c_390_n 4.45536e-19 $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_200 N_A_257_147#_c_218_n N_A_257_243#_c_391_n 0.00150324f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_201 N_A_257_147#_M1016_g N_A_257_243#_c_392_n 0.00279659f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_202 N_A_257_147#_c_216_n N_A_257_243#_c_392_n 0.00685679f $X=4.71 $Y=0.615
+ $X2=0 $Y2=0
cc_203 N_A_257_147#_M1016_g N_A_257_243#_c_393_n 0.00229895f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_204 N_A_257_147#_c_213_n N_A_257_243#_c_393_n 0.00616579f $X=4.315 $Y=1.105
+ $X2=0 $Y2=0
cc_205 N_A_257_147#_c_214_n N_A_257_243#_c_393_n 0.0131915f $X=4.335 $Y=1.275
+ $X2=0 $Y2=0
cc_206 N_A_257_147#_c_215_n N_A_257_243#_c_393_n 0.00905906f $X=4.335 $Y=1.495
+ $X2=0 $Y2=0
cc_207 N_A_257_147#_c_219_n N_A_257_243#_c_393_n 0.00379592f $X=4.08 $Y=1.19
+ $X2=0 $Y2=0
cc_208 N_A_257_147#_c_224_n N_A_257_243#_c_393_n 0.0104611f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_209 N_A_257_147#_c_226_n N_A_257_243#_c_393_n 2.87747e-19 $X=4.375 $Y=1.53
+ $X2=0 $Y2=0
cc_210 N_A_257_147#_c_228_n N_A_257_243#_c_393_n 0.00364961f $X=4.08 $Y=1.325
+ $X2=0 $Y2=0
cc_211 N_A_257_147#_c_224_n N_A_257_243#_c_405_n 0.00296332f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_212 N_A_257_147#_c_214_n N_A_257_243#_c_432_n 0.00348195f $X=4.335 $Y=1.275
+ $X2=0 $Y2=0
cc_213 N_A_257_147#_c_215_n N_A_257_243#_c_432_n 0.00667477f $X=4.335 $Y=1.495
+ $X2=0 $Y2=0
cc_214 N_A_257_147#_c_219_n N_A_257_243#_c_432_n 0.00199715f $X=4.08 $Y=1.19
+ $X2=0 $Y2=0
cc_215 N_A_257_147#_c_224_n N_A_257_243#_c_432_n 0.00814639f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_216 N_A_257_147#_c_226_n N_A_257_243#_c_432_n 3.27004e-19 $X=4.375 $Y=1.53
+ $X2=0 $Y2=0
cc_217 N_A_257_147#_c_228_n N_A_257_243#_c_432_n 0.00245924f $X=4.08 $Y=1.325
+ $X2=0 $Y2=0
cc_218 N_A_257_147#_c_224_n N_A_257_243#_c_394_n 0.068469f $X=4.23 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_257_147#_c_211_n N_A_257_243#_c_395_n 0.00155066f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_220 N_A_257_147#_c_224_n N_A_257_243#_c_395_n 0.0132091f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_221 N_A_257_147#_M1016_g N_A_257_243#_c_396_n 0.00449775f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_222 N_A_257_147#_c_213_n N_A_257_243#_c_396_n 0.0056501f $X=4.315 $Y=1.105
+ $X2=0 $Y2=0
cc_223 N_A_257_147#_c_214_n N_A_257_243#_c_396_n 0.00254727f $X=4.335 $Y=1.275
+ $X2=0 $Y2=0
cc_224 N_A_257_147#_c_216_n N_A_257_243#_c_396_n 0.00142728f $X=4.71 $Y=0.615
+ $X2=0 $Y2=0
cc_225 N_A_257_147#_c_219_n N_A_257_243#_c_396_n 0.00107245f $X=4.08 $Y=1.19
+ $X2=0 $Y2=0
cc_226 N_A_257_147#_c_224_n N_A_257_243#_c_396_n 0.0151647f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_227 N_A_257_147#_M1016_g N_A_257_243#_c_397_n 0.0055766f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_228 N_A_257_147#_c_213_n N_A_257_243#_c_397_n 0.00974359f $X=4.315 $Y=1.105
+ $X2=0 $Y2=0
cc_229 N_A_257_147#_c_214_n N_A_257_243#_c_397_n 0.00522313f $X=4.335 $Y=1.275
+ $X2=0 $Y2=0
cc_230 N_A_257_147#_c_216_n N_A_257_243#_c_397_n 0.00132323f $X=4.71 $Y=0.615
+ $X2=0 $Y2=0
cc_231 N_A_257_147#_c_219_n N_A_257_243#_c_397_n 0.00134732f $X=4.08 $Y=1.19
+ $X2=0 $Y2=0
cc_232 N_A_257_147#_c_224_n N_A_257_243#_c_397_n 9.74566e-19 $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_233 N_A_257_147#_c_211_n N_A_257_243#_c_398_n 0.00708004f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_234 N_A_257_147#_c_212_n N_A_257_243#_c_398_n 0.0165261f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_235 N_A_257_147#_c_224_n N_A_257_243#_c_398_n 8.52878e-19 $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_236 N_A_257_147#_c_211_n N_A_257_243#_c_399_n 0.0242697f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_237 N_A_257_147#_c_212_n N_A_257_243#_c_399_n 2.60953e-19 $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_238 N_A_257_147#_c_224_n N_A_257_243#_c_399_n 0.00446365f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_239 N_A_257_147#_M1005_g N_A_257_243#_c_400_n 0.0107241f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_240 N_A_257_147#_c_224_n N_A_465_315#_M1000_d 3.75899e-19 $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_241 N_A_257_147#_M1009_g N_A_465_315#_M1018_g 0.0155568f $X=1.84 $Y=2.275
+ $X2=0 $Y2=0
cc_242 N_A_257_147#_c_224_n N_A_465_315#_M1012_g 0.00428067f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_243 N_A_257_147#_c_216_n N_A_465_315#_M1014_g 4.79422e-19 $X=4.71 $Y=0.615
+ $X2=0 $Y2=0
cc_244 N_A_257_147#_c_224_n N_A_465_315#_c_516_n 0.0228159f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_245 N_A_257_147#_M1016_g N_A_465_315#_c_511_n 4.75033e-19 $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_246 N_A_257_147#_c_224_n N_A_465_315#_c_511_n 0.0271467f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_247 N_A_257_147#_c_228_n N_A_465_315#_c_530_n 0.00446021f $X=4.08 $Y=1.325
+ $X2=0 $Y2=0
cc_248 N_A_257_147#_M1007_d N_A_465_315#_c_518_n 0.00483989f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_249 N_A_257_147#_c_214_n N_A_465_315#_c_518_n 0.00128309f $X=4.335 $Y=1.275
+ $X2=0 $Y2=0
cc_250 N_A_257_147#_c_215_n N_A_465_315#_c_518_n 0.0178907f $X=4.335 $Y=1.495
+ $X2=0 $Y2=0
cc_251 N_A_257_147#_c_222_n N_A_465_315#_c_518_n 0.0316717f $X=4.845 $Y=1.66
+ $X2=0 $Y2=0
cc_252 N_A_257_147#_c_224_n N_A_465_315#_c_518_n 0.0132019f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_253 N_A_257_147#_c_226_n N_A_465_315#_c_518_n 0.00170504f $X=4.375 $Y=1.53
+ $X2=0 $Y2=0
cc_254 N_A_257_147#_c_228_n N_A_465_315#_c_518_n 0.0145602f $X=4.08 $Y=1.325
+ $X2=0 $Y2=0
cc_255 N_A_257_147#_c_222_n N_A_465_315#_c_519_n 0.0122409f $X=4.845 $Y=1.66
+ $X2=0 $Y2=0
cc_256 N_A_257_147#_c_224_n N_A_465_315#_c_520_n 0.0039188f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_257 N_A_257_147#_c_227_n N_A_465_315#_c_520_n 0.00753208f $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_258 N_A_257_147#_c_224_n N_A_465_315#_c_541_n 0.00517255f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_259 N_A_257_147#_c_228_n N_A_465_315#_c_542_n 0.00322985f $X=4.08 $Y=1.325
+ $X2=0 $Y2=0
cc_260 N_A_257_147#_c_222_n N_A_465_315#_c_521_n 0.00984522f $X=4.845 $Y=1.66
+ $X2=0 $Y2=0
cc_261 N_A_257_147#_c_222_n N_A_465_315#_c_522_n 5.47076e-19 $X=4.845 $Y=1.66
+ $X2=0 $Y2=0
cc_262 N_A_257_147#_c_224_n N_A_287_413#_M1000_g 0.0075269f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_263 N_A_257_147#_M1005_g N_A_287_413#_c_648_n 0.00581419f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_264 N_A_257_147#_c_211_n N_A_287_413#_c_648_n 0.0249382f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_265 N_A_257_147#_c_212_n N_A_287_413#_c_648_n 9.8177e-19 $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_266 N_A_257_147#_c_218_n N_A_287_413#_c_648_n 0.00398233f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_267 N_A_257_147#_M1009_g N_A_287_413#_c_652_n 0.0131252f $X=1.84 $Y=2.275
+ $X2=0 $Y2=0
cc_268 N_A_257_147#_c_224_n N_A_287_413#_c_652_n 0.00594058f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_269 N_A_257_147#_c_236_n N_A_287_413#_c_652_n 0.00121651f $X=1.76 $Y=1.53
+ $X2=0 $Y2=0
cc_270 N_A_257_147#_c_225_n N_A_287_413#_c_652_n 0.0302261f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_271 N_A_257_147#_c_227_n N_A_287_413#_c_652_n 6.45937e-19 $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_272 N_A_257_147#_c_224_n N_A_287_413#_c_643_n 0.0205826f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_273 N_A_257_147#_c_236_n N_A_287_413#_c_643_n 5.20192e-19 $X=1.76 $Y=1.53
+ $X2=0 $Y2=0
cc_274 N_A_257_147#_c_225_n N_A_287_413#_c_643_n 0.0436285f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_275 N_A_257_147#_c_227_n N_A_287_413#_c_643_n 0.00709868f $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_276 N_A_257_147#_c_211_n N_A_287_413#_c_639_n 0.00602675f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_277 N_A_257_147#_c_218_n N_A_287_413#_c_639_n 0.0146898f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_278 N_A_257_147#_c_224_n N_A_287_413#_c_639_n 0.00783084f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_279 N_A_257_147#_c_224_n N_A_287_413#_c_640_n 0.00746407f $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_280 N_A_257_147#_c_224_n N_A_287_413#_c_641_n 3.55037e-19 $X=4.23 $Y=1.53
+ $X2=0 $Y2=0
cc_281 N_A_257_147#_M1016_g N_CLK_c_736_n 0.00418129f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_282 N_A_257_147#_c_213_n N_CLK_c_736_n 0.00385476f $X=4.315 $Y=1.105 $X2=0
+ $Y2=0
cc_283 N_A_257_147#_c_214_n N_CLK_c_736_n 0.00171427f $X=4.335 $Y=1.275 $X2=0
+ $Y2=0
cc_284 N_A_257_147#_c_219_n N_CLK_c_736_n 0.012847f $X=4.08 $Y=1.19 $X2=0 $Y2=0
cc_285 N_A_257_147#_M1016_g N_CLK_c_739_n 0.019901f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_286 N_A_257_147#_c_216_n N_CLK_c_739_n 0.00707977f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_287 N_A_257_147#_c_213_n N_CLK_c_740_n 0.00700455f $X=4.315 $Y=1.105 $X2=0
+ $Y2=0
cc_288 N_A_257_147#_c_214_n N_CLK_c_740_n 2.58523e-19 $X=4.335 $Y=1.275 $X2=0
+ $Y2=0
cc_289 N_A_257_147#_c_222_n N_CLK_c_740_n 9.73222e-19 $X=4.845 $Y=1.66 $X2=0
+ $Y2=0
cc_290 N_A_257_147#_c_216_n N_CLK_c_740_n 0.0200908f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_291 N_A_257_147#_c_217_n N_CLK_c_740_n 0.00136651f $X=4.68 $Y=0.465 $X2=0
+ $Y2=0
cc_292 N_A_257_147#_c_226_n N_CLK_c_740_n 0.00109922f $X=4.375 $Y=1.53 $X2=0
+ $Y2=0
cc_293 N_A_257_147#_c_222_n N_CLK_c_741_n 0.00555242f $X=4.845 $Y=1.66 $X2=0
+ $Y2=0
cc_294 N_A_257_147#_c_215_n N_CLK_c_742_n 4.8674e-19 $X=4.335 $Y=1.495 $X2=0
+ $Y2=0
cc_295 N_A_257_147#_c_222_n N_CLK_c_742_n 0.00777662f $X=4.845 $Y=1.66 $X2=0
+ $Y2=0
cc_296 N_A_257_147#_c_226_n N_CLK_c_742_n 4.65417e-19 $X=4.375 $Y=1.53 $X2=0
+ $Y2=0
cc_297 N_A_257_147#_c_215_n N_CLK_c_747_n 0.00400264f $X=4.335 $Y=1.495 $X2=0
+ $Y2=0
cc_298 N_A_257_147#_c_222_n N_CLK_c_747_n 0.016003f $X=4.845 $Y=1.66 $X2=0 $Y2=0
cc_299 N_A_257_147#_c_226_n N_CLK_c_747_n 0.00159708f $X=4.375 $Y=1.53 $X2=0
+ $Y2=0
cc_300 N_A_257_147#_c_228_n N_CLK_c_747_n 0.0376094f $X=4.08 $Y=1.325 $X2=0
+ $Y2=0
cc_301 N_A_257_147#_c_213_n N_CLK_c_744_n 0.00940108f $X=4.315 $Y=1.105 $X2=0
+ $Y2=0
cc_302 N_A_257_147#_c_214_n N_CLK_c_744_n 0.0110934f $X=4.335 $Y=1.275 $X2=0
+ $Y2=0
cc_303 N_A_257_147#_c_215_n N_CLK_c_744_n 0.00281426f $X=4.335 $Y=1.495 $X2=0
+ $Y2=0
cc_304 N_A_257_147#_c_222_n N_CLK_c_744_n 0.0171599f $X=4.845 $Y=1.66 $X2=0
+ $Y2=0
cc_305 N_A_257_147#_c_216_n N_CLK_c_744_n 0.00864905f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_306 N_A_257_147#_c_217_n N_A_1020_47#_c_827_n 0.0196051f $X=4.68 $Y=0.465
+ $X2=0 $Y2=0
cc_307 N_A_257_147#_c_216_n N_A_1020_47#_c_819_n 0.0108704f $X=4.71 $Y=0.615
+ $X2=0 $Y2=0
cc_308 N_A_257_147#_c_224_n N_VPWR_M1018_d 0.0020643f $X=4.23 $Y=1.53 $X2=0
+ $Y2=0
cc_309 N_A_257_147#_c_215_n N_VPWR_M1001_d 0.00463165f $X=4.335 $Y=1.495 $X2=0
+ $Y2=0
cc_310 N_A_257_147#_c_222_n N_VPWR_M1001_d 4.52908e-19 $X=4.845 $Y=1.66 $X2=0
+ $Y2=0
cc_311 N_A_257_147#_c_224_n N_VPWR_M1001_d 4.60476e-19 $X=4.23 $Y=1.53 $X2=0
+ $Y2=0
cc_312 N_A_257_147#_c_228_n N_VPWR_c_906_n 0.0233072f $X=4.08 $Y=1.325 $X2=0
+ $Y2=0
cc_313 N_A_257_147#_M1009_g N_VPWR_c_909_n 0.00357877f $X=1.84 $Y=2.275 $X2=0
+ $Y2=0
cc_314 N_A_257_147#_M1009_g N_VPWR_c_910_n 0.00145256f $X=1.84 $Y=2.275 $X2=0
+ $Y2=0
cc_315 N_A_257_147#_c_224_n N_VPWR_c_910_n 7.31718e-19 $X=4.23 $Y=1.53 $X2=0
+ $Y2=0
cc_316 N_A_257_147#_M1009_g N_VPWR_c_898_n 0.00579685f $X=1.84 $Y=2.275 $X2=0
+ $Y2=0
cc_317 N_A_257_147#_c_225_n N_VPWR_c_898_n 0.00150144f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_318 N_A_257_147#_M1005_g N_A_27_47#_c_1002_n 0.0029712f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_319 N_A_257_147#_c_211_n N_A_27_47#_c_1002_n 0.0067219f $X=1.45 $Y=0.87 $X2=0
+ $Y2=0
cc_320 N_A_257_147#_c_212_n N_A_27_47#_c_1002_n 4.43441e-19 $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_321 N_A_257_147#_M1005_g N_A_27_47#_c_1025_n 0.00382934f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_322 N_A_257_147#_c_216_n N_VGND_M1016_d 0.00164398f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_323 N_A_257_147#_M1005_g N_VGND_c_1082_n 0.00109585f $X=1.375 $Y=0.415 $X2=0
+ $Y2=0
cc_324 N_A_257_147#_M1016_g N_VGND_c_1084_n 0.00853729f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_325 N_A_257_147#_c_214_n N_VGND_c_1084_n 0.00117442f $X=4.335 $Y=1.275 $X2=0
+ $Y2=0
cc_326 N_A_257_147#_c_216_n N_VGND_c_1084_n 0.013843f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_327 N_A_257_147#_M1005_g N_VGND_c_1088_n 0.00456464f $X=1.375 $Y=0.415 $X2=0
+ $Y2=0
cc_328 N_A_257_147#_c_212_n N_VGND_c_1088_n 2.64403e-19 $X=1.45 $Y=0.87 $X2=0
+ $Y2=0
cc_329 N_A_257_147#_M1016_g N_VGND_c_1089_n 0.0046653f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_330 N_A_257_147#_c_216_n N_VGND_c_1094_n 0.00258611f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_331 N_A_257_147#_c_217_n N_VGND_c_1094_n 0.0151508f $X=4.68 $Y=0.465 $X2=0
+ $Y2=0
cc_332 N_A_257_147#_M1020_d N_VGND_c_1096_n 0.00227267f $X=4.545 $Y=0.235 $X2=0
+ $Y2=0
cc_333 N_A_257_147#_M1005_g N_VGND_c_1096_n 0.00806939f $X=1.375 $Y=0.415 $X2=0
+ $Y2=0
cc_334 N_A_257_147#_M1016_g N_VGND_c_1096_n 0.00669841f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_335 N_A_257_147#_c_212_n N_VGND_c_1096_n 3.49206e-19 $X=1.45 $Y=0.87 $X2=0
+ $Y2=0
cc_336 N_A_257_147#_c_216_n N_VGND_c_1096_n 0.00553659f $X=4.71 $Y=0.615 $X2=0
+ $Y2=0
cc_337 N_A_257_147#_c_217_n N_VGND_c_1096_n 0.00864204f $X=4.68 $Y=0.465 $X2=0
+ $Y2=0
cc_338 N_A_257_243#_c_394_n N_A_465_315#_M1006_d 5.81953e-19 $X=3.77 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_339 N_A_257_243#_c_391_n N_A_465_315#_M1012_g 0.00692236f $X=1.9 $Y=1.215
+ $X2=0 $Y2=0
cc_340 N_A_257_243#_c_394_n N_A_465_315#_M1012_g 0.00342271f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_341 N_A_257_243#_c_398_n N_A_465_315#_M1012_g 0.0115616f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_342 N_A_257_243#_c_399_n N_A_465_315#_M1012_g 7.79891e-19 $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_343 N_A_257_243#_c_400_n N_A_465_315#_M1012_g 0.0139526f $X=1.96 $Y=0.705
+ $X2=0 $Y2=0
cc_344 N_A_257_243#_c_392_n N_A_465_315#_c_511_n 0.100963f $X=3.84 $Y=0.465
+ $X2=0 $Y2=0
cc_345 N_A_257_243#_c_405_n N_A_465_315#_c_511_n 0.00461785f $X=3.745 $Y=1.66
+ $X2=0 $Y2=0
cc_346 N_A_257_243#_c_394_n N_A_465_315#_c_511_n 0.0208446f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_347 N_A_257_243#_c_396_n N_A_465_315#_c_511_n 2.9182e-19 $X=3.915 $Y=0.85
+ $X2=0 $Y2=0
cc_348 N_A_257_243#_M1001_s N_A_465_315#_c_518_n 0.00483614f $X=3.75 $Y=1.515
+ $X2=0 $Y2=0
cc_349 N_A_257_243#_c_405_n N_A_465_315#_c_518_n 0.0134309f $X=3.745 $Y=1.66
+ $X2=0 $Y2=0
cc_350 N_A_257_243#_c_432_n N_A_465_315#_c_518_n 0.0159566f $X=3.875 $Y=1.66
+ $X2=0 $Y2=0
cc_351 N_A_257_243#_c_405_n N_A_465_315#_c_542_n 0.00982836f $X=3.745 $Y=1.66
+ $X2=0 $Y2=0
cc_352 N_A_257_243#_c_394_n N_A_287_413#_c_637_n 0.00847687f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_353 N_A_257_243#_c_405_n N_A_287_413#_M1000_g 5.08874e-19 $X=3.745 $Y=1.66
+ $X2=0 $Y2=0
cc_354 N_A_257_243#_c_389_n N_A_287_413#_c_648_n 7.07243e-19 $X=1.825 $Y=1.29
+ $X2=0 $Y2=0
cc_355 N_A_257_243#_c_394_n N_A_287_413#_c_648_n 0.00173863f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_356 N_A_257_243#_c_395_n N_A_287_413#_c_648_n 0.0020338f $X=2.22 $Y=0.85
+ $X2=0 $Y2=0
cc_357 N_A_257_243#_c_398_n N_A_287_413#_c_648_n 0.00258224f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_358 N_A_257_243#_c_399_n N_A_287_413#_c_648_n 0.0175669f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_359 N_A_257_243#_c_400_n N_A_287_413#_c_648_n 0.0128508f $X=1.96 $Y=0.705
+ $X2=0 $Y2=0
cc_360 N_A_257_243#_M1021_g N_A_287_413#_c_652_n 0.00300964f $X=1.36 $Y=2.275
+ $X2=0 $Y2=0
cc_361 N_A_257_243#_M1021_g N_A_287_413#_c_643_n 6.3244e-19 $X=1.36 $Y=2.275
+ $X2=0 $Y2=0
cc_362 N_A_257_243#_c_394_n N_A_287_413#_c_638_n 0.0162752f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_363 N_A_257_243#_c_395_n N_A_287_413#_c_638_n 0.00275249f $X=2.22 $Y=0.85
+ $X2=0 $Y2=0
cc_364 N_A_257_243#_c_398_n N_A_287_413#_c_638_n 7.44567e-19 $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_365 N_A_257_243#_c_399_n N_A_287_413#_c_638_n 0.0205672f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_366 N_A_257_243#_c_400_n N_A_287_413#_c_638_n 0.00302624f $X=1.96 $Y=0.705
+ $X2=0 $Y2=0
cc_367 N_A_257_243#_c_391_n N_A_287_413#_c_639_n 0.00377955f $X=1.9 $Y=1.215
+ $X2=0 $Y2=0
cc_368 N_A_257_243#_c_394_n N_A_287_413#_c_639_n 0.00154998f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_369 N_A_257_243#_c_395_n N_A_287_413#_c_639_n 0.00160742f $X=2.22 $Y=0.85
+ $X2=0 $Y2=0
cc_370 N_A_257_243#_c_398_n N_A_287_413#_c_639_n 0.00153556f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_371 N_A_257_243#_c_399_n N_A_287_413#_c_639_n 0.0128543f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_372 N_A_257_243#_c_394_n N_A_287_413#_c_640_n 0.0106635f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_373 N_A_257_243#_c_394_n N_A_287_413#_c_641_n 0.0044627f $X=3.77 $Y=0.85
+ $X2=0 $Y2=0
cc_374 N_A_257_243#_M1021_g N_VPWR_c_909_n 0.00577801f $X=1.36 $Y=2.275 $X2=0
+ $Y2=0
cc_375 N_A_257_243#_M1021_g N_VPWR_c_898_n 0.0103326f $X=1.36 $Y=2.275 $X2=0
+ $Y2=0
cc_376 N_A_257_243#_c_394_n N_VGND_M1012_d 4.25819e-19 $X=3.77 $Y=0.85 $X2=0
+ $Y2=0
cc_377 N_A_257_243#_c_394_n N_VGND_c_1083_n 0.0140576f $X=3.77 $Y=0.85 $X2=0
+ $Y2=0
cc_378 N_A_257_243#_c_400_n N_VGND_c_1088_n 0.00357877f $X=1.96 $Y=0.705 $X2=0
+ $Y2=0
cc_379 N_A_257_243#_c_392_n N_VGND_c_1089_n 0.0244536f $X=3.84 $Y=0.465 $X2=0
+ $Y2=0
cc_380 N_A_257_243#_M1016_s N_VGND_c_1096_n 0.00182676f $X=3.715 $Y=0.235 $X2=0
+ $Y2=0
cc_381 N_A_257_243#_c_392_n N_VGND_c_1096_n 0.00625164f $X=3.84 $Y=0.465 $X2=0
+ $Y2=0
cc_382 N_A_257_243#_c_394_n N_VGND_c_1096_n 0.0724491f $X=3.77 $Y=0.85 $X2=0
+ $Y2=0
cc_383 N_A_257_243#_c_395_n N_VGND_c_1096_n 0.014828f $X=2.22 $Y=0.85 $X2=0
+ $Y2=0
cc_384 N_A_257_243#_c_396_n N_VGND_c_1096_n 0.0152609f $X=3.915 $Y=0.85 $X2=0
+ $Y2=0
cc_385 N_A_257_243#_c_397_n N_VGND_c_1096_n 6.43573e-19 $X=3.915 $Y=0.85 $X2=0
+ $Y2=0
cc_386 N_A_257_243#_c_400_n N_VGND_c_1096_n 0.00589934f $X=1.96 $Y=0.705 $X2=0
+ $Y2=0
cc_387 N_A_465_315#_M1012_g N_A_287_413#_c_637_n 0.0188679f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_388 N_A_465_315#_c_511_n N_A_287_413#_c_637_n 0.0293052f $X=3.32 $Y=0.42
+ $X2=0 $Y2=0
cc_389 N_A_465_315#_M1018_g N_A_287_413#_M1000_g 0.0129074f $X=2.43 $Y=2.275
+ $X2=0 $Y2=0
cc_390 N_A_465_315#_M1012_g N_A_287_413#_M1000_g 0.00670688f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_391 N_A_465_315#_c_516_n N_A_287_413#_M1000_g 0.014093f $X=3.185 $Y=1.77
+ $X2=0 $Y2=0
cc_392 N_A_465_315#_c_520_n N_A_287_413#_M1000_g 0.00808806f $X=2.46 $Y=1.74
+ $X2=0 $Y2=0
cc_393 N_A_465_315#_c_541_n N_A_287_413#_M1000_g 2.06052e-19 $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_394 N_A_465_315#_c_542_n N_A_287_413#_M1000_g 0.00982347f $X=3.295 $Y=1.86
+ $X2=0 $Y2=0
cc_395 N_A_465_315#_M1012_g N_A_287_413#_c_648_n 0.00893118f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_396 N_A_465_315#_M1018_g N_A_287_413#_c_652_n 0.00282173f $X=2.43 $Y=2.275
+ $X2=0 $Y2=0
cc_397 N_A_465_315#_M1018_g N_A_287_413#_c_643_n 0.00426352f $X=2.43 $Y=2.275
+ $X2=0 $Y2=0
cc_398 N_A_465_315#_M1012_g N_A_287_413#_c_643_n 0.00550388f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_399 N_A_465_315#_c_520_n N_A_287_413#_c_643_n 0.00271662f $X=2.46 $Y=1.74
+ $X2=0 $Y2=0
cc_400 N_A_465_315#_c_541_n N_A_287_413#_c_643_n 0.0255746f $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_401 N_A_465_315#_M1012_g N_A_287_413#_c_638_n 0.0114396f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_465_315#_M1012_g N_A_287_413#_c_639_n 0.00791638f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_465_315#_c_520_n N_A_287_413#_c_639_n 0.00300149f $X=2.46 $Y=1.74
+ $X2=0 $Y2=0
cc_404 N_A_465_315#_c_541_n N_A_287_413#_c_639_n 0.00700208f $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_405 N_A_465_315#_M1012_g N_A_287_413#_c_640_n 0.00928658f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_406 N_A_465_315#_c_516_n N_A_287_413#_c_640_n 0.0171291f $X=3.185 $Y=1.77
+ $X2=0 $Y2=0
cc_407 N_A_465_315#_c_511_n N_A_287_413#_c_640_n 0.0310043f $X=3.32 $Y=0.42
+ $X2=0 $Y2=0
cc_408 N_A_465_315#_c_541_n N_A_287_413#_c_640_n 0.00230595f $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_409 N_A_465_315#_M1012_g N_A_287_413#_c_641_n 0.0213485f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_465_315#_c_516_n N_A_287_413#_c_641_n 0.00123339f $X=3.185 $Y=1.77
+ $X2=0 $Y2=0
cc_411 N_A_465_315#_M1014_g N_CLK_M1015_g 0.0696057f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_A_465_315#_M1014_g N_CLK_M1022_g 0.00642463f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_465_315#_c_522_n N_CLK_M1022_g 0.0375236f $X=5.575 $Y=1.52 $X2=0
+ $Y2=0
cc_414 N_A_465_315#_M1014_g N_CLK_c_740_n 0.0166168f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_465_315#_M1014_g N_CLK_c_741_n 0.01681f $X=5.435 $Y=0.445 $X2=0 $Y2=0
cc_416 N_A_465_315#_c_518_n N_CLK_c_741_n 0.00524792f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_417 N_A_465_315#_c_521_n N_CLK_c_741_n 0.0352231f $X=5.485 $Y=1.52 $X2=0
+ $Y2=0
cc_418 N_A_465_315#_c_522_n N_CLK_c_741_n 0.00488951f $X=5.575 $Y=1.52 $X2=0
+ $Y2=0
cc_419 N_A_465_315#_M1014_g N_CLK_c_747_n 0.00137667f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_420 N_A_465_315#_c_518_n N_CLK_c_747_n 0.0130735f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_421 N_A_465_315#_c_519_n N_CLK_c_747_n 0.00320853f $X=5.335 $Y=1.915 $X2=0
+ $Y2=0
cc_422 N_A_465_315#_c_521_n N_CLK_c_747_n 0.00137462f $X=5.485 $Y=1.52 $X2=0
+ $Y2=0
cc_423 N_A_465_315#_c_522_n N_CLK_c_747_n 0.00332804f $X=5.575 $Y=1.52 $X2=0
+ $Y2=0
cc_424 N_A_465_315#_M1014_g N_CLK_c_744_n 3.32747e-19 $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_425 N_A_465_315#_M1014_g N_A_1020_47#_c_818_n 0.0112069f $X=5.435 $Y=0.445
+ $X2=0 $Y2=0
cc_426 N_A_465_315#_M1008_g N_A_1020_47#_c_820_n 9.63993e-19 $X=5.575 $Y=2.165
+ $X2=0 $Y2=0
cc_427 N_A_465_315#_c_519_n N_A_1020_47#_c_820_n 0.0143305f $X=5.335 $Y=1.915
+ $X2=0 $Y2=0
cc_428 N_A_465_315#_c_521_n N_A_1020_47#_c_820_n 0.0144034f $X=5.485 $Y=1.52
+ $X2=0 $Y2=0
cc_429 N_A_465_315#_c_522_n N_A_1020_47#_c_820_n 0.002146f $X=5.575 $Y=1.52
+ $X2=0 $Y2=0
cc_430 N_A_465_315#_c_516_n N_VPWR_M1018_d 0.00488989f $X=3.185 $Y=1.77 $X2=0
+ $Y2=0
cc_431 N_A_465_315#_c_518_n N_VPWR_M1001_d 0.00612262f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_432 N_A_465_315#_c_518_n N_VPWR_M1008_s 0.00399258f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_433 N_A_465_315#_c_519_n N_VPWR_M1008_s 7.75292e-19 $X=5.335 $Y=1.915 $X2=0
+ $Y2=0
cc_434 N_A_465_315#_c_530_n N_VPWR_c_904_n 0.0176738f $X=3.32 $Y=2.205 $X2=0
+ $Y2=0
cc_435 N_A_465_315#_c_518_n N_VPWR_c_904_n 0.114438f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_436 N_A_465_315#_c_530_n N_VPWR_c_905_n 0.0133789f $X=3.32 $Y=2.205 $X2=0
+ $Y2=0
cc_437 N_A_465_315#_c_518_n N_VPWR_c_905_n 0.00215449f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_438 N_A_465_315#_c_518_n N_VPWR_c_906_n 0.0216591f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_439 N_A_465_315#_M1008_g N_VPWR_c_907_n 0.0046653f $X=5.575 $Y=2.165 $X2=0
+ $Y2=0
cc_440 N_A_465_315#_M1018_g N_VPWR_c_909_n 7.6274e-19 $X=2.43 $Y=2.275 $X2=0
+ $Y2=0
cc_441 N_A_465_315#_M1018_g N_VPWR_c_910_n 0.0247949f $X=2.43 $Y=2.275 $X2=0
+ $Y2=0
cc_442 N_A_465_315#_c_520_n N_VPWR_c_910_n 0.0022365f $X=2.46 $Y=1.74 $X2=0
+ $Y2=0
cc_443 N_A_465_315#_c_541_n N_VPWR_c_910_n 0.044273f $X=2.545 $Y=1.74 $X2=0
+ $Y2=0
cc_444 N_A_465_315#_M1008_g N_VPWR_c_911_n 0.00882421f $X=5.575 $Y=2.165 $X2=0
+ $Y2=0
cc_445 N_A_465_315#_c_521_n N_VPWR_c_911_n 8.53981e-19 $X=5.485 $Y=1.52 $X2=0
+ $Y2=0
cc_446 N_A_465_315#_c_522_n N_VPWR_c_911_n 4.82886e-19 $X=5.575 $Y=1.52 $X2=0
+ $Y2=0
cc_447 N_A_465_315#_M1000_d N_VPWR_c_898_n 0.00223109f $X=3.185 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_A_465_315#_M1018_g N_VPWR_c_898_n 0.002381f $X=2.43 $Y=2.275 $X2=0
+ $Y2=0
cc_449 N_A_465_315#_M1008_g N_VPWR_c_898_n 0.00794739f $X=5.575 $Y=2.165 $X2=0
+ $Y2=0
cc_450 N_A_465_315#_c_516_n N_VPWR_c_898_n 0.00508158f $X=3.185 $Y=1.77 $X2=0
+ $Y2=0
cc_451 N_A_465_315#_c_530_n N_VPWR_c_898_n 0.00839556f $X=3.32 $Y=2.205 $X2=0
+ $Y2=0
cc_452 N_A_465_315#_c_518_n N_VPWR_c_898_n 0.0139993f $X=5.18 $Y=2 $X2=0 $Y2=0
cc_453 N_A_465_315#_c_520_n N_VPWR_c_898_n 6.86139e-19 $X=2.46 $Y=1.74 $X2=0
+ $Y2=0
cc_454 N_A_465_315#_c_541_n N_VPWR_c_898_n 0.00214472f $X=2.545 $Y=1.74 $X2=0
+ $Y2=0
cc_455 N_A_465_315#_M1012_g N_VGND_c_1083_n 0.00849127f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_456 N_A_465_315#_c_511_n N_VGND_c_1083_n 0.0156967f $X=3.32 $Y=0.42 $X2=0
+ $Y2=0
cc_457 N_A_465_315#_M1012_g N_VGND_c_1088_n 0.00486707f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_465_315#_c_511_n N_VGND_c_1089_n 0.0133789f $X=3.32 $Y=0.42 $X2=0
+ $Y2=0
cc_459 N_A_465_315#_M1014_g N_VGND_c_1094_n 0.00365142f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_465_315#_M1014_g N_VGND_c_1095_n 0.00928177f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_461 N_A_465_315#_M1006_d N_VGND_c_1096_n 0.00204319f $X=3.185 $Y=0.235 $X2=0
+ $Y2=0
cc_462 N_A_465_315#_M1012_g N_VGND_c_1096_n 0.00673447f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_463 N_A_465_315#_M1014_g N_VGND_c_1096_n 0.00559219f $X=5.435 $Y=0.445 $X2=0
+ $Y2=0
cc_464 N_A_465_315#_c_511_n N_VGND_c_1096_n 0.00399922f $X=3.32 $Y=0.42 $X2=0
+ $Y2=0
cc_465 N_A_287_413#_M1000_g N_VPWR_c_904_n 0.00239902f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_466 N_A_287_413#_M1000_g N_VPWR_c_905_n 0.00468308f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_467 N_A_287_413#_c_652_n N_VPWR_c_909_n 0.0463617f $X=2.035 $Y=2.295 $X2=0
+ $Y2=0
cc_468 N_A_287_413#_M1000_g N_VPWR_c_910_n 0.00514863f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_A_287_413#_c_652_n N_VPWR_c_910_n 0.0295853f $X=2.035 $Y=2.295 $X2=0
+ $Y2=0
cc_470 N_A_287_413#_c_643_n N_VPWR_c_910_n 0.00379592f $X=2.12 $Y=2.125 $X2=0
+ $Y2=0
cc_471 N_A_287_413#_M1021_d N_VPWR_c_898_n 0.00263412f $X=1.435 $Y=2.065 $X2=0
+ $Y2=0
cc_472 N_A_287_413#_M1000_g N_VPWR_c_898_n 0.00805978f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_287_413#_c_652_n N_VPWR_c_898_n 0.0285676f $X=2.035 $Y=2.295 $X2=0
+ $Y2=0
cc_474 N_A_287_413#_c_648_n N_A_27_47#_c_1025_n 0.0219377f $X=2.33 $Y=0.395
+ $X2=0 $Y2=0
cc_475 N_A_287_413#_c_652_n A_383_413# 0.00832946f $X=2.035 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_476 N_A_287_413#_c_643_n A_383_413# 0.00151526f $X=2.12 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_477 N_A_287_413#_c_637_n N_VGND_c_1083_n 0.00734556f $X=3.11 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_287_413#_c_648_n N_VGND_c_1083_n 0.0231479f $X=2.33 $Y=0.395 $X2=0
+ $Y2=0
cc_479 N_A_287_413#_c_638_n N_VGND_c_1083_n 0.0210362f $X=2.415 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_287_413#_c_640_n N_VGND_c_1083_n 0.022345f $X=2.93 $Y=1.16 $X2=0
+ $Y2=0
cc_481 N_A_287_413#_c_641_n N_VGND_c_1083_n 0.00484825f $X=3.11 $Y=1.16 $X2=0
+ $Y2=0
cc_482 N_A_287_413#_c_648_n N_VGND_c_1088_n 0.0673769f $X=2.33 $Y=0.395 $X2=0
+ $Y2=0
cc_483 N_A_287_413#_c_637_n N_VGND_c_1089_n 0.00585385f $X=3.11 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_A_287_413#_M1005_d N_VGND_c_1096_n 0.00299551f $X=1.45 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_287_413#_c_637_n N_VGND_c_1096_n 0.00794139f $X=3.11 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_A_287_413#_c_648_n N_VGND_c_1096_n 0.0299006f $X=2.33 $Y=0.395 $X2=0
+ $Y2=0
cc_487 N_A_287_413#_c_648_n A_395_47# 0.00874765f $X=2.33 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_488 N_A_287_413#_c_638_n A_395_47# 0.00160798f $X=2.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_489 N_CLK_M1015_g N_A_1020_47#_c_816_n 0.0160282f $X=5.795 $Y=0.445 $X2=0
+ $Y2=0
cc_490 N_CLK_c_743_n N_A_1020_47#_c_816_n 0.00278662f $X=5.995 $Y=1.05 $X2=0
+ $Y2=0
cc_491 N_CLK_M1022_g N_A_1020_47#_M1013_g 0.035715f $X=5.995 $Y=2.165 $X2=0
+ $Y2=0
cc_492 N_CLK_M1015_g N_A_1020_47#_c_818_n 0.0109898f $X=5.795 $Y=0.445 $X2=0
+ $Y2=0
cc_493 N_CLK_c_741_n N_A_1020_47#_c_818_n 0.0552543f $X=5.885 $Y=1.05 $X2=0
+ $Y2=0
cc_494 N_CLK_c_743_n N_A_1020_47#_c_818_n 0.00537215f $X=5.995 $Y=1.05 $X2=0
+ $Y2=0
cc_495 N_CLK_c_739_n N_A_1020_47#_c_819_n 4.25479e-19 $X=4.66 $Y=0.73 $X2=0
+ $Y2=0
cc_496 N_CLK_c_740_n N_A_1020_47#_c_819_n 6.3229e-19 $X=4.66 $Y=0.88 $X2=0 $Y2=0
cc_497 N_CLK_c_741_n N_A_1020_47#_c_819_n 0.0181374f $X=5.885 $Y=1.05 $X2=0
+ $Y2=0
cc_498 N_CLK_M1022_g N_A_1020_47#_c_820_n 0.0268601f $X=5.995 $Y=2.165 $X2=0
+ $Y2=0
cc_499 N_CLK_c_741_n N_A_1020_47#_c_820_n 0.045368f $X=5.885 $Y=1.05 $X2=0 $Y2=0
cc_500 N_CLK_c_743_n N_A_1020_47#_c_820_n 0.00644546f $X=5.995 $Y=1.05 $X2=0
+ $Y2=0
cc_501 N_CLK_M1015_g N_A_1020_47#_c_821_n 0.00235168f $X=5.795 $Y=0.445 $X2=0
+ $Y2=0
cc_502 N_CLK_c_741_n N_A_1020_47#_c_821_n 0.00294772f $X=5.885 $Y=1.05 $X2=0
+ $Y2=0
cc_503 N_CLK_c_743_n N_A_1020_47#_c_821_n 0.001185f $X=5.995 $Y=1.05 $X2=0 $Y2=0
cc_504 N_CLK_c_741_n N_A_1020_47#_c_822_n 2.88786e-19 $X=5.885 $Y=1.05 $X2=0
+ $Y2=0
cc_505 N_CLK_c_743_n N_A_1020_47#_c_822_n 0.0202296f $X=5.995 $Y=1.05 $X2=0
+ $Y2=0
cc_506 N_CLK_M1022_g N_VPWR_c_901_n 0.00166155f $X=5.995 $Y=2.165 $X2=0 $Y2=0
cc_507 N_CLK_c_747_n N_VPWR_c_906_n 0.024098f $X=4.715 $Y=1.325 $X2=0 $Y2=0
cc_508 N_CLK_M1022_g N_VPWR_c_907_n 0.00424239f $X=5.995 $Y=2.165 $X2=0 $Y2=0
cc_509 N_CLK_M1022_g N_VPWR_c_911_n 5.79077e-19 $X=5.995 $Y=2.165 $X2=0 $Y2=0
cc_510 N_CLK_M1022_g N_VPWR_c_898_n 0.00576116f $X=5.995 $Y=2.165 $X2=0 $Y2=0
cc_511 N_CLK_c_739_n N_VGND_c_1084_n 0.00809304f $X=4.66 $Y=0.73 $X2=0 $Y2=0
cc_512 N_CLK_c_739_n N_VGND_c_1094_n 0.00337001f $X=4.66 $Y=0.73 $X2=0 $Y2=0
cc_513 N_CLK_c_740_n N_VGND_c_1094_n 0.00229357f $X=4.66 $Y=0.88 $X2=0 $Y2=0
cc_514 N_CLK_M1015_g N_VGND_c_1095_n 0.0188261f $X=5.795 $Y=0.445 $X2=0 $Y2=0
cc_515 N_CLK_c_739_n N_VGND_c_1096_n 0.0053254f $X=4.66 $Y=0.73 $X2=0 $Y2=0
cc_516 N_CLK_c_740_n N_VGND_c_1096_n 0.00262886f $X=4.66 $Y=0.88 $X2=0 $Y2=0
cc_517 N_A_1020_47#_c_820_n N_VPWR_M1022_d 0.00224468f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_518 N_A_1020_47#_M1013_g N_VPWR_c_901_n 0.00533931f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_519 N_A_1020_47#_M1019_g N_VPWR_c_901_n 6.03273e-19 $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_520 N_A_1020_47#_c_820_n N_VPWR_c_901_n 0.0180293f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_521 N_A_1020_47#_M1019_g N_VPWR_c_903_n 0.0031814f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_522 N_A_1020_47#_c_820_n N_VPWR_c_907_n 0.0145632f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_523 N_A_1020_47#_M1013_g N_VPWR_c_908_n 0.00564095f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_524 N_A_1020_47#_M1019_g N_VPWR_c_908_n 0.0054895f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_525 N_A_1020_47#_M1008_d N_VPWR_c_898_n 0.00411223f $X=5.65 $Y=1.845 $X2=0
+ $Y2=0
cc_526 N_A_1020_47#_M1013_g N_VPWR_c_898_n 0.00950335f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_527 N_A_1020_47#_M1019_g N_VPWR_c_898_n 0.010667f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_528 N_A_1020_47#_c_820_n N_VPWR_c_898_n 0.013348f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_529 N_A_1020_47#_c_816_n N_GCLK_c_1052_n 0.00121413f $X=6.47 $Y=0.995 $X2=0
+ $Y2=0
cc_530 N_A_1020_47#_c_817_n N_GCLK_c_1052_n 0.00621583f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_1020_47#_c_820_n N_GCLK_c_1052_n 0.00420505f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_532 N_A_1020_47#_c_821_n N_GCLK_c_1052_n 0.00847884f $X=6.315 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_A_1020_47#_c_822_n N_GCLK_c_1052_n 0.00528944f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_534 N_A_1020_47#_c_817_n N_GCLK_c_1061_n 0.00269264f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_535 N_A_1020_47#_c_822_n N_GCLK_c_1061_n 0.00103776f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_536 N_A_1020_47#_M1019_g N_GCLK_c_1063_n 0.00259971f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_537 N_A_1020_47#_c_822_n N_GCLK_c_1063_n 0.00105578f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_538 N_A_1020_47#_M1013_g N_GCLK_c_1054_n 0.00121211f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_539 N_A_1020_47#_M1019_g N_GCLK_c_1054_n 0.00769664f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_540 N_A_1020_47#_c_820_n N_GCLK_c_1054_n 0.00954314f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_541 N_A_1020_47#_c_822_n N_GCLK_c_1054_n 0.00193313f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_542 N_A_1020_47#_c_820_n N_GCLK_c_1069_n 0.0203737f $X=5.785 $Y=2.085 $X2=0
+ $Y2=0
cc_543 N_A_1020_47#_c_822_n N_GCLK_c_1069_n 0.00775129f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_544 N_A_1020_47#_M1019_g GCLK 0.0101586f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_545 N_A_1020_47#_c_822_n GCLK 0.0197662f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_546 N_A_1020_47#_c_817_n N_GCLK_c_1073_n 0.00550796f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_547 N_A_1020_47#_c_818_n N_VGND_M1015_d 0.006707f $X=6.23 $Y=0.7 $X2=0 $Y2=0
cc_548 N_A_1020_47#_c_821_n N_VGND_M1015_d 0.00134384f $X=6.315 $Y=0.995 $X2=0
+ $Y2=0
cc_549 N_A_1020_47#_c_817_n N_VGND_c_1086_n 0.00318017f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_550 N_A_1020_47#_c_816_n N_VGND_c_1090_n 0.00564095f $X=6.47 $Y=0.995 $X2=0
+ $Y2=0
cc_551 N_A_1020_47#_c_817_n N_VGND_c_1090_n 0.0054895f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_552 N_A_1020_47#_c_827_n N_VGND_c_1094_n 0.0141623f $X=5.225 $Y=0.46 $X2=0
+ $Y2=0
cc_553 N_A_1020_47#_c_818_n N_VGND_c_1094_n 0.00272823f $X=6.23 $Y=0.7 $X2=0
+ $Y2=0
cc_554 N_A_1020_47#_c_816_n N_VGND_c_1095_n 0.00995471f $X=6.47 $Y=0.995 $X2=0
+ $Y2=0
cc_555 N_A_1020_47#_c_817_n N_VGND_c_1095_n 4.79177e-19 $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_556 N_A_1020_47#_c_818_n N_VGND_c_1095_n 0.051428f $X=6.23 $Y=0.7 $X2=0 $Y2=0
cc_557 N_A_1020_47#_c_822_n N_VGND_c_1095_n 3.22676e-19 $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_558 N_A_1020_47#_M1014_s N_VGND_c_1096_n 0.00225325f $X=5.1 $Y=0.235 $X2=0
+ $Y2=0
cc_559 N_A_1020_47#_c_816_n N_VGND_c_1096_n 0.00937895f $X=6.47 $Y=0.995 $X2=0
+ $Y2=0
cc_560 N_A_1020_47#_c_817_n N_VGND_c_1096_n 0.0106281f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_561 N_A_1020_47#_c_827_n N_VGND_c_1096_n 0.00795901f $X=5.225 $Y=0.46 $X2=0
+ $Y2=0
cc_562 N_A_1020_47#_c_818_n N_VGND_c_1096_n 0.00875485f $X=6.23 $Y=0.7 $X2=0
+ $Y2=0
cc_563 N_A_1020_47#_c_818_n A_1102_47# 9.80231e-19 $X=6.23 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_564 N_VPWR_c_898_n A_109_369# 0.00168634f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_565 N_VPWR_c_898_n N_A_27_47#_M1003_d 0.00386882f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_566 N_VPWR_c_900_n N_A_27_47#_c_1001_n 0.0101554f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_567 N_VPWR_c_909_n N_A_27_47#_c_1012_n 0.0098369f $X=2.375 $Y=2.44 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_898_n N_A_27_47#_c_1012_n 0.00639994f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_909_n N_A_27_47#_c_1020_n 0.033302f $X=2.375 $Y=2.44 $X2=0 $Y2=0
cc_570 N_VPWR_c_898_n N_A_27_47#_c_1020_n 0.0209902f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_571 N_VPWR_c_898_n A_383_413# 0.00809303f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_572 N_VPWR_c_898_n N_GCLK_M1013_s 0.00307068f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_573 N_VPWR_c_908_n GCLK 0.0157287f $X=7.01 $Y=2.72 $X2=0 $Y2=0
cc_574 N_VPWR_c_898_n GCLK 0.0102114f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_575 N_VPWR_c_903_n GCLK 0.022003f $X=7.1 $Y=1.66 $X2=0 $Y2=0
cc_576 A_109_369# N_A_27_47#_c_1001_n 0.00276145f $X=0.545 $Y=1.845 $X2=0 $Y2=0
cc_577 A_109_369# N_A_27_47#_c_1012_n 8.01918e-19 $X=0.545 $Y=1.845 $X2=0 $Y2=0
cc_578 A_109_369# N_A_27_47#_c_1020_n 6.12987e-19 $X=0.545 $Y=1.845 $X2=0.215
+ $Y2=2
cc_579 N_A_27_47#_c_1002_n N_VGND_M1023_d 7.33468e-19 $X=1.015 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_580 N_A_27_47#_c_1003_n N_VGND_M1023_d 8.45526e-19 $X=0.685 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_581 N_A_27_47#_c_1003_n N_VGND_c_1082_n 0.0158273f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_582 N_A_27_47#_c_1000_n N_VGND_c_1087_n 0.0172026f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_583 N_A_27_47#_c_1003_n N_VGND_c_1087_n 0.00258611f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_584 N_A_27_47#_c_1002_n N_VGND_c_1088_n 0.00256355f $X=1.015 $Y=0.7 $X2=0
+ $Y2=0
cc_585 N_A_27_47#_c_1025_n N_VGND_c_1088_n 0.0120906f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_586 N_A_27_47#_M1023_s N_VGND_c_1096_n 0.00226128f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_587 N_A_27_47#_M1010_d N_VGND_c_1096_n 0.00617083f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_588 N_A_27_47#_c_1000_n N_VGND_c_1096_n 0.00977915f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_589 N_A_27_47#_c_1002_n N_VGND_c_1096_n 0.00427891f $X=1.015 $Y=0.7 $X2=0
+ $Y2=0
cc_590 N_A_27_47#_c_1003_n N_VGND_c_1096_n 0.00582244f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_591 N_A_27_47#_c_1025_n N_VGND_c_1096_n 0.00681108f $X=1.1 $Y=0.42 $X2=0
+ $Y2=0
cc_592 GCLK N_VGND_c_1086_n 0.022003f $X=7.105 $Y=1.105 $X2=0 $Y2=0
cc_593 N_GCLK_c_1073_n N_VGND_c_1090_n 0.0156348f $X=6.68 $Y=0.42 $X2=0 $Y2=0
cc_594 N_GCLK_M1002_s N_VGND_c_1096_n 0.0030199f $X=6.545 $Y=0.235 $X2=0 $Y2=0
cc_595 N_GCLK_c_1073_n N_VGND_c_1096_n 0.0101215f $X=6.68 $Y=0.42 $X2=0 $Y2=0
cc_596 N_VGND_c_1096_n A_395_47# 0.00299863f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_597 N_VGND_c_1095_n A_1102_47# 0.00105937f $X=6.4 $Y=0.18 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__bufinv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.265000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  4.295000 0.255000  4.545000 0.260000 ;
        RECT  4.295000 0.260000  4.625000 0.735000 ;
        RECT  4.295000 0.735000 10.955000 0.905000 ;
        RECT  4.295000 1.445000 10.955000 1.615000 ;
        RECT  4.295000 1.615000  4.625000 2.465000 ;
        RECT  5.135000 0.260000  5.465000 0.735000 ;
        RECT  5.135000 1.615000  5.465000 2.465000 ;
        RECT  5.215000 0.255000  5.385000 0.260000 ;
        RECT  5.975000 0.260000  6.305000 0.735000 ;
        RECT  5.975000 1.615000  6.305000 2.465000 ;
        RECT  6.055000 0.255000  6.225000 0.260000 ;
        RECT  6.815000 0.260000  7.145000 0.735000 ;
        RECT  6.815000 1.615000  7.145000 2.465000 ;
        RECT  7.655000 0.260000  7.985000 0.735000 ;
        RECT  7.655000 1.615000  7.985000 2.465000 ;
        RECT  8.495000 0.260000  8.825000 0.735000 ;
        RECT  8.495000 1.615000  8.825000 2.465000 ;
        RECT  9.335000 0.260000  9.665000 0.735000 ;
        RECT  9.335000 1.615000  9.665000 2.465000 ;
        RECT 10.175000 0.260000 10.505000 0.735000 ;
        RECT 10.175000 1.615000 10.505000 2.465000 ;
        RECT 10.680000 0.905000 10.955000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.595000  0.085000  0.765000 0.565000 ;
        RECT  1.435000  0.085000  1.605000 0.565000 ;
        RECT  2.275000  0.085000  2.445000 0.565000 ;
        RECT  3.115000  0.085000  3.285000 0.565000 ;
        RECT  3.955000  0.085000  4.125000 0.565000 ;
        RECT  4.795000  0.085000  4.965000 0.565000 ;
        RECT  5.635000  0.085000  5.805000 0.565000 ;
        RECT  6.475000  0.085000  6.645000 0.565000 ;
        RECT  7.315000  0.085000  7.485000 0.565000 ;
        RECT  8.155000  0.085000  8.325000 0.565000 ;
        RECT  8.995000  0.085000  9.165000 0.565000 ;
        RECT  9.835000  0.085000 10.005000 0.565000 ;
        RECT 10.675000  0.085000 10.845000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.040000 2.805000 ;
        RECT  0.595000 1.785000  0.765000 2.635000 ;
        RECT  1.435000 1.785000  1.605000 2.635000 ;
        RECT  2.275000 1.835000  2.445000 2.635000 ;
        RECT  3.115000 1.835000  3.285000 2.635000 ;
        RECT  3.955000 1.835000  4.125000 2.635000 ;
        RECT  4.795000 1.835000  4.965000 2.635000 ;
        RECT  5.635000 1.835000  5.805000 2.635000 ;
        RECT  6.475000 1.835000  6.645000 2.635000 ;
        RECT  7.315000 1.835000  7.485000 2.635000 ;
        RECT  8.155000 1.835000  8.325000 2.635000 ;
        RECT  8.995000 1.835000  9.165000 2.635000 ;
        RECT  9.835000 1.835000 10.005000 2.635000 ;
        RECT 10.675000 1.835000 10.845000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.260000  0.425000 0.735000 ;
      RECT 0.095000 0.735000  1.605000 0.905000 ;
      RECT 0.095000 1.445000  1.605000 1.615000 ;
      RECT 0.095000 1.615000  0.425000 2.465000 ;
      RECT 0.935000 0.260000  1.265000 0.735000 ;
      RECT 0.935000 1.615000  1.265000 2.465000 ;
      RECT 1.435000 0.905000  1.605000 1.075000 ;
      RECT 1.435000 1.075000  3.745000 1.275000 ;
      RECT 1.435000 1.275000  1.605000 1.445000 ;
      RECT 1.775000 0.260000  2.105000 0.735000 ;
      RECT 1.775000 0.735000  4.125000 0.905000 ;
      RECT 1.775000 1.445000  4.125000 1.615000 ;
      RECT 1.775000 1.615000  2.105000 2.465000 ;
      RECT 2.615000 0.260000  2.945000 0.735000 ;
      RECT 2.615000 1.615000  2.945000 2.465000 ;
      RECT 3.455000 0.260000  3.785000 0.735000 ;
      RECT 3.455000 1.615000  3.785000 2.465000 ;
      RECT 3.950000 0.905000  4.125000 1.075000 ;
      RECT 3.950000 1.075000 10.510000 1.275000 ;
      RECT 3.950000 1.275000  4.125000 1.445000 ;
  END
END sky130_fd_sc_hd__bufinv_16

* File: sky130_fd_sc_hd__or3_2.spice.SKY130_FD_SC_HD__OR3_2.pxi
* Created: Thu Aug 27 14:43:24 2020
* 
x_PM_SKY130_FD_SC_HD__OR3_2%C N_C_M1001_g N_C_M1005_g C N_C_c_61_n
+ PM_SKY130_FD_SC_HD__OR3_2%C
x_PM_SKY130_FD_SC_HD__OR3_2%B N_B_M1002_g N_B_M1009_g N_B_c_86_n N_B_c_87_n B B
+ N_B_c_89_n N_B_c_90_n PM_SKY130_FD_SC_HD__OR3_2%B
x_PM_SKY130_FD_SC_HD__OR3_2%A N_A_M1008_g N_A_M1007_g A A A N_A_c_128_n
+ N_A_c_129_n N_A_c_130_n PM_SKY130_FD_SC_HD__OR3_2%A
x_PM_SKY130_FD_SC_HD__OR3_2%A_30_53# N_A_30_53#_M1001_s N_A_30_53#_M1009_d
+ N_A_30_53#_M1005_s N_A_30_53#_c_179_n N_A_30_53#_M1004_g N_A_30_53#_M1000_g
+ N_A_30_53#_c_180_n N_A_30_53#_M1006_g N_A_30_53#_M1003_g N_A_30_53#_c_181_n
+ N_A_30_53#_c_182_n N_A_30_53#_c_183_n N_A_30_53#_c_191_n N_A_30_53#_c_278_p
+ N_A_30_53#_c_184_n N_A_30_53#_c_210_n N_A_30_53#_c_192_n N_A_30_53#_c_193_n
+ N_A_30_53#_c_185_n N_A_30_53#_c_194_n N_A_30_53#_c_186_n N_A_30_53#_c_187_n
+ N_A_30_53#_c_188_n PM_SKY130_FD_SC_HD__OR3_2%A_30_53#
x_PM_SKY130_FD_SC_HD__OR3_2%VPWR N_VPWR_M1007_d N_VPWR_M1003_d N_VPWR_c_294_n
+ N_VPWR_c_295_n N_VPWR_c_296_n VPWR N_VPWR_c_297_n N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_293_n PM_SKY130_FD_SC_HD__OR3_2%VPWR
x_PM_SKY130_FD_SC_HD__OR3_2%X N_X_M1004_s N_X_M1000_s N_X_c_328_n N_X_c_330_n
+ N_X_c_326_n X PM_SKY130_FD_SC_HD__OR3_2%X
x_PM_SKY130_FD_SC_HD__OR3_2%VGND N_VGND_M1001_d N_VGND_M1008_d N_VGND_M1006_d
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n VGND
+ N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n
+ N_VGND_c_360_n PM_SKY130_FD_SC_HD__OR3_2%VGND
cc_1 VNB N_C_M1001_g 0.0346235f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.475
cc_2 VNB C 0.0151697f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_C_c_61_n 0.0367867f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_4 VNB N_B_M1002_g 0.0163726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_B_c_86_n 0.013575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_B_c_87_n 0.0110772f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_7 VNB N_A_M1008_g 0.0266374f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.475
cc_8 VNB N_A_c_128_n 0.0206834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_c_129_n 0.00216296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_130_n 0.00336902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_30_53#_c_179_n 0.0164401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_30_53#_c_180_n 0.0207347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_30_53#_c_181_n 0.0135183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_30_53#_c_182_n 0.00380274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_30_53#_c_183_n 0.00916336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_30_53#_c_184_n 0.00106516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_30_53#_c_185_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_30_53#_c_186_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_30_53#_c_187_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_30_53#_c_188_n 0.0464346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_293_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_326_n 7.68963e-19 $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_23 VNB N_VGND_c_351_n 0.00101984f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_24 VNB N_VGND_c_352_n 5.60747e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_353_n 0.0104904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_354_n 0.036417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_355_n 0.0152668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_356_n 0.0115649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_357_n 0.0171221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_358_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_359_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_360_n 0.165754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_C_M1005_g 0.025409f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.695
cc_34 VPB C 0.00431076f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_35 VPB N_C_c_61_n 0.0101292f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_36 VPB N_B_M1002_g 0.0242436f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_B_c_89_n 0.0370191f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_38 VPB N_B_c_90_n 0.0354382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_M1007_g 0.0214023f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.695
cc_40 VPB A 0.00148181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_c_128_n 0.00403484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_c_129_n 0.00322575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_30_53#_M1000_g 0.0209283f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_44 VPB N_A_30_53#_M1003_g 0.0238856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_30_53#_c_191_n 0.00292112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_30_53#_c_192_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_30_53#_c_193_n 0.0209903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_30_53#_c_194_n 0.00139593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_30_53#_c_188_n 0.00736414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_294_n 0.0120872f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_51 VPB N_VPWR_c_295_n 0.0104612f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_52 VPB N_VPWR_c_296_n 0.0504714f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_53 VPB N_VPWR_c_297_n 0.0381055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_298_n 0.018077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_299_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_293_n 0.0566157f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_X_c_326_n 0.00111849f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_58 C N_B_M1002_g 2.5296e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_59 N_C_c_61_n N_B_M1002_g 0.0395944f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_60 N_C_M1001_g N_B_c_86_n 0.0136742f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_61 N_C_M1001_g N_B_c_87_n 0.0395944f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_62 N_C_M1005_g N_B_c_90_n 0.00441056f $X=0.485 $Y=1.695 $X2=0 $Y2=0
cc_63 N_C_M1005_g A 0.00430965f $X=0.485 $Y=1.695 $X2=0 $Y2=0
cc_64 C N_A_c_130_n 0.0279382f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_65 N_C_c_61_n N_A_c_130_n 0.00270522f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_66 N_C_M1001_g N_A_30_53#_c_182_n 0.0163896f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_67 C N_A_30_53#_c_182_n 0.00546144f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_68 N_C_c_61_n N_A_30_53#_c_182_n 3.50292e-19 $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_69 C N_A_30_53#_c_183_n 0.0212035f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_70 N_C_c_61_n N_A_30_53#_c_183_n 0.00184772f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_71 N_C_M1005_g N_A_30_53#_c_191_n 0.0104454f $X=0.485 $Y=1.695 $X2=0 $Y2=0
cc_72 N_C_M1005_g N_A_30_53#_c_193_n 0.00733639f $X=0.485 $Y=1.695 $X2=0 $Y2=0
cc_73 C N_A_30_53#_c_193_n 0.0239899f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_74 N_C_c_61_n N_A_30_53#_c_193_n 0.00205394f $X=0.485 $Y=1.16 $X2=0 $Y2=0
cc_75 N_C_M1001_g N_VGND_c_351_n 0.00953333f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_76 N_C_M1001_g N_VGND_c_355_n 0.00322006f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_77 N_C_M1001_g N_VGND_c_360_n 0.00466042f $X=0.485 $Y=0.475 $X2=0 $Y2=0
cc_78 N_B_M1002_g N_A_M1008_g 0.0033853f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_79 N_B_c_86_n N_A_M1008_g 0.0187947f $X=0.875 $Y=0.76 $X2=0 $Y2=0
cc_80 N_B_M1002_g N_A_M1007_g 0.0246267f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_81 N_B_c_90_n N_A_M1007_g 9.37151e-19 $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_82 N_B_M1002_g A 0.00791433f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_83 N_B_M1002_g N_A_c_128_n 0.0167622f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_84 N_B_M1002_g N_A_c_129_n 0.00970058f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_85 N_B_c_87_n N_A_c_129_n 0.00177283f $X=0.875 $Y=0.91 $X2=0 $Y2=0
cc_86 N_B_M1002_g N_A_c_130_n 0.00470079f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_87 N_B_c_86_n N_A_30_53#_c_182_n 0.00683722f $X=0.875 $Y=0.76 $X2=0 $Y2=0
cc_88 N_B_c_87_n N_A_30_53#_c_182_n 0.00604526f $X=0.875 $Y=0.91 $X2=0 $Y2=0
cc_89 N_B_M1002_g N_A_30_53#_c_191_n 0.0104077f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_90 N_B_c_89_n N_A_30_53#_c_191_n 0.00120401f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_91 N_B_c_90_n N_A_30_53#_c_191_n 0.0489918f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_92 N_B_c_90_n N_A_30_53#_c_210_n 3.54753e-19 $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_93 N_B_M1002_g N_A_30_53#_c_193_n 6.80151e-19 $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_94 N_B_c_90_n N_A_30_53#_c_193_n 0.0268584f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_95 N_B_M1002_g N_A_30_53#_c_194_n 0.00286901f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_96 N_B_c_90_n N_A_30_53#_c_194_n 0.0137296f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_97 N_B_M1002_g N_VPWR_c_294_n 0.00249809f $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_98 N_B_c_89_n N_VPWR_c_294_n 7.14013e-19 $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_99 N_B_c_90_n N_VPWR_c_294_n 0.0251801f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_100 N_B_c_89_n N_VPWR_c_297_n 0.00736312f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_101 N_B_c_90_n N_VPWR_c_297_n 0.0598896f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_102 N_B_c_89_n N_VPWR_c_293_n 0.0106165f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_103 N_B_c_90_n N_VPWR_c_293_n 0.0435145f $X=0.905 $Y=2.28 $X2=0 $Y2=0
cc_104 N_B_c_86_n N_VGND_c_351_n 0.00679416f $X=0.875 $Y=0.76 $X2=0 $Y2=0
cc_105 N_B_c_87_n N_VGND_c_351_n 2.19529e-19 $X=0.875 $Y=0.91 $X2=0 $Y2=0
cc_106 N_B_c_86_n N_VGND_c_352_n 5.25642e-19 $X=0.875 $Y=0.76 $X2=0 $Y2=0
cc_107 N_B_c_86_n N_VGND_c_356_n 0.00322006f $X=0.875 $Y=0.76 $X2=0 $Y2=0
cc_108 N_B_c_86_n N_VGND_c_360_n 0.00390029f $X=0.875 $Y=0.76 $X2=0 $Y2=0
cc_109 N_A_M1008_g N_A_30_53#_c_179_n 0.0172443f $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_110 N_A_M1007_g N_A_30_53#_M1000_g 0.0189524f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_111 N_A_c_129_n N_A_30_53#_c_182_n 0.0148461f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_c_130_n N_A_30_53#_c_182_n 0.0183663f $X=0.717 $Y=1.325 $X2=0 $Y2=0
cc_113 N_A_M1007_g N_A_30_53#_c_191_n 2.12667e-19 $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_114 A N_A_30_53#_c_191_n 0.0122114f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_115 N_A_c_129_n N_A_30_53#_c_191_n 0.00875823f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_M1008_g N_A_30_53#_c_184_n 0.0116406f $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_117 N_A_c_128_n N_A_30_53#_c_184_n 0.00220162f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_c_129_n N_A_30_53#_c_184_n 0.0166868f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_M1007_g N_A_30_53#_c_210_n 0.0117152f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_120 N_A_c_129_n N_A_30_53#_c_210_n 0.0104093f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_M1007_g N_A_30_53#_c_192_n 0.0034529f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_122 N_A_c_128_n N_A_30_53#_c_185_n 5.77159e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_129_n N_A_30_53#_c_185_n 0.0146254f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_M1007_g N_A_30_53#_c_194_n 0.00969506f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_125 A N_A_30_53#_c_194_n 0.00603332f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_126 N_A_c_128_n N_A_30_53#_c_194_n 0.00156816f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_129_n N_A_30_53#_c_194_n 0.0112884f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_c_128_n N_A_30_53#_c_186_n 0.00186332f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_c_129_n N_A_30_53#_c_186_n 0.0271506f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_M1008_g N_A_30_53#_c_187_n 0.0034529f $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_131 N_A_c_128_n N_A_30_53#_c_188_n 0.0203649f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_c_129_n N_A_30_53#_c_188_n 3.51645e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_133 A A_112_297# 0.00106198f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_134 N_A_M1007_g N_VPWR_c_294_n 0.00294311f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_135 N_A_M1007_g N_VPWR_c_297_n 0.00264561f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_136 N_A_M1007_g N_VPWR_c_293_n 0.00333991f $X=1.325 $Y=1.695 $X2=0 $Y2=0
cc_137 N_A_M1008_g N_VGND_c_351_n 5.2354e-19 $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_138 N_A_M1008_g N_VGND_c_352_n 0.00709299f $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_139 N_A_M1008_g N_VGND_c_356_n 0.00322006f $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_140 N_A_M1008_g N_VGND_c_360_n 0.00390029f $X=1.325 $Y=0.475 $X2=0 $Y2=0
cc_141 N_A_30_53#_c_191_n A_112_297# 0.0010205f $X=1.1 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_142 N_A_30_53#_c_191_n A_184_297# 0.0024109f $X=1.1 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_30_53#_c_194_n A_184_297# 0.0048682f $X=1.185 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_144 N_A_30_53#_c_210_n N_VPWR_M1007_d 0.00526233f $X=1.6 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A_30_53#_M1000_g N_VPWR_c_294_n 0.00348231f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_30_53#_c_210_n N_VPWR_c_294_n 0.0190361f $X=1.6 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A_30_53#_c_194_n N_VPWR_c_294_n 0.00579452f $X=1.185 $Y=1.58 $X2=0
+ $Y2=0
cc_148 N_A_30_53#_c_188_n N_VPWR_c_294_n 2.11345e-19 $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_30_53#_M1003_g N_VPWR_c_296_n 0.00736854f $X=2.235 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_30_53#_M1000_g N_VPWR_c_298_n 0.00585385f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_30_53#_M1003_g N_VPWR_c_298_n 0.00503406f $X=2.235 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_30_53#_M1000_g N_VPWR_c_293_n 0.0118387f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_30_53#_M1003_g N_VPWR_c_293_n 0.0096815f $X=2.235 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_30_53#_c_180_n N_X_c_328_n 0.00536146f $X=2.235 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_30_53#_c_188_n N_X_c_328_n 0.00259703f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_30_53#_M1003_g N_X_c_330_n 0.00294462f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_30_53#_c_188_n N_X_c_330_n 0.00288868f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_30_53#_c_179_n N_X_c_326_n 0.00151661f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_30_53#_M1000_g N_X_c_326_n 0.00115345f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_30_53#_c_180_n N_X_c_326_n 0.0069941f $X=2.235 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_30_53#_M1003_g N_X_c_326_n 0.00632068f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_30_53#_c_184_n N_X_c_326_n 0.00352178f $X=1.6 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_30_53#_c_192_n N_X_c_326_n 0.00841218f $X=1.685 $Y=1.495 $X2=0 $Y2=0
cc_164 N_A_30_53#_c_186_n N_X_c_326_n 0.0232251f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_30_53#_c_187_n N_X_c_326_n 0.00836616f $X=1.737 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_30_53#_c_188_n N_X_c_326_n 0.0230606f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_30_53#_M1003_g X 0.0119134f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_30_53#_c_182_n N_VGND_M1001_d 0.00160115f $X=1.03 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_30_53#_c_184_n N_VGND_M1008_d 0.00482895f $X=1.6 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_30_53#_c_187_n N_VGND_M1008_d 6.98847e-19 $X=1.737 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_30_53#_c_182_n N_VGND_c_351_n 0.0160613f $X=1.03 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_30_53#_c_179_n N_VGND_c_352_n 0.0079064f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_30_53#_c_180_n N_VGND_c_352_n 9.49203e-19 $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_174 N_A_30_53#_c_184_n N_VGND_c_352_n 0.020701f $X=1.6 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_30_53#_c_188_n N_VGND_c_352_n 2.33671e-19 $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_A_30_53#_c_180_n N_VGND_c_354_n 0.00674522f $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_30_53#_c_181_n N_VGND_c_355_n 0.0131002f $X=0.275 $Y=0.47 $X2=0 $Y2=0
cc_178 N_A_30_53#_c_182_n N_VGND_c_355_n 0.00232396f $X=1.03 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_30_53#_c_182_n N_VGND_c_356_n 0.00232396f $X=1.03 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_30_53#_c_278_p N_VGND_c_356_n 0.00846569f $X=1.115 $Y=0.47 $X2=0
+ $Y2=0
cc_181 N_A_30_53#_c_184_n N_VGND_c_356_n 0.00232396f $X=1.6 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_30_53#_c_179_n N_VGND_c_357_n 0.00524631f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_30_53#_c_180_n N_VGND_c_357_n 0.00513402f $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_30_53#_c_184_n N_VGND_c_357_n 3.34073e-19 $X=1.6 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_30_53#_c_179_n N_VGND_c_360_n 0.00851181f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_30_53#_c_180_n N_VGND_c_360_n 0.00968945f $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_30_53#_c_181_n N_VGND_c_360_n 0.00942308f $X=0.275 $Y=0.47 $X2=0
+ $Y2=0
cc_188 N_A_30_53#_c_182_n N_VGND_c_360_n 0.00970544f $X=1.03 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_30_53#_c_278_p N_VGND_c_360_n 0.00625722f $X=1.115 $Y=0.47 $X2=0
+ $Y2=0
cc_190 N_A_30_53#_c_184_n N_VGND_c_360_n 0.00637905f $X=1.6 $Y=0.74 $X2=0 $Y2=0
cc_191 N_VPWR_c_293_n N_X_M1000_s 0.00393857f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_296_n N_X_c_326_n 0.0783202f $X=2.47 $Y=1.62 $X2=0 $Y2=0
cc_193 N_VPWR_c_298_n X 0.0168871f $X=2.385 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_c_293_n X 0.0102668f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_296_n N_VGND_c_354_n 0.0124587f $X=2.47 $Y=1.62 $X2=0 $Y2=0
cc_196 N_X_c_328_n N_VGND_c_354_n 0.0261408f $X=2.13 $Y=0.587 $X2=0 $Y2=0
cc_197 N_X_c_326_n N_VGND_c_354_n 0.011394f $X=2.077 $Y=1.495 $X2=0 $Y2=0
cc_198 N_X_c_328_n N_VGND_c_357_n 0.00796253f $X=2.13 $Y=0.587 $X2=0 $Y2=0
cc_199 N_X_M1004_s N_VGND_c_360_n 0.00409985f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_200 N_X_c_328_n N_VGND_c_360_n 0.00913686f $X=2.13 $Y=0.587 $X2=0 $Y2=0

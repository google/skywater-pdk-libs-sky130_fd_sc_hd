# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__xor3_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__xor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.525000 1.075000 8.935000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 0.995000 7.875000 1.445000 ;
        RECT 7.705000 1.445000 8.285000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.880000 0.995000 3.515000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.350000 0.765000 0.660000 ;
        RECT 0.595000 0.660000 1.605000 0.830000 ;
        RECT 0.595000 0.830000 1.535000 0.925000 ;
        RECT 0.695000 1.440000 1.420000 1.455000 ;
        RECT 0.695000 1.455000 1.705000 2.045000 ;
        RECT 0.695000 2.045000 0.865000 2.465000 ;
        RECT 1.105000 0.925000 1.420000 1.440000 ;
        RECT 1.435000 0.350000 1.605000 0.660000 ;
        RECT 1.535000 2.045000 1.705000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.175000  0.085000  0.345000 0.545000 ;
        RECT 0.935000  0.085000  1.265000 0.465000 ;
        RECT 1.855000  0.085000  2.025000 0.525000 ;
        RECT 4.950000  0.085000  5.120000 0.885000 ;
        RECT 8.995000  0.085000  9.165000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
        RECT 9.805000 -0.085000 9.975000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.275000 2.135000  0.445000 2.635000 ;
        RECT 1.035000 2.215000  1.365000 2.635000 ;
        RECT 1.875000 2.215000  2.205000 2.635000 ;
        RECT 4.705000 2.235000  5.035000 2.635000 ;
        RECT 8.915000 2.275000  9.245000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
        RECT 9.805000 2.635000 9.975000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.820000 0.965000 2.045000 1.325000 ;
      RECT 1.875000 0.695000 2.365000 0.865000 ;
      RECT 1.875000 0.865000 2.045000 0.965000 ;
      RECT 1.875000 1.325000 2.045000 1.875000 ;
      RECT 1.875000 1.875000 2.545000 2.045000 ;
      RECT 2.195000 0.255000 3.760000 0.425000 ;
      RECT 2.195000 0.425000 2.365000 0.695000 ;
      RECT 2.370000 1.535000 3.855000 1.705000 ;
      RECT 2.375000 2.045000 2.545000 2.235000 ;
      RECT 2.375000 2.235000 3.915000 2.405000 ;
      RECT 2.540000 0.595000 2.710000 1.535000 ;
      RECT 2.890000 1.895000 4.195000 2.065000 ;
      RECT 2.990000 0.655000 4.100000 0.825000 ;
      RECT 3.410000 0.425000 3.760000 0.455000 ;
      RECT 3.685000 0.995000 4.055000 1.325000 ;
      RECT 3.685000 1.325000 3.855000 1.535000 ;
      RECT 3.930000 0.255000 4.780000 0.425000 ;
      RECT 3.930000 0.425000 4.100000 0.655000 ;
      RECT 4.025000 1.525000 4.555000 1.695000 ;
      RECT 4.025000 1.695000 4.195000 1.895000 ;
      RECT 4.130000 2.235000 4.535000 2.405000 ;
      RECT 4.270000 0.595000 4.440000 1.375000 ;
      RECT 4.270000 1.375000 4.555000 1.525000 ;
      RECT 4.365000 1.895000 5.540000 2.065000 ;
      RECT 4.365000 2.065000 4.535000 2.235000 ;
      RECT 4.610000 0.425000 4.780000 1.035000 ;
      RECT 4.610000 1.035000 4.865000 1.040000 ;
      RECT 4.610000 1.040000 4.880000 1.045000 ;
      RECT 4.610000 1.045000 4.890000 1.050000 ;
      RECT 4.610000 1.050000 4.895000 1.205000 ;
      RECT 4.725000 1.205000 4.895000 1.895000 ;
      RECT 5.125000 1.445000 5.540000 1.715000 ;
      RECT 5.300000 0.415000 5.540000 1.445000 ;
      RECT 5.370000 2.065000 5.540000 2.275000 ;
      RECT 5.370000 2.275000 8.465000 2.445000 ;
      RECT 5.715000 0.265000 6.130000 0.485000 ;
      RECT 5.715000 0.485000 5.935000 0.595000 ;
      RECT 5.715000 0.595000 5.885000 2.105000 ;
      RECT 6.075000 0.720000 6.470000 0.825000 ;
      RECT 6.075000 0.825000 6.275000 0.890000 ;
      RECT 6.075000 0.890000 6.245000 2.275000 ;
      RECT 6.105000 0.655000 6.470000 0.720000 ;
      RECT 6.300000 0.320000 6.470000 0.655000 ;
      RECT 6.415000 1.445000 7.195000 1.615000 ;
      RECT 6.415000 1.615000 6.830000 2.045000 ;
      RECT 6.430000 0.995000 6.855000 1.270000 ;
      RECT 6.640000 0.630000 6.855000 0.995000 ;
      RECT 7.025000 0.255000 8.170000 0.425000 ;
      RECT 7.025000 0.425000 7.195000 1.445000 ;
      RECT 7.365000 0.595000 7.535000 1.935000 ;
      RECT 7.365000 1.935000 9.675000 2.105000 ;
      RECT 7.705000 0.425000 8.170000 0.465000 ;
      RECT 8.045000 0.730000 8.250000 0.945000 ;
      RECT 8.045000 0.945000 8.355000 1.275000 ;
      RECT 8.455000 1.495000 9.275000 1.705000 ;
      RECT 8.495000 0.295000 8.785000 0.735000 ;
      RECT 8.495000 0.735000 9.275000 0.750000 ;
      RECT 8.535000 0.750000 9.275000 0.905000 ;
      RECT 9.105000 0.905000 9.275000 0.995000 ;
      RECT 9.105000 0.995000 9.335000 1.325000 ;
      RECT 9.105000 1.325000 9.275000 1.495000 ;
      RECT 9.190000 1.875000 9.675000 1.935000 ;
      RECT 9.415000 0.255000 9.675000 0.585000 ;
      RECT 9.415000 2.105000 9.675000 2.465000 ;
      RECT 9.505000 0.585000 9.675000 1.875000 ;
    LAYER mcon ;
      RECT 4.385000 1.445000 4.555000 1.615000 ;
      RECT 5.305000 0.765000 5.475000 0.935000 ;
      RECT 5.765000 0.425000 5.935000 0.595000 ;
      RECT 6.685000 0.765000 6.855000 0.935000 ;
      RECT 6.685000 1.445000 6.855000 1.615000 ;
      RECT 8.065000 0.765000 8.235000 0.935000 ;
      RECT 8.525000 0.425000 8.695000 0.595000 ;
    LAYER met1 ;
      RECT 4.325000 1.415000 4.615000 1.460000 ;
      RECT 4.325000 1.460000 6.915000 1.600000 ;
      RECT 4.325000 1.600000 4.615000 1.645000 ;
      RECT 5.245000 0.735000 5.535000 0.780000 ;
      RECT 5.245000 0.780000 8.295000 0.920000 ;
      RECT 5.245000 0.920000 5.535000 0.965000 ;
      RECT 5.705000 0.395000 5.995000 0.440000 ;
      RECT 5.705000 0.440000 8.755000 0.580000 ;
      RECT 5.705000 0.580000 5.995000 0.625000 ;
      RECT 6.625000 0.735000 6.915000 0.780000 ;
      RECT 6.625000 0.920000 6.915000 0.965000 ;
      RECT 6.625000 1.415000 6.915000 1.460000 ;
      RECT 6.625000 1.600000 6.915000 1.645000 ;
      RECT 8.005000 0.735000 8.295000 0.780000 ;
      RECT 8.005000 0.920000 8.295000 0.965000 ;
      RECT 8.465000 0.395000 8.755000 0.440000 ;
      RECT 8.465000 0.580000 8.755000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_4
END LIBRARY

* File: sky130_fd_sc_hd__o21ai_2.pxi.spice
* Created: Thu Aug 27 14:35:45 2020
* 
x_PM_SKY130_FD_SC_HD__O21AI_2%A1 N_A1_c_55_n N_A1_M1009_g N_A1_M1003_g
+ N_A1_M1008_g N_A1_M1011_g N_A1_c_62_n N_A1_c_56_n N_A1_c_57_n A1 A1
+ N_A1_c_58_n PM_SKY130_FD_SC_HD__O21AI_2%A1
x_PM_SKY130_FD_SC_HD__O21AI_2%A2 N_A2_c_130_n N_A2_M1000_g N_A2_M1005_g
+ N_A2_c_131_n N_A2_M1004_g N_A2_M1010_g A2 N_A2_c_132_n N_A2_c_133_n
+ PM_SKY130_FD_SC_HD__O21AI_2%A2
x_PM_SKY130_FD_SC_HD__O21AI_2%B1 N_B1_c_183_n N_B1_M1002_g N_B1_M1001_g
+ N_B1_c_185_n N_B1_c_186_n N_B1_M1007_g N_B1_M1006_g N_B1_c_187_n B1 B1
+ N_B1_c_189_n PM_SKY130_FD_SC_HD__O21AI_2%B1
x_PM_SKY130_FD_SC_HD__O21AI_2%VPWR N_VPWR_M1003_s N_VPWR_M1008_s N_VPWR_M1006_d
+ N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n
+ VPWR N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_231_n
+ PM_SKY130_FD_SC_HD__O21AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O21AI_2%A_112_297# N_A_112_297#_M1003_d
+ N_A_112_297#_M1010_d N_A_112_297#_c_286_n N_A_112_297#_c_287_n
+ N_A_112_297#_c_293_n N_A_112_297#_c_295_n
+ PM_SKY130_FD_SC_HD__O21AI_2%A_112_297#
x_PM_SKY130_FD_SC_HD__O21AI_2%Y N_Y_M1002_d N_Y_M1005_s N_Y_M1001_s N_Y_c_323_n
+ Y Y Y Y N_Y_c_305_n N_Y_c_302_n N_Y_c_310_n PM_SKY130_FD_SC_HD__O21AI_2%Y
x_PM_SKY130_FD_SC_HD__O21AI_2%A_29_47# N_A_29_47#_M1009_d N_A_29_47#_M1000_d
+ N_A_29_47#_M1011_d N_A_29_47#_M1007_s N_A_29_47#_c_338_n N_A_29_47#_c_344_n
+ N_A_29_47#_c_339_n N_A_29_47#_c_349_n N_A_29_47#_c_340_n N_A_29_47#_c_355_n
+ N_A_29_47#_c_356_n N_A_29_47#_c_375_n N_A_29_47#_c_341_n N_A_29_47#_c_342_n
+ PM_SKY130_FD_SC_HD__O21AI_2%A_29_47#
x_PM_SKY130_FD_SC_HD__O21AI_2%VGND N_VGND_M1009_s N_VGND_M1004_s N_VGND_c_411_n
+ N_VGND_c_412_n VGND N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n PM_SKY130_FD_SC_HD__O21AI_2%VGND
cc_1 VNB N_A1_c_55_n 0.0662345f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.96
cc_2 VNB N_A1_c_56_n 0.00492907f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_3 VNB N_A1_c_57_n 0.0234542f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_4 VNB N_A1_c_58_n 0.0175595f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.995
cc_5 VNB N_A2_c_130_n 0.0163913f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.96
cc_6 VNB N_A2_c_131_n 0.0173283f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=1.325
cc_7 VNB N_A2_c_132_n 0.00529918f $X=-0.19 $Y=-0.24 $X2=1.847 $Y2=1.53
cc_8 VNB N_A2_c_133_n 0.0341549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_183_n 0.0145588f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.96
cc_10 VNB N_B1_M1001_g 0.00684821f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.985
cc_11 VNB N_B1_c_185_n 0.0117721f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=1.325
cc_12 VNB N_B1_c_186_n 0.0178464f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=1.985
cc_13 VNB N_B1_c_187_n 0.00685304f $X=-0.19 $Y=-0.24 $X2=1.847 $Y2=1.16
cc_14 VNB B1 0.0205286f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_15 VNB N_B1_c_189_n 0.0355749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_231_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_302_n 0.00295442f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_18 VNB N_A_29_47#_c_338_n 0.018052f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.53
cc_19 VNB N_A_29_47#_c_339_n 0.00909933f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_20 VNB N_A_29_47#_c_340_n 0.00429425f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_21 VNB N_A_29_47#_c_341_n 0.00126312f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_22 VNB N_A_29_47#_c_342_n 0.0136468f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.132
cc_23 VNB N_VGND_c_411_n 0.0047158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_412_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.53
cc_25 VNB N_VGND_c_413_n 0.0185988f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_26 VNB N_VGND_c_414_n 0.0381669f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_27 VNB N_VGND_c_415_n 0.181368f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_28 VNB N_VGND_c_416_n 0.0210524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_417_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.325
cc_30 VPB N_A1_c_55_n 0.00826134f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.96
cc_31 VPB N_A1_M1003_g 0.0235373f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_32 VPB N_A1_M1008_g 0.0185491f $X=-0.19 $Y=1.305 $X2=1.845 $Y2=1.985
cc_33 VPB N_A1_c_62_n 0.00778906f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.53
cc_34 VPB N_A1_c_56_n 0.00301297f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_35 VPB N_A1_c_57_n 0.00631455f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_36 VPB A1 0.00518033f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_37 VPB A1 0.00726806f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.445
cc_38 VPB N_A2_M1005_g 0.0186077f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_39 VPB N_A2_M1010_g 0.0193374f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=0.56
cc_40 VPB N_A2_c_133_n 0.00611931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B1_M1001_g 0.0204212f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_42 VPB N_B1_M1006_g 0.0238197f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.53
cc_43 VPB B1 0.00656808f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_44 VPB N_B1_c_189_n 0.010139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_232_n 0.0106587f $X=-0.19 $Y=1.305 $X2=1.845 $Y2=1.985
cc_46 VPB N_VPWR_c_233_n 0.0305655f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=0.995
cc_47 VPB N_VPWR_c_234_n 0.00227295f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.53
cc_48 VPB N_VPWR_c_235_n 0.00997098f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_49 VPB N_VPWR_c_236_n 0.0380928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_237_n 0.0333972f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.445
cc_51 VPB N_VPWR_c_238_n 0.0143915f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.132
cc_52 VPB N_VPWR_c_239_n 0.00519461f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.445
cc_53 VPB N_VPWR_c_231_n 0.0434267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_Y_c_302_n 0.00367686f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_55 N_A1_c_55_n N_A2_c_130_n 0.0255609f $X=0.485 $Y=0.96 $X2=-0.19 $Y2=-0.24
cc_56 N_A1_M1003_g N_A2_M1005_g 0.0267552f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A1_c_62_n N_A2_M1005_g 0.0149806f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_58 A1 N_A2_M1005_g 5.96887e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A1_c_58_n N_A2_c_131_n 0.0211228f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A1_M1008_g N_A2_M1010_g 0.032548f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A1_c_62_n N_A2_M1010_g 0.0101073f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_62 N_A1_c_55_n N_A2_c_132_n 0.00157245f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_63 N_A1_c_62_n N_A2_c_132_n 0.0573639f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_64 N_A1_c_56_n N_A2_c_132_n 0.0164124f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A1_c_57_n N_A2_c_132_n 2.11058e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_66 A1 N_A2_c_132_n 0.0166956f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A1_c_55_n N_A2_c_133_n 0.022502f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_68 N_A1_c_62_n N_A2_c_133_n 0.0040428f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_69 N_A1_c_56_n N_A2_c_133_n 0.0052341f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A1_c_57_n N_A2_c_133_n 0.0162104f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_71 A1 N_A2_c_133_n 5.80215e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_72 N_A1_c_58_n N_B1_c_183_n 0.0117405f $X=1.865 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_73 N_A1_M1008_g N_B1_M1001_g 0.0359212f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A1_c_56_n N_B1_c_187_n 0.00488621f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A1_c_57_n N_B1_c_187_n 0.021305f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_76 A1 N_VPWR_M1003_s 0.00289981f $X=0.14 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_77 N_A1_c_56_n N_VPWR_M1008_s 0.00277374f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A1_c_55_n N_VPWR_c_233_n 0.00107824f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_79 N_A1_M1003_g N_VPWR_c_233_n 0.013399f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_80 A1 N_VPWR_c_233_n 0.0227573f $X=0.14 $Y=1.445 $X2=0 $Y2=0
cc_81 N_A1_M1008_g N_VPWR_c_234_n 0.00764053f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A1_M1003_g N_VPWR_c_237_n 0.00486043f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A1_M1008_g N_VPWR_c_237_n 0.00411597f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A1_M1003_g N_VPWR_c_231_n 0.00825064f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A1_M1008_g N_VPWR_c_231_n 0.00500252f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A1_c_62_n N_A_112_297#_M1003_d 0.00176461f $X=1.6 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A1_c_62_n N_A_112_297#_M1010_d 0.00162243f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_88 N_A1_c_56_n N_A_112_297#_M1010_d 0.00154655f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A1_c_62_n N_A_112_297#_c_286_n 0.0135055f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_90 N_A1_c_62_n N_Y_M1005_s 0.00176891f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_91 N_A1_M1008_g N_Y_c_305_n 0.0131497f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A1_c_56_n N_Y_c_305_n 0.0296112f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A1_c_57_n N_Y_c_305_n 5.23705e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A1_c_56_n N_Y_c_302_n 0.0239848f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A1_c_57_n N_Y_c_302_n 4.57631e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A1_M1008_g N_Y_c_310_n 7.08948e-19 $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A1_c_62_n N_Y_c_310_n 0.0319158f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_98 N_A1_c_55_n N_A_29_47#_c_338_n 0.00614277f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_99 N_A1_c_55_n N_A_29_47#_c_344_n 0.0101054f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_100 N_A1_c_62_n N_A_29_47#_c_344_n 0.00381797f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_101 A1 N_A_29_47#_c_344_n 0.00101523f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A1_c_55_n N_A_29_47#_c_339_n 0.0081483f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_103 A1 N_A_29_47#_c_339_n 0.0242892f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A1_c_55_n N_A_29_47#_c_349_n 5.21391e-19 $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_105 N_A1_c_58_n N_A_29_47#_c_349_n 6.10472e-19 $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A1_c_62_n N_A_29_47#_c_340_n 0.00480305f $X=1.6 $Y=1.53 $X2=0 $Y2=0
cc_107 N_A1_c_56_n N_A_29_47#_c_340_n 0.032123f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A1_c_57_n N_A_29_47#_c_340_n 0.00424827f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A1_c_58_n N_A_29_47#_c_340_n 0.0101432f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A1_c_58_n N_A_29_47#_c_355_n 0.00224274f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A1_c_58_n N_A_29_47#_c_356_n 0.00475971f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_c_55_n N_VGND_c_411_n 0.00267631f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_113 N_A1_c_58_n N_VGND_c_412_n 0.00534468f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A1_c_58_n N_VGND_c_414_n 0.0042335f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A1_c_55_n N_VGND_c_415_n 0.00675612f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_116 N_A1_c_58_n N_VGND_c_415_n 0.00625656f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A1_c_55_n N_VGND_c_416_n 0.00424868f $X=0.485 $Y=0.96 $X2=0 $Y2=0
cc_118 N_A2_M1005_g N_VPWR_c_233_n 0.00107483f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A2_M1010_g N_VPWR_c_234_n 9.48926e-19 $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A2_M1005_g N_VPWR_c_237_n 0.00357877f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A2_M1010_g N_VPWR_c_237_n 0.00357877f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A2_M1005_g N_VPWR_c_231_n 0.00530427f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A2_M1010_g N_VPWR_c_231_n 0.00546392f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A2_M1005_g N_A_112_297#_c_287_n 0.0121906f $X=0.915 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A2_M1010_g N_A_112_297#_c_287_n 0.00837827f $X=1.345 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A2_M1010_g N_Y_c_305_n 0.00867291f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A2_M1010_g N_Y_c_310_n 0.0041292f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A2_c_130_n N_A_29_47#_c_338_n 5.21391e-19 $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_130_n N_A_29_47#_c_344_n 0.00883087f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_132_n N_A_29_47#_c_344_n 0.0208462f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A2_c_133_n N_A_29_47#_c_344_n 0.00154684f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A2_c_130_n N_A_29_47#_c_349_n 0.00614277f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_131_n N_A_29_47#_c_349_n 0.00692975f $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A2_c_131_n N_A_29_47#_c_340_n 0.0093975f $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A2_c_132_n N_A_29_47#_c_340_n 0.00781738f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A2_c_131_n N_A_29_47#_c_356_n 4.90982e-19 $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A2_c_130_n N_A_29_47#_c_341_n 7.36376e-19 $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A2_c_131_n N_A_29_47#_c_341_n 7.36376e-19 $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_132_n N_A_29_47#_c_341_n 0.019141f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A2_c_133_n N_A_29_47#_c_341_n 0.00253097f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_c_130_n N_VGND_c_411_n 0.00267631f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_131_n N_VGND_c_412_n 0.00384786f $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A2_c_130_n N_VGND_c_413_n 0.00424868f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A2_c_131_n N_VGND_c_413_n 0.00424868f $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A2_c_130_n N_VGND_c_415_n 0.00581418f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A2_c_131_n N_VGND_c_415_n 0.00616657f $X=1.345 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B1_M1001_g N_VPWR_c_234_n 0.00170542f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B1_M1001_g N_VPWR_c_236_n 6.89506e-19 $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B1_M1006_g N_VPWR_c_236_n 0.0156754f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_150 B1 N_VPWR_c_236_n 0.0255942f $X=2.9 $Y=0.765 $X2=0 $Y2=0
cc_151 N_B1_c_189_n N_VPWR_c_236_n 0.00174034f $X=2.745 $Y=1.142 $X2=0 $Y2=0
cc_152 N_B1_M1001_g N_VPWR_c_238_n 0.00441055f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B1_M1006_g N_VPWR_c_238_n 0.00564095f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B1_M1001_g N_VPWR_c_231_n 0.00604582f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B1_M1006_g N_VPWR_c_231_n 0.00953074f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B1_M1001_g N_Y_c_305_n 0.0160158f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B1_c_183_n N_Y_c_302_n 0.0018621f $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_158 N_B1_M1001_g N_Y_c_302_n 0.00312743f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B1_c_185_n N_Y_c_302_n 0.0144006f $X=2.67 $Y=1.062 $X2=0 $Y2=0
cc_160 N_B1_c_186_n N_Y_c_302_n 5.61747e-19 $X=2.745 $Y=0.96 $X2=0 $Y2=0
cc_161 B1 N_Y_c_302_n 0.0427649f $X=2.9 $Y=0.765 $X2=0 $Y2=0
cc_162 N_B1_c_189_n N_Y_c_302_n 0.0041517f $X=2.745 $Y=1.142 $X2=0 $Y2=0
cc_163 B1 N_A_29_47#_M1007_s 0.00248682f $X=2.9 $Y=0.765 $X2=0 $Y2=0
cc_164 N_B1_c_183_n N_A_29_47#_c_340_n 0.00296067f $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_165 N_B1_c_183_n N_A_29_47#_c_355_n 5.89792e-19 $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_166 N_B1_c_183_n N_A_29_47#_c_356_n 0.0042062f $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_167 N_B1_c_186_n N_A_29_47#_c_356_n 4.72667e-19 $X=2.745 $Y=0.96 $X2=0 $Y2=0
cc_168 N_B1_c_183_n N_A_29_47#_c_375_n 0.0105206f $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_169 N_B1_c_185_n N_A_29_47#_c_375_n 3.28898e-19 $X=2.67 $Y=1.062 $X2=0 $Y2=0
cc_170 N_B1_c_186_n N_A_29_47#_c_375_n 0.0124922f $X=2.745 $Y=0.96 $X2=0 $Y2=0
cc_171 N_B1_c_183_n N_A_29_47#_c_342_n 5.00002e-19 $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_172 N_B1_c_186_n N_A_29_47#_c_342_n 0.00334667f $X=2.745 $Y=0.96 $X2=0 $Y2=0
cc_173 B1 N_A_29_47#_c_342_n 0.0207723f $X=2.9 $Y=0.765 $X2=0 $Y2=0
cc_174 N_B1_c_189_n N_A_29_47#_c_342_n 0.00118211f $X=2.745 $Y=1.142 $X2=0 $Y2=0
cc_175 N_B1_c_183_n N_VGND_c_414_n 0.00357842f $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_176 N_B1_c_186_n N_VGND_c_414_n 0.00359389f $X=2.745 $Y=0.96 $X2=0 $Y2=0
cc_177 N_B1_c_183_n N_VGND_c_415_n 0.00530424f $X=2.315 $Y=0.96 $X2=0 $Y2=0
cc_178 N_B1_c_186_n N_VGND_c_415_n 0.00617523f $X=2.745 $Y=0.96 $X2=0 $Y2=0
cc_179 B1 N_VGND_c_415_n 8.28511e-19 $X=2.9 $Y=0.765 $X2=0 $Y2=0
cc_180 N_VPWR_c_231_n N_A_112_297#_M1003_d 0.00375981f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_181 N_VPWR_c_231_n N_A_112_297#_M1010_d 0.00308454f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_237_n N_A_112_297#_c_287_n 0.0385283f $X=1.91 $Y=2.72 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_231_n N_A_112_297#_c_287_n 0.0245637f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_237_n N_A_112_297#_c_293_n 0.0135892f $X=1.91 $Y=2.72 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_231_n N_A_112_297#_c_293_n 0.00847259f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_237_n N_A_112_297#_c_295_n 0.0124917f $X=1.91 $Y=2.72 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_231_n N_A_112_297#_c_295_n 0.00710224f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_231_n N_Y_M1005_s 0.00224864f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_c_231_n N_Y_M1001_s 0.00325133f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_238_n N_Y_c_323_n 0.0140505f $X=2.815 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_231_n N_Y_c_323_n 0.00897324f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_M1008_s N_Y_c_305_n 0.00694363f $X=1.92 $Y=1.485 $X2=0 $Y2=0
cc_193 N_VPWR_c_234_n N_Y_c_305_n 0.0140852f $X=2.075 $Y=2.34 $X2=0 $Y2=0
cc_194 N_VPWR_c_237_n N_Y_c_305_n 0.00217464f $X=1.91 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_238_n N_Y_c_305_n 0.0020229f $X=2.815 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_231_n N_Y_c_305_n 0.0102471f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_197 N_A_112_297#_c_287_n N_Y_M1005_s 0.003328f $X=1.525 $Y=2.38 $X2=0.485
+ $Y2=0.56
cc_198 N_A_112_297#_M1010_d N_Y_c_305_n 0.00510373f $X=1.42 $Y=1.485 $X2=0 $Y2=0
cc_199 N_A_112_297#_c_287_n N_Y_c_305_n 0.00623241f $X=1.525 $Y=2.38 $X2=0 $Y2=0
cc_200 N_A_112_297#_c_295_n N_Y_c_305_n 0.0138908f $X=1.61 $Y=2.3 $X2=0 $Y2=0
cc_201 N_A_112_297#_c_287_n N_Y_c_310_n 0.0135861f $X=1.525 $Y=2.38 $X2=0 $Y2=0
cc_202 N_Y_M1002_d N_A_29_47#_c_375_n 0.0032157f $X=2.39 $Y=0.235 $X2=0 $Y2=0
cc_203 N_Y_c_302_n N_A_29_47#_c_375_n 0.0126484f $X=2.53 $Y=0.76 $X2=0 $Y2=0
cc_204 N_Y_M1002_d N_VGND_c_415_n 0.00224864f $X=2.39 $Y=0.235 $X2=0 $Y2=0
cc_205 N_A_29_47#_c_344_n N_VGND_M1009_s 0.00350645f $X=0.965 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A_29_47#_c_340_n N_VGND_M1004_s 0.00795142f $X=1.935 $Y=0.8 $X2=0 $Y2=0
cc_207 N_A_29_47#_c_344_n N_VGND_c_411_n 0.0129597f $X=0.965 $Y=0.8 $X2=0 $Y2=0
cc_208 N_A_29_47#_c_349_n N_VGND_c_412_n 0.0169695f $X=1.13 $Y=0.4 $X2=0 $Y2=0
cc_209 N_A_29_47#_c_340_n N_VGND_c_412_n 0.0131159f $X=1.935 $Y=0.8 $X2=0 $Y2=0
cc_210 N_A_29_47#_c_355_n N_VGND_c_412_n 0.0102296f $X=2.1 $Y=0.425 $X2=0 $Y2=0
cc_211 N_A_29_47#_c_356_n N_VGND_c_412_n 0.00676824f $X=2.1 $Y=0.715 $X2=0 $Y2=0
cc_212 N_A_29_47#_c_344_n N_VGND_c_413_n 0.00213388f $X=0.965 $Y=0.8 $X2=0 $Y2=0
cc_213 N_A_29_47#_c_349_n N_VGND_c_413_n 0.0188428f $X=1.13 $Y=0.4 $X2=0 $Y2=0
cc_214 N_A_29_47#_c_340_n N_VGND_c_413_n 0.00285904f $X=1.935 $Y=0.8 $X2=0 $Y2=0
cc_215 N_A_29_47#_c_340_n N_VGND_c_414_n 0.0030068f $X=1.935 $Y=0.8 $X2=0 $Y2=0
cc_216 N_A_29_47#_c_355_n N_VGND_c_414_n 0.0189784f $X=2.1 $Y=0.425 $X2=0 $Y2=0
cc_217 N_A_29_47#_c_375_n N_VGND_c_414_n 0.0311267f $X=2.815 $Y=0.34 $X2=0 $Y2=0
cc_218 N_A_29_47#_c_342_n N_VGND_c_414_n 0.0188277f $X=2.97 $Y=0.34 $X2=0 $Y2=0
cc_219 N_A_29_47#_M1009_d N_VGND_c_415_n 0.00213418f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_A_29_47#_M1000_d N_VGND_c_415_n 0.00223231f $X=0.99 $Y=0.235 $X2=0
+ $Y2=0
cc_221 N_A_29_47#_M1011_d N_VGND_c_415_n 0.00223231f $X=1.96 $Y=0.235 $X2=0
+ $Y2=0
cc_222 N_A_29_47#_M1007_s N_VGND_c_415_n 0.00213418f $X=2.82 $Y=0.235 $X2=0
+ $Y2=0
cc_223 N_A_29_47#_c_338_n N_VGND_c_415_n 0.0124245f $X=0.27 $Y=0.4 $X2=0 $Y2=0
cc_224 N_A_29_47#_c_344_n N_VGND_c_415_n 0.00889701f $X=0.965 $Y=0.8 $X2=0 $Y2=0
cc_225 N_A_29_47#_c_349_n N_VGND_c_415_n 0.0122425f $X=1.13 $Y=0.4 $X2=0 $Y2=0
cc_226 N_A_29_47#_c_340_n N_VGND_c_415_n 0.0119492f $X=1.935 $Y=0.8 $X2=0 $Y2=0
cc_227 N_A_29_47#_c_355_n N_VGND_c_415_n 0.0123102f $X=2.1 $Y=0.425 $X2=0 $Y2=0
cc_228 N_A_29_47#_c_375_n N_VGND_c_415_n 0.0192538f $X=2.815 $Y=0.34 $X2=0 $Y2=0
cc_229 N_A_29_47#_c_342_n N_VGND_c_415_n 0.0115692f $X=2.97 $Y=0.34 $X2=0 $Y2=0
cc_230 N_A_29_47#_c_338_n N_VGND_c_416_n 0.0209424f $X=0.27 $Y=0.4 $X2=0 $Y2=0
cc_231 N_A_29_47#_c_344_n N_VGND_c_416_n 0.00213388f $X=0.965 $Y=0.8 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 1.355000 2.775000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.180000 0.305000 9.530000 0.725000 ;
        RECT 9.180000 0.725000 9.560000 0.790000 ;
        RECT 9.180000 0.790000 9.610000 0.825000 ;
        RECT 9.200000 1.505000 9.610000 1.540000 ;
        RECT 9.200000 1.540000 9.530000 2.465000 ;
        RECT 9.355000 1.430000 9.610000 1.505000 ;
        RECT 9.390000 0.825000 9.610000 1.430000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 0.265000 10.940000 0.795000 ;
        RECT 10.685000 1.445000 10.940000 2.325000 ;
        RECT 10.730000 0.795000 10.940000 1.445000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.055000 3.995000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.750000 3.235000 0.785000 ;
        RECT 1.760000 0.785000 2.010000 0.810000 ;
        RECT 1.760000 0.810000 1.990000 0.820000 ;
        RECT 1.760000 0.820000 1.975000 0.835000 ;
        RECT 1.760000 0.835000 1.970000 0.840000 ;
        RECT 1.760000 0.840000 1.965000 0.850000 ;
        RECT 1.760000 0.850000 1.960000 0.855000 ;
        RECT 1.760000 0.855000 1.955000 0.860000 ;
        RECT 1.760000 0.860000 1.950000 0.870000 ;
        RECT 1.760000 0.870000 1.945000 0.875000 ;
        RECT 1.760000 0.875000 1.940000 0.880000 ;
        RECT 1.760000 0.880000 1.930000 1.685000 ;
        RECT 1.790000 0.735000 3.235000 0.750000 ;
        RECT 1.805000 0.725000 3.235000 0.735000 ;
        RECT 1.820000 0.715000 3.235000 0.725000 ;
        RECT 1.830000 0.705000 3.235000 0.715000 ;
        RECT 1.840000 0.690000 3.235000 0.705000 ;
        RECT 1.860000 0.655000 3.235000 0.690000 ;
        RECT 1.875000 0.615000 3.235000 0.655000 ;
        RECT 2.455000 0.305000 2.630000 0.615000 ;
        RECT 3.065000 0.785000 3.235000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.420000  0.255000  1.705000 0.585000 ;
      RECT  1.420000  0.585000  1.590000 1.860000 ;
      RECT  1.420000  1.860000  3.230000 2.075000 ;
      RECT  1.420000  2.075000  1.705000 2.445000 ;
      RECT  1.875000  2.245000  2.205000 2.635000 ;
      RECT  1.955000  0.085000  2.285000 0.445000 ;
      RECT  2.100000  0.955000  2.445000 1.125000 ;
      RECT  2.100000  1.125000  2.270000 1.860000 ;
      RECT  2.675000  2.245000  3.570000 2.415000 ;
      RECT  2.800000  0.275000  3.575000 0.445000 ;
      RECT  3.060000  1.355000  3.255000 1.685000 ;
      RECT  3.060000  1.685000  3.230000 1.860000 ;
      RECT  3.400000  1.825000  4.335000 1.995000 ;
      RECT  3.400000  1.995000  3.570000 2.245000 ;
      RECT  3.405000  0.445000  3.575000 0.715000 ;
      RECT  3.405000  0.715000  4.335000 0.885000 ;
      RECT  3.740000  2.165000  3.910000 2.635000 ;
      RECT  3.745000  0.085000  3.945000 0.545000 ;
      RECT  4.165000  0.365000  4.515000 0.535000 ;
      RECT  4.165000  0.535000  4.335000 0.715000 ;
      RECT  4.165000  0.885000  4.335000 1.825000 ;
      RECT  4.165000  1.995000  4.335000 2.070000 ;
      RECT  4.165000  2.070000  4.450000 2.440000 ;
      RECT  4.505000  0.705000  5.085000 1.035000 ;
      RECT  4.505000  1.035000  4.745000 1.905000 ;
      RECT  4.645000  2.190000  5.715000 2.360000 ;
      RECT  4.685000  0.365000  5.425000 0.535000 ;
      RECT  4.935000  1.655000  5.375000 2.010000 ;
      RECT  5.255000  0.535000  5.425000 1.315000 ;
      RECT  5.255000  1.315000  6.055000 1.485000 ;
      RECT  5.545000  1.485000  6.055000 1.575000 ;
      RECT  5.545000  1.575000  5.715000 2.190000 ;
      RECT  5.595000  0.765000  6.395000 1.065000 ;
      RECT  5.595000  1.065000  5.765000 1.095000 ;
      RECT  5.675000  0.085000  6.045000 0.585000 ;
      RECT  5.885000  1.245000  6.055000 1.315000 ;
      RECT  5.885000  1.835000  6.055000 2.635000 ;
      RECT  6.225000  0.365000  6.685000 0.535000 ;
      RECT  6.225000  0.535000  6.395000 0.765000 ;
      RECT  6.225000  1.065000  6.395000 2.135000 ;
      RECT  6.225000  2.135000  6.475000 2.465000 ;
      RECT  6.565000  0.705000  7.115000 1.035000 ;
      RECT  6.565000  1.245000  6.755000 1.965000 ;
      RECT  6.700000  2.165000  7.585000 2.335000 ;
      RECT  6.915000  0.365000  7.455000 0.535000 ;
      RECT  6.925000  1.035000  7.115000 1.575000 ;
      RECT  6.925000  1.575000  7.245000 1.905000 ;
      RECT  7.285000  0.535000  7.455000 0.995000 ;
      RECT  7.285000  0.995000  8.315000 1.325000 ;
      RECT  7.285000  1.325000  7.585000 1.405000 ;
      RECT  7.415000  1.405000  7.585000 2.165000 ;
      RECT  7.700000  0.085000  8.070000 0.615000 ;
      RECT  7.755000  1.575000  8.670000 1.905000 ;
      RECT  7.765000  2.135000  8.070000 2.635000 ;
      RECT  8.340000  0.300000  8.670000 0.825000 ;
      RECT  8.380000  1.905000  8.670000 2.455000 ;
      RECT  8.485000  0.825000  8.670000 0.995000 ;
      RECT  8.485000  0.995000  9.220000 1.325000 ;
      RECT  8.485000  1.325000  8.670000 1.575000 ;
      RECT  8.840000  0.085000  9.010000 0.695000 ;
      RECT  8.840000  1.625000  9.010000 2.635000 ;
      RECT  9.700000  0.345000  9.950000 0.620000 ;
      RECT  9.700000  1.685000 10.030000 2.425000 ;
      RECT  9.780000  0.620000  9.950000 0.995000 ;
      RECT  9.780000  0.995000 10.560000 1.325000 ;
      RECT  9.780000  1.325000 10.030000 1.685000 ;
      RECT 10.185000  0.085000 10.515000 0.805000 ;
      RECT 10.210000  1.495000 10.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.015000  0.765000  1.185000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  0.765000  4.915000 0.935000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.165000  1.785000  5.335000 1.955000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.575000  1.785000  6.745000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  0.765000  6.755000 0.935000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 6.805000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 0.955000 0.735000 1.245000 0.780000 ;
      RECT 0.955000 0.780000 6.815000 0.920000 ;
      RECT 0.955000 0.920000 1.245000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.105000 1.755000 5.395000 1.800000 ;
      RECT 5.105000 1.940000 5.395000 1.985000 ;
      RECT 6.515000 1.755000 6.805000 1.800000 ;
      RECT 6.515000 1.940000 6.805000 1.985000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxbp_1
END LIBRARY

* File: sky130_fd_sc_hd__a22o_4.pxi.spice
* Created: Tue Sep  1 18:53:28 2020
* 
x_PM_SKY130_FD_SC_HD__A22O_4%A_96_21# N_A_96_21#_M1001_s N_A_96_21#_M1014_d
+ N_A_96_21#_M1013_d N_A_96_21#_M1010_d N_A_96_21#_c_111_n N_A_96_21#_M1000_g
+ N_A_96_21#_M1003_g N_A_96_21#_c_112_n N_A_96_21#_M1004_g N_A_96_21#_M1006_g
+ N_A_96_21#_c_113_n N_A_96_21#_M1005_g N_A_96_21#_M1007_g N_A_96_21#_c_114_n
+ N_A_96_21#_M1017_g N_A_96_21#_M1019_g N_A_96_21#_c_115_n N_A_96_21#_c_116_n
+ N_A_96_21#_c_117_n N_A_96_21#_c_118_n N_A_96_21#_c_132_n N_A_96_21#_c_133_n
+ N_A_96_21#_c_144_p N_A_96_21#_c_119_n N_A_96_21#_c_120_n N_A_96_21#_c_121_n
+ N_A_96_21#_c_145_p N_A_96_21#_c_122_n N_A_96_21#_c_123_n N_A_96_21#_c_147_p
+ N_A_96_21#_c_124_n N_A_96_21#_c_125_n N_A_96_21#_c_126_n
+ PM_SKY130_FD_SC_HD__A22O_4%A_96_21#
x_PM_SKY130_FD_SC_HD__A22O_4%B2 N_B2_c_277_n N_B2_M1022_g N_B2_M1013_g
+ N_B2_c_278_n N_B2_M1023_g N_B2_M1021_g N_B2_c_285_n N_B2_c_279_n N_B2_c_280_n
+ B2 N_B2_c_281_n N_B2_c_282_n PM_SKY130_FD_SC_HD__A22O_4%B2
x_PM_SKY130_FD_SC_HD__A22O_4%B1 N_B1_c_362_n N_B1_M1001_g N_B1_M1009_g
+ N_B1_c_363_n N_B1_M1018_g N_B1_M1010_g B1 N_B1_c_365_n
+ PM_SKY130_FD_SC_HD__A22O_4%B1
x_PM_SKY130_FD_SC_HD__A22O_4%A2 N_A2_c_405_n N_A2_M1012_g N_A2_M1002_g
+ N_A2_c_406_n N_A2_M1016_g N_A2_M1008_g N_A2_c_407_n N_A2_c_408_n N_A2_c_417_n
+ N_A2_c_418_n N_A2_c_409_n N_A2_c_410_n A2 N_A2_c_411_n A2
+ PM_SKY130_FD_SC_HD__A22O_4%A2
x_PM_SKY130_FD_SC_HD__A22O_4%A1 N_A1_c_490_n N_A1_M1014_g N_A1_M1011_g
+ N_A1_c_491_n N_A1_M1015_g N_A1_M1020_g A1 N_A1_c_492_n
+ PM_SKY130_FD_SC_HD__A22O_4%A1
x_PM_SKY130_FD_SC_HD__A22O_4%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1019_d
+ N_VPWR_M1002_d N_VPWR_M1020_d N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_536_n
+ N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n
+ N_VPWR_c_542_n N_VPWR_c_543_n VPWR N_VPWR_c_544_n N_VPWR_c_545_n
+ N_VPWR_c_546_n N_VPWR_c_533_n N_VPWR_c_548_n N_VPWR_c_549_n
+ PM_SKY130_FD_SC_HD__A22O_4%VPWR
x_PM_SKY130_FD_SC_HD__A22O_4%X N_X_M1000_d N_X_M1005_d N_X_M1003_s N_X_M1007_s
+ N_X_c_630_n N_X_c_631_n N_X_c_635_n N_X_c_636_n N_X_c_644_n N_X_c_676_n
+ N_X_c_637_n N_X_c_632_n N_X_c_659_n N_X_c_680_n N_X_c_633_n N_X_c_638_n X
+ PM_SKY130_FD_SC_HD__A22O_4%X
x_PM_SKY130_FD_SC_HD__A22O_4%A_484_297# N_A_484_297#_M1013_s
+ N_A_484_297#_M1009_s N_A_484_297#_M1021_s N_A_484_297#_M1011_s
+ N_A_484_297#_M1008_s N_A_484_297#_c_704_n N_A_484_297#_c_708_n
+ N_A_484_297#_c_723_n N_A_484_297#_c_718_n N_A_484_297#_c_748_n
+ N_A_484_297#_c_727_n N_A_484_297#_c_701_n N_A_484_297#_c_753_n
+ N_A_484_297#_c_711_n N_A_484_297#_c_712_n N_A_484_297#_c_733_n
+ PM_SKY130_FD_SC_HD__A22O_4%A_484_297#
x_PM_SKY130_FD_SC_HD__A22O_4%VGND N_VGND_M1000_s N_VGND_M1004_s N_VGND_M1017_s
+ N_VGND_M1023_s N_VGND_M1016_d N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n N_VGND_c_767_n
+ N_VGND_c_768_n N_VGND_c_769_n VGND N_VGND_c_770_n N_VGND_c_771_n
+ N_VGND_c_772_n N_VGND_c_773_n N_VGND_c_774_n PM_SKY130_FD_SC_HD__A22O_4%VGND
x_PM_SKY130_FD_SC_HD__A22O_4%A_566_47# N_A_566_47#_M1022_d N_A_566_47#_M1018_d
+ N_A_566_47#_c_857_n PM_SKY130_FD_SC_HD__A22O_4%A_566_47#
x_PM_SKY130_FD_SC_HD__A22O_4%A_918_47# N_A_918_47#_M1012_s N_A_918_47#_M1015_s
+ N_A_918_47#_c_872_n N_A_918_47#_c_877_n N_A_918_47#_c_870_n
+ PM_SKY130_FD_SC_HD__A22O_4%A_918_47#
cc_1 VNB N_A_96_21#_c_111_n 0.0191784f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_2 VNB N_A_96_21#_c_112_n 0.0157977f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_3 VNB N_A_96_21#_c_113_n 0.0157964f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.995
cc_4 VNB N_A_96_21#_c_114_n 0.0190654f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.995
cc_5 VNB N_A_96_21#_c_115_n 6.30857e-19 $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.175
cc_6 VNB N_A_96_21#_c_116_n 6.59699e-19 $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=1.785
cc_7 VNB N_A_96_21#_c_117_n 0.00475766f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=1.075
cc_8 VNB N_A_96_21#_c_118_n 2.79314e-19 $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=0.82
cc_9 VNB N_A_96_21#_c_119_n 0.00129702f $X=-0.19 $Y=-0.24 $X2=3.475 $Y2=0.775
cc_10 VNB N_A_96_21#_c_120_n 4.62713e-19 $X=-0.19 $Y=-0.24 $X2=3.3 $Y2=0.775
cc_11 VNB N_A_96_21#_c_121_n 0.00424408f $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=1.175
cc_12 VNB N_A_96_21#_c_122_n 0.0119901f $X=-0.19 $Y=-0.24 $X2=3.17 $Y2=0.775
cc_13 VNB N_A_96_21#_c_123_n 4.16442e-19 $X=-0.19 $Y=-0.24 $X2=3.605 $Y2=0.775
cc_14 VNB N_A_96_21#_c_124_n 0.00219468f $X=-0.19 $Y=-0.24 $X2=5.145 $Y2=0.73
cc_15 VNB N_A_96_21#_c_125_n 0.0137328f $X=-0.19 $Y=-0.24 $X2=4.935 $Y2=0.775
cc_16 VNB N_A_96_21#_c_126_n 0.0689431f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.16
cc_17 VNB N_B2_c_277_n 0.0198931f $X=-0.19 $Y=-0.24 $X2=3.25 $Y2=0.235
cc_18 VNB N_B2_c_278_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B2_c_279_n 0.00349181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B2_c_280_n 0.0193014f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_21 VNB N_B2_c_281_n 0.0241314f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_22 VNB N_B2_c_282_n 0.00590555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B1_c_362_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=3.25 $Y2=0.235
cc_24 VNB N_B1_c_363_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB B1 0.00141292f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_26 VNB N_B1_c_365_n 0.0299865f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_27 VNB N_A2_c_405_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=3.25 $Y2=0.235
cc_28 VNB N_A2_c_406_n 0.0218917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A2_c_407_n 0.00358835f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.985
cc_30 VNB N_A2_c_408_n 0.0192902f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.985
cc_31 VNB N_A2_c_409_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.325
cc_32 VNB N_A2_c_410_n 0.00191001f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_33 VNB N_A2_c_411_n 0.0280032f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_34 VNB A2 0.032006f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.995
cc_35 VNB N_A1_c_490_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=3.25 $Y2=0.235
cc_36 VNB N_A1_c_491_n 0.0161504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A1_c_492_n 0.0313079f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_38 VNB N_VPWR_c_533_n 0.269736f $X=-0.19 $Y=-0.24 $X2=4.935 $Y2=0.82
cc_39 VNB N_X_c_630_n 0.0014432f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_40 VNB N_X_c_631_n 0.00986769f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_41 VNB N_X_c_632_n 0.00440603f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_42 VNB N_X_c_633_n 0.00222466f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_43 VNB X 0.0213229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_760_n 0.00419326f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.985
cc_45 VNB N_VGND_c_761_n 0.0169505f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_46 VNB N_VGND_c_762_n 0.0130399f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_47 VNB N_VGND_c_763_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_48 VNB N_VGND_c_764_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_49 VNB N_VGND_c_765_n 0.00668678f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.985
cc_50 VNB N_VGND_c_766_n 0.0365907f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.56
cc_51 VNB N_VGND_c_767_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.56
cc_52 VNB N_VGND_c_768_n 0.0369054f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.985
cc_53 VNB N_VGND_c_769_n 0.00326621f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.985
cc_54 VNB N_VGND_c_770_n 0.0139174f $X=-0.19 $Y=-0.24 $X2=3.385 $Y2=0.775
cc_55 VNB N_VGND_c_771_n 0.324107f $X=-0.19 $Y=-0.24 $X2=3.385 $Y2=0.73
cc_56 VNB N_VGND_c_772_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_773_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=1.96
cc_58 VNB N_VGND_c_774_n 0.0202712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_918_47#_c_870_n 0.00245731f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_60 VPB N_A_96_21#_M1003_g 0.0219695f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_61 VPB N_A_96_21#_M1006_g 0.0181176f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_62 VPB N_A_96_21#_M1007_g 0.0181312f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.985
cc_63 VPB N_A_96_21#_M1019_g 0.0218481f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.985
cc_64 VPB N_A_96_21#_c_116_n 0.00822582f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=1.785
cc_65 VPB N_A_96_21#_c_132_n 0.010722f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.87
cc_66 VPB N_A_96_21#_c_133_n 0.00201536f $X=-0.19 $Y=1.305 $X2=2.23 $Y2=1.87
cc_67 VPB N_A_96_21#_c_126_n 0.0103574f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.16
cc_68 VPB N_B2_M1013_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_B2_M1021_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_70 VPB N_B2_c_285_n 0.00732858f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_71 VPB N_B2_c_279_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_B2_c_280_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.995
cc_73 VPB N_B2_c_281_n 0.00475082f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_74 VPB N_B2_c_282_n 0.00311667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B1_M1009_g 0.0183531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_B1_M1010_g 0.0183545f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_77 VPB N_B1_c_365_n 0.00400363f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_78 VPB N_A2_M1002_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A2_M1008_g 0.0245822f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_80 VPB N_A2_c_407_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_81 VPB N_A2_c_408_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_82 VPB N_A2_c_417_n 0.00789162f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.995
cc_83 VPB N_A2_c_418_n 2.50157e-19 $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_84 VPB N_A2_c_409_n 0.00130531f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.325
cc_85 VPB N_A2_c_411_n 0.00538302f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=0.56
cc_86 VPB N_A1_M1011_g 0.0183373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A1_M1020_g 0.0183337f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_88 VPB N_A1_c_492_n 0.00400351f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_89 VPB N_VPWR_c_534_n 0.0140014f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.325
cc_90 VPB N_VPWR_c_535_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_91 VPB N_VPWR_c_536_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_92 VPB N_VPWR_c_537_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_538_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.325
cc_94 VPB N_VPWR_c_539_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=0.995
cc_95 VPB N_VPWR_c_540_n 0.0584886f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.325
cc_96 VPB N_VPWR_c_541_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.985
cc_97 VPB N_VPWR_c_542_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_543_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.175
cc_99 VPB N_VPWR_c_544_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_100 VPB N_VPWR_c_545_n 0.0163782f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=1.275
cc_101 VPB N_VPWR_c_546_n 0.0241f $X=-0.19 $Y=1.305 $X2=3.385 $Y2=0.73
cc_102 VPB N_VPWR_c_533_n 0.0603204f $X=-0.19 $Y=1.305 $X2=4.935 $Y2=0.82
cc_103 VPB N_VPWR_c_548_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.965 $Y2=1.96
cc_104 VPB N_VPWR_c_549_n 0.0047828f $X=-0.19 $Y=1.305 $X2=3.605 $Y2=0.775
cc_105 VPB N_X_c_635_n 0.00152588f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_106 VPB N_X_c_636_n 0.0124376f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.325
cc_107 VPB N_X_c_637_n 0.00471275f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=0.995
cc_108 VPB N_X_c_638_n 0.00204415f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_109 VPB X 0.00756106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_484_297#_c_701_n 0.00338184f $X=-0.19 $Y=1.305 $X2=1.815
+ $Y2=0.995
cc_111 N_A_96_21#_c_117_n N_B2_c_277_n 0.0024189f $X=2.085 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_96_21#_c_120_n N_B2_c_277_n 4.8408e-19 $X=3.3 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_96_21#_c_122_n N_B2_c_277_n 0.0139498f $X=3.17 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_96_21#_c_116_n N_B2_M1013_g 0.00590249f $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_115 N_A_96_21#_c_132_n N_B2_M1013_g 0.0113813f $X=2.84 $Y=1.87 $X2=0 $Y2=0
cc_116 N_A_96_21#_c_123_n N_B2_c_278_n 4.88987e-19 $X=3.605 $Y=0.775 $X2=0 $Y2=0
cc_117 N_A_96_21#_c_125_n N_B2_c_278_n 0.0122419f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_118 N_A_96_21#_M1013_d N_B2_c_285_n 0.00124334f $X=2.83 $Y=1.485 $X2=0 $Y2=0
cc_119 N_A_96_21#_M1010_d N_B2_c_285_n 0.00164852f $X=3.67 $Y=1.485 $X2=0 $Y2=0
cc_120 N_A_96_21#_c_144_p N_B2_c_285_n 0.0315971f $X=3.68 $Y=1.87 $X2=0 $Y2=0
cc_121 N_A_96_21#_c_145_p N_B2_c_285_n 0.00677369f $X=2.965 $Y=1.87 $X2=0 $Y2=0
cc_122 N_A_96_21#_c_122_n N_B2_c_285_n 0.0112883f $X=3.17 $Y=0.775 $X2=0 $Y2=0
cc_123 N_A_96_21#_c_147_p N_B2_c_285_n 0.0122128f $X=3.805 $Y=1.87 $X2=0 $Y2=0
cc_124 N_A_96_21#_c_125_n N_B2_c_279_n 0.0254297f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_125 N_A_96_21#_c_125_n N_B2_c_280_n 0.00295599f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_126 N_A_96_21#_c_116_n N_B2_c_281_n 2.32165e-19 $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_127 N_A_96_21#_c_117_n N_B2_c_281_n 0.00245123f $X=2.085 $Y=1.075 $X2=0 $Y2=0
cc_128 N_A_96_21#_c_121_n N_B2_c_281_n 0.00100933f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_129 N_A_96_21#_c_122_n N_B2_c_281_n 0.00295599f $X=3.17 $Y=0.775 $X2=0 $Y2=0
cc_130 N_A_96_21#_M1013_d N_B2_c_282_n 0.00104582f $X=2.83 $Y=1.485 $X2=0 $Y2=0
cc_131 N_A_96_21#_c_116_n N_B2_c_282_n 0.0269082f $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_132 N_A_96_21#_c_132_n N_B2_c_282_n 0.0273041f $X=2.84 $Y=1.87 $X2=0 $Y2=0
cc_133 N_A_96_21#_c_121_n N_B2_c_282_n 0.0169378f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_134 N_A_96_21#_c_145_p N_B2_c_282_n 0.00564423f $X=2.965 $Y=1.87 $X2=0 $Y2=0
cc_135 N_A_96_21#_c_122_n N_B2_c_282_n 0.0424183f $X=3.17 $Y=0.775 $X2=0 $Y2=0
cc_136 N_A_96_21#_c_126_n N_B2_c_282_n 0.00131745f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_96_21#_c_120_n N_B1_c_362_n 0.00570524f $X=3.3 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_96_21#_c_122_n N_B1_c_362_n 0.00541406f $X=3.17 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_139 N_A_96_21#_c_144_p N_B1_M1009_g 0.00924026f $X=3.68 $Y=1.87 $X2=0 $Y2=0
cc_140 N_A_96_21#_c_123_n N_B1_c_363_n 0.00595698f $X=3.605 $Y=0.775 $X2=0 $Y2=0
cc_141 N_A_96_21#_c_125_n N_B1_c_363_n 0.00487822f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_142 N_A_96_21#_c_144_p N_B1_M1010_g 0.00924026f $X=3.68 $Y=1.87 $X2=0 $Y2=0
cc_143 N_A_96_21#_c_122_n B1 0.0400898f $X=3.17 $Y=0.775 $X2=0 $Y2=0
cc_144 N_A_96_21#_c_119_n N_B1_c_365_n 0.00224214f $X=3.475 $Y=0.775 $X2=0 $Y2=0
cc_145 N_A_96_21#_c_124_n N_A2_c_405_n 4.80264e-19 $X=5.145 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_96_21#_c_125_n N_A2_c_405_n 0.0122419f $X=4.935 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_96_21#_c_125_n N_A2_c_407_n 0.0254297f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_148 N_A_96_21#_c_125_n N_A2_c_408_n 0.00295599f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_149 N_A_96_21#_c_125_n N_A2_c_417_n 0.0071189f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_150 N_A_96_21#_c_124_n N_A1_c_490_n 0.0054298f $X=5.145 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_96_21#_c_125_n N_A1_c_490_n 0.00582863f $X=4.935 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_96_21#_c_124_n N_A1_c_491_n 0.00381649f $X=5.145 $Y=0.73 $X2=0 $Y2=0
cc_153 N_A_96_21#_c_125_n A1 0.0300382f $X=4.935 $Y=0.775 $X2=0 $Y2=0
cc_154 N_A_96_21#_c_124_n N_A1_c_492_n 0.00224214f $X=5.145 $Y=0.73 $X2=0 $Y2=0
cc_155 N_A_96_21#_c_116_n N_VPWR_M1019_d 0.0033596f $X=2.065 $Y=1.785 $X2=0
+ $Y2=0
cc_156 N_A_96_21#_c_133_n N_VPWR_M1019_d 0.00410134f $X=2.23 $Y=1.87 $X2=0 $Y2=0
cc_157 N_A_96_21#_M1003_g N_VPWR_c_535_n 0.00338128f $X=0.555 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_96_21#_M1006_g N_VPWR_c_536_n 0.00157837f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_96_21#_M1007_g N_VPWR_c_536_n 0.00157837f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_96_21#_M1019_g N_VPWR_c_537_n 0.00338128f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_96_21#_c_133_n N_VPWR_c_537_n 0.0176408f $X=2.23 $Y=1.87 $X2=0 $Y2=0
cc_162 N_A_96_21#_M1003_g N_VPWR_c_544_n 0.00585385f $X=0.555 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_96_21#_M1006_g N_VPWR_c_544_n 0.00585385f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_96_21#_M1007_g N_VPWR_c_545_n 0.00585385f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_96_21#_M1019_g N_VPWR_c_545_n 0.00585385f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_96_21#_M1013_d N_VPWR_c_533_n 0.00215227f $X=2.83 $Y=1.485 $X2=0
+ $Y2=0
cc_167 N_A_96_21#_M1010_d N_VPWR_c_533_n 0.0021603f $X=3.67 $Y=1.485 $X2=0 $Y2=0
cc_168 N_A_96_21#_M1003_g N_VPWR_c_533_n 0.0114631f $X=0.555 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_96_21#_M1006_g N_VPWR_c_533_n 0.0104367f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_96_21#_M1007_g N_VPWR_c_533_n 0.0104367f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_96_21#_M1019_g N_VPWR_c_533_n 0.0117628f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_96_21#_c_132_n N_VPWR_c_533_n 0.00780718f $X=2.84 $Y=1.87 $X2=0 $Y2=0
cc_173 N_A_96_21#_c_133_n N_VPWR_c_533_n 0.00435471f $X=2.23 $Y=1.87 $X2=0 $Y2=0
cc_174 N_A_96_21#_c_144_p N_VPWR_c_533_n 0.00127799f $X=3.68 $Y=1.87 $X2=0 $Y2=0
cc_175 N_A_96_21#_c_111_n N_X_c_630_n 0.0111411f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_96_21#_c_115_n N_X_c_630_n 0.00410208f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_177 N_A_96_21#_M1003_g N_X_c_635_n 0.015729f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_96_21#_c_115_n N_X_c_635_n 0.00686379f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_179 N_A_96_21#_c_111_n N_X_c_644_n 0.0108342f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_96_21#_c_112_n N_X_c_644_n 0.00621819f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_96_21#_c_113_n N_X_c_644_n 5.19281e-19 $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_96_21#_M1006_g N_X_c_637_n 0.0133439f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_96_21#_M1007_g N_X_c_637_n 0.0133089f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_96_21#_M1019_g N_X_c_637_n 3.45391e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_96_21#_c_115_n N_X_c_637_n 0.0618991f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_186 N_A_96_21#_c_116_n N_X_c_637_n 0.00344747f $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_187 N_A_96_21#_c_126_n N_X_c_637_n 0.00436768f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_96_21#_c_112_n N_X_c_632_n 0.00870364f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_96_21#_c_113_n N_X_c_632_n 0.0098365f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_96_21#_c_114_n N_X_c_632_n 0.00298809f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_96_21#_c_115_n N_X_c_632_n 0.0626515f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_192 N_A_96_21#_c_118_n N_X_c_632_n 0.00808484f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_193 N_A_96_21#_c_126_n N_X_c_632_n 0.00452472f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_96_21#_c_112_n N_X_c_659_n 5.22228e-19 $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_96_21#_c_113_n N_X_c_659_n 0.00630972f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_96_21#_c_114_n N_X_c_659_n 0.0109565f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_96_21#_c_111_n N_X_c_633_n 0.00113258f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_96_21#_c_112_n N_X_c_633_n 0.00113258f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_96_21#_c_115_n N_X_c_633_n 0.0265057f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_200 N_A_96_21#_c_126_n N_X_c_633_n 0.00230227f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_96_21#_c_115_n N_X_c_638_n 0.0203891f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_202 N_A_96_21#_c_126_n N_X_c_638_n 0.00222737f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_96_21#_c_111_n X 0.0198998f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_96_21#_c_115_n X 0.0164324f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_205 N_A_96_21#_c_132_n N_A_484_297#_M1013_s 0.00496426f $X=2.84 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_206 N_A_96_21#_c_144_p N_A_484_297#_M1009_s 0.00317012f $X=3.68 $Y=1.87 $X2=0
+ $Y2=0
cc_207 N_A_96_21#_M1013_d N_A_484_297#_c_704_n 0.00310345f $X=2.83 $Y=1.485
+ $X2=0 $Y2=0
cc_208 N_A_96_21#_c_132_n N_A_484_297#_c_704_n 0.00506389f $X=2.84 $Y=1.87 $X2=0
+ $Y2=0
cc_209 N_A_96_21#_c_144_p N_A_484_297#_c_704_n 0.00506389f $X=3.68 $Y=1.87 $X2=0
+ $Y2=0
cc_210 N_A_96_21#_c_145_p N_A_484_297#_c_704_n 0.0112088f $X=2.965 $Y=1.87 $X2=0
+ $Y2=0
cc_211 N_A_96_21#_M1010_d N_A_484_297#_c_708_n 0.00312348f $X=3.67 $Y=1.485
+ $X2=0 $Y2=0
cc_212 N_A_96_21#_c_144_p N_A_484_297#_c_708_n 0.00506389f $X=3.68 $Y=1.87 $X2=0
+ $Y2=0
cc_213 N_A_96_21#_c_147_p N_A_484_297#_c_708_n 0.0112811f $X=3.805 $Y=1.87 $X2=0
+ $Y2=0
cc_214 N_A_96_21#_c_132_n N_A_484_297#_c_711_n 0.0150802f $X=2.84 $Y=1.87 $X2=0
+ $Y2=0
cc_215 N_A_96_21#_c_144_p N_A_484_297#_c_712_n 0.0116461f $X=3.68 $Y=1.87 $X2=0
+ $Y2=0
cc_216 N_A_96_21#_c_118_n N_VGND_M1017_s 0.00546399f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_217 N_A_96_21#_c_122_n N_VGND_M1017_s 0.00639474f $X=3.17 $Y=0.775 $X2=0
+ $Y2=0
cc_218 N_A_96_21#_c_125_n N_VGND_M1023_s 0.00306523f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_219 N_A_96_21#_c_111_n N_VGND_c_760_n 0.00316354f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_96_21#_c_111_n N_VGND_c_761_n 0.00423737f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_96_21#_c_112_n N_VGND_c_761_n 0.00423737f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_96_21#_c_112_n N_VGND_c_763_n 0.00146448f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_96_21#_c_113_n N_VGND_c_763_n 0.00146339f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_96_21#_c_125_n N_VGND_c_764_n 0.0125492f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_225 N_A_96_21#_c_122_n N_VGND_c_766_n 0.00194318f $X=3.17 $Y=0.775 $X2=0
+ $Y2=0
cc_226 N_A_96_21#_c_125_n N_VGND_c_766_n 0.0025354f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_227 N_A_96_21#_c_125_n N_VGND_c_768_n 0.00239348f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_228 N_A_96_21#_M1001_s N_VGND_c_771_n 0.00216833f $X=3.25 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_96_21#_M1014_d N_VGND_c_771_n 0.00216833f $X=5.01 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_A_96_21#_c_111_n N_VGND_c_771_n 0.00674307f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_96_21#_c_112_n N_VGND_c_771_n 0.00571669f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_96_21#_c_113_n N_VGND_c_771_n 0.0057163f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_96_21#_c_114_n N_VGND_c_771_n 0.0108251f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_96_21#_c_118_n N_VGND_c_771_n 0.00127084f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_235 N_A_96_21#_c_122_n N_VGND_c_771_n 0.00619164f $X=3.17 $Y=0.775 $X2=0
+ $Y2=0
cc_236 N_A_96_21#_c_125_n N_VGND_c_771_n 0.0121714f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_237 N_A_96_21#_c_113_n N_VGND_c_773_n 0.00423334f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_96_21#_c_114_n N_VGND_c_773_n 0.00541359f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_96_21#_c_114_n N_VGND_c_774_n 0.00335921f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_96_21#_c_118_n N_VGND_c_774_n 0.0232224f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_241 N_A_96_21#_c_122_n N_VGND_c_774_n 0.0291799f $X=3.17 $Y=0.775 $X2=0 $Y2=0
cc_242 N_A_96_21#_c_122_n N_A_566_47#_M1022_d 0.00195168f $X=3.17 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_243 N_A_96_21#_c_125_n N_A_566_47#_M1018_d 0.00195168f $X=4.935 $Y=0.775
+ $X2=0 $Y2=0
cc_244 N_A_96_21#_M1001_s N_A_566_47#_c_857_n 0.00305026f $X=3.25 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_96_21#_c_120_n N_A_566_47#_c_857_n 0.0224636f $X=3.3 $Y=0.775 $X2=0
+ $Y2=0
cc_246 N_A_96_21#_c_122_n N_A_566_47#_c_857_n 0.0121378f $X=3.17 $Y=0.775 $X2=0
+ $Y2=0
cc_247 N_A_96_21#_c_125_n N_A_566_47#_c_857_n 0.011913f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_248 N_A_96_21#_c_125_n N_A_918_47#_M1012_s 0.00195168f $X=4.935 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_249 N_A_96_21#_M1014_d N_A_918_47#_c_872_n 0.00305026f $X=5.01 $Y=0.235 $X2=0
+ $Y2=0
cc_250 N_A_96_21#_c_124_n N_A_918_47#_c_872_n 0.0183915f $X=5.145 $Y=0.73 $X2=0
+ $Y2=0
cc_251 N_A_96_21#_c_125_n N_A_918_47#_c_872_n 0.0123626f $X=4.935 $Y=0.775 $X2=0
+ $Y2=0
cc_252 N_A_96_21#_c_124_n N_A_918_47#_c_870_n 0.0105248f $X=5.145 $Y=0.73 $X2=0
+ $Y2=0
cc_253 N_B2_c_277_n N_B1_c_362_n 0.0268717f $X=2.755 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_254 N_B2_M1013_g N_B1_M1009_g 0.0428045f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B2_c_285_n N_B1_M1009_g 0.00991308f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_256 N_B2_c_278_n N_B1_c_363_n 0.0268673f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B2_M1021_g N_B1_M1010_g 0.0428494f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B2_c_285_n N_B1_M1010_g 0.0102793f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_259 N_B2_c_285_n B1 0.0391837f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_260 N_B2_c_279_n B1 0.0172311f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B2_c_280_n B1 6.66616e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_262 N_B2_c_281_n B1 2.07818e-19 $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B2_c_282_n B1 0.0169874f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B2_c_285_n N_B1_c_365_n 0.00214031f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_265 N_B2_c_279_n N_B1_c_365_n 0.00458063f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B2_c_280_n N_B1_c_365_n 0.0223771f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B2_c_281_n N_B1_c_365_n 0.0223106f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B2_c_282_n N_B1_c_365_n 0.00592594f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B2_c_278_n N_A2_c_405_n 0.0207366f $X=4.015 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_270 N_B2_M1021_g N_A2_M1002_g 0.02101f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B2_c_285_n N_A2_M1002_g 5.77655e-19 $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_272 N_B2_c_279_n N_A2_M1002_g 3.59226e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B2_M1021_g N_A2_c_407_n 3.59226e-19 $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B2_c_279_n N_A2_c_407_n 0.0307171f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_275 N_B2_c_280_n N_A2_c_407_n 7.80994e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B2_c_279_n N_A2_c_408_n 7.80994e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_277 N_B2_c_280_n N_A2_c_408_n 0.0197715f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_278 N_B2_M1021_g N_A2_c_418_n 5.77655e-19 $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B2_c_285_n N_A2_c_418_n 0.0154679f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_280 N_B2_M1013_g N_VPWR_c_537_n 0.00214938f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B2_M1013_g N_VPWR_c_540_n 0.00357877f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B2_M1021_g N_VPWR_c_540_n 0.00357877f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_283 N_B2_M1013_g N_VPWR_c_533_n 0.00657948f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B2_M1021_g N_VPWR_c_533_n 0.00546478f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B2_c_282_n N_A_484_297#_M1013_s 0.00407272f $X=2.755 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_286 N_B2_c_285_n N_A_484_297#_M1009_s 0.00166235f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_287 N_B2_c_285_n N_A_484_297#_M1021_s 0.00151125f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_288 N_B2_M1013_g N_A_484_297#_c_704_n 0.00851673f $X=2.755 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_B2_M1021_g N_A_484_297#_c_708_n 0.0121306f $X=4.015 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_B2_c_285_n N_A_484_297#_c_718_n 0.00292685f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_291 N_B2_c_278_n N_VGND_c_764_n 0.00512705f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_277_n N_VGND_c_766_n 0.0042294f $X=2.755 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B2_c_278_n N_VGND_c_766_n 0.0042294f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B2_c_277_n N_VGND_c_771_n 0.00709599f $X=2.755 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B2_c_278_n N_VGND_c_771_n 0.00609665f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B2_c_277_n N_VGND_c_774_n 0.00481673f $X=2.755 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B2_c_277_n N_A_566_47#_c_857_n 0.00315446f $X=2.755 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_B2_c_278_n N_A_566_47#_c_857_n 0.00329629f $X=4.015 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_B1_M1009_g N_VPWR_c_540_n 0.00357877f $X=3.175 $Y=1.985 $X2=0 $Y2=0
cc_300 N_B1_M1010_g N_VPWR_c_540_n 0.00357877f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_301 N_B1_M1009_g N_VPWR_c_533_n 0.00525341f $X=3.175 $Y=1.985 $X2=0 $Y2=0
cc_302 N_B1_M1010_g N_VPWR_c_533_n 0.00525341f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_303 N_B1_M1009_g N_A_484_297#_c_704_n 0.00851673f $X=3.175 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_B1_M1010_g N_A_484_297#_c_708_n 0.00851673f $X=3.595 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_B1_c_362_n N_VGND_c_766_n 0.00357877f $X=3.175 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B1_c_363_n N_VGND_c_766_n 0.00357877f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_c_362_n N_VGND_c_771_n 0.00525237f $X=3.175 $Y=0.995 $X2=0 $Y2=0
cc_308 N_B1_c_363_n N_VGND_c_771_n 0.00525237f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B1_c_362_n N_A_566_47#_c_857_n 0.00917157f $X=3.175 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_B1_c_363_n N_A_566_47#_c_857_n 0.00915387f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_A2_c_405_n N_A1_c_490_n 0.0268761f $X=4.515 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_312 N_A2_M1002_g N_A1_M1011_g 0.0432836f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A2_c_417_n N_A1_M1011_g 0.0108086f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_314 N_A2_c_406_n N_A1_c_491_n 0.012379f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_M1008_g N_A1_M1020_g 0.042557f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A2_c_417_n N_A1_M1020_g 0.0113924f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_317 N_A2_c_407_n A1 0.0133594f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A2_c_408_n A1 2.2122e-19 $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A2_c_417_n A1 0.0349894f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_320 N_A2_c_410_n A1 0.0172564f $X=5.735 $Y=1.175 $X2=0 $Y2=0
cc_321 N_A2_c_411_n A1 2.00336e-19 $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A2_c_407_n N_A1_c_492_n 0.00527477f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A2_c_408_n N_A1_c_492_n 0.022397f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A2_c_417_n N_A1_c_492_n 0.00214031f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_325 N_A2_c_409_n N_A1_c_492_n 0.00362491f $X=5.65 $Y=1.445 $X2=0 $Y2=0
cc_326 N_A2_c_410_n N_A1_c_492_n 0.00144374f $X=5.735 $Y=1.175 $X2=0 $Y2=0
cc_327 N_A2_c_411_n N_A1_c_492_n 0.0222902f $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A2_c_417_n N_VPWR_M1002_d 0.00130005f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_329 N_A2_c_418_n N_VPWR_M1002_d 3.52503e-19 $X=4.68 $Y=1.53 $X2=0 $Y2=0
cc_330 N_A2_c_417_n N_VPWR_M1020_d 0.00167975f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_331 N_A2_M1002_g N_VPWR_c_538_n 0.00302074f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A2_M1008_g N_VPWR_c_539_n 0.00302074f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A2_M1002_g N_VPWR_c_540_n 0.00585385f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A2_M1008_g N_VPWR_c_546_n 0.00585385f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A2_M1002_g N_VPWR_c_533_n 0.0061234f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A2_M1008_g N_VPWR_c_533_n 0.00700792f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A2_c_418_n N_A_484_297#_M1021_s 0.00151125f $X=4.68 $Y=1.53 $X2=0 $Y2=0
cc_338 N_A2_c_417_n N_A_484_297#_M1011_s 0.00165831f $X=5.565 $Y=1.53 $X2=0
+ $Y2=0
cc_339 N_A2_M1002_g N_A_484_297#_c_723_n 0.0095558f $X=4.515 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A2_c_417_n N_A_484_297#_c_723_n 0.0190307f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_341 N_A2_c_418_n N_A_484_297#_c_723_n 0.013811f $X=4.68 $Y=1.53 $X2=0 $Y2=0
cc_342 N_A2_c_418_n N_A_484_297#_c_718_n 0.00292685f $X=4.68 $Y=1.53 $X2=0 $Y2=0
cc_343 N_A2_M1008_g N_A_484_297#_c_727_n 0.01084f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A2_c_417_n N_A_484_297#_c_727_n 0.0245652f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_345 A2 N_A_484_297#_c_727_n 0.00397033f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_346 N_A2_M1008_g N_A_484_297#_c_701_n 6.58332e-19 $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_347 N_A2_c_417_n N_A_484_297#_c_701_n 0.00786716f $X=5.565 $Y=1.53 $X2=0
+ $Y2=0
cc_348 A2 N_A_484_297#_c_701_n 0.0166332f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_349 N_A2_c_417_n N_A_484_297#_c_733_n 0.0126919f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_350 N_A2_c_405_n N_VGND_c_764_n 0.00518302f $X=4.515 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A2_c_406_n N_VGND_c_765_n 0.00460417f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A2_c_411_n N_VGND_c_765_n 2.29969e-19 $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_353 A2 N_VGND_c_765_n 0.0137431f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_354 N_A2_c_405_n N_VGND_c_768_n 0.0042294f $X=4.515 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A2_c_406_n N_VGND_c_768_n 0.00539841f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_356 N_A2_c_405_n N_VGND_c_771_n 0.00607156f $X=4.515 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A2_c_406_n N_VGND_c_771_n 0.0105876f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A2_c_405_n N_A_918_47#_c_872_n 0.00324504f $X=4.515 $Y=0.995 $X2=0
+ $Y2=0
cc_359 N_A2_c_406_n N_A_918_47#_c_877_n 0.00266812f $X=5.775 $Y=0.995 $X2=0
+ $Y2=0
cc_360 N_A2_c_406_n N_A_918_47#_c_870_n 0.00511693f $X=5.775 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A2_c_417_n N_A_918_47#_c_870_n 0.00310205f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_362 N_A2_c_410_n N_A_918_47#_c_870_n 0.0139065f $X=5.735 $Y=1.175 $X2=0 $Y2=0
cc_363 N_A2_c_411_n N_A_918_47#_c_870_n 0.00152613f $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_364 N_A1_M1011_g N_VPWR_c_538_n 0.00157837f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A1_M1020_g N_VPWR_c_539_n 0.00157837f $X=5.355 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A1_M1011_g N_VPWR_c_542_n 0.00585385f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A1_M1020_g N_VPWR_c_542_n 0.00585385f $X=5.355 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A1_M1011_g N_VPWR_c_533_n 0.00591203f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A1_M1020_g N_VPWR_c_533_n 0.00591203f $X=5.355 $Y=1.985 $X2=0 $Y2=0
cc_370 N_A1_M1011_g N_A_484_297#_c_723_n 0.00956194f $X=4.935 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_A1_M1020_g N_A_484_297#_c_727_n 0.00956194f $X=5.355 $Y=1.985 $X2=0
+ $Y2=0
cc_372 N_A1_c_490_n N_VGND_c_768_n 0.00357877f $X=4.935 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A1_c_491_n N_VGND_c_768_n 0.00357877f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A1_c_490_n N_VGND_c_771_n 0.00525237f $X=4.935 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A1_c_491_n N_VGND_c_771_n 0.00525237f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A1_c_490_n N_A_918_47#_c_872_n 0.00918928f $X=4.935 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A1_c_491_n N_A_918_47#_c_872_n 0.0111772f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_378 A1 N_A_918_47#_c_872_n 0.00209698f $X=5.225 $Y=1.105 $X2=0 $Y2=0
cc_379 N_VPWR_c_533_n N_X_M1003_s 0.00284632f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_c_533_n N_X_M1007_s 0.00284632f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_M1003_d N_X_c_635_n 6.05749e-19 $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_382 N_VPWR_c_535_n N_X_c_635_n 0.00365338f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_383 N_VPWR_M1003_d N_X_c_636_n 0.00347536f $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_384 N_VPWR_c_535_n N_X_c_636_n 0.011469f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_385 N_VPWR_c_544_n N_X_c_676_n 0.0142343f $X=1.06 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_c_533_n N_X_c_676_n 0.00955092f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_M1006_d N_X_c_637_n 0.00169858f $X=1.05 $Y=1.485 $X2=0 $Y2=0
cc_388 N_VPWR_c_536_n N_X_c_637_n 0.0121607f $X=1.185 $Y=1.99 $X2=0 $Y2=0
cc_389 N_VPWR_c_545_n N_X_c_680_n 0.0142343f $X=1.9 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_533_n N_X_c_680_n 0.00955092f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_533_n N_A_484_297#_M1013_s 0.00207714f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_392 N_VPWR_c_533_n N_A_484_297#_M1009_s 0.00213597f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_533_n N_A_484_297#_M1021_s 0.00284453f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_533_n N_A_484_297#_M1011_s 0.00223619f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_533_n N_A_484_297#_M1008_s 0.00349344f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_540_n N_A_484_297#_c_704_n 0.0329893f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_533_n N_A_484_297#_c_704_n 0.0204667f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_540_n N_A_484_297#_c_708_n 0.0529483f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_533_n N_A_484_297#_c_708_n 0.0331756f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_M1002_d N_A_484_297#_c_723_n 0.00325521f $X=4.59 $Y=1.485 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_538_n N_A_484_297#_c_723_n 0.0123301f $X=4.725 $Y=2.3 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_533_n N_A_484_297#_c_723_n 0.0109281f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_542_n N_A_484_297#_c_748_n 0.0142343f $X=5.44 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_533_n N_A_484_297#_c_748_n 0.00955092f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_M1020_d N_A_484_297#_c_727_n 0.00325404f $X=5.43 $Y=1.485 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_539_n N_A_484_297#_c_727_n 0.0123301f $X=5.565 $Y=2.3 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_533_n N_A_484_297#_c_727_n 0.012579f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_546_n N_A_484_297#_c_753_n 0.0142403f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_533_n N_A_484_297#_c_753_n 0.00781266f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_537_n N_A_484_297#_c_711_n 0.0186128f $X=2.025 $Y=2.3 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_540_n N_A_484_297#_c_711_n 0.0151494f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_533_n N_A_484_297#_c_711_n 0.00938745f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_540_n N_A_484_297#_c_712_n 0.0137033f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_533_n N_A_484_297#_c_712_n 0.00938745f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_X_c_630_n N_VGND_M1000_s 5.40298e-19 $X=0.6 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_416 N_X_c_631_n N_VGND_M1000_s 0.00329182f $X=0.37 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_417 N_X_c_632_n N_VGND_M1004_s 0.00162089f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_418 N_X_c_630_n N_VGND_c_760_n 0.00402428f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_419 N_X_c_631_n N_VGND_c_760_n 0.00920832f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_420 N_X_c_644_n N_VGND_c_761_n 0.017716f $X=0.765 $Y=0.39 $X2=0 $Y2=0
cc_421 N_X_c_632_n N_VGND_c_761_n 0.00198695f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_422 N_X_c_630_n N_VGND_c_762_n 0.0019947f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_423 N_X_c_631_n N_VGND_c_762_n 0.00293744f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_424 N_X_c_632_n N_VGND_c_763_n 0.0122559f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_425 N_X_M1000_d N_VGND_c_771_n 0.00215535f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_426 N_X_M1005_d N_VGND_c_771_n 0.00215201f $X=1.47 $Y=0.235 $X2=0 $Y2=0
cc_427 N_X_c_630_n N_VGND_c_771_n 0.00407016f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_428 N_X_c_631_n N_VGND_c_771_n 0.00542613f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_429 N_X_c_644_n N_VGND_c_771_n 0.0121406f $X=0.765 $Y=0.39 $X2=0 $Y2=0
cc_430 N_X_c_632_n N_VGND_c_771_n 0.00835832f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_431 N_X_c_659_n N_VGND_c_771_n 0.0122069f $X=1.605 $Y=0.39 $X2=0 $Y2=0
cc_432 N_X_c_632_n N_VGND_c_773_n 0.00198695f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_433 N_X_c_659_n N_VGND_c_773_n 0.0188551f $X=1.605 $Y=0.39 $X2=0 $Y2=0
cc_434 N_VGND_c_771_n N_A_566_47#_M1022_d 0.00215227f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_435 N_VGND_c_771_n N_A_566_47#_M1018_d 0.00215227f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_764_n N_A_566_47#_c_857_n 0.0142796f $X=4.27 $Y=0.39 $X2=0 $Y2=0
cc_437 N_VGND_c_766_n N_A_566_47#_c_857_n 0.0646671f $X=4.185 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_771_n N_A_566_47#_c_857_n 0.0418989f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_771_n N_A_918_47#_M1012_s 0.00215227f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_440 N_VGND_c_771_n N_A_918_47#_M1015_s 0.00215206f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_c_764_n N_A_918_47#_c_872_n 0.014815f $X=4.27 $Y=0.39 $X2=0 $Y2=0
cc_442 N_VGND_c_768_n N_A_918_47#_c_872_n 0.0504977f $X=5.9 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_771_n N_A_918_47#_c_872_n 0.0327385f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_c_768_n N_A_918_47#_c_877_n 0.0151965f $X=5.9 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_771_n N_A_918_47#_c_877_n 0.00940324f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_765_n N_A_918_47#_c_870_n 0.0154056f $X=5.985 $Y=0.39 $X2=0
+ $Y2=0

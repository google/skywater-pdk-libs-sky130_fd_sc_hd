* File: sky130_fd_sc_hd__clkbuf_1.spice
* Created: Tue Sep  1 19:00:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkbuf_1.pex.spice"
.subckt sky130_fd_sc_hd__clkbuf_1  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_75_212#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0754 AS=0.1352 PD=0.81 PS=1.56 NRD=1.152 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1001 N_A_75_212#_M1001_d N_A_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0754 PD=1.56 PS=0.81 NRD=0 NRS=1.152 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_VPWR_M1000_d N_A_75_212#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.79
+ AD=0.11455 AS=0.2054 PD=1.08 PS=2.1 NRD=1.2411 NRS=0 M=1 R=5.26667 SA=75000.2
+ SB=75000.6 A=0.1185 P=1.88 MULT=1
MM1002 N_A_75_212#_M1002_d N_A_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.79
+ AD=0.2054 AS=0.11455 PD=2.1 PS=1.08 NRD=0 NRS=1.2411 M=1 R=5.26667 SA=75000.6
+ SB=75000.2 A=0.1185 P=1.88 MULT=1
DX4_noxref VNB VPB NWDIODE A=2.8248 P=6.73
*
.include "sky130_fd_sc_hd__clkbuf_1.pxi.spice"
*
.ends
*
*

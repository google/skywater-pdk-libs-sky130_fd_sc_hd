* File: sky130_fd_sc_hd__sdfxtp_2.pex.spice
* Created: Thu Aug 27 14:47:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%CLK 1 2 3 5 6 8 11 13 14
c42 1 0 2.71124e-20 $X=0.31 $Y=1.325
r43 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.16 $X2=0.27
+ $Y2=1.53
r44 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r45 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.475 $Y2=1.665
r46 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=1.665
r47 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=2.135
r48 3 18 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r49 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r50 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r51 1 18 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r52 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_27_47# 1 2 9 13 17 19 20 25 29 31 35 39
+ 43 44 45 49 50 52 55 56 57 58 59 60 69 75 78 79 80 82 86
c247 86 0 1.77381e-19 $X=6.695 $Y=1.41
c248 52 0 8.70797e-20 $X=0.76 $Y=1.235
c249 50 0 1.81794e-19 $X=0.73 $Y=1.795
c250 45 0 3.29888e-20 $X=0.615 $Y=1.88
c251 29 0 4.21632e-20 $X=6.7 $Y=2.275
c252 19 0 1.57835e-19 $X=5.01 $Y=1.32
r253 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.41
+ $X2=6.695 $Y2=1.575
r254 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.695
+ $Y=1.41 $X2=6.695 $Y2=1.41
r255 82 85 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.695 $Y=1.32
+ $X2=6.695 $Y2=1.41
r256 78 81 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.74
+ $X2=5.145 $Y2=1.905
r257 78 80 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.74
+ $X2=5.145 $Y2=1.575
r258 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=1.74 $X2=5.145 $Y2=1.74
r259 74 75 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=0.89 $Y=1.235
+ $X2=0.895 $Y2=1.235
r260 70 86 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.705 $Y=1.87
+ $X2=6.705 $Y2=1.41
r261 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.705 $Y=1.87
+ $X2=6.705 $Y2=1.87
r262 66 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r263 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=1.87
+ $X2=0.725 $Y2=1.87
r264 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r265 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.56 $Y=1.87
+ $X2=6.705 $Y2=1.87
r266 59 60 1.39232 $w=1.4e-07 $l=1.125e-06 $layer=MET1_cond $X=6.56 $Y=1.87
+ $X2=5.435 $Y2=1.87
r267 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.87 $Y=1.87
+ $X2=0.725 $Y2=1.87
r268 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r269 57 58 5.29083 $w=1.4e-07 $l=4.275e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=0.87 $Y2=1.87
r270 53 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r271 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r272 50 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r273 50 52 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r274 49 56 6.0623 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=0.97
r275 49 52 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=1.235
r276 47 56 9.38461 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=0.805
+ $X2=0.712 $Y2=0.97
r277 46 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r278 45 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r279 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.35 $Y2=1.88
r280 43 47 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.712 $Y2=0.805
r281 43 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r282 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r283 37 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r284 33 35 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.345 $Y=1.245
+ $X2=7.345 $Y2=0.415
r285 32 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.83 $Y=1.32
+ $X2=6.695 $Y2=1.32
r286 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.27 $Y=1.32
+ $X2=7.345 $Y2=1.245
r287 31 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.27 $Y=1.32
+ $X2=6.83 $Y2=1.32
r288 29 87 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.7 $Y=2.275 $X2=6.7
+ $Y2=1.575
r289 25 81 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.085 $Y=2.275
+ $X2=5.085 $Y2=1.905
r290 21 80 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.085 $Y=1.395
+ $X2=5.085 $Y2=1.575
r291 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.01 $Y=1.32
+ $X2=5.085 $Y2=1.395
r292 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=5.01 $Y=1.32
+ $X2=4.7 $Y2=1.32
r293 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.625 $Y=1.245
+ $X2=4.7 $Y2=1.32
r294 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.625 $Y=1.245
+ $X2=4.625 $Y2=0.415
r295 11 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=1.235
r296 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=2.135
r297 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r298 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r299 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r300 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%SCE 3 9 11 15 19 22 25 26 28 29 30 34 35 38
+ 39 42
c120 30 0 1.66251e-19 $X=3.08 $Y=0.7
c121 9 0 5.27825e-20 $X=1.85 $Y=0.445
r122 43 44 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.865 $Y=1.58
+ $X2=1.865 $Y2=1.655
r123 37 39 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.51
r124 37 38 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.7
r125 35 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=0.95
+ $X2=3.165 $Y2=0.785
r126 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=0.95 $X2=3.165 $Y2=0.95
r127 32 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=0.785
+ $X2=3.165 $Y2=0.95
r128 31 38 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.65 $Y=0.7
+ $X2=2.562 $Y2=0.7
r129 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.08 $Y=0.7
+ $X2=3.165 $Y2=0.785
r130 30 31 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.08 $Y=0.7
+ $X2=2.65 $Y2=0.7
r131 28 38 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=2.562 $Y2=0.7
r132 28 29 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=1.95 $Y2=0.7
r133 26 43 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.865 $Y=1.52
+ $X2=1.865 $Y2=1.58
r134 26 42 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.865 $Y=1.52
+ $X2=1.865 $Y2=1.385
r135 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=1.52 $X2=1.865 $Y2=1.52
r136 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=0.785
+ $X2=1.95 $Y2=0.7
r137 23 25 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.865 $Y=0.785
+ $X2=1.865 $Y2=1.52
r138 22 42 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.845 $Y=0.83
+ $X2=1.845 $Y2=1.385
r139 21 22 21.5285 $w=1.55e-07 $l=4.5e-08 $layer=POLY_cond $X=1.847 $Y=0.785
+ $X2=1.847 $Y2=0.83
r140 19 46 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.225 $Y=0.445
+ $X2=3.225 $Y2=0.785
r141 13 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.26 $Y=1.655
+ $X2=2.26 $Y2=2.165
r142 12 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.58
+ $X2=1.865 $Y2=1.58
r143 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.185 $Y=1.58
+ $X2=2.26 $Y2=1.655
r144 11 12 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.185 $Y=1.58
+ $X2=2.03 $Y2=1.58
r145 9 21 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.85 $Y=0.445
+ $X2=1.85 $Y2=0.785
r146 3 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.835 $Y=2.165
+ $X2=1.835 $Y2=1.655
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_299_47# 1 2 9 13 16 19 21 24 25 28 32 34
+ 38 39 41 43 44
c128 41 0 7.46557e-20 $X=2.205 $Y=1.967
c129 24 0 1.60762e-19 $X=2.205 $Y=1.86
r130 44 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.185 $Y=1.52
+ $X2=3.185 $Y2=1.685
r131 43 46 9.59627 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.172 $Y=1.52
+ $X2=3.172 $Y2=1.685
r132 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.52 $X2=3.185 $Y2=1.52
r133 39 48 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.295 $Y=1.04
+ $X2=2.295 $Y2=0.905
r134 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.04 $X2=2.295 $Y2=1.04
r135 35 38 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.205 $Y=1.04
+ $X2=2.295 $Y2=1.04
r136 29 32 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.52 $Y=0.36
+ $X2=1.64 $Y2=0.36
r137 28 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.16 $Y=1.86
+ $X2=3.16 $Y2=1.685
r138 26 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=1.967
+ $X2=2.205 $Y2=1.967
r139 25 28 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.075 $Y=1.967
+ $X2=3.16 $Y2=1.86
r140 25 26 42.0776 $w=2.13e-07 $l=7.85e-07 $layer=LI1_cond $X=3.075 $Y=1.967
+ $X2=2.29 $Y2=1.967
r141 24 41 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.205 $Y=1.86
+ $X2=2.205 $Y2=1.967
r142 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=1.125
+ $X2=2.205 $Y2=1.04
r143 23 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.205 $Y=1.125
+ $X2=2.205 $Y2=1.86
r144 22 34 1.46632 $w=2.15e-07 $l=1.38e-07 $layer=LI1_cond $X=1.71 $Y=1.967
+ $X2=1.572 $Y2=1.967
r145 21 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=1.967
+ $X2=2.205 $Y2=1.967
r146 21 22 21.9768 $w=2.13e-07 $l=4.1e-07 $layer=LI1_cond $X=2.12 $Y=1.967
+ $X2=1.71 $Y2=1.967
r147 17 34 5.02022 $w=2.22e-07 $l=1.08e-07 $layer=LI1_cond $X=1.572 $Y=2.075
+ $X2=1.572 $Y2=1.967
r148 17 19 4.1907 $w=2.73e-07 $l=1e-07 $layer=LI1_cond $X=1.572 $Y=2.075
+ $X2=1.572 $Y2=2.175
r149 16 34 5.02022 $w=2.22e-07 $l=1.30434e-07 $layer=LI1_cond $X=1.52 $Y=1.86
+ $X2=1.572 $Y2=1.967
r150 15 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.445
+ $X2=1.52 $Y2=0.36
r151 15 16 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.52 $Y=0.445
+ $X2=1.52 $Y2=1.86
r152 13 52 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.14 $Y=2.165
+ $X2=3.14 $Y2=1.685
r153 9 48 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.355 $Y=0.445
+ $X2=2.355 $Y2=0.905
r154 2 19 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.845 $X2=1.625 $Y2=2.175
r155 1 32 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.64 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%D 3 7 9 12 13
r49 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.52
+ $X2=2.705 $Y2=1.685
r50 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.52
+ $X2=2.705 $Y2=1.355
r51 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.52 $X2=2.705 $Y2=1.52
r52 9 13 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.59 $Y=1.52
+ $X2=2.705 $Y2=1.52
r53 7 14 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.745 $Y=0.445
+ $X2=2.745 $Y2=1.355
r54 3 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.72 $Y=2.165
+ $X2=2.72 $Y2=1.685
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%SCD 3 7 9 10 14
c48 3 0 1.66251e-19 $X=3.605 $Y=0.445
r49 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.355
+ $X2=3.665 $Y2=1.52
r50 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.355
+ $X2=3.665 $Y2=1.19
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.665
+ $Y=1.355 $X2=3.665 $Y2=1.355
r52 10 15 4.27171 $w=4.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.775 $Y=1.53
+ $X2=3.775 $Y2=1.355
r53 9 15 4.02761 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.775 $Y=1.19
+ $X2=3.775 $Y2=1.355
r54 7 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.605 $Y=2.165
+ $X2=3.605 $Y2=1.52
r55 3 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.605 $Y=0.445
+ $X2=3.605 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_193_47# 1 2 9 13 14 16 19 23 24 27 30 33
+ 37 38 40 41 42 43 46 52 59 60 61 66
c217 66 0 1.77381e-19 $X=6.925 $Y=0.87
c218 42 0 1.57835e-19 $X=6.57 $Y=0.85
c219 40 0 5.27825e-20 $X=4.685 $Y=0.85
r220 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.925
+ $Y=0.87 $X2=6.925 $Y2=0.87
r221 63 66 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.83 $Y=0.87
+ $X2=6.925 $Y2=0.87
r222 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.045 $Y=0.87
+ $X2=5.045 $Y2=0.705
r223 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.045
+ $Y=0.87 $X2=5.045 $Y2=0.87
r224 53 67 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.715 $Y=0.87
+ $X2=6.925 $Y2=0.87
r225 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.715 $Y=0.85
+ $X2=6.715 $Y2=0.85
r226 50 60 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.83 $Y=0.87
+ $X2=5.045 $Y2=0.87
r227 50 80 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.83 $Y=0.87
+ $X2=4.67 $Y2=0.87
r228 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0.85
+ $X2=4.83 $Y2=0.85
r229 46 75 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.132 $Y=0.85
+ $X2=1.132 $Y2=1.96
r230 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.135 $Y=0.85
+ $X2=1.135 $Y2=0.85
r231 43 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=0.85
+ $X2=4.83 $Y2=0.85
r232 42 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.57 $Y=0.85
+ $X2=6.715 $Y2=0.85
r233 42 43 1.97401 $w=1.4e-07 $l=1.595e-06 $layer=MET1_cond $X=6.57 $Y=0.85
+ $X2=4.975 $Y2=0.85
r234 41 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.28 $Y=0.85
+ $X2=1.135 $Y2=0.85
r235 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=4.83 $Y2=0.85
r236 40 41 4.2141 $w=1.4e-07 $l=3.405e-06 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=1.28 $Y2=0.85
r237 38 69 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=7.205 $Y=1.74
+ $X2=7.12 $Y2=1.74
r238 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.205
+ $Y=1.74 $X2=7.205 $Y2=1.74
r239 34 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.065 $Y=1.74
+ $X2=7.205 $Y2=1.74
r240 33 67 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.97 $Y=0.87
+ $X2=6.925 $Y2=0.87
r241 32 46 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=1.132 $Y=0.715
+ $X2=1.132 $Y2=0.85
r242 30 32 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.13 $Y=0.51
+ $X2=1.13 $Y2=0.715
r243 27 34 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.065 $Y=1.575
+ $X2=7.065 $Y2=1.74
r244 26 33 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.065 $Y=1.035
+ $X2=6.97 $Y2=0.87
r245 26 27 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.065 $Y=1.035
+ $X2=7.065 $Y2=1.575
r246 24 57 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.635 $Y=1.74
+ $X2=4.635 $Y2=1.875
r247 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.74 $X2=4.635 $Y2=1.74
r248 21 80 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.67 $Y=1.035
+ $X2=4.67 $Y2=0.87
r249 21 23 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.67 $Y=1.035
+ $X2=4.67 $Y2=1.74
r250 17 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.12 $Y=1.875
+ $X2=7.12 $Y2=1.74
r251 17 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.12 $Y=1.875
+ $X2=7.12 $Y2=2.275
r252 14 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.83 $Y=0.705
+ $X2=6.83 $Y2=0.87
r253 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.83 $Y=0.705
+ $X2=6.83 $Y2=0.415
r254 13 61 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.105 $Y=0.415
+ $X2=5.105 $Y2=0.705
r255 9 57 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.62 $Y=2.275 $X2=4.62
+ $Y2=1.875
r256 2 75 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.815 $X2=1.105 $Y2=1.96
r257 1 30 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_1098_183# 1 2 9 13 15 18 21 23 29 30 32
+ 33 36
r95 35 36 5.54023 $w=2.61e-07 $l=3e-08 $layer=POLY_cond $X=5.565 $Y=0.93
+ $X2=5.595 $Y2=0.93
r96 32 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=2.3
+ $X2=6.395 $Y2=2.135
r97 27 36 24.0077 $w=2.61e-07 $l=1.3e-07 $layer=POLY_cond $X=5.725 $Y=0.93
+ $X2=5.595 $Y2=0.93
r98 26 29 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=0.93
+ $X2=5.81 $Y2=0.93
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=0.93 $X2=5.725 $Y2=0.93
r100 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.44 $Y=0.45
+ $X2=6.565 $Y2=0.45
r101 19 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.355 $Y=1.065
+ $X2=6.355 $Y2=0.915
r102 19 33 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.355 $Y=1.065
+ $X2=6.355 $Y2=2.135
r103 18 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.355 $Y=0.765
+ $X2=6.355 $Y2=0.915
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.355 $Y=0.535
+ $X2=6.44 $Y2=0.45
r105 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.355 $Y=0.535
+ $X2=6.355 $Y2=0.765
r106 15 30 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.915
+ $X2=6.355 $Y2=0.915
r107 15 29 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.27 $Y=0.915
+ $X2=5.81 $Y2=0.915
r108 11 36 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.595 $Y=0.795
+ $X2=5.595 $Y2=0.93
r109 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.595 $Y=0.795
+ $X2=5.595 $Y2=0.445
r110 7 35 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.565 $Y=1.065
+ $X2=5.565 $Y2=0.93
r111 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.565 $Y=1.065
+ $X2=5.565 $Y2=2.275
r112 2 32 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.735 $X2=6.435 $Y2=2.3
r113 1 23 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.4
+ $Y=0.235 $X2=6.565 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_939_413# 1 2 8 11 13 15 18 20 21 22 26 31
+ 33 35
c109 31 0 1.42307e-19 $X=5.385 $Y=1.315
r110 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.015
+ $Y=1.41 $X2=6.015 $Y2=1.41
r111 35 37 17.1405 $w=2.42e-07 $l=3.4e-07 $layer=LI1_cond $X=5.675 $Y=1.41
+ $X2=6.015 $Y2=1.41
r112 32 35 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=1.575
+ $X2=5.675 $Y2=1.41
r113 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.675 $Y=1.575
+ $X2=5.675 $Y2=2.19
r114 31 35 14.6198 $w=2.42e-07 $l=2.9e-07 $layer=LI1_cond $X=5.385 $Y=1.41
+ $X2=5.675 $Y2=1.41
r115 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.385 $Y=0.535
+ $X2=5.385 $Y2=1.315
r116 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.3 $Y=0.45
+ $X2=5.385 $Y2=0.535
r117 26 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.3 $Y=0.45
+ $X2=4.895 $Y2=0.45
r118 22 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.59 $Y=2.275
+ $X2=5.675 $Y2=2.19
r119 22 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.59 $Y=2.275
+ $X2=4.855 $Y2=2.275
r120 20 38 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.15 $Y=1.41
+ $X2=6.015 $Y2=1.41
r121 20 21 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.15 $Y=1.41
+ $X2=6.225 $Y2=1.41
r122 16 18 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.225 $Y=1.025
+ $X2=6.325 $Y2=1.025
r123 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.325 $Y=0.95
+ $X2=6.325 $Y2=1.025
r124 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.325 $Y=0.95
+ $X2=6.325 $Y2=0.555
r125 9 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.225 $Y=1.545
+ $X2=6.225 $Y2=1.41
r126 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.225 $Y=1.545
+ $X2=6.225 $Y2=2.11
r127 8 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.225 $Y=1.275
+ $X2=6.225 $Y2=1.41
r128 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.225 $Y=1.1
+ $X2=6.225 $Y2=1.025
r129 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.225 $Y=1.1
+ $X2=6.225 $Y2=1.275
r130 2 24 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=2.065 $X2=4.855 $Y2=2.275
r131 1 28 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.235 $X2=4.895 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_1526_315# 1 2 9 13 15 17 20 22 24 27 29
+ 32 36 39 41 44 48 52 53 62
c99 62 0 1.11165e-19 $X=9.635 $Y=1.16
r100 61 62 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=9.215 $Y=1.16
+ $X2=9.635 $Y2=1.16
r101 54 56 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.705 $Y=1.74
+ $X2=7.82 $Y2=1.74
r102 48 50 17.5434 $w=3.48e-07 $l=4.4e-07 $layer=LI1_cond $X=8.56 $Y=0.385
+ $X2=8.56 $Y2=0.825
r103 45 61 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.18 $Y=1.16
+ $X2=9.215 $Y2=1.16
r104 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.18
+ $Y=1.16 $X2=9.18 $Y2=1.16
r105 42 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=1.16
+ $X2=8.65 $Y2=1.16
r106 42 44 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.735 $Y=1.16
+ $X2=9.18 $Y2=1.16
r107 41 52 7.13466 $w=2.2e-07 $l=1.88348e-07 $layer=LI1_cond $X=8.65 $Y=1.575
+ $X2=8.6 $Y2=1.74
r108 40 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.65 $Y=1.325
+ $X2=8.65 $Y2=1.16
r109 40 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.65 $Y=1.325
+ $X2=8.65 $Y2=1.575
r110 39 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.65 $Y=0.995
+ $X2=8.65 $Y2=1.16
r111 39 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.65 $Y=0.995
+ $X2=8.65 $Y2=0.825
r112 34 52 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=8.6 $Y=1.905
+ $X2=8.6 $Y2=1.74
r113 34 36 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.6 $Y=1.905
+ $X2=8.6 $Y2=2.29
r114 32 56 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.885 $Y=1.74
+ $X2=7.82 $Y2=1.74
r115 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.885
+ $Y=1.74 $X2=7.885 $Y2=1.74
r116 29 52 0.067832 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=8.465 $Y=1.74
+ $X2=8.6 $Y2=1.74
r117 29 31 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=8.465 $Y=1.74
+ $X2=7.885 $Y2=1.74
r118 25 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.635 $Y=1.325
+ $X2=9.635 $Y2=1.16
r119 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.635 $Y=1.325
+ $X2=9.635 $Y2=1.985
r120 22 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.635 $Y=0.995
+ $X2=9.635 $Y2=1.16
r121 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.635 $Y=0.995
+ $X2=9.635 $Y2=0.56
r122 18 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.215 $Y=1.325
+ $X2=9.215 $Y2=1.16
r123 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.215 $Y=1.325
+ $X2=9.215 $Y2=1.985
r124 15 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.215 $Y=0.995
+ $X2=9.215 $Y2=1.16
r125 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.215 $Y=0.995
+ $X2=9.215 $Y2=0.56
r126 11 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.82 $Y=1.575
+ $X2=7.82 $Y2=1.74
r127 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.82 $Y=1.575
+ $X2=7.82 $Y2=0.445
r128 7 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1.905
+ $X2=7.705 $Y2=1.74
r129 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.705 $Y=1.905
+ $X2=7.705 $Y2=2.275
r130 2 52 600 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=1.485 $X2=8.55 $Y2=1.68
r131 2 36 600 $w=1.7e-07 $l=8.65246e-07 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=1.485 $X2=8.55 $Y2=2.29
r132 1 48 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=8.425
+ $Y=0.235 $X2=8.55 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_1355_413# 1 2 7 9 12 14 15 16 20 27 30 33
+ 34
c88 30 0 1.11165e-19 $X=8.31 $Y=1.16
c89 27 0 4.21632e-20 $X=7.545 $Y=2.165
c90 15 0 1.26335e-19 $X=8.76 $Y=1.16
r91 33 35 11.5578 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=7.48 $Y=1.16
+ $X2=7.48 $Y2=1.405
r92 33 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.48 $Y=1.16
+ $X2=7.48 $Y2=0.995
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.31
+ $Y=1.16 $X2=8.31 $Y2=1.16
r94 28 33 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.63 $Y=1.16
+ $X2=7.48 $Y2=1.16
r95 28 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.63 $Y=1.16
+ $X2=8.31 $Y2=1.16
r96 27 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.545 $Y=2.165
+ $X2=7.545 $Y2=1.405
r97 24 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.415 $Y=0.535
+ $X2=7.415 $Y2=0.995
r98 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.33 $Y=0.45
+ $X2=7.415 $Y2=0.535
r99 20 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.33 $Y=0.45
+ $X2=7.125 $Y2=0.45
r100 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.46 $Y=2.25
+ $X2=7.545 $Y2=2.165
r101 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.46 $Y=2.25
+ $X2=6.91 $Y2=2.25
r102 14 31 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=8.685 $Y=1.16
+ $X2=8.31 $Y2=1.16
r103 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.685 $Y=1.16
+ $X2=8.76 $Y2=1.16
r104 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=1.325
+ $X2=8.76 $Y2=1.16
r105 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.76 $Y=1.325
+ $X2=8.76 $Y2=1.985
r106 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=0.995
+ $X2=8.76 $Y2=1.16
r107 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.76 $Y=0.995
+ $X2=8.76 $Y2=0.56
r108 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=2.065 $X2=6.91 $Y2=2.25
r109 1 22 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=6.905
+ $Y=0.235 $X2=7.125 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 42 46 48
+ 50 55 56 57 59 64 69 81 88 94 97 100 103 106 110
c163 110 0 1.81794e-19 $X=9.89 $Y=2.72
c164 2 0 2.35417e-19 $X=1.91 $Y=1.845
c165 1 0 3.29888e-20 $X=0.55 $Y=1.815
r166 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r167 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r168 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r169 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r170 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r171 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r172 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r173 92 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r174 92 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r175 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r176 89 106 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=9.08 $Y=2.72
+ $X2=8.992 $Y2=2.72
r177 89 91 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.08 $Y=2.72
+ $X2=9.43 $Y2=2.72
r178 88 109 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=9.775 $Y=2.72
+ $X2=9.947 $Y2=2.72
r179 88 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.775 $Y=2.72
+ $X2=9.43 $Y2=2.72
r180 87 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r181 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r182 84 87 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r183 83 86 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r184 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r185 81 103 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.81 $Y=2.72
+ $X2=7.962 $Y2=2.72
r186 81 86 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.81 $Y=2.72
+ $X2=7.59 $Y2=2.72
r187 80 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r188 80 101 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r189 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r190 77 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=3.84 $Y2=2.72
r191 77 79 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r192 76 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r193 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r194 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r195 73 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r196 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r197 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r198 70 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.045 $Y2=2.72
r199 70 72 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.53 $Y2=2.72
r200 69 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.84 $Y2=2.72
r201 69 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.45 $Y2=2.72
r202 68 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r203 68 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r204 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r205 65 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=0.685 $Y2=2.72
r206 65 67 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r207 64 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=2.045 $Y2=2.72
r208 64 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=1.61 $Y2=2.72
r209 59 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.685 $Y2=2.72
r210 59 61 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r211 57 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r212 57 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r213 55 79 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=5.75 $Y2=2.72
r214 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=6.015 $Y2=2.72
r215 54 83 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.1 $Y=2.72
+ $X2=6.21 $Y2=2.72
r216 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.1 $Y=2.72
+ $X2=6.015 $Y2=2.72
r217 50 53 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.86 $Y=1.63
+ $X2=9.86 $Y2=2.31
r218 48 109 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=9.86 $Y=2.635
+ $X2=9.947 $Y2=2.72
r219 48 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.86 $Y=2.635
+ $X2=9.86 $Y2=2.31
r220 44 106 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=8.992 $Y=2.635
+ $X2=8.992 $Y2=2.72
r221 44 46 53.5532 $w=1.73e-07 $l=8.45e-07 $layer=LI1_cond $X=8.992 $Y=2.635
+ $X2=8.992 $Y2=1.79
r222 43 103 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.115 $Y=2.72
+ $X2=7.962 $Y2=2.72
r223 42 106 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=8.905 $Y=2.72
+ $X2=8.992 $Y2=2.72
r224 42 43 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.905 $Y=2.72
+ $X2=8.115 $Y2=2.72
r225 38 103 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.962 $Y=2.635
+ $X2=7.962 $Y2=2.72
r226 38 40 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=7.962 $Y=2.635
+ $X2=7.962 $Y2=2.3
r227 34 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=2.635
+ $X2=6.015 $Y2=2.72
r228 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.015 $Y=2.635
+ $X2=6.015 $Y2=2
r229 30 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=2.635
+ $X2=3.84 $Y2=2.72
r230 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.84 $Y=2.635
+ $X2=3.84 $Y2=2.33
r231 26 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.72
r232 26 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.33
r233 22 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.72
r234 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.22
r235 7 53 400 $w=1.7e-07 $l=8.9687e-07 $layer=licon1_PDIFF $count=1 $X=9.71
+ $Y=1.485 $X2=9.86 $Y2=2.31
r236 7 50 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.71
+ $Y=1.485 $X2=9.86 $Y2=1.63
r237 6 46 300 $w=1.7e-07 $l=3.74566e-07 $layer=licon1_PDIFF $count=2 $X=8.835
+ $Y=1.485 $X2=8.99 $Y2=1.79
r238 5 40 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=2.065 $X2=8.025 $Y2=2.3
r239 4 36 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=5.64
+ $Y=2.065 $X2=6.015 $Y2=2
r240 3 32 600 $w=1.7e-07 $l=5.59308e-07 $layer=licon1_PDIFF $count=1 $X=3.68
+ $Y=1.845 $X2=3.84 $Y2=2.33
r241 2 28 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.845 $X2=2.045 $Y2=2.33
r242 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.815 $X2=0.685 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%A_559_369# 1 2 3 4 13 17 22 24 25 26 27 28
+ 30 32 36 38 39
r111 39 41 21.3062 $w=2.09e-07 $l=3.65e-07 $layer=LI1_cond $X=4.327 $Y=1.91
+ $X2=4.327 $Y2=2.275
r112 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.295 $Y=0.45
+ $X2=4.395 $Y2=0.45
r113 32 39 5.42244 $w=2.09e-07 $l=9.97246e-08 $layer=LI1_cond $X=4.295 $Y=1.825
+ $X2=4.327 $Y2=1.91
r114 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=0.865
+ $X2=4.295 $Y2=0.78
r115 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.295 $Y=0.865
+ $X2=4.295 $Y2=1.825
r116 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=0.695
+ $X2=4.295 $Y2=0.78
r117 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=0.535
+ $X2=4.295 $Y2=0.45
r118 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.295 $Y=0.535
+ $X2=4.295 $Y2=0.695
r119 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=0.78
+ $X2=4.295 $Y2=0.78
r120 27 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.21 $Y=0.78
+ $X2=3.59 $Y2=0.78
r121 25 39 1.94907 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.21 $Y=1.91
+ $X2=4.327 $Y2=1.91
r122 25 26 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.21 $Y=1.91
+ $X2=3.585 $Y2=1.91
r123 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=0.695
+ $X2=3.59 $Y2=0.78
r124 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.505 $Y=0.445
+ $X2=3.505 $Y2=0.695
r125 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=1.995
+ $X2=3.585 $Y2=1.91
r126 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.5 $Y=1.995
+ $X2=3.5 $Y2=2.245
r127 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=0.36
+ $X2=3.505 $Y2=0.445
r128 17 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.42 $Y=0.36
+ $X2=3.01 $Y2=0.36
r129 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=2.33
+ $X2=3.5 $Y2=2.245
r130 13 15 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.415 $Y=2.33
+ $X2=2.93 $Y2=2.33
r131 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=2.065 $X2=4.36 $Y2=2.275
r132 3 15 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.845 $X2=2.93 $Y2=2.33
r133 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.235 $X2=4.395 $Y2=0.45
r134 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=3.01 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%Q 1 2 11 12 13 14 15 27
c31 12 0 1.26335e-19 $X=9.432 $Y=1.505
r32 15 24 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=9.432 $Y=2.21
+ $X2=9.432 $Y2=2.31
r33 14 15 11.3574 $w=3.43e-07 $l=3.4e-07 $layer=LI1_cond $X=9.432 $Y=1.87
+ $X2=9.432 $Y2=2.21
r34 13 31 13.323 $w=3.43e-07 $l=3.1e-07 $layer=LI1_cond $X=9.432 $Y=0.51
+ $X2=9.432 $Y2=0.82
r35 13 27 3.84148 $w=3.43e-07 $l=1.15e-07 $layer=LI1_cond $X=9.432 $Y=0.51
+ $X2=9.432 $Y2=0.395
r36 12 31 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=9.52 $Y=1.505
+ $X2=9.52 $Y2=0.82
r37 11 12 7.14324 $w=3.43e-07 $l=1.25e-07 $layer=LI1_cond $X=9.432 $Y=1.63
+ $X2=9.432 $Y2=1.505
r38 9 14 6.447 $w=3.43e-07 $l=1.93e-07 $layer=LI1_cond $X=9.432 $Y=1.677
+ $X2=9.432 $Y2=1.87
r39 9 11 1.56999 $w=3.43e-07 $l=4.7e-08 $layer=LI1_cond $X=9.432 $Y=1.677
+ $X2=9.432 $Y2=1.63
r40 2 24 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=1.485 $X2=9.425 $Y2=2.31
r41 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=1.485 $X2=9.425 $Y2=1.63
r42 1 27 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=9.29
+ $Y=0.235 $X2=9.425 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_2%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 44 48
+ 50 52 54 56 61 66 74 82 88 91 94 97 100 103 107
c163 107 0 2.71124e-20 $X=9.89 $Y=0
r164 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r165 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r166 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r167 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r168 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r169 95 98 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r170 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r171 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r172 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r173 86 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r174 86 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r175 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r176 83 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=0 $X2=8.99
+ $Y2=0
r177 83 85 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.075 $Y=0
+ $X2=9.43 $Y2=0
r178 82 106 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=9.775 $Y=0
+ $X2=9.947 $Y2=0
r179 82 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.775 $Y=0 $X2=9.43
+ $Y2=0
r180 81 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r181 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r182 78 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r183 78 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r184 77 80 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=7.59
+ $Y2=0
r185 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r186 75 97 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=5.905
+ $Y2=0
r187 75 77 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=6.21
+ $Y2=0
r188 74 100 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.93 $Y2=0
r189 74 80 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.59 $Y2=0
r190 73 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r191 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r192 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r193 70 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r194 69 72 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r195 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r196 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.14
+ $Y2=0
r197 67 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r198 66 94 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.86
+ $Y2=0
r199 66 72 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.45
+ $Y2=0
r200 65 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r201 65 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r202 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r203 62 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r204 62 64 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r205 61 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.14
+ $Y2=0
r206 61 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r207 56 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r208 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r209 54 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r210 54 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r211 50 106 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.947 $Y2=0
r212 50 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0.395
r213 46 103 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=0.085
+ $X2=8.99 $Y2=0
r214 46 48 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.99 $Y=0.085
+ $X2=8.99 $Y2=0.53
r215 45 100 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=7.93 $Y2=0
r216 44 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=0 $X2=8.99
+ $Y2=0
r217 44 45 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.905 $Y=0
+ $X2=8.115 $Y2=0
r218 40 100 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r219 40 42 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.45
r220 36 97 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0.085
+ $X2=5.905 $Y2=0
r221 36 38 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.905 $Y=0.085
+ $X2=5.905 $Y2=0.42
r222 35 94 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.86
+ $Y2=0
r223 34 97 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.72 $Y=0 $X2=5.905
+ $Y2=0
r224 34 35 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=5.72 $Y=0 $X2=3.96
+ $Y2=0
r225 30 94 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0
r226 30 32 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0.36
r227 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r228 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.36
r229 22 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r230 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r231 7 52 91 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=2 $X=9.71
+ $Y=0.235 $X2=9.86 $Y2=0.395
r232 6 48 182 $w=1.7e-07 $l=3.64349e-07 $layer=licon1_NDIFF $count=1 $X=8.835
+ $Y=0.235 $X2=8.99 $Y2=0.53
r233 5 42 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=7.895
+ $Y=0.235 $X2=8.03 $Y2=0.45
r234 4 38 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=5.67
+ $Y=0.235 $X2=5.975 $Y2=0.42
r235 3 32 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.68
+ $Y=0.235 $X2=3.845 $Y2=0.36
r236 2 28 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.14 $Y2=0.36
r237 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__sedfxbp_1.spice
* Created: Tue Sep  1 19:31:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sedfxbp_1.pex.spice"
.subckt sky130_fd_sc_hd__sedfxbp_1  VNB VPB CLK D DE SCD SCE VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1042 N_VGND_M1042_d N_CLK_M1042_g N_A_27_47#_M1042_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_193_47#_M1024_d N_A_27_47#_M1024_g N_VGND_M1042_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_381_47# N_D_M1004_g N_A_299_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_DE_M1005_g A_381_47# VNB NSHORT L=0.15 W=0.42 AD=0.1092
+ AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_DE_M1039_g N_A_423_343#_M1039_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.1092 PD=0.71 PS=1.36 NRD=1.428 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1025 A_729_47# N_A_423_343#_M1025_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0609 PD=0.78 PS=0.71 NRD=35.712 NRS=1.428 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1043 N_A_299_47#_M1043_d N_A_791_264#_M1043_g A_729_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0756 PD=0.69 PS=0.78 NRD=0 NRS=35.712 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_A_915_47#_M1035_d N_A_885_21#_M1035_g N_A_299_47#_M1043_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_SCE_M1008_g N_A_885_21#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1026 A_1226_119# N_SCD_M1026_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1012 N_A_915_47#_M1012_d N_SCE_M1012_g A_1226_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.242469 AS=0.0441 PD=1.62077 PS=0.63 NRD=1.428 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1029 N_A_1446_413#_M1029_d N_A_27_47#_M1029_g N_A_915_47#_M1012_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0522 AS=0.207831 PD=0.65 PS=1.38923 NRD=0 NRS=34.992 M=1
+ R=2.4 SA=75000.6 SB=75001.8 A=0.054 P=1.02 MULT=1
MM1014 A_1561_47# N_A_193_47#_M1014_g N_A_1446_413#_M1029_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0700615 AS=0.0522 PD=0.738462 PS=0.65 NRD=46.536 NRS=4.992 M=1
+ R=2.4 SA=75001 SB=75001.3 A=0.054 P=1.02 MULT=1
MM1021 N_VGND_M1021_d N_A_1610_159#_M1021_g A_1561_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0958472 AS=0.0817385 PD=0.859811 PS=0.861538 NRD=0 NRS=39.888 M=1 R=2.8
+ SA=75001.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1006 N_A_1610_159#_M1006_d N_A_1446_413#_M1006_g N_VGND_M1021_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.146053 PD=1.8 PS=1.31019 NRD=0 NRS=30.936 M=1
+ R=4.26667 SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1040 A_1974_47# N_A_1610_159#_M1040_g N_VGND_M1040_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0730154 AS=0.1092 PD=0.813077 PS=1.36 NRD=33.948 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1028 N_A_2051_413#_M1028_d N_A_193_47#_M1028_g A_1974_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0684 AS=0.0625846 PD=0.74 PS=0.696923 NRD=3.324 NRS=39.612 M=1
+ R=2.4 SA=75000.7 SB=75001.7 A=0.054 P=1.02 MULT=1
MM1030 A_2177_47# N_A_27_47#_M1030_g N_A_2051_413#_M1028_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0684 PD=0.687692 PS=0.74 NRD=38.076 NRS=30 M=1 R=2.4
+ SA=75001.2 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1002 N_VGND_M1002_d N_A_791_264#_M1002_g A_2177_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.0710769 PD=0.773271 PS=0.802308 NRD=17.136 NRS=32.628 M=1
+ R=2.8 SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_Q_N_M1003_d N_A_791_264#_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.121799 PD=1.82 PS=1.19673 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1038_d N_A_2051_413#_M1038_g N_A_791_264#_M1038_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=17.136 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1041 N_Q_M1041_d N_A_2051_413#_M1041_g N_VGND_M1038_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.121799 PD=1.86 PS=1.19673 NRD=0.912 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_27_47#_M1016_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1031 A_381_369# N_D_M1031_g N_A_299_47#_M1031_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1664 PD=0.85 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.5 A=0.096 P=1.58 MULT=1
MM1033 N_VPWR_M1033_d N_A_423_343#_M1033_g A_381_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1664 AS=0.0672 PD=1.8 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_VPWR_M1013_d N_DE_M1013_g N_A_423_343#_M1013_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0928 AS=0.1664 PD=0.93 PS=1.8 NRD=1.5366 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1017 A_729_369# N_DE_M1017_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.0928 PD=1 PS=0.93 NRD=38.4741 NRS=1.5366 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1036 N_A_299_47#_M1036_d N_A_791_264#_M1036_g A_729_369# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0992 AS=0.1152 PD=0.95 PS=1 NRD=0 NRS=38.4741 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1015 N_A_915_47#_M1015_d N_SCE_M1015_g N_A_299_47#_M1036_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1984 AS=0.0992 PD=1.9 PS=0.95 NRD=13.8491 NRS=10.7562 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_SCE_M1034_g N_A_885_21#_M1034_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1264 AS=0.1696 PD=1.035 PS=1.81 NRD=16.9223 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1023 A_1231_369# N_SCD_M1023_g N_VPWR_M1034_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1056 AS=0.1264 PD=0.97 PS=1.035 NRD=33.8446 NRS=18.4589 M=1 R=4.26667
+ SA=75000.7 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1032 N_A_915_47#_M1032_d N_A_885_21#_M1032_g A_1231_369# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.161992 AS=0.1056 PD=1.31019 PS=0.97 NRD=19.9955 NRS=33.8446 M=1
+ R=4.26667 SA=75001.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 N_A_1446_413#_M1011_d N_A_193_47#_M1011_g N_A_915_47#_M1032_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06405 AS=0.106308 PD=0.725 PS=0.859811 NRD=4.6886
+ NRS=48.068 M=1 R=2.8 SA=75001.8 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1018 A_1537_413# N_A_27_47#_M1018_g N_A_1446_413#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07665 AS=0.06405 PD=0.785 PS=0.725 NRD=59.7895 NRS=7.0329 M=1
+ R=2.8 SA=75002.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1610_159#_M1009_g A_1537_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.128423 AS=0.07665 PD=0.904615 PS=0.785 NRD=97.318 NRS=59.7895 M=1
+ R=2.8 SA=75002.8 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1019 N_A_1610_159#_M1019_d N_A_1446_413#_M1019_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=0.75 AD=0.195 AS=0.229327 PD=2.02 PS=1.61538 NRD=0 NRS=6.5601 M=1 R=5
+ SA=75002.1 SB=75000.2 A=0.1125 P=1.8 MULT=1
MM1037 A_1960_413# N_A_1610_159#_M1037_g N_VPWR_M1037_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06405 AS=0.1092 PD=0.725 PS=1.36 NRD=45.7237 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1027 N_A_2051_413#_M1027_d N_A_27_47#_M1027_g A_1960_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.06405 PD=0.69 PS=0.725 NRD=0 NRS=45.7237 M=1 R=2.8
+ SA=75000.6 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1020 A_2135_413# N_A_193_47#_M1020_g N_A_2051_413#_M1027_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0882 AS=0.0567 PD=0.84 PS=0.69 NRD=72.693 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_791_264#_M1010_g A_2135_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.0882 PD=0.789718 PS=0.84 NRD=29.3136 NRS=72.693 M=1 R=2.8
+ SA=75001.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_Q_N_M1001_d N_A_791_264#_M1001_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.205282 PD=2.52 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_A_2051_413#_M1022_g N_A_791_264#_M1022_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.120195 AS=0.1728 PD=1.04195 PS=1.82 NRD=18.4589 NRS=1.5366
+ M=1 R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1007 N_Q_M1007_d N_A_2051_413#_M1007_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.187805 PD=2.56 PS=1.62805 NRD=0.9653 NRS=0 M=1 R=6.66667
+ SA=75000.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX44_noxref VNB VPB NWDIODE A=23.1962 P=32.75
c_149 VNB 0 1.01407e-19 $X=0.145 $Y=-0.085
c_282 VPB 0 1.40584e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__sedfxbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__bufbuf_16.spice
* Created: Thu Aug 27 14:10:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__bufbuf_16.pex.spice"
.subckt sky130_fd_sc_hd__bufbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1049 N_A_109_47#_M1049_d N_A_M1049_g N_VGND_M1049_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_215_47#_M1006_d N_A_109_47#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75010.3 A=0.0975 P=1.6 MULT=1
MM1007 N_A_215_47#_M1007_d N_A_109_47#_M1007_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75009.8 A=0.0975 P=1.6 MULT=1
MM1011 N_A_215_47#_M1007_d N_A_109_47#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75009.4 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1011_s N_A_215_47#_M1010_g N_A_549_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75009 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_215_47#_M1012_g N_A_549_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75008.6 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1012_d N_A_215_47#_M1020_g N_A_549_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75008.2 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A_215_47#_M1021_g N_A_549_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75007.7 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1021_d N_A_215_47#_M1023_g N_A_549_47#_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1033 N_VGND_M1033_d N_A_215_47#_M1033_g N_A_549_47#_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1033_d N_A_549_47#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75006.5 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_549_47#_M1009_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1009_d N_A_549_47#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.8
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A_549_47#_M1018_g N_X_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.2
+ SB=75005.2 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1018_d N_A_549_47#_M1026_g N_X_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.6
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1027_d N_A_549_47#_M1027_g N_X_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.1
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1028 N_VGND_M1027_d N_A_549_47#_M1028_g N_X_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.5
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1029 N_VGND_M1029_d N_A_549_47#_M1029_g N_X_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.9
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1035 N_VGND_M1029_d N_A_549_47#_M1035_g N_X_M1035_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.3
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1038_d N_A_549_47#_M1038_g N_X_M1035_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.7
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1040 N_VGND_M1038_d N_A_549_47#_M1040_g N_X_M1040_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1041 N_VGND_M1041_d N_A_549_47#_M1041_g N_X_M1040_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1042 N_VGND_M1041_d N_A_549_47#_M1042_g N_X_M1042_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1043 N_VGND_M1043_d N_A_549_47#_M1043_g N_X_M1042_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1046 N_VGND_M1043_d N_A_549_47#_M1046_g N_X_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1051 N_VGND_M1051_d N_A_549_47#_M1051_g N_X_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75010.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1032 N_A_109_47#_M1032_d N_A_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_109_47#_M1003_g N_A_215_47#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75010.3 A=0.15 P=2.3 MULT=1
MM1034 N_VPWR_M1003_d N_A_109_47#_M1034_g N_A_215_47#_M1034_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75009.8 A=0.15 P=2.3 MULT=1
MM1044 N_VPWR_M1044_d N_A_109_47#_M1044_g N_A_215_47#_M1034_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75009.4 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1044_d N_A_215_47#_M1013_g N_A_549_47#_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75009 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_215_47#_M1014_g N_A_549_47#_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75008.6 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1014_d N_A_215_47#_M1019_g N_A_549_47#_M1019_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75008.2 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_A_215_47#_M1024_g N_A_549_47#_M1019_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75007.7 A=0.15 P=2.3 MULT=1
MM1025 N_VPWR_M1024_d N_A_215_47#_M1025_g N_A_549_47#_M1025_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75007.3 A=0.15 P=2.3 MULT=1
MM1045 N_VPWR_M1045_d N_A_215_47#_M1045_g N_A_549_47#_M1025_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75006.9 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_549_47#_M1001_g N_VPWR_M1045_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75006.5 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1001_d N_A_549_47#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75006.1 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1004_d N_A_549_47#_M1004_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8
+ SB=75005.6 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1004_d N_A_549_47#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1008_d N_A_549_47#_M1008_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.6
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1015 N_X_M1008_d N_A_549_47#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.1
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1016 N_X_M1016_d N_A_549_47#_M1016_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.5
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1022 N_X_M1016_d N_A_549_47#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.9
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1030 N_X_M1030_d N_A_549_47#_M1030_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.3
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1031 N_X_M1030_d N_A_549_47#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.7
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1036 N_X_M1036_d N_A_549_47#_M1036_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1037 N_X_M1036_d N_A_549_47#_M1037_g N_VPWR_M1037_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1039 N_X_M1039_d N_A_549_47#_M1039_g N_VPWR_M1037_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1047 N_X_M1039_d N_A_549_47#_M1047_g N_VPWR_M1047_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1048 N_X_M1048_d N_A_549_47#_M1048_g N_VPWR_M1047_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1050 N_X_M1048_d N_A_549_47#_M1050_g N_VPWR_M1050_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75010.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX52_noxref VNB VPB NWDIODE A=19.8057 P=27.89
*
.include "sky130_fd_sc_hd__bufbuf_16.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdfxbp_2.pxi.spice
* Created: Tue Sep  1 19:31:09 2020
* 
x_PM_SKY130_FD_SC_HD__SDFXBP_2%CLK N_CLK_c_246_n N_CLK_c_250_n N_CLK_c_247_n
+ N_CLK_M1037_g N_CLK_c_251_n N_CLK_M1012_g N_CLK_c_252_n CLK
+ PM_SKY130_FD_SC_HD__SDFXBP_2%CLK
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_27_47# N_A_27_47#_M1037_s N_A_27_47#_M1012_s
+ N_A_27_47#_M1027_g N_A_27_47#_M1036_g N_A_27_47#_M1024_g N_A_27_47#_c_290_n
+ N_A_27_47#_c_291_n N_A_27_47#_M1000_g N_A_27_47#_M1018_g N_A_27_47#_c_292_n
+ N_A_27_47#_M1023_g N_A_27_47#_c_525_p N_A_27_47#_c_294_n N_A_27_47#_c_295_n
+ N_A_27_47#_c_307_n N_A_27_47#_c_296_n N_A_27_47#_c_413_p N_A_27_47#_c_308_n
+ N_A_27_47#_c_309_n N_A_27_47#_c_297_n N_A_27_47#_c_310_n N_A_27_47#_c_311_n
+ N_A_27_47#_c_312_n N_A_27_47#_c_313_n N_A_27_47#_c_314_n N_A_27_47#_c_298_n
+ N_A_27_47#_c_316_n N_A_27_47#_c_317_n N_A_27_47#_c_318_n N_A_27_47#_c_299_n
+ N_A_27_47#_c_300_n PM_SKY130_FD_SC_HD__SDFXBP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%SCE N_SCE_M1030_g N_SCE_M1039_g N_SCE_M1026_g
+ N_SCE_M1021_g N_SCE_c_537_n N_SCE_c_547_n N_SCE_c_538_n N_SCE_c_559_p
+ N_SCE_c_539_n N_SCE_c_540_n N_SCE_c_541_n N_SCE_c_542_n SCE
+ PM_SKY130_FD_SC_HD__SDFXBP_2%SCE
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_299_47# N_A_299_47#_M1039_s N_A_299_47#_M1030_s
+ N_A_299_47#_M1016_g N_A_299_47#_M1007_g N_A_299_47#_c_646_n
+ N_A_299_47#_c_653_n N_A_299_47#_c_661_n N_A_299_47#_c_647_n
+ N_A_299_47#_c_663_n N_A_299_47#_c_655_n N_A_299_47#_c_648_n
+ N_A_299_47#_c_656_n N_A_299_47#_c_649_n N_A_299_47#_c_650_n
+ N_A_299_47#_c_668_n N_A_299_47#_c_657_n N_A_299_47#_c_658_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%A_299_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%D N_D_M1010_g N_D_M1017_g D N_D_c_774_n
+ N_D_c_775_n PM_SKY130_FD_SC_HD__SDFXBP_2%D
x_PM_SKY130_FD_SC_HD__SDFXBP_2%SCD N_SCD_M1011_g N_SCD_M1004_g SCD N_SCD_c_822_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%SCD
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_193_47# N_A_193_47#_M1027_d N_A_193_47#_M1036_d
+ N_A_193_47#_M1015_g N_A_193_47#_M1020_g N_A_193_47#_c_868_n
+ N_A_193_47#_M1022_g N_A_193_47#_M1008_g N_A_193_47#_c_869_n
+ N_A_193_47#_c_885_n N_A_193_47#_c_870_n N_A_193_47#_c_871_n
+ N_A_193_47#_c_872_n N_A_193_47#_c_887_n N_A_193_47#_c_888_n
+ N_A_193_47#_c_873_n N_A_193_47#_c_874_n N_A_193_47#_c_875_n
+ N_A_193_47#_c_1007_p N_A_193_47#_c_876_n N_A_193_47#_c_877_n
+ N_A_193_47#_c_878_n N_A_193_47#_c_879_n N_A_193_47#_c_880_n
+ N_A_193_47#_c_881_n PM_SKY130_FD_SC_HD__SDFXBP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_1097_183# N_A_1097_183#_M1001_d
+ N_A_1097_183#_M1033_d N_A_1097_183#_M1013_g N_A_1097_183#_M1034_g
+ N_A_1097_183#_c_1085_n N_A_1097_183#_c_1111_n N_A_1097_183#_c_1131_p
+ N_A_1097_183#_c_1112_n N_A_1097_183#_c_1086_n N_A_1097_183#_c_1087_n
+ N_A_1097_183#_c_1099_n N_A_1097_183#_c_1088_n N_A_1097_183#_c_1089_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%A_1097_183#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_938_413# N_A_938_413#_M1024_d
+ N_A_938_413#_M1015_d N_A_938_413#_c_1178_n N_A_938_413#_M1033_g
+ N_A_938_413#_c_1179_n N_A_938_413#_M1001_g N_A_938_413#_c_1180_n
+ N_A_938_413#_c_1181_n N_A_938_413#_c_1182_n N_A_938_413#_c_1196_n
+ N_A_938_413#_c_1222_n N_A_938_413#_c_1183_n N_A_938_413#_c_1188_n
+ N_A_938_413#_c_1184_n PM_SKY130_FD_SC_HD__SDFXBP_2%A_938_413#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_1525_315# N_A_1525_315#_M1032_s
+ N_A_1525_315#_M1035_s N_A_1525_315#_M1031_g N_A_1525_315#_M1003_g
+ N_A_1525_315#_c_1287_n N_A_1525_315#_M1028_g N_A_1525_315#_M1005_g
+ N_A_1525_315#_c_1288_n N_A_1525_315#_M1029_g N_A_1525_315#_M1019_g
+ N_A_1525_315#_c_1289_n N_A_1525_315#_c_1290_n N_A_1525_315#_c_1291_n
+ N_A_1525_315#_c_1292_n N_A_1525_315#_M1025_g N_A_1525_315#_M1038_g
+ N_A_1525_315#_c_1304_n N_A_1525_315#_c_1305_n N_A_1525_315#_c_1306_n
+ N_A_1525_315#_c_1307_n N_A_1525_315#_c_1308_n N_A_1525_315#_c_1293_n
+ N_A_1525_315#_c_1309_n N_A_1525_315#_c_1294_n N_A_1525_315#_c_1295_n
+ N_A_1525_315#_c_1311_n N_A_1525_315#_c_1326_p
+ PM_SKY130_FD_SC_HD__SDFXBP_2%A_1525_315#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_1354_413# N_A_1354_413#_M1022_d
+ N_A_1354_413#_M1018_d N_A_1354_413#_c_1422_n N_A_1354_413#_M1032_g
+ N_A_1354_413#_M1035_g N_A_1354_413#_c_1423_n N_A_1354_413#_c_1424_n
+ N_A_1354_413#_c_1434_n N_A_1354_413#_c_1437_n N_A_1354_413#_c_1431_n
+ N_A_1354_413#_c_1425_n N_A_1354_413#_c_1426_n N_A_1354_413#_c_1427_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%A_1354_413#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_2049_47# N_A_2049_47#_M1025_s
+ N_A_2049_47#_M1038_s N_A_2049_47#_c_1509_n N_A_2049_47#_M1006_g
+ N_A_2049_47#_M1002_g N_A_2049_47#_c_1510_n N_A_2049_47#_M1009_g
+ N_A_2049_47#_M1014_g N_A_2049_47#_c_1511_n N_A_2049_47#_c_1516_n
+ N_A_2049_47#_c_1512_n N_A_2049_47#_c_1532_n N_A_2049_47#_c_1513_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%A_2049_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%VPWR N_VPWR_M1012_d N_VPWR_M1030_d N_VPWR_M1004_d
+ N_VPWR_M1013_d N_VPWR_M1031_d N_VPWR_M1035_d N_VPWR_M1019_d N_VPWR_M1038_d
+ N_VPWR_M1014_d N_VPWR_c_1579_n N_VPWR_c_1580_n N_VPWR_c_1581_n N_VPWR_c_1582_n
+ N_VPWR_c_1583_n N_VPWR_c_1584_n N_VPWR_c_1585_n N_VPWR_c_1586_n
+ N_VPWR_c_1587_n N_VPWR_c_1588_n N_VPWR_c_1589_n N_VPWR_c_1590_n
+ N_VPWR_c_1591_n N_VPWR_c_1592_n N_VPWR_c_1593_n VPWR N_VPWR_c_1594_n
+ N_VPWR_c_1595_n N_VPWR_c_1596_n N_VPWR_c_1597_n N_VPWR_c_1598_n
+ N_VPWR_c_1599_n N_VPWR_c_1600_n N_VPWR_c_1601_n N_VPWR_c_1602_n
+ N_VPWR_c_1603_n N_VPWR_c_1604_n N_VPWR_c_1605_n N_VPWR_c_1578_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%VPWR
x_PM_SKY130_FD_SC_HD__SDFXBP_2%A_560_369# N_A_560_369#_M1017_d
+ N_A_560_369#_M1024_s N_A_560_369#_M1010_d N_A_560_369#_M1015_s
+ N_A_560_369#_c_1782_n N_A_560_369#_c_1794_n N_A_560_369#_c_1806_n
+ N_A_560_369#_c_1771_n N_A_560_369#_c_1778_n N_A_560_369#_c_1779_n
+ N_A_560_369#_c_1772_n N_A_560_369#_c_1773_n N_A_560_369#_c_1774_n
+ N_A_560_369#_c_1775_n N_A_560_369#_c_1776_n N_A_560_369#_c_1777_n
+ N_A_560_369#_c_1781_n PM_SKY130_FD_SC_HD__SDFXBP_2%A_560_369#
x_PM_SKY130_FD_SC_HD__SDFXBP_2%Q N_Q_M1028_s N_Q_M1005_s N_Q_c_1895_n
+ N_Q_c_1892_n N_Q_c_1893_n Q N_Q_c_1911_n PM_SKY130_FD_SC_HD__SDFXBP_2%Q
x_PM_SKY130_FD_SC_HD__SDFXBP_2%Q_N N_Q_N_M1006_s N_Q_N_M1002_s N_Q_N_c_1933_n
+ N_Q_N_c_1934_n Q_N Q_N PM_SKY130_FD_SC_HD__SDFXBP_2%Q_N
x_PM_SKY130_FD_SC_HD__SDFXBP_2%VGND N_VGND_M1037_d N_VGND_M1039_d N_VGND_M1011_d
+ N_VGND_M1034_d N_VGND_M1003_d N_VGND_M1032_d N_VGND_M1029_d N_VGND_M1025_d
+ N_VGND_M1009_d N_VGND_c_1951_n N_VGND_c_1952_n N_VGND_c_1953_n N_VGND_c_1954_n
+ N_VGND_c_1955_n N_VGND_c_1956_n N_VGND_c_1957_n N_VGND_c_1958_n
+ N_VGND_c_1959_n N_VGND_c_1960_n N_VGND_c_1961_n N_VGND_c_1962_n VGND
+ N_VGND_c_1963_n N_VGND_c_1964_n N_VGND_c_1965_n N_VGND_c_1966_n
+ N_VGND_c_1967_n N_VGND_c_1968_n N_VGND_c_1969_n N_VGND_c_1970_n
+ N_VGND_c_1971_n N_VGND_c_1972_n N_VGND_c_1973_n N_VGND_c_1974_n
+ N_VGND_c_1975_n N_VGND_c_1976_n N_VGND_c_1977_n N_VGND_c_1978_n
+ PM_SKY130_FD_SC_HD__SDFXBP_2%VGND
cc_1 VNB N_CLK_c_246_n 0.0573151f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_247_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0185843f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_4 VNB N_A_27_47#_M1027_g 0.0381832f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1024_g 0.052087f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_6 VNB N_A_27_47#_c_290_n 0.0136466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_291_n 0.00249911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_292_n 0.0158261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1023_g 0.043789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_294_n 0.00319094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_295_n 0.00642096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_296_n 8.11193e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_297_n 0.00238722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_298_n 0.0228343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_299_n 0.00980602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_300_n 0.00148891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SCE_M1039_g 0.0506961f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_18 VNB N_SCE_M1021_g 0.016865f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_19 VNB N_SCE_c_537_n 0.00457617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_538_n 0.00290318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_539_n 0.00348269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_540_n 0.00118673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_541_n 0.0272673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_542_n 0.00148358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_299_47#_M1016_g 0.0216917f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_26 VNB N_A_299_47#_c_646_n 0.0137707f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_27 VNB N_A_299_47#_c_647_n 0.00262794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_299_47#_c_648_n 0.00249039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_299_47#_c_649_n 0.00285099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_299_47#_c_650_n 0.0299041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_D_M1017_g 0.0443856f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_32 VNB N_SCD_M1011_g 0.0447042f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_33 VNB SCD 0.0130762f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_34 VNB N_SCD_c_822_n 0.0127645f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_868_n 0.0180432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_869_n 0.00330396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_870_n 0.00369255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_871_n 0.00403969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_872_n 0.00632811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_873_n 0.0486971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_193_47#_c_874_n 0.00572932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_193_47#_c_875_n 0.0103972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_193_47#_c_876_n 0.0114429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_193_47#_c_877_n 6.97704e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_193_47#_c_878_n 0.0266741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_193_47#_c_879_n 0.005674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_880_n 0.0176138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_881_n 0.0285203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1097_183#_M1013_g 0.0146965f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_50 VNB N_A_1097_183#_M1034_g 0.0210316f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_51 VNB N_A_1097_183#_c_1085_n 0.00354578f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_52 VNB N_A_1097_183#_c_1086_n 0.00364457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1097_183#_c_1087_n 0.00130588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1097_183#_c_1088_n 0.00302393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1097_183#_c_1089_n 0.0338642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_938_413#_c_1178_n 0.0118275f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_57 VNB N_A_938_413#_c_1179_n 0.0158415f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_58 VNB N_A_938_413#_c_1180_n 0.0152351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_938_413#_c_1181_n 0.00913873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_938_413#_c_1182_n 8.51874e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_938_413#_c_1183_n 0.0118261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_938_413#_c_1184_n 0.00180949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1525_315#_M1003_g 0.0478726f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.105
cc_64 VNB N_A_1525_315#_c_1287_n 0.016402f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_65 VNB N_A_1525_315#_c_1288_n 0.0193862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1525_315#_c_1289_n 0.0451281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1525_315#_c_1290_n 0.030097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1525_315#_c_1291_n 0.0304242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1525_315#_c_1292_n 0.0179157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1525_315#_c_1293_n 0.00160611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1525_315#_c_1294_n 0.00373683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1525_315#_c_1295_n 0.00820384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1354_413#_c_1422_n 0.0203674f $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=2.135
cc_74 VNB N_A_1354_413#_c_1423_n 0.0412143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1354_413#_c_1424_n 0.00807206f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_76 VNB N_A_1354_413#_c_1425_n 0.00923861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1354_413#_c_1426_n 0.00584041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1354_413#_c_1427_n 0.00344545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_2049_47#_c_1509_n 0.0167328f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_80 VNB N_A_2049_47#_c_1510_n 0.0197001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_2049_47#_c_1511_n 0.00788325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_2049_47#_c_1512_n 0.00338009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_2049_47#_c_1513_n 0.0503595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VPWR_c_1578_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_560_369#_c_1771_n 2.29256e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_560_369#_c_1772_n 0.0115446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_560_369#_c_1773_n 0.00220658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_560_369#_c_1774_n 0.00348474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_560_369#_c_1775_n 0.00913814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_560_369#_c_1776_n 0.00243436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_560_369#_c_1777_n 0.00182555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_Q_c_1892_n 9.91593e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_Q_c_1893_n 3.20153e-19 $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_94 VNB Q_N 0.00103626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1951_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1952_n 0.00281433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1953_n 0.00486519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1954_n 0.0457659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1955_n 0.0058544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1956_n 0.00237946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1957_n 0.0217892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1958_n 0.00423032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1959_n 0.00898265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1960_n 0.00428548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1961_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1962_n 0.00964018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1963_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1964_n 0.0289225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1965_n 0.0346138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1966_n 0.0430904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1967_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1968_n 0.0204144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1969_n 0.0153766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1970_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1971_n 0.00512961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1972_n 0.00381885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1973_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1974_n 0.00513917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1975_n 0.00365128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1976_n 0.00442067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1977_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1978_n 0.570034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VPB N_CLK_c_246_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_124 VPB N_CLK_c_250_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_125 VPB N_CLK_c_251_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.74
cc_126 VPB N_CLK_c_252_n 0.0235707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_127 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.105
cc_128 VPB N_A_27_47#_M1036_g 0.03676f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.105
cc_129 VPB N_A_27_47#_c_290_n 0.0143056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_291_n 0.0052612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_M1000_g 0.0191311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_M1018_g 0.033754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_292_n 0.0210291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_307_n 0.00185683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_308_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_309_n 0.00356676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_310_n 0.0567661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_311_n 0.00130301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_312_n 0.00139996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_313_n 9.17012e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_314_n 0.00536377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_298_n 0.0115869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_316_n 0.0266783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_317_n 0.00853708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_318_n 0.0106236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_299_n 0.020895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_300_n 0.00437972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_SCE_M1030_g 0.0236254f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_149 VPB N_SCE_M1039_g 0.00509704f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.135
cc_150 VPB N_SCE_M1026_g 0.0196072f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_151 VPB N_SCE_c_537_n 0.00116063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_SCE_c_547_n 0.0437017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_299_47#_M1007_g 0.0184813f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.105
cc_154 VPB N_A_299_47#_c_646_n 0.010521f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_155 VPB N_A_299_47#_c_653_n 0.00406887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_299_47#_c_647_n 0.00417171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_299_47#_c_655_n 0.00158406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_299_47#_c_656_n 0.00180574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_299_47#_c_657_n 0.0014433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_299_47#_c_658_n 0.027856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_D_M1010_g 0.0192049f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_162 VPB N_D_M1017_g 0.00360779f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.135
cc_163 VPB N_D_c_774_n 0.0271103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_D_c_775_n 0.00449122f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.105
cc_165 VPB N_SCD_M1004_g 0.0328806f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.135
cc_166 VPB SCD 0.0103452f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_167 VPB N_SCD_c_822_n 0.018616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_193_47#_M1015_g 0.024991f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_169 VPB N_A_193_47#_M1008_g 0.0221869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_193_47#_c_869_n 0.00462988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_193_47#_c_885_n 0.0328226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_193_47#_c_870_n 0.00311128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_193_47#_c_887_n 0.00568216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_193_47#_c_888_n 0.0266658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_193_47#_c_876_n 0.0173137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1097_183#_M1013_g 0.049805f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_177 VPB N_A_1097_183#_c_1088_n 0.00255179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_938_413#_M1033_g 0.0226707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_179 VPB N_A_938_413#_c_1181_n 0.0189969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_938_413#_c_1182_n 0.00681499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_938_413#_c_1188_n 0.00161138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_938_413#_c_1184_n 0.00887906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1525_315#_M1031_g 0.025189f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_184 VPB N_A_1525_315#_M1003_g 0.0178898f $X=-0.19 $Y=1.305 $X2=0.155
+ $Y2=1.105
cc_185 VPB N_A_1525_315#_M1005_g 0.0190109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1525_315#_M1019_g 0.0222885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1525_315#_c_1289_n 0.0234771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1525_315#_c_1290_n 0.00739451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1525_315#_c_1291_n 5.42563e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1525_315#_M1038_g 0.0252846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1525_315#_c_1304_n 0.0126982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1525_315#_c_1305_n 0.0137898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1525_315#_c_1306_n 0.0118556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1525_315#_c_1307_n 0.0408358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_1525_315#_c_1308_n 0.00754758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1525_315#_c_1309_n 0.00234285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1525_315#_c_1294_n 0.00373683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1525_315#_c_1311_n 9.71818e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1354_413#_M1035_g 0.0235713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1354_413#_c_1423_n 0.0157151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1354_413#_c_1424_n 5.11281e-19 $X=-0.19 $Y=1.305 $X2=0.33
+ $Y2=1.16
cc_202 VPB N_A_1354_413#_c_1431_n 0.0126796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1354_413#_c_1425_n 0.00365405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1354_413#_c_1426_n 0.0050339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_2049_47#_M1002_g 0.0195085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_2049_47#_M1014_g 0.022964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_2049_47#_c_1516_n 0.0122047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_2049_47#_c_1512_n 0.00405051f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_2049_47#_c_1513_n 0.00886788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1579_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1580_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1581_n 0.00470486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1582_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1583_n 0.00548955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1584_n 0.0218906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1585_n 0.00474144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1586_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1587_n 0.00499301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1588_n 0.0111867f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1589_n 0.0105994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1590_n 0.0517085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1591_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1592_n 0.0190118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1593_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1594_n 0.0156572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1595_n 0.0255003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1596_n 0.0378453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1597_n 0.0449606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1598_n 0.0219039f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1599_n 0.0158909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1600_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1601_n 0.00436214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1602_n 0.00324297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1603_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1604_n 0.00343636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1605_n 0.00459796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1578_n 0.0730545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_560_369#_c_1778_n 0.00823319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_A_560_369#_c_1779_n 0.00155557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_560_369#_c_1775_n 0.0110678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_560_369#_c_1781_n 0.00997623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_Q_c_1892_n 0.0017899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB Q_N 0.00211514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 N_CLK_c_246_n N_A_27_47#_M1027_g 0.0049062f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_245 N_CLK_c_247_n N_A_27_47#_M1027_g 0.0187731f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_246 CLK N_A_27_47#_M1027_g 3.14819e-19 $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_247 N_CLK_c_250_n N_A_27_47#_M1036_g 0.00531917f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_248 N_CLK_c_252_n N_A_27_47#_M1036_g 0.0276478f $X=0.475 $Y=1.665 $X2=0 $Y2=0
cc_249 CLK N_A_27_47#_M1036_g 5.73308e-19 $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_250 N_CLK_c_246_n N_A_27_47#_c_294_n 0.00761961f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_251 N_CLK_c_247_n N_A_27_47#_c_294_n 0.00668648f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_252 CLK N_A_27_47#_c_294_n 0.00774265f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_253 N_CLK_c_246_n N_A_27_47#_c_295_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_254 CLK N_A_27_47#_c_295_n 0.0144574f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_255 N_CLK_c_251_n N_A_27_47#_c_307_n 0.0128144f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_256 N_CLK_c_252_n N_A_27_47#_c_307_n 0.0013816f $X=0.475 $Y=1.665 $X2=0 $Y2=0
cc_257 CLK N_A_27_47#_c_307_n 0.00728212f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_258 N_CLK_c_246_n N_A_27_47#_c_296_n 3.98708e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_259 CLK N_A_27_47#_c_296_n 0.0516739f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_260 N_CLK_c_246_n N_A_27_47#_c_308_n 2.90926e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_261 N_CLK_c_250_n N_A_27_47#_c_308_n 7.09762e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_262 N_CLK_c_252_n N_A_27_47#_c_308_n 0.00440146f $X=0.475 $Y=1.665 $X2=0
+ $Y2=0
cc_263 N_CLK_c_246_n N_A_27_47#_c_309_n 2.26313e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_264 N_CLK_c_251_n N_A_27_47#_c_309_n 2.17882e-19 $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_265 N_CLK_c_252_n N_A_27_47#_c_309_n 0.00358837f $X=0.475 $Y=1.665 $X2=0
+ $Y2=0
cc_266 CLK N_A_27_47#_c_309_n 0.0153364f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_267 N_CLK_c_246_n N_A_27_47#_c_297_n 0.00381855f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_268 N_CLK_c_251_n N_A_27_47#_c_311_n 0.00100908f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_269 N_CLK_c_246_n N_A_27_47#_c_298_n 0.0169285f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_270 CLK N_A_27_47#_c_298_n 0.00161876f $X=0.155 $Y=1.105 $X2=0 $Y2=0
cc_271 N_CLK_c_251_n N_VPWR_c_1579_n 0.00946555f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_272 N_CLK_c_251_n N_VPWR_c_1594_n 0.00332278f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_273 N_CLK_c_251_n N_VPWR_c_1578_n 0.00485269f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_274 N_CLK_c_247_n N_VGND_c_1951_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_275 N_CLK_c_246_n N_VGND_c_1963_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_276 N_CLK_c_247_n N_VGND_c_1963_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_277 N_CLK_c_247_n N_VGND_c_1978_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_310_n N_SCE_M1030_g 0.00319643f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_310_n N_SCE_M1026_g 0.00116169f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_310_n N_SCE_c_537_n 0.00414929f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_310_n N_SCE_c_547_n 0.00341967f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_310_n N_A_299_47#_M1007_g 7.69535e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_310_n N_A_299_47#_c_646_n 0.0120648f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_310_n N_A_299_47#_c_661_n 0.0163793f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_310_n N_A_299_47#_c_647_n 0.00933005f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_310_n N_A_299_47#_c_663_n 0.0369342f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_310_n N_A_299_47#_c_655_n 0.0113096f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1027_g N_A_299_47#_c_648_n 9.61905e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_310_n N_A_299_47#_c_656_n 0.0130054f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_310_n N_A_299_47#_c_650_n 0.00287433f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_310_n N_A_299_47#_c_668_n 0.0046527f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_310_n N_A_299_47#_c_657_n 7.81108e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_310_n N_A_299_47#_c_658_n 0.0016565f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_310_n N_D_M1010_g 0.00219328f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_310_n N_D_c_774_n 0.00308822f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_310_n N_D_c_775_n 0.0085184f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_310_n N_SCD_M1004_g 0.00188492f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_310_n SCD 0.0127788f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_310_n N_A_193_47#_M1036_d 6.81311e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_310_n N_A_193_47#_M1015_g 0.00371812f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_316_n N_A_193_47#_M1015_g 0.014411f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_317_n N_A_193_47#_M1015_g 9.60176e-19 $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_M1023_g N_A_193_47#_c_868_n 0.0144677f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_M1018_g N_A_193_47#_M1008_g 0.0175056f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_314_n N_A_193_47#_M1008_g 0.00136781f $X=6.71 $Y=1.87 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_300_n N_A_193_47#_M1008_g 5.16255e-19 $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1024_g N_A_193_47#_c_869_n 0.00772368f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_290_n N_A_193_47#_c_869_n 0.00687115f $X=5.005 $Y=1.32 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_291_n N_A_193_47#_c_869_n 0.00418731f $X=4.695 $Y=1.32 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_310_n N_A_193_47#_c_869_n 0.0139192f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_313_n N_A_193_47#_c_869_n 2.15174e-19 $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_316_n N_A_193_47#_c_869_n 7.29366e-19 $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_317_n N_A_193_47#_c_869_n 0.0168988f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_318_n N_A_193_47#_c_869_n 0.00604391f $X=5.14 $Y=1.575 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_291_n N_A_193_47#_c_885_n 0.0162569f $X=4.695 $Y=1.32 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_310_n N_A_193_47#_c_885_n 0.00545515f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_316_n N_A_193_47#_c_885_n 0.0174998f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_317_n N_A_193_47#_c_885_n 0.00118389f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_292_n N_A_193_47#_c_870_n 0.0117161f $X=7.265 $Y=1.32 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_M1023_g N_A_193_47#_c_870_n 0.00430042f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_299_n N_A_193_47#_c_870_n 0.00402309f $X=6.69 $Y=1.32 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_300_n N_A_193_47#_c_870_n 0.0234373f $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1027_g N_A_193_47#_c_871_n 0.00136529f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_294_n N_A_193_47#_c_871_n 0.00442897f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1023_g N_A_193_47#_c_872_n 0.0020279f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_299_n N_A_193_47#_c_872_n 0.00222109f $X=6.69 $Y=1.32 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_300_n N_A_193_47#_c_872_n 0.0119224f $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_M1018_g N_A_193_47#_c_887_n 0.00117691f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_292_n N_A_193_47#_c_887_n 0.00338756f $X=7.265 $Y=1.32 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_314_n N_A_193_47#_c_887_n 0.00513984f $X=6.71 $Y=1.87 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_300_n N_A_193_47#_c_887_n 0.0245563f $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_M1018_g N_A_193_47#_c_888_n 0.0130792f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_292_n N_A_193_47#_c_888_n 0.0212127f $X=7.265 $Y=1.32 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_300_n N_A_193_47#_c_888_n 6.54911e-19 $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_M1024_g N_A_193_47#_c_873_n 0.00225641f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_M1027_g N_A_193_47#_c_874_n 0.00662116f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_294_n N_A_193_47#_c_874_n 0.0022123f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_297_n N_A_193_47#_c_874_n 0.00516669f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_299_n N_A_193_47#_c_875_n 5.41218e-19 $X=6.69 $Y=1.32 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1027_g N_A_193_47#_c_876_n 0.00851768f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_294_n N_A_193_47#_c_876_n 0.0055484f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_296_n N_A_193_47#_c_876_n 0.0597663f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_413_p N_A_193_47#_c_876_n 0.00826639f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_297_n N_A_193_47#_c_876_n 0.00884862f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_310_n N_A_193_47#_c_876_n 0.0247251f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_311_n N_A_193_47#_c_876_n 0.00246357f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_298_n N_A_193_47#_c_876_n 0.0174894f $X=0.895 $Y=1.235 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_299_n N_A_193_47#_c_877_n 6.19017e-19 $X=6.69 $Y=1.32 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_300_n N_A_193_47#_c_877_n 0.00125233f $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_M1024_g N_A_193_47#_c_878_n 0.0213105f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_290_n N_A_193_47#_c_878_n 0.0174066f $X=5.005 $Y=1.32 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_316_n N_A_193_47#_c_878_n 5.43883e-19 $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_317_n N_A_193_47#_c_878_n 4.76262e-19 $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_M1024_g N_A_193_47#_c_879_n 0.0116468f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_290_n N_A_193_47#_c_879_n 0.00587088f $X=5.005 $Y=1.32 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_317_n N_A_193_47#_c_879_n 0.00398178f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_M1024_g N_A_193_47#_c_880_n 0.0102604f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1023_g N_A_193_47#_c_881_n 0.0193601f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_299_n N_A_193_47#_c_881_n 0.020308f $X=6.69 $Y=1.32 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_312_n N_A_1097_183#_M1033_d 0.00523078f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_290_n N_A_1097_183#_M1013_g 0.0113457f $X=5.005 $Y=1.32
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_M1000_g N_A_1097_183#_M1013_g 0.0276008f $X=5.08 $Y=2.275
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_312_n N_A_1097_183#_M1013_g 0.00281129f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_313_n N_A_1097_183#_M1013_g 0.00148824f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_316_n N_A_1097_183#_M1013_g 0.0206011f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_317_n N_A_1097_183#_M1013_g 0.0022f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_312_n N_A_1097_183#_c_1099_n 0.00261642f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_M1018_g N_A_1097_183#_c_1088_n 0.00455971f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_312_n N_A_1097_183#_c_1088_n 0.0193938f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_314_n N_A_1097_183#_c_1088_n 0.00311096f $X=6.71 $Y=1.87
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_299_n N_A_1097_183#_c_1088_n 0.00225153f $X=6.69 $Y=1.32
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_300_n N_A_1097_183#_c_1088_n 0.0517157f $X=6.69 $Y=1.41
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_299_n N_A_938_413#_c_1178_n 0.0158005f $X=6.69 $Y=1.32 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_300_n N_A_938_413#_c_1178_n 3.03019e-19 $X=6.69 $Y=1.41
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_M1018_g N_A_938_413#_M1033_g 0.0247799f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_312_n N_A_938_413#_M1033_g 0.00700233f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_300_n N_A_938_413#_M1033_g 8.29633e-19 $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_312_n N_A_938_413#_c_1181_n 0.00109659f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_M1000_g N_A_938_413#_c_1196_n 0.00859863f $X=5.08 $Y=2.275
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_310_n N_A_938_413#_c_1196_n 0.00699281f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_312_n N_A_938_413#_c_1196_n 0.00369623f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_313_n N_A_938_413#_c_1196_n 0.00172439f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_316_n N_A_938_413#_c_1196_n 5.38487e-19 $X=5.14 $Y=1.74
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_317_n N_A_938_413#_c_1196_n 0.0252832f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1024_g N_A_938_413#_c_1183_n 9.86268e-19 $X=4.62 $Y=0.415
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_290_n N_A_938_413#_c_1183_n 8.14452e-19 $X=5.005 $Y=1.32
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_M1000_g N_A_938_413#_c_1188_n 9.97608e-19 $X=5.08 $Y=2.275
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_312_n N_A_938_413#_c_1188_n 0.0183205f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_313_n N_A_938_413#_c_1188_n 0.00258875f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_316_n N_A_938_413#_c_1188_n 7.00613e-19 $X=5.14 $Y=1.74
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_317_n N_A_938_413#_c_1188_n 0.0250097f $X=5.14 $Y=1.74 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_290_n N_A_938_413#_c_1184_n 0.00225879f $X=5.005 $Y=1.32
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_312_n N_A_938_413#_c_1184_n 0.0173913f $X=6.565 $Y=1.87
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_313_n N_A_938_413#_c_1184_n 0.00179088f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_317_n N_A_938_413#_c_1184_n 0.00980238f $X=5.14 $Y=1.74
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_318_n N_A_938_413#_c_1184_n 4.44848e-19 $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_M1023_g N_A_1525_315#_M1003_g 0.0463015f $X=7.34 $Y=0.415
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_M1018_g N_A_1354_413#_c_1434_n 0.00281529f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_314_n N_A_1354_413#_c_1434_n 0.00241029f $X=6.71 $Y=1.87
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_300_n N_A_1354_413#_c_1434_n 0.0022468f $X=6.69 $Y=1.41
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_M1023_g N_A_1354_413#_c_1437_n 0.00800808f $X=7.34 $Y=0.415
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_314_n N_A_1354_413#_c_1431_n 0.00230468f $X=6.71 $Y=1.87
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_300_n N_A_1354_413#_c_1431_n 9.59883e-19 $X=6.69 $Y=1.41
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_M1023_g N_A_1354_413#_c_1425_n 3.1587e-19 $X=7.34 $Y=0.415
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_292_n N_A_1354_413#_c_1426_n 0.00558094f $X=7.265 $Y=1.32
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_M1023_g N_A_1354_413#_c_1426_n 0.0061466f $X=7.34 $Y=0.415
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_M1023_g N_A_1354_413#_c_1427_n 0.0110507f $X=7.34 $Y=0.415
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_413_p N_VPWR_M1012_d 6.91013e-19 $X=0.73 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_409 N_A_27_47#_c_311_n N_VPWR_M1012_d 0.0017551f $X=0.875 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_410 N_A_27_47#_c_312_n N_VPWR_M1013_d 0.00678497f $X=6.565 $Y=1.87 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_M1036_g N_VPWR_c_1579_n 0.00937841f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_307_n N_VPWR_c_1579_n 0.0030205f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_413_p N_VPWR_c_1579_n 0.0133497f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_309_n N_VPWR_c_1579_n 0.012721f $X=0.265 $Y=1.96 $X2=0 $Y2=0
cc_415 N_A_27_47#_c_311_n N_VPWR_c_1579_n 0.00324852f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_310_n N_VPWR_c_1580_n 0.00123614f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_310_n N_VPWR_c_1581_n 8.00522e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_312_n N_VPWR_c_1582_n 0.00950843f $X=6.565 $Y=1.87 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_M1000_g N_VPWR_c_1590_n 0.0037886f $X=5.08 $Y=2.275 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_307_n N_VPWR_c_1594_n 0.0018545f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_309_n N_VPWR_c_1594_n 0.0120313f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1036_g N_VPWR_c_1595_n 0.00442511f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_M1018_g N_VPWR_c_1597_n 0.00430107f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_300_n N_VPWR_c_1597_n 0.00157744f $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_M1036_g N_VPWR_c_1578_n 0.0053417f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_M1000_g N_VPWR_c_1578_n 0.00557377f $X=5.08 $Y=2.275 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_M1018_g N_VPWR_c_1578_n 0.0057371f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_307_n N_VPWR_c_1578_n 0.00405127f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_309_n N_VPWR_c_1578_n 0.00646745f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_310_n N_VPWR_c_1578_n 0.198964f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_431 N_A_27_47#_c_311_n N_VPWR_c_1578_n 0.014581f $X=0.875 $Y=1.87 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_312_n N_VPWR_c_1578_n 0.0535471f $X=6.565 $Y=1.87 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_313_n N_VPWR_c_1578_n 0.0147031f $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_314_n N_VPWR_c_1578_n 0.0159163f $X=6.71 $Y=1.87 $X2=0 $Y2=0
cc_435 N_A_27_47#_c_300_n N_VPWR_c_1578_n 0.00100625f $X=6.69 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_310_n N_A_560_369#_c_1782_n 0.00584375f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_310_n N_A_560_369#_c_1778_n 0.022293f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_310_n N_A_560_369#_c_1779_n 0.0102354f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_M1024_g N_A_560_369#_c_1774_n 0.0044467f $X=4.62 $Y=0.415
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_M1024_g N_A_560_369#_c_1775_n 0.00902644f $X=4.62 $Y=0.415
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_310_n N_A_560_369#_c_1775_n 0.0104876f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_M1024_g N_A_560_369#_c_1776_n 0.00178202f $X=4.62 $Y=0.415
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_M1024_g N_A_560_369#_c_1777_n 0.00164257f $X=4.62 $Y=0.415
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_310_n N_A_560_369#_c_1781_n 0.0126037f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_317_n N_A_560_369#_c_1781_n 0.00314032f $X=5.14 $Y=1.74
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_310_n A_644_369# 0.00134881f $X=5.145 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_447 N_A_27_47#_c_294_n N_VGND_M1037_d 0.00166329f $X=0.615 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_448 N_A_27_47#_M1027_g N_VGND_c_1951_n 0.0100209f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_294_n N_VGND_c_1951_n 0.0150403f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_296_n N_VGND_c_1951_n 0.00108069f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_298_n N_VGND_c_1951_n 5.70216e-19 $X=0.895 $Y=1.235 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_M1024_g N_VGND_c_1953_n 0.00344097f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1024_g N_VGND_c_1954_n 0.00431421f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_M1023_g N_VGND_c_1956_n 0.00230753f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_525_p N_VGND_c_1963_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_294_n N_VGND_c_1963_n 0.00243651f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_M1027_g N_VGND_c_1964_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_M1023_g N_VGND_c_1966_n 0.00379696f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_M1037_s N_VGND_c_1978_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_M1027_g N_VGND_c_1978_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_M1024_g N_VGND_c_1978_n 0.00721503f $X=4.62 $Y=0.415 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_M1023_g N_VGND_c_1978_n 0.00575728f $X=7.34 $Y=0.415 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_525_p N_VGND_c_1978_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_294_n N_VGND_c_1978_n 0.00564532f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_465 N_SCE_M1039_g N_A_299_47#_M1016_g 0.0204373f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_466 N_SCE_c_537_n N_A_299_47#_M1016_g 0.00147314f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_467 N_SCE_c_538_n N_A_299_47#_M1016_g 0.0107276f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_468 N_SCE_M1030_g N_A_299_47#_c_646_n 0.00433634f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_469 N_SCE_M1039_g N_A_299_47#_c_646_n 0.0181395f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_470 N_SCE_c_537_n N_A_299_47#_c_646_n 0.0621897f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_471 N_SCE_c_547_n N_A_299_47#_c_646_n 0.00715683f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_472 N_SCE_c_559_p N_A_299_47#_c_646_n 0.0130375f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_473 N_SCE_M1030_g N_A_299_47#_c_661_n 0.0125417f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_474 N_SCE_c_537_n N_A_299_47#_c_661_n 0.0103251f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_475 N_SCE_c_547_n N_A_299_47#_c_661_n 0.0039772f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_476 N_SCE_M1030_g N_A_299_47#_c_647_n 0.00142881f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_477 N_SCE_M1039_g N_A_299_47#_c_647_n 0.00145274f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_478 N_SCE_M1026_g N_A_299_47#_c_647_n 0.00581038f $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_479 N_SCE_c_537_n N_A_299_47#_c_647_n 0.0405813f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_480 N_SCE_c_547_n N_A_299_47#_c_647_n 0.00894616f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_481 N_SCE_M1026_g N_A_299_47#_c_663_n 0.00531583f $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_482 N_SCE_M1039_g N_A_299_47#_c_648_n 0.00239556f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_483 N_SCE_c_559_p N_A_299_47#_c_648_n 0.00168685f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_484 N_SCE_c_547_n N_A_299_47#_c_656_n 2.83838e-19 $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_485 N_SCE_M1039_g N_A_299_47#_c_649_n 5.26825e-19 $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_SCE_c_537_n N_A_299_47#_c_649_n 0.0134242f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_487 N_SCE_c_547_n N_A_299_47#_c_649_n 3.95711e-19 $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_488 N_SCE_c_538_n N_A_299_47#_c_649_n 0.0208599f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_489 N_SCE_c_540_n N_A_299_47#_c_649_n 0.00389077f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_490 N_SCE_M1039_g N_A_299_47#_c_650_n 0.0174183f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_491 N_SCE_c_537_n N_A_299_47#_c_650_n 0.00156762f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_492 N_SCE_c_547_n N_A_299_47#_c_650_n 0.00745174f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_493 N_SCE_c_538_n N_A_299_47#_c_650_n 0.00319888f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_494 N_SCE_M1026_g N_A_299_47#_c_668_n 0.00695809f $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_495 N_SCE_c_540_n N_A_299_47#_c_657_n 0.00959271f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_496 N_SCE_c_541_n N_A_299_47#_c_657_n 3.983e-19 $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_497 N_SCE_c_540_n N_A_299_47#_c_658_n 2.12418e-19 $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_498 N_SCE_c_541_n N_A_299_47#_c_658_n 0.0144723f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_499 N_SCE_M1026_g N_D_M1010_g 0.0370747f $X=2.255 $Y=2.165 $X2=0 $Y2=0
cc_500 N_SCE_M1021_g N_D_M1017_g 0.0137065f $X=3.23 $Y=0.445 $X2=0 $Y2=0
cc_501 N_SCE_c_539_n N_D_M1017_g 0.0126031f $X=3.085 $Y=0.7 $X2=0 $Y2=0
cc_502 N_SCE_c_540_n N_D_M1017_g 0.00203037f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_503 N_SCE_c_541_n N_D_M1017_g 0.0213831f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_504 N_SCE_M1039_g N_D_c_774_n 3.44894e-19 $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_505 N_SCE_c_547_n N_D_c_774_n 0.0112854f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_506 N_SCE_c_539_n N_D_c_774_n 8.44684e-19 $X=3.085 $Y=0.7 $X2=0 $Y2=0
cc_507 N_SCE_c_542_n N_D_c_774_n 0.0011605f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_508 N_SCE_c_547_n N_D_c_775_n 0.00125504f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_509 N_SCE_c_539_n N_D_c_775_n 0.00197762f $X=3.085 $Y=0.7 $X2=0 $Y2=0
cc_510 N_SCE_c_542_n N_D_c_775_n 0.00315365f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_511 N_SCE_M1021_g N_SCD_M1011_g 0.0572953f $X=3.23 $Y=0.445 $X2=0 $Y2=0
cc_512 N_SCE_c_540_n N_SCD_M1011_g 0.00138865f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_513 N_SCE_c_540_n SCD 0.00392926f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_514 N_SCE_c_541_n SCD 2.85078e-19 $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_515 N_SCE_M1039_g N_A_193_47#_c_873_n 0.00255572f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_516 N_SCE_M1021_g N_A_193_47#_c_873_n 5.27825e-19 $X=3.23 $Y=0.445 $X2=0
+ $Y2=0
cc_517 N_SCE_c_537_n N_A_193_47#_c_873_n 0.0167276f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_518 N_SCE_c_547_n N_A_193_47#_c_873_n 0.0049774f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_519 N_SCE_c_538_n N_A_193_47#_c_873_n 0.0166296f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_520 N_SCE_c_559_p N_A_193_47#_c_873_n 0.00356182f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_521 N_SCE_c_539_n N_A_193_47#_c_873_n 0.0205248f $X=3.085 $Y=0.7 $X2=0 $Y2=0
cc_522 N_SCE_c_540_n N_A_193_47#_c_873_n 0.0108868f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_523 N_SCE_c_541_n N_A_193_47#_c_873_n 0.0037338f $X=3.17 $Y=0.95 $X2=0 $Y2=0
cc_524 N_SCE_c_542_n N_A_193_47#_c_873_n 0.00735012f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_525 N_SCE_M1030_g N_A_193_47#_c_876_n 0.00160127f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_526 N_SCE_M1030_g N_VPWR_c_1580_n 0.0086701f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_527 N_SCE_M1026_g N_VPWR_c_1580_n 0.00953157f $X=2.255 $Y=2.165 $X2=0 $Y2=0
cc_528 N_SCE_M1030_g N_VPWR_c_1595_n 0.00340533f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_529 N_SCE_M1026_g N_VPWR_c_1596_n 0.00340456f $X=2.255 $Y=2.165 $X2=0 $Y2=0
cc_530 N_SCE_M1030_g N_VPWR_c_1578_n 0.00515557f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_531 N_SCE_M1026_g N_VPWR_c_1578_n 0.00392879f $X=2.255 $Y=2.165 $X2=0 $Y2=0
cc_532 N_SCE_c_539_n N_A_560_369#_M1017_d 0.00218892f $X=3.085 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_533 N_SCE_M1026_g N_A_560_369#_c_1782_n 5.73988e-19 $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_534 N_SCE_M1021_g N_A_560_369#_c_1794_n 0.00763758f $X=3.23 $Y=0.445 $X2=0
+ $Y2=0
cc_535 N_SCE_c_539_n N_A_560_369#_c_1794_n 0.0207306f $X=3.085 $Y=0.7 $X2=0
+ $Y2=0
cc_536 N_SCE_c_541_n N_A_560_369#_c_1794_n 2.32966e-19 $X=3.17 $Y=0.95 $X2=0
+ $Y2=0
cc_537 N_SCE_M1021_g N_A_560_369#_c_1771_n 0.00405684f $X=3.23 $Y=0.445 $X2=0
+ $Y2=0
cc_538 N_SCE_c_539_n N_A_560_369#_c_1771_n 0.00630259f $X=3.085 $Y=0.7 $X2=0
+ $Y2=0
cc_539 N_SCE_M1021_g N_A_560_369#_c_1773_n 9.7798e-19 $X=3.23 $Y=0.445 $X2=0
+ $Y2=0
cc_540 N_SCE_c_539_n N_A_560_369#_c_1773_n 0.00793437f $X=3.085 $Y=0.7 $X2=0
+ $Y2=0
cc_541 N_SCE_c_540_n N_A_560_369#_c_1773_n 0.00554533f $X=3.17 $Y=0.95 $X2=0
+ $Y2=0
cc_542 N_SCE_c_538_n N_VGND_M1039_d 0.00250602f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_543 N_SCE_M1039_g N_VGND_c_1952_n 0.00411511f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_544 N_SCE_c_538_n N_VGND_c_1952_n 0.0185636f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_545 N_SCE_M1039_g N_VGND_c_1964_n 0.00409976f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_546 N_SCE_c_559_p N_VGND_c_1964_n 0.00251644f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_547 N_SCE_M1021_g N_VGND_c_1965_n 0.00362032f $X=3.23 $Y=0.445 $X2=0 $Y2=0
cc_548 N_SCE_c_538_n N_VGND_c_1965_n 0.00263191f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_549 N_SCE_c_539_n N_VGND_c_1965_n 0.00274476f $X=3.085 $Y=0.7 $X2=0 $Y2=0
cc_550 SCE N_VGND_c_1965_n 0.00782706f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_551 N_SCE_M1039_g N_VGND_c_1978_n 0.00687529f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_552 N_SCE_M1021_g N_VGND_c_1978_n 0.00526606f $X=3.23 $Y=0.445 $X2=0 $Y2=0
cc_553 N_SCE_c_538_n N_VGND_c_1978_n 0.00307132f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_554 N_SCE_c_559_p N_VGND_c_1978_n 0.00183549f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_555 N_SCE_c_539_n N_VGND_c_1978_n 0.00232388f $X=3.085 $Y=0.7 $X2=0 $Y2=0
cc_556 SCE N_VGND_c_1978_n 0.00302552f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_557 SCE A_487_47# 0.00226988f $X=2.475 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_558 N_A_299_47#_M1007_g N_D_M1010_g 0.028319f $X=3.145 $Y=2.165 $X2=0 $Y2=0
cc_559 N_A_299_47#_c_647_n N_D_M1010_g 0.00113649f $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_560 N_A_299_47#_c_663_n N_D_M1010_g 0.0119158f $X=3.08 $Y=1.967 $X2=0 $Y2=0
cc_561 N_A_299_47#_c_655_n N_D_M1010_g 0.00126571f $X=3.165 $Y=1.86 $X2=0 $Y2=0
cc_562 N_A_299_47#_M1016_g N_D_M1017_g 0.0412183f $X=2.36 $Y=0.445 $X2=0 $Y2=0
cc_563 N_A_299_47#_c_647_n N_D_M1017_g 0.00512253f $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_564 N_A_299_47#_c_649_n N_D_M1017_g 6.95345e-19 $X=2.3 $Y=1.04 $X2=0 $Y2=0
cc_565 N_A_299_47#_c_650_n N_D_M1017_g 0.0168474f $X=2.3 $Y=1.04 $X2=0 $Y2=0
cc_566 N_A_299_47#_c_647_n N_D_c_774_n 6.06547e-19 $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_567 N_A_299_47#_c_663_n N_D_c_774_n 0.00290918f $X=3.08 $Y=1.967 $X2=0 $Y2=0
cc_568 N_A_299_47#_c_657_n N_D_c_774_n 0.0011165f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_569 N_A_299_47#_c_658_n N_D_c_774_n 0.0197807f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_570 N_A_299_47#_c_647_n N_D_c_775_n 0.0254462f $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_571 N_A_299_47#_c_663_n N_D_c_775_n 0.0199968f $X=3.08 $Y=1.967 $X2=0 $Y2=0
cc_572 N_A_299_47#_c_649_n N_D_c_775_n 2.73452e-19 $X=2.3 $Y=1.04 $X2=0 $Y2=0
cc_573 N_A_299_47#_c_657_n N_D_c_775_n 0.0157256f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_574 N_A_299_47#_c_658_n N_D_c_775_n 0.00104184f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_575 N_A_299_47#_M1007_g N_SCD_M1004_g 0.0359024f $X=3.145 $Y=2.165 $X2=0
+ $Y2=0
cc_576 N_A_299_47#_c_663_n N_SCD_M1004_g 2.17192e-19 $X=3.08 $Y=1.967 $X2=0
+ $Y2=0
cc_577 N_A_299_47#_c_655_n N_SCD_M1004_g 0.002483f $X=3.165 $Y=1.86 $X2=0 $Y2=0
cc_578 N_A_299_47#_c_657_n SCD 0.0159098f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_579 N_A_299_47#_c_658_n SCD 0.00104233f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_580 N_A_299_47#_c_657_n N_SCD_c_822_n 3.53677e-19 $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_581 N_A_299_47#_c_658_n N_SCD_c_822_n 0.0204284f $X=3.19 $Y=1.52 $X2=0 $Y2=0
cc_582 N_A_299_47#_c_646_n N_A_193_47#_c_871_n 0.0978547f $X=1.52 $Y=1.86 $X2=0
+ $Y2=0
cc_583 N_A_299_47#_c_648_n N_A_193_47#_c_871_n 0.00751783f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_584 N_A_299_47#_M1016_g N_A_193_47#_c_873_n 0.00170787f $X=2.36 $Y=0.445
+ $X2=0 $Y2=0
cc_585 N_A_299_47#_c_646_n N_A_193_47#_c_873_n 0.0181188f $X=1.52 $Y=1.86 $X2=0
+ $Y2=0
cc_586 N_A_299_47#_c_648_n N_A_193_47#_c_873_n 0.00465031f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_587 N_A_299_47#_c_649_n N_A_193_47#_c_873_n 0.00873594f $X=2.3 $Y=1.04 $X2=0
+ $Y2=0
cc_588 N_A_299_47#_c_650_n N_A_193_47#_c_873_n 0.00457609f $X=2.3 $Y=1.04 $X2=0
+ $Y2=0
cc_589 N_A_299_47#_c_657_n N_A_193_47#_c_873_n 0.00166362f $X=3.19 $Y=1.52 $X2=0
+ $Y2=0
cc_590 N_A_299_47#_c_658_n N_A_193_47#_c_873_n 6.70678e-19 $X=3.19 $Y=1.52 $X2=0
+ $Y2=0
cc_591 N_A_299_47#_c_646_n N_A_193_47#_c_874_n 0.00264809f $X=1.52 $Y=1.86 $X2=0
+ $Y2=0
cc_592 N_A_299_47#_c_653_n N_A_193_47#_c_876_n 0.0272627f $X=1.625 $Y=2.175
+ $X2=0 $Y2=0
cc_593 N_A_299_47#_c_656_n N_A_193_47#_c_876_n 0.0158132f $X=1.572 $Y=1.967
+ $X2=0 $Y2=0
cc_594 N_A_299_47#_c_661_n N_VPWR_M1030_d 0.00416053f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_595 N_A_299_47#_c_661_n N_VPWR_c_1580_n 0.0128774f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_596 N_A_299_47#_c_668_n N_VPWR_c_1580_n 0.00214536f $X=2.205 $Y=1.967 $X2=0
+ $Y2=0
cc_597 N_A_299_47#_c_653_n N_VPWR_c_1595_n 0.0168466f $X=1.625 $Y=2.175 $X2=0
+ $Y2=0
cc_598 N_A_299_47#_c_661_n N_VPWR_c_1595_n 0.00240758f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_599 N_A_299_47#_M1007_g N_VPWR_c_1596_n 0.00368123f $X=3.145 $Y=2.165 $X2=0
+ $Y2=0
cc_600 N_A_299_47#_c_663_n N_VPWR_c_1596_n 0.00604259f $X=3.08 $Y=1.967 $X2=0
+ $Y2=0
cc_601 N_A_299_47#_c_668_n N_VPWR_c_1596_n 0.00138725f $X=2.205 $Y=1.967 $X2=0
+ $Y2=0
cc_602 N_A_299_47#_M1030_s N_VPWR_c_1578_n 0.00184114f $X=1.5 $Y=1.845 $X2=0
+ $Y2=0
cc_603 N_A_299_47#_M1007_g N_VPWR_c_1578_n 0.00535446f $X=3.145 $Y=2.165 $X2=0
+ $Y2=0
cc_604 N_A_299_47#_c_653_n N_VPWR_c_1578_n 0.00494372f $X=1.625 $Y=2.175 $X2=0
+ $Y2=0
cc_605 N_A_299_47#_c_661_n N_VPWR_c_1578_n 0.00247958f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_606 N_A_299_47#_c_663_n N_VPWR_c_1578_n 0.00555531f $X=3.08 $Y=1.967 $X2=0
+ $Y2=0
cc_607 N_A_299_47#_c_668_n N_VPWR_c_1578_n 0.00120782f $X=2.205 $Y=1.967 $X2=0
+ $Y2=0
cc_608 N_A_299_47#_c_663_n A_466_369# 0.00555859f $X=3.08 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_609 N_A_299_47#_c_663_n N_A_560_369#_M1010_d 0.00427378f $X=3.08 $Y=1.967
+ $X2=0 $Y2=0
cc_610 N_A_299_47#_M1007_g N_A_560_369#_c_1782_n 0.00811134f $X=3.145 $Y=2.165
+ $X2=0 $Y2=0
cc_611 N_A_299_47#_c_663_n N_A_560_369#_c_1782_n 0.0265702f $X=3.08 $Y=1.967
+ $X2=0 $Y2=0
cc_612 N_A_299_47#_c_658_n N_A_560_369#_c_1782_n 0.0012413f $X=3.19 $Y=1.52
+ $X2=0 $Y2=0
cc_613 N_A_299_47#_M1007_g N_A_560_369#_c_1806_n 0.00367162f $X=3.145 $Y=2.165
+ $X2=0 $Y2=0
cc_614 N_A_299_47#_M1007_g N_A_560_369#_c_1779_n 5.41855e-19 $X=3.145 $Y=2.165
+ $X2=0 $Y2=0
cc_615 N_A_299_47#_c_663_n N_A_560_369#_c_1779_n 0.00683183f $X=3.08 $Y=1.967
+ $X2=0 $Y2=0
cc_616 N_A_299_47#_c_655_n N_A_560_369#_c_1779_n 0.00221463f $X=3.165 $Y=1.86
+ $X2=0 $Y2=0
cc_617 N_A_299_47#_c_648_n N_VGND_c_1951_n 0.002159f $X=1.64 $Y=0.36 $X2=0 $Y2=0
cc_618 N_A_299_47#_M1016_g N_VGND_c_1952_n 0.00745268f $X=2.36 $Y=0.445 $X2=0
+ $Y2=0
cc_619 N_A_299_47#_c_648_n N_VGND_c_1964_n 0.0193961f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_620 N_A_299_47#_M1016_g N_VGND_c_1965_n 0.00365142f $X=2.36 $Y=0.445 $X2=0
+ $Y2=0
cc_621 N_A_299_47#_M1039_s N_VGND_c_1978_n 0.00186585f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_622 N_A_299_47#_M1016_g N_VGND_c_1978_n 0.00396023f $X=2.36 $Y=0.445 $X2=0
+ $Y2=0
cc_623 N_A_299_47#_c_648_n N_VGND_c_1978_n 0.00613328f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_624 N_D_M1017_g N_SCD_M1011_g 0.00367381f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_625 N_D_M1017_g N_A_193_47#_c_873_n 0.00435815f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_626 N_D_c_774_n N_A_193_47#_c_873_n 0.00255857f $X=2.71 $Y=1.52 $X2=0 $Y2=0
cc_627 N_D_c_775_n N_A_193_47#_c_873_n 0.00706402f $X=2.71 $Y=1.52 $X2=0 $Y2=0
cc_628 N_D_M1010_g N_VPWR_c_1580_n 0.00181754f $X=2.725 $Y=2.165 $X2=0 $Y2=0
cc_629 N_D_M1010_g N_VPWR_c_1596_n 0.00385655f $X=2.725 $Y=2.165 $X2=0 $Y2=0
cc_630 N_D_M1010_g N_VPWR_c_1578_n 0.00548378f $X=2.725 $Y=2.165 $X2=0 $Y2=0
cc_631 N_D_M1010_g N_A_560_369#_c_1782_n 0.00619595f $X=2.725 $Y=2.165 $X2=0
+ $Y2=0
cc_632 N_D_M1017_g N_A_560_369#_c_1794_n 0.00166377f $X=2.75 $Y=0.445 $X2=0
+ $Y2=0
cc_633 N_D_M1017_g N_VGND_c_1952_n 0.00138865f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_634 N_D_M1017_g N_VGND_c_1965_n 0.0042011f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_635 N_D_M1017_g N_VGND_c_1978_n 0.00560912f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_636 N_SCD_M1011_g N_A_193_47#_c_873_n 0.00245438f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_637 SCD N_A_193_47#_c_873_n 0.0132488f $X=3.855 $Y=1.105 $X2=0 $Y2=0
cc_638 N_SCD_M1004_g N_VPWR_c_1581_n 0.00615911f $X=3.61 $Y=2.165 $X2=0 $Y2=0
cc_639 N_SCD_M1004_g N_VPWR_c_1596_n 0.00412211f $X=3.61 $Y=2.165 $X2=0 $Y2=0
cc_640 N_SCD_M1004_g N_VPWR_c_1578_n 0.00690372f $X=3.61 $Y=2.165 $X2=0 $Y2=0
cc_641 N_SCD_M1004_g N_A_560_369#_c_1782_n 0.00495708f $X=3.61 $Y=2.165 $X2=0
+ $Y2=0
cc_642 N_SCD_M1011_g N_A_560_369#_c_1794_n 0.00446703f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_643 N_SCD_M1004_g N_A_560_369#_c_1806_n 0.00677278f $X=3.61 $Y=2.165 $X2=0
+ $Y2=0
cc_644 N_SCD_M1011_g N_A_560_369#_c_1771_n 0.00629065f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_645 N_SCD_M1004_g N_A_560_369#_c_1778_n 0.00857009f $X=3.61 $Y=2.165 $X2=0
+ $Y2=0
cc_646 SCD N_A_560_369#_c_1778_n 0.0313936f $X=3.855 $Y=1.105 $X2=0 $Y2=0
cc_647 N_SCD_c_822_n N_A_560_369#_c_1778_n 5.47858e-19 $X=3.67 $Y=1.355 $X2=0
+ $Y2=0
cc_648 N_SCD_M1004_g N_A_560_369#_c_1779_n 0.00253324f $X=3.61 $Y=2.165 $X2=0
+ $Y2=0
cc_649 SCD N_A_560_369#_c_1779_n 0.00365006f $X=3.855 $Y=1.105 $X2=0 $Y2=0
cc_650 N_SCD_M1011_g N_A_560_369#_c_1772_n 0.00825679f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_651 SCD N_A_560_369#_c_1772_n 0.0308767f $X=3.855 $Y=1.105 $X2=0 $Y2=0
cc_652 N_SCD_c_822_n N_A_560_369#_c_1772_n 5.22795e-19 $X=3.67 $Y=1.355 $X2=0
+ $Y2=0
cc_653 N_SCD_M1011_g N_A_560_369#_c_1773_n 0.00228451f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_654 SCD N_A_560_369#_c_1773_n 0.00395813f $X=3.855 $Y=1.105 $X2=0 $Y2=0
cc_655 N_SCD_M1011_g N_A_560_369#_c_1774_n 0.0022162f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_656 N_SCD_M1011_g N_A_560_369#_c_1775_n 0.00407065f $X=3.61 $Y=0.445 $X2=0
+ $Y2=0
cc_657 N_SCD_M1004_g N_A_560_369#_c_1775_n 0.00427612f $X=3.61 $Y=2.165 $X2=0
+ $Y2=0
cc_658 SCD N_A_560_369#_c_1775_n 0.0508929f $X=3.855 $Y=1.105 $X2=0 $Y2=0
cc_659 N_SCD_c_822_n N_A_560_369#_c_1775_n 0.00137588f $X=3.67 $Y=1.355 $X2=0
+ $Y2=0
cc_660 N_SCD_M1004_g N_A_560_369#_c_1781_n 0.00286352f $X=3.61 $Y=2.165 $X2=0
+ $Y2=0
cc_661 N_SCD_M1011_g N_VGND_c_1953_n 0.00562907f $X=3.61 $Y=0.445 $X2=0 $Y2=0
cc_662 N_SCD_M1011_g N_VGND_c_1965_n 0.00404961f $X=3.61 $Y=0.445 $X2=0 $Y2=0
cc_663 N_SCD_M1011_g N_VGND_c_1978_n 0.00665506f $X=3.61 $Y=0.445 $X2=0 $Y2=0
cc_664 N_A_193_47#_c_872_n N_A_1097_183#_M1001_d 0.00133652f $X=6.965 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_665 N_A_193_47#_c_875_n N_A_1097_183#_M1001_d 0.00107859f $X=6.58 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_666 N_A_193_47#_c_877_n N_A_1097_183#_M1001_d 5.46694e-19 $X=6.725 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_667 N_A_193_47#_c_875_n N_A_1097_183#_M1034_g 0.00208483f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_668 N_A_193_47#_c_880_n N_A_1097_183#_M1034_g 0.013781f $X=5.04 $Y=0.705
+ $X2=0 $Y2=0
cc_669 N_A_193_47#_c_875_n N_A_1097_183#_c_1085_n 0.0221014f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_670 N_A_193_47#_c_877_n N_A_1097_183#_c_1111_n 8.79173e-19 $X=6.725 $Y=0.85
+ $X2=0 $Y2=0
cc_671 N_A_193_47#_c_872_n N_A_1097_183#_c_1112_n 0.00716698f $X=6.965 $Y=0.87
+ $X2=0 $Y2=0
cc_672 N_A_193_47#_c_875_n N_A_1097_183#_c_1112_n 0.00405538f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_673 N_A_193_47#_c_877_n N_A_1097_183#_c_1112_n 0.0012409f $X=6.725 $Y=0.85
+ $X2=0 $Y2=0
cc_674 N_A_193_47#_c_875_n N_A_1097_183#_c_1086_n 0.00899288f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_675 N_A_193_47#_c_870_n N_A_1097_183#_c_1087_n 0.00114045f $X=7.06 $Y=1.575
+ $X2=0 $Y2=0
cc_676 N_A_193_47#_c_872_n N_A_1097_183#_c_1087_n 0.0187423f $X=6.965 $Y=0.87
+ $X2=0 $Y2=0
cc_677 N_A_193_47#_c_875_n N_A_1097_183#_c_1087_n 0.0176435f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_678 N_A_193_47#_c_877_n N_A_1097_183#_c_1087_n 0.00182243f $X=6.725 $Y=0.85
+ $X2=0 $Y2=0
cc_679 N_A_193_47#_c_881_n N_A_1097_183#_c_1087_n 5.82389e-19 $X=6.92 $Y=0.87
+ $X2=0 $Y2=0
cc_680 N_A_193_47#_c_870_n N_A_1097_183#_c_1088_n 0.00620052f $X=7.06 $Y=1.575
+ $X2=0 $Y2=0
cc_681 N_A_193_47#_c_875_n N_A_1097_183#_c_1089_n 0.00299829f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_682 N_A_193_47#_c_878_n N_A_1097_183#_c_1089_n 0.0179412f $X=5.04 $Y=0.87
+ $X2=0 $Y2=0
cc_683 N_A_193_47#_c_870_n N_A_938_413#_c_1178_n 6.31337e-19 $X=7.06 $Y=1.575
+ $X2=0 $Y2=0
cc_684 N_A_193_47#_c_868_n N_A_938_413#_c_1179_n 0.00957285f $X=6.825 $Y=0.705
+ $X2=0 $Y2=0
cc_685 N_A_193_47#_c_872_n N_A_938_413#_c_1179_n 0.00100831f $X=6.965 $Y=0.87
+ $X2=0 $Y2=0
cc_686 N_A_193_47#_c_870_n N_A_938_413#_c_1180_n 3.37852e-19 $X=7.06 $Y=1.575
+ $X2=0 $Y2=0
cc_687 N_A_193_47#_c_881_n N_A_938_413#_c_1180_n 0.00957285f $X=6.92 $Y=0.87
+ $X2=0 $Y2=0
cc_688 N_A_193_47#_M1015_g N_A_938_413#_c_1196_n 0.00169093f $X=4.615 $Y=2.275
+ $X2=0 $Y2=0
cc_689 N_A_193_47#_c_869_n N_A_938_413#_c_1196_n 0.00286257f $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_690 N_A_193_47#_c_885_n N_A_938_413#_c_1196_n 6.94615e-19 $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_691 N_A_193_47#_c_875_n N_A_938_413#_c_1222_n 0.00505066f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_692 N_A_193_47#_c_1007_p N_A_938_413#_c_1222_n 0.00102631f $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_693 N_A_193_47#_c_878_n N_A_938_413#_c_1222_n 0.00256542f $X=5.04 $Y=0.87
+ $X2=0 $Y2=0
cc_694 N_A_193_47#_c_879_n N_A_938_413#_c_1222_n 0.0237558f $X=5.04 $Y=0.87
+ $X2=0 $Y2=0
cc_695 N_A_193_47#_c_880_n N_A_938_413#_c_1222_n 0.00840911f $X=5.04 $Y=0.705
+ $X2=0 $Y2=0
cc_696 N_A_193_47#_c_869_n N_A_938_413#_c_1183_n 0.00981359f $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_697 N_A_193_47#_c_875_n N_A_938_413#_c_1183_n 0.0188221f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_698 N_A_193_47#_c_1007_p N_A_938_413#_c_1183_n 4.71298e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_699 N_A_193_47#_c_879_n N_A_938_413#_c_1183_n 0.023986f $X=5.04 $Y=0.87 $X2=0
+ $Y2=0
cc_700 N_A_193_47#_c_880_n N_A_938_413#_c_1183_n 0.00604394f $X=5.04 $Y=0.705
+ $X2=0 $Y2=0
cc_701 N_A_193_47#_c_869_n N_A_938_413#_c_1184_n 0.00649323f $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_702 N_A_193_47#_c_875_n N_A_938_413#_c_1184_n 0.00803733f $X=6.58 $Y=0.85
+ $X2=0 $Y2=0
cc_703 N_A_193_47#_M1008_g N_A_1525_315#_c_1307_n 0.018025f $X=7.115 $Y=2.275
+ $X2=0 $Y2=0
cc_704 N_A_193_47#_c_888_n N_A_1525_315#_c_1307_n 0.0119764f $X=7.2 $Y=1.74
+ $X2=0 $Y2=0
cc_705 N_A_193_47#_M1008_g N_A_1354_413#_c_1434_n 0.00974744f $X=7.115 $Y=2.275
+ $X2=0 $Y2=0
cc_706 N_A_193_47#_c_887_n N_A_1354_413#_c_1434_n 0.012999f $X=7.2 $Y=1.74 $X2=0
+ $Y2=0
cc_707 N_A_193_47#_c_888_n N_A_1354_413#_c_1434_n 0.00300896f $X=7.2 $Y=1.74
+ $X2=0 $Y2=0
cc_708 N_A_193_47#_c_872_n N_A_1354_413#_c_1437_n 0.0153172f $X=6.965 $Y=0.87
+ $X2=0 $Y2=0
cc_709 N_A_193_47#_c_881_n N_A_1354_413#_c_1437_n 8.54271e-19 $X=6.92 $Y=0.87
+ $X2=0 $Y2=0
cc_710 N_A_193_47#_M1008_g N_A_1354_413#_c_1431_n 0.0046302f $X=7.115 $Y=2.275
+ $X2=0 $Y2=0
cc_711 N_A_193_47#_c_870_n N_A_1354_413#_c_1431_n 0.00868218f $X=7.06 $Y=1.575
+ $X2=0 $Y2=0
cc_712 N_A_193_47#_c_887_n N_A_1354_413#_c_1431_n 0.024681f $X=7.2 $Y=1.74 $X2=0
+ $Y2=0
cc_713 N_A_193_47#_c_888_n N_A_1354_413#_c_1431_n 0.00187857f $X=7.2 $Y=1.74
+ $X2=0 $Y2=0
cc_714 N_A_193_47#_c_870_n N_A_1354_413#_c_1426_n 0.0272384f $X=7.06 $Y=1.575
+ $X2=0 $Y2=0
cc_715 N_A_193_47#_c_888_n N_A_1354_413#_c_1426_n 0.00102186f $X=7.2 $Y=1.74
+ $X2=0 $Y2=0
cc_716 N_A_193_47#_c_868_n N_A_1354_413#_c_1427_n 8.96907e-19 $X=6.825 $Y=0.705
+ $X2=0 $Y2=0
cc_717 N_A_193_47#_c_872_n N_A_1354_413#_c_1427_n 0.0255918f $X=6.965 $Y=0.87
+ $X2=0 $Y2=0
cc_718 N_A_193_47#_c_877_n N_A_1354_413#_c_1427_n 8.3858e-19 $X=6.725 $Y=0.85
+ $X2=0 $Y2=0
cc_719 N_A_193_47#_c_881_n N_A_1354_413#_c_1427_n 3.08898e-19 $X=6.92 $Y=0.87
+ $X2=0 $Y2=0
cc_720 N_A_193_47#_c_876_n N_VPWR_c_1579_n 0.0127357f $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_721 N_A_193_47#_c_876_n N_VPWR_c_1580_n 5.63902e-19 $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_722 N_A_193_47#_M1015_g N_VPWR_c_1581_n 0.00265717f $X=4.615 $Y=2.275 $X2=0
+ $Y2=0
cc_723 N_A_193_47#_M1015_g N_VPWR_c_1590_n 0.005785f $X=4.615 $Y=2.275 $X2=0
+ $Y2=0
cc_724 N_A_193_47#_c_876_n N_VPWR_c_1595_n 0.015988f $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_725 N_A_193_47#_M1008_g N_VPWR_c_1597_n 0.00383564f $X=7.115 $Y=2.275 $X2=0
+ $Y2=0
cc_726 N_A_193_47#_M1015_g N_VPWR_c_1578_n 0.00734982f $X=4.615 $Y=2.275 $X2=0
+ $Y2=0
cc_727 N_A_193_47#_M1008_g N_VPWR_c_1578_n 0.00579176f $X=7.115 $Y=2.275 $X2=0
+ $Y2=0
cc_728 N_A_193_47#_c_869_n N_VPWR_c_1578_n 0.00189161f $X=4.63 $Y=1.74 $X2=0
+ $Y2=0
cc_729 N_A_193_47#_c_885_n N_VPWR_c_1578_n 3.04586e-19 $X=4.63 $Y=1.74 $X2=0
+ $Y2=0
cc_730 N_A_193_47#_c_876_n N_VPWR_c_1578_n 0.00409094f $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_731 N_A_193_47#_c_873_n N_A_560_369#_c_1794_n 0.00537221f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_732 N_A_193_47#_c_873_n N_A_560_369#_c_1772_n 0.021391f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_733 N_A_193_47#_c_873_n N_A_560_369#_c_1773_n 0.00971398f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_734 N_A_193_47#_c_869_n N_A_560_369#_c_1775_n 0.058581f $X=4.63 $Y=1.74 $X2=0
+ $Y2=0
cc_735 N_A_193_47#_c_885_n N_A_560_369#_c_1775_n 0.0052844f $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_736 N_A_193_47#_c_873_n N_A_560_369#_c_1775_n 0.0123751f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_737 N_A_193_47#_c_1007_p N_A_560_369#_c_1775_n 2.40577e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_738 N_A_193_47#_c_879_n N_A_560_369#_c_1775_n 0.0125023f $X=5.04 $Y=0.87
+ $X2=0 $Y2=0
cc_739 N_A_193_47#_c_873_n N_A_560_369#_c_1776_n 0.00506513f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_740 N_A_193_47#_c_879_n N_A_560_369#_c_1776_n 6.01474e-19 $X=5.04 $Y=0.87
+ $X2=0 $Y2=0
cc_741 N_A_193_47#_c_873_n N_A_560_369#_c_1777_n 0.00562077f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_742 N_A_193_47#_c_1007_p N_A_560_369#_c_1777_n 2.71985e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_743 N_A_193_47#_c_879_n N_A_560_369#_c_1777_n 0.0122401f $X=5.04 $Y=0.87
+ $X2=0 $Y2=0
cc_744 N_A_193_47#_M1015_g N_A_560_369#_c_1781_n 0.00485506f $X=4.615 $Y=2.275
+ $X2=0 $Y2=0
cc_745 N_A_193_47#_c_869_n N_A_560_369#_c_1781_n 0.00558861f $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_746 N_A_193_47#_c_885_n N_A_560_369#_c_1781_n 0.00162985f $X=4.63 $Y=1.74
+ $X2=0 $Y2=0
cc_747 N_A_193_47#_c_873_n N_VGND_c_1952_n 0.00118059f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_748 N_A_193_47#_c_873_n N_VGND_c_1953_n 8.73533e-19 $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_749 N_A_193_47#_c_879_n N_VGND_c_1954_n 0.00254426f $X=5.04 $Y=0.87 $X2=0
+ $Y2=0
cc_750 N_A_193_47#_c_880_n N_VGND_c_1954_n 0.0037981f $X=5.04 $Y=0.705 $X2=0
+ $Y2=0
cc_751 N_A_193_47#_c_875_n N_VGND_c_1955_n 0.00197288f $X=6.58 $Y=0.85 $X2=0
+ $Y2=0
cc_752 N_A_193_47#_c_871_n N_VGND_c_1964_n 0.0100142f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_753 N_A_193_47#_c_868_n N_VGND_c_1966_n 0.00435108f $X=6.825 $Y=0.705 $X2=0
+ $Y2=0
cc_754 N_A_193_47#_c_872_n N_VGND_c_1966_n 0.00341023f $X=6.965 $Y=0.87 $X2=0
+ $Y2=0
cc_755 N_A_193_47#_c_881_n N_VGND_c_1966_n 8.04624e-19 $X=6.92 $Y=0.87 $X2=0
+ $Y2=0
cc_756 N_A_193_47#_M1027_d N_VGND_c_1978_n 0.00281453f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_757 N_A_193_47#_c_868_n N_VGND_c_1978_n 0.00619334f $X=6.825 $Y=0.705 $X2=0
+ $Y2=0
cc_758 N_A_193_47#_c_871_n N_VGND_c_1978_n 0.00380969f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_759 N_A_193_47#_c_872_n N_VGND_c_1978_n 0.00383201f $X=6.965 $Y=0.87 $X2=0
+ $Y2=0
cc_760 N_A_193_47#_c_873_n N_VGND_c_1978_n 0.156876f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_A_193_47#_c_874_n N_VGND_c_1978_n 0.0151167f $X=1.28 $Y=0.85 $X2=0
+ $Y2=0
cc_762 N_A_193_47#_c_875_n N_VGND_c_1978_n 0.0737651f $X=6.58 $Y=0.85 $X2=0
+ $Y2=0
cc_763 N_A_193_47#_c_1007_p N_VGND_c_1978_n 0.0146285f $X=4.975 $Y=0.85 $X2=0
+ $Y2=0
cc_764 N_A_193_47#_c_877_n N_VGND_c_1978_n 0.0146952f $X=6.725 $Y=0.85 $X2=0
+ $Y2=0
cc_765 N_A_193_47#_c_879_n N_VGND_c_1978_n 0.00247273f $X=5.04 $Y=0.87 $X2=0
+ $Y2=0
cc_766 N_A_193_47#_c_880_n N_VGND_c_1978_n 0.00563926f $X=5.04 $Y=0.705 $X2=0
+ $Y2=0
cc_767 N_A_193_47#_c_881_n N_VGND_c_1978_n 0.00134095f $X=6.92 $Y=0.87 $X2=0
+ $Y2=0
cc_768 N_A_1097_183#_c_1088_n N_A_938_413#_c_1178_n 0.00595764f $X=6.39 $Y=2.135
+ $X2=0 $Y2=0
cc_769 N_A_1097_183#_M1013_g N_A_938_413#_M1033_g 0.0139082f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_770 N_A_1097_183#_c_1099_n N_A_938_413#_M1033_g 0.00378805f $X=6.43 $Y=2.3
+ $X2=0 $Y2=0
cc_771 N_A_1097_183#_c_1088_n N_A_938_413#_M1033_g 0.0122998f $X=6.39 $Y=2.135
+ $X2=0 $Y2=0
cc_772 N_A_1097_183#_M1034_g N_A_938_413#_c_1179_n 0.0109128f $X=5.59 $Y=0.445
+ $X2=0 $Y2=0
cc_773 N_A_1097_183#_c_1085_n N_A_938_413#_c_1179_n 0.00351053f $X=6.265
+ $Y=0.915 $X2=0 $Y2=0
cc_774 N_A_1097_183#_c_1111_n N_A_938_413#_c_1179_n 0.00675936f $X=6.35 $Y=0.765
+ $X2=0 $Y2=0
cc_775 N_A_1097_183#_c_1131_p N_A_938_413#_c_1179_n 0.004701f $X=6.435 $Y=0.45
+ $X2=0 $Y2=0
cc_776 N_A_1097_183#_c_1087_n N_A_938_413#_c_1179_n 0.00333126f $X=6.35 $Y=0.915
+ $X2=0 $Y2=0
cc_777 N_A_1097_183#_c_1089_n N_A_938_413#_c_1179_n 0.00500517f $X=5.59 $Y=0.93
+ $X2=0 $Y2=0
cc_778 N_A_1097_183#_M1013_g N_A_938_413#_c_1180_n 0.00398999f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_779 N_A_1097_183#_c_1085_n N_A_938_413#_c_1180_n 0.00996228f $X=6.265
+ $Y=0.915 $X2=0 $Y2=0
cc_780 N_A_1097_183#_c_1086_n N_A_938_413#_c_1180_n 2.46578e-19 $X=5.805 $Y=0.93
+ $X2=0 $Y2=0
cc_781 N_A_1097_183#_c_1087_n N_A_938_413#_c_1180_n 0.00234347f $X=6.35 $Y=0.915
+ $X2=0 $Y2=0
cc_782 N_A_1097_183#_c_1088_n N_A_938_413#_c_1180_n 0.00394884f $X=6.39 $Y=2.135
+ $X2=0 $Y2=0
cc_783 N_A_1097_183#_c_1089_n N_A_938_413#_c_1180_n 0.00573363f $X=5.59 $Y=0.93
+ $X2=0 $Y2=0
cc_784 N_A_1097_183#_M1013_g N_A_938_413#_c_1181_n 0.0173592f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_785 N_A_1097_183#_c_1085_n N_A_938_413#_c_1181_n 0.00400764f $X=6.265
+ $Y=0.915 $X2=0 $Y2=0
cc_786 N_A_1097_183#_c_1089_n N_A_938_413#_c_1181_n 0.00238133f $X=5.59 $Y=0.93
+ $X2=0 $Y2=0
cc_787 N_A_1097_183#_c_1088_n N_A_938_413#_c_1182_n 0.00611615f $X=6.39 $Y=2.135
+ $X2=0 $Y2=0
cc_788 N_A_1097_183#_M1013_g N_A_938_413#_c_1196_n 0.0101048f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_789 N_A_1097_183#_M1034_g N_A_938_413#_c_1183_n 0.00441151f $X=5.59 $Y=0.445
+ $X2=0 $Y2=0
cc_790 N_A_1097_183#_c_1086_n N_A_938_413#_c_1183_n 0.0243525f $X=5.805 $Y=0.93
+ $X2=0 $Y2=0
cc_791 N_A_1097_183#_c_1089_n N_A_938_413#_c_1183_n 0.0095167f $X=5.59 $Y=0.93
+ $X2=0 $Y2=0
cc_792 N_A_1097_183#_M1013_g N_A_938_413#_c_1188_n 0.0153783f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_793 N_A_1097_183#_c_1088_n N_A_938_413#_c_1188_n 0.00754007f $X=6.39 $Y=2.135
+ $X2=0 $Y2=0
cc_794 N_A_1097_183#_M1013_g N_A_938_413#_c_1184_n 0.0138593f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_795 N_A_1097_183#_c_1085_n N_A_938_413#_c_1184_n 0.0186614f $X=6.265 $Y=0.915
+ $X2=0 $Y2=0
cc_796 N_A_1097_183#_c_1086_n N_A_938_413#_c_1184_n 0.0112018f $X=5.805 $Y=0.93
+ $X2=0 $Y2=0
cc_797 N_A_1097_183#_c_1088_n N_A_938_413#_c_1184_n 0.0245884f $X=6.39 $Y=2.135
+ $X2=0 $Y2=0
cc_798 N_A_1097_183#_c_1089_n N_A_938_413#_c_1184_n 0.00213749f $X=5.59 $Y=0.93
+ $X2=0 $Y2=0
cc_799 N_A_1097_183#_c_1099_n N_A_1354_413#_c_1434_n 0.0109209f $X=6.43 $Y=2.3
+ $X2=0 $Y2=0
cc_800 N_A_1097_183#_M1013_g N_VPWR_c_1582_n 0.0057281f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_801 N_A_1097_183#_c_1088_n N_VPWR_c_1582_n 0.0237f $X=6.39 $Y=2.135 $X2=0
+ $Y2=0
cc_802 N_A_1097_183#_M1013_g N_VPWR_c_1590_n 0.00378797f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_803 N_A_1097_183#_c_1099_n N_VPWR_c_1597_n 0.015079f $X=6.43 $Y=2.3 $X2=0
+ $Y2=0
cc_804 N_A_1097_183#_M1033_d N_VPWR_c_1578_n 0.00285796f $X=6.295 $Y=1.735 $X2=0
+ $Y2=0
cc_805 N_A_1097_183#_M1013_g N_VPWR_c_1578_n 0.00596544f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_806 N_A_1097_183#_c_1099_n N_VPWR_c_1578_n 0.00439826f $X=6.43 $Y=2.3 $X2=0
+ $Y2=0
cc_807 N_A_1097_183#_c_1085_n N_VGND_M1034_d 0.00306998f $X=6.265 $Y=0.915 $X2=0
+ $Y2=0
cc_808 N_A_1097_183#_M1034_g N_VGND_c_1954_n 0.00585385f $X=5.59 $Y=0.445 $X2=0
+ $Y2=0
cc_809 N_A_1097_183#_M1034_g N_VGND_c_1955_n 0.00603751f $X=5.59 $Y=0.445 $X2=0
+ $Y2=0
cc_810 N_A_1097_183#_c_1111_n N_VGND_c_1955_n 0.00354103f $X=6.35 $Y=0.765 $X2=0
+ $Y2=0
cc_811 N_A_1097_183#_c_1131_p N_VGND_c_1955_n 0.013122f $X=6.435 $Y=0.45 $X2=0
+ $Y2=0
cc_812 N_A_1097_183#_c_1086_n N_VGND_c_1955_n 0.0258565f $X=5.805 $Y=0.93 $X2=0
+ $Y2=0
cc_813 N_A_1097_183#_c_1089_n N_VGND_c_1955_n 0.00122075f $X=5.59 $Y=0.93 $X2=0
+ $Y2=0
cc_814 N_A_1097_183#_c_1131_p N_VGND_c_1966_n 0.00594819f $X=6.435 $Y=0.45 $X2=0
+ $Y2=0
cc_815 N_A_1097_183#_c_1112_n N_VGND_c_1966_n 0.0100275f $X=6.56 $Y=0.45 $X2=0
+ $Y2=0
cc_816 N_A_1097_183#_M1001_d N_VGND_c_1978_n 0.00246943f $X=6.395 $Y=0.235 $X2=0
+ $Y2=0
cc_817 N_A_1097_183#_M1034_g N_VGND_c_1978_n 0.0070154f $X=5.59 $Y=0.445 $X2=0
+ $Y2=0
cc_818 N_A_1097_183#_c_1085_n N_VGND_c_1978_n 0.0042145f $X=6.265 $Y=0.915 $X2=0
+ $Y2=0
cc_819 N_A_1097_183#_c_1131_p N_VGND_c_1978_n 0.00261981f $X=6.435 $Y=0.45 $X2=0
+ $Y2=0
cc_820 N_A_1097_183#_c_1112_n N_VGND_c_1978_n 0.00442918f $X=6.56 $Y=0.45 $X2=0
+ $Y2=0
cc_821 N_A_1097_183#_c_1086_n N_VGND_c_1978_n 0.00269026f $X=5.805 $Y=0.93 $X2=0
+ $Y2=0
cc_822 N_A_938_413#_c_1196_n N_VPWR_M1013_d 0.00236303f $X=5.585 $Y=2.275 $X2=0
+ $Y2=0
cc_823 N_A_938_413#_c_1188_n N_VPWR_M1013_d 0.00412006f $X=5.67 $Y=2.19 $X2=0
+ $Y2=0
cc_824 N_A_938_413#_M1033_g N_VPWR_c_1582_n 0.00314007f $X=6.22 $Y=2.11 $X2=0
+ $Y2=0
cc_825 N_A_938_413#_c_1181_n N_VPWR_c_1582_n 9.53331e-19 $X=6.145 $Y=1.41 $X2=0
+ $Y2=0
cc_826 N_A_938_413#_c_1196_n N_VPWR_c_1582_n 0.0138309f $X=5.585 $Y=2.275 $X2=0
+ $Y2=0
cc_827 N_A_938_413#_c_1188_n N_VPWR_c_1582_n 0.0252361f $X=5.67 $Y=2.19 $X2=0
+ $Y2=0
cc_828 N_A_938_413#_c_1184_n N_VPWR_c_1582_n 0.00741701f $X=5.67 $Y=1.41 $X2=0
+ $Y2=0
cc_829 N_A_938_413#_c_1196_n N_VPWR_c_1590_n 0.0359536f $X=5.585 $Y=2.275 $X2=0
+ $Y2=0
cc_830 N_A_938_413#_M1033_g N_VPWR_c_1597_n 0.00541359f $X=6.22 $Y=2.11 $X2=0
+ $Y2=0
cc_831 N_A_938_413#_M1015_d N_VPWR_c_1578_n 0.00217001f $X=4.69 $Y=2.065 $X2=0
+ $Y2=0
cc_832 N_A_938_413#_M1033_g N_VPWR_c_1578_n 0.00665748f $X=6.22 $Y=2.11 $X2=0
+ $Y2=0
cc_833 N_A_938_413#_c_1196_n N_VPWR_c_1578_n 0.0161661f $X=5.585 $Y=2.275 $X2=0
+ $Y2=0
cc_834 N_A_938_413#_c_1196_n A_1031_413# 0.0045944f $X=5.585 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_835 N_A_938_413#_c_1222_n N_VGND_c_1954_n 0.0255873f $X=5.295 $Y=0.45 $X2=0
+ $Y2=0
cc_836 N_A_938_413#_c_1179_n N_VGND_c_1955_n 0.00816054f $X=6.32 $Y=0.95 $X2=0
+ $Y2=0
cc_837 N_A_938_413#_c_1179_n N_VGND_c_1966_n 0.00407056f $X=6.32 $Y=0.95 $X2=0
+ $Y2=0
cc_838 N_A_938_413#_M1024_d N_VGND_c_1978_n 0.00228142f $X=4.695 $Y=0.235 $X2=0
+ $Y2=0
cc_839 N_A_938_413#_c_1179_n N_VGND_c_1978_n 0.00620172f $X=6.32 $Y=0.95 $X2=0
+ $Y2=0
cc_840 N_A_938_413#_c_1222_n N_VGND_c_1978_n 0.0113221f $X=5.295 $Y=0.45 $X2=0
+ $Y2=0
cc_841 N_A_938_413#_c_1222_n A_1035_47# 0.00455507f $X=5.295 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_842 N_A_938_413#_c_1183_n A_1035_47# 0.00200718f $X=5.38 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_843 N_A_1525_315#_c_1287_n N_A_1354_413#_c_1422_n 0.0203579f $X=9.21 $Y=0.995
+ $X2=0 $Y2=0
cc_844 N_A_1525_315#_c_1293_n N_A_1354_413#_c_1422_n 0.00487327f $X=8.632
+ $Y=0.995 $X2=0 $Y2=0
cc_845 N_A_1525_315#_c_1295_n N_A_1354_413#_c_1422_n 0.00674772f $X=8.56
+ $Y=0.385 $X2=0 $Y2=0
cc_846 N_A_1525_315#_M1005_g N_A_1354_413#_M1035_g 0.0206926f $X=9.21 $Y=1.985
+ $X2=0 $Y2=0
cc_847 N_A_1525_315#_c_1308_n N_A_1354_413#_M1035_g 0.00599733f $X=8.56 $Y=2.34
+ $X2=0 $Y2=0
cc_848 N_A_1525_315#_c_1309_n N_A_1354_413#_M1035_g 0.00717661f $X=8.632
+ $Y=1.575 $X2=0 $Y2=0
cc_849 N_A_1525_315#_c_1311_n N_A_1354_413#_M1035_g 0.00383694f $X=8.56 $Y=1.66
+ $X2=0 $Y2=0
cc_850 N_A_1525_315#_M1003_g N_A_1354_413#_c_1423_n 0.0164567f $X=7.815 $Y=0.445
+ $X2=0 $Y2=0
cc_851 N_A_1525_315#_c_1306_n N_A_1354_413#_c_1423_n 0.00567751f $X=8.395
+ $Y=1.74 $X2=0 $Y2=0
cc_852 N_A_1525_315#_c_1295_n N_A_1354_413#_c_1423_n 0.00747686f $X=8.56
+ $Y=0.385 $X2=0 $Y2=0
cc_853 N_A_1525_315#_c_1311_n N_A_1354_413#_c_1423_n 0.00591375f $X=8.56 $Y=1.66
+ $X2=0 $Y2=0
cc_854 N_A_1525_315#_c_1326_p N_A_1354_413#_c_1423_n 0.0168258f $X=8.632 $Y=1.16
+ $X2=0 $Y2=0
cc_855 N_A_1525_315#_c_1290_n N_A_1354_413#_c_1424_n 0.0216171f $X=9.705 $Y=1.16
+ $X2=0 $Y2=0
cc_856 N_A_1525_315#_c_1294_n N_A_1354_413#_c_1424_n 0.0180498f $X=9.19 $Y=1.16
+ $X2=0 $Y2=0
cc_857 N_A_1525_315#_c_1326_p N_A_1354_413#_c_1424_n 9.32228e-19 $X=8.632
+ $Y=1.16 $X2=0 $Y2=0
cc_858 N_A_1525_315#_M1031_g N_A_1354_413#_c_1434_n 0.00194535f $X=7.7 $Y=2.275
+ $X2=0 $Y2=0
cc_859 N_A_1525_315#_M1003_g N_A_1354_413#_c_1437_n 0.00114979f $X=7.815
+ $Y=0.445 $X2=0 $Y2=0
cc_860 N_A_1525_315#_c_1306_n N_A_1354_413#_c_1431_n 0.0262086f $X=8.395 $Y=1.74
+ $X2=0 $Y2=0
cc_861 N_A_1525_315#_c_1307_n N_A_1354_413#_c_1431_n 0.00865902f $X=7.88 $Y=1.74
+ $X2=0 $Y2=0
cc_862 N_A_1525_315#_M1003_g N_A_1354_413#_c_1425_n 0.0181285f $X=7.815 $Y=0.445
+ $X2=0 $Y2=0
cc_863 N_A_1525_315#_c_1306_n N_A_1354_413#_c_1425_n 0.0343168f $X=8.395 $Y=1.74
+ $X2=0 $Y2=0
cc_864 N_A_1525_315#_c_1307_n N_A_1354_413#_c_1425_n 0.00739167f $X=7.88 $Y=1.74
+ $X2=0 $Y2=0
cc_865 N_A_1525_315#_c_1295_n N_A_1354_413#_c_1425_n 7.42989e-19 $X=8.56
+ $Y=0.385 $X2=0 $Y2=0
cc_866 N_A_1525_315#_c_1326_p N_A_1354_413#_c_1425_n 0.0277655f $X=8.632 $Y=1.16
+ $X2=0 $Y2=0
cc_867 N_A_1525_315#_M1003_g N_A_1354_413#_c_1426_n 0.00880678f $X=7.815
+ $Y=0.445 $X2=0 $Y2=0
cc_868 N_A_1525_315#_M1003_g N_A_1354_413#_c_1427_n 0.00779225f $X=7.815
+ $Y=0.445 $X2=0 $Y2=0
cc_869 N_A_1525_315#_c_1291_n N_A_2049_47#_c_1509_n 0.00317818f $X=10.525
+ $Y=1.325 $X2=0 $Y2=0
cc_870 N_A_1525_315#_c_1292_n N_A_2049_47#_c_1509_n 0.0140671f $X=10.58 $Y=0.73
+ $X2=0 $Y2=0
cc_871 N_A_1525_315#_c_1304_n N_A_2049_47#_M1002_g 0.00474627f $X=10.552
+ $Y=1.515 $X2=0 $Y2=0
cc_872 N_A_1525_315#_c_1305_n N_A_2049_47#_M1002_g 0.0181632f $X=10.552 $Y=1.665
+ $X2=0 $Y2=0
cc_873 N_A_1525_315#_c_1288_n N_A_2049_47#_c_1511_n 0.00507334f $X=9.63 $Y=0.995
+ $X2=0 $Y2=0
cc_874 N_A_1525_315#_c_1291_n N_A_2049_47#_c_1511_n 0.00936266f $X=10.525
+ $Y=1.325 $X2=0 $Y2=0
cc_875 N_A_1525_315#_c_1292_n N_A_2049_47#_c_1511_n 0.00172958f $X=10.58 $Y=0.73
+ $X2=0 $Y2=0
cc_876 N_A_1525_315#_M1019_g N_A_2049_47#_c_1516_n 0.00606518f $X=9.63 $Y=1.985
+ $X2=0 $Y2=0
cc_877 N_A_1525_315#_M1038_g N_A_2049_47#_c_1516_n 0.0120617f $X=10.58 $Y=2.165
+ $X2=0 $Y2=0
cc_878 N_A_1525_315#_c_1304_n N_A_2049_47#_c_1516_n 0.00799512f $X=10.552
+ $Y=1.515 $X2=0 $Y2=0
cc_879 N_A_1525_315#_c_1305_n N_A_2049_47#_c_1516_n 0.00666896f $X=10.552
+ $Y=1.665 $X2=0 $Y2=0
cc_880 N_A_1525_315#_c_1291_n N_A_2049_47#_c_1512_n 0.0133342f $X=10.525
+ $Y=1.325 $X2=0 $Y2=0
cc_881 N_A_1525_315#_c_1305_n N_A_2049_47#_c_1512_n 0.00159098f $X=10.552
+ $Y=1.665 $X2=0 $Y2=0
cc_882 N_A_1525_315#_c_1289_n N_A_2049_47#_c_1532_n 0.0245362f $X=10.45 $Y=1.16
+ $X2=0 $Y2=0
cc_883 N_A_1525_315#_c_1291_n N_A_2049_47#_c_1532_n 0.00652717f $X=10.525
+ $Y=1.325 $X2=0 $Y2=0
cc_884 N_A_1525_315#_c_1291_n N_A_2049_47#_c_1513_n 0.0178735f $X=10.525
+ $Y=1.325 $X2=0 $Y2=0
cc_885 N_A_1525_315#_M1031_g N_VPWR_c_1583_n 0.0115962f $X=7.7 $Y=2.275 $X2=0
+ $Y2=0
cc_886 N_A_1525_315#_c_1306_n N_VPWR_c_1583_n 0.0182102f $X=8.395 $Y=1.74 $X2=0
+ $Y2=0
cc_887 N_A_1525_315#_c_1307_n N_VPWR_c_1583_n 0.0049226f $X=7.88 $Y=1.74 $X2=0
+ $Y2=0
cc_888 N_A_1525_315#_c_1308_n N_VPWR_c_1583_n 0.0179808f $X=8.56 $Y=2.34 $X2=0
+ $Y2=0
cc_889 N_A_1525_315#_c_1308_n N_VPWR_c_1584_n 0.0197786f $X=8.56 $Y=2.34 $X2=0
+ $Y2=0
cc_890 N_A_1525_315#_M1005_g N_VPWR_c_1585_n 0.00655352f $X=9.21 $Y=1.985 $X2=0
+ $Y2=0
cc_891 N_A_1525_315#_c_1290_n N_VPWR_c_1585_n 4.10671e-19 $X=9.705 $Y=1.16 $X2=0
+ $Y2=0
cc_892 N_A_1525_315#_c_1294_n N_VPWR_c_1585_n 0.0100037f $X=9.19 $Y=1.16 $X2=0
+ $Y2=0
cc_893 N_A_1525_315#_M1019_g N_VPWR_c_1586_n 0.0109361f $X=9.63 $Y=1.985 $X2=0
+ $Y2=0
cc_894 N_A_1525_315#_c_1289_n N_VPWR_c_1586_n 0.00543326f $X=10.45 $Y=1.16 $X2=0
+ $Y2=0
cc_895 N_A_1525_315#_M1038_g N_VPWR_c_1586_n 0.00401192f $X=10.58 $Y=2.165 $X2=0
+ $Y2=0
cc_896 N_A_1525_315#_c_1305_n N_VPWR_c_1586_n 2.01664e-19 $X=10.552 $Y=1.665
+ $X2=0 $Y2=0
cc_897 N_A_1525_315#_c_1305_n N_VPWR_c_1587_n 0.0119616f $X=10.552 $Y=1.665
+ $X2=0 $Y2=0
cc_898 N_A_1525_315#_M1005_g N_VPWR_c_1592_n 0.00542757f $X=9.21 $Y=1.985 $X2=0
+ $Y2=0
cc_899 N_A_1525_315#_M1019_g N_VPWR_c_1592_n 0.00542757f $X=9.63 $Y=1.985 $X2=0
+ $Y2=0
cc_900 N_A_1525_315#_M1031_g N_VPWR_c_1597_n 0.00585385f $X=7.7 $Y=2.275 $X2=0
+ $Y2=0
cc_901 N_A_1525_315#_M1038_g N_VPWR_c_1598_n 0.00542953f $X=10.58 $Y=2.165 $X2=0
+ $Y2=0
cc_902 N_A_1525_315#_M1035_s N_VPWR_c_1578_n 0.00209642f $X=8.435 $Y=1.485 $X2=0
+ $Y2=0
cc_903 N_A_1525_315#_M1031_g N_VPWR_c_1578_n 0.0124099f $X=7.7 $Y=2.275 $X2=0
+ $Y2=0
cc_904 N_A_1525_315#_M1005_g N_VPWR_c_1578_n 0.00968319f $X=9.21 $Y=1.985 $X2=0
+ $Y2=0
cc_905 N_A_1525_315#_M1019_g N_VPWR_c_1578_n 0.0108549f $X=9.63 $Y=1.985 $X2=0
+ $Y2=0
cc_906 N_A_1525_315#_M1038_g N_VPWR_c_1578_n 0.0111168f $X=10.58 $Y=2.165 $X2=0
+ $Y2=0
cc_907 N_A_1525_315#_c_1306_n N_VPWR_c_1578_n 0.0121091f $X=8.395 $Y=1.74 $X2=0
+ $Y2=0
cc_908 N_A_1525_315#_c_1307_n N_VPWR_c_1578_n 7.75814e-19 $X=7.88 $Y=1.74 $X2=0
+ $Y2=0
cc_909 N_A_1525_315#_c_1308_n N_VPWR_c_1578_n 0.0123666f $X=8.56 $Y=2.34 $X2=0
+ $Y2=0
cc_910 N_A_1525_315#_M1005_g N_Q_c_1895_n 0.0105686f $X=9.21 $Y=1.985 $X2=0
+ $Y2=0
cc_911 N_A_1525_315#_M1019_g N_Q_c_1895_n 0.0112795f $X=9.63 $Y=1.985 $X2=0
+ $Y2=0
cc_912 N_A_1525_315#_c_1309_n N_Q_c_1895_n 0.00124581f $X=8.632 $Y=1.575 $X2=0
+ $Y2=0
cc_913 N_A_1525_315#_c_1311_n N_Q_c_1895_n 0.00156787f $X=8.56 $Y=1.66 $X2=0
+ $Y2=0
cc_914 N_A_1525_315#_c_1287_n N_Q_c_1892_n 0.00216579f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_915 N_A_1525_315#_M1005_g N_Q_c_1892_n 0.00477172f $X=9.21 $Y=1.985 $X2=0
+ $Y2=0
cc_916 N_A_1525_315#_c_1288_n N_Q_c_1892_n 0.00302688f $X=9.63 $Y=0.995 $X2=0
+ $Y2=0
cc_917 N_A_1525_315#_M1019_g N_Q_c_1892_n 0.00724125f $X=9.63 $Y=1.985 $X2=0
+ $Y2=0
cc_918 N_A_1525_315#_c_1290_n N_Q_c_1892_n 0.0215544f $X=9.705 $Y=1.16 $X2=0
+ $Y2=0
cc_919 N_A_1525_315#_c_1309_n N_Q_c_1892_n 0.00100004f $X=8.632 $Y=1.575 $X2=0
+ $Y2=0
cc_920 N_A_1525_315#_c_1294_n N_Q_c_1892_n 0.026582f $X=9.19 $Y=1.16 $X2=0 $Y2=0
cc_921 N_A_1525_315#_c_1287_n N_Q_c_1893_n 0.0024123f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_922 N_A_1525_315#_c_1288_n N_Q_c_1893_n 0.0031371f $X=9.63 $Y=0.995 $X2=0
+ $Y2=0
cc_923 N_A_1525_315#_c_1290_n N_Q_c_1893_n 0.00212054f $X=9.705 $Y=1.16 $X2=0
+ $Y2=0
cc_924 N_A_1525_315#_c_1294_n N_Q_c_1893_n 0.00157529f $X=9.19 $Y=1.16 $X2=0
+ $Y2=0
cc_925 N_A_1525_315#_c_1295_n N_Q_c_1893_n 0.00105214f $X=8.56 $Y=0.385 $X2=0
+ $Y2=0
cc_926 N_A_1525_315#_c_1287_n N_Q_c_1911_n 0.00652062f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_927 N_A_1525_315#_c_1288_n N_Q_c_1911_n 0.00717234f $X=9.63 $Y=0.995 $X2=0
+ $Y2=0
cc_928 N_A_1525_315#_c_1295_n N_Q_c_1911_n 0.00281621f $X=8.56 $Y=0.385 $X2=0
+ $Y2=0
cc_929 N_A_1525_315#_M1003_g N_VGND_c_1956_n 0.0215676f $X=7.815 $Y=0.445 $X2=0
+ $Y2=0
cc_930 N_A_1525_315#_c_1295_n N_VGND_c_1956_n 0.0198494f $X=8.56 $Y=0.385 $X2=0
+ $Y2=0
cc_931 N_A_1525_315#_c_1295_n N_VGND_c_1957_n 0.0181097f $X=8.56 $Y=0.385 $X2=0
+ $Y2=0
cc_932 N_A_1525_315#_c_1287_n N_VGND_c_1958_n 0.001944f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_933 N_A_1525_315#_c_1290_n N_VGND_c_1958_n 6.02862e-19 $X=9.705 $Y=1.16 $X2=0
+ $Y2=0
cc_934 N_A_1525_315#_c_1294_n N_VGND_c_1958_n 0.0103606f $X=9.19 $Y=1.16 $X2=0
+ $Y2=0
cc_935 N_A_1525_315#_c_1288_n N_VGND_c_1959_n 0.00501847f $X=9.63 $Y=0.995 $X2=0
+ $Y2=0
cc_936 N_A_1525_315#_c_1289_n N_VGND_c_1959_n 0.0072715f $X=10.45 $Y=1.16 $X2=0
+ $Y2=0
cc_937 N_A_1525_315#_c_1292_n N_VGND_c_1959_n 0.00478714f $X=10.58 $Y=0.73 $X2=0
+ $Y2=0
cc_938 N_A_1525_315#_c_1292_n N_VGND_c_1960_n 0.00667732f $X=10.58 $Y=0.73 $X2=0
+ $Y2=0
cc_939 N_A_1525_315#_c_1287_n N_VGND_c_1967_n 0.00541359f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_940 N_A_1525_315#_c_1288_n N_VGND_c_1967_n 0.00541359f $X=9.63 $Y=0.995 $X2=0
+ $Y2=0
cc_941 N_A_1525_315#_c_1291_n N_VGND_c_1968_n 0.00105583f $X=10.525 $Y=1.325
+ $X2=0 $Y2=0
cc_942 N_A_1525_315#_c_1292_n N_VGND_c_1968_n 0.00585385f $X=10.58 $Y=0.73 $X2=0
+ $Y2=0
cc_943 N_A_1525_315#_M1032_s N_VGND_c_1978_n 0.00212021f $X=8.435 $Y=0.235 $X2=0
+ $Y2=0
cc_944 N_A_1525_315#_M1003_g N_VGND_c_1978_n 9.61436e-19 $X=7.815 $Y=0.445 $X2=0
+ $Y2=0
cc_945 N_A_1525_315#_c_1287_n N_VGND_c_1978_n 0.00965588f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_946 N_A_1525_315#_c_1288_n N_VGND_c_1978_n 0.0099975f $X=9.63 $Y=0.995 $X2=0
+ $Y2=0
cc_947 N_A_1525_315#_c_1291_n N_VGND_c_1978_n 0.00138273f $X=10.525 $Y=1.325
+ $X2=0 $Y2=0
cc_948 N_A_1525_315#_c_1292_n N_VGND_c_1978_n 0.0122138f $X=10.58 $Y=0.73 $X2=0
+ $Y2=0
cc_949 N_A_1525_315#_c_1295_n N_VGND_c_1978_n 0.0134083f $X=8.56 $Y=0.385 $X2=0
+ $Y2=0
cc_950 N_A_1354_413#_M1035_g N_VPWR_c_1583_n 0.00211737f $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_951 N_A_1354_413#_M1035_g N_VPWR_c_1584_n 0.00541763f $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_952 N_A_1354_413#_M1035_g N_VPWR_c_1585_n 0.00321253f $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_953 N_A_1354_413#_c_1434_n N_VPWR_c_1597_n 0.0273845f $X=7.455 $Y=2.25 $X2=0
+ $Y2=0
cc_954 N_A_1354_413#_M1018_d N_VPWR_c_1578_n 0.00217593f $X=6.77 $Y=2.065 $X2=0
+ $Y2=0
cc_955 N_A_1354_413#_M1035_g N_VPWR_c_1578_n 0.0109823f $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_956 N_A_1354_413#_c_1434_n N_VPWR_c_1578_n 0.0274677f $X=7.455 $Y=2.25 $X2=0
+ $Y2=0
cc_957 N_A_1354_413#_c_1434_n A_1438_413# 0.0105858f $X=7.455 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_958 N_A_1354_413#_c_1431_n A_1438_413# 0.00184879f $X=7.54 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_959 N_A_1354_413#_M1035_g N_Q_c_1895_n 4.53355e-19 $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_960 N_A_1354_413#_c_1422_n N_Q_c_1911_n 3.39217e-19 $X=8.77 $Y=0.995 $X2=0
+ $Y2=0
cc_961 N_A_1354_413#_c_1422_n N_VGND_c_1956_n 0.00262644f $X=8.77 $Y=0.995 $X2=0
+ $Y2=0
cc_962 N_A_1354_413#_c_1437_n N_VGND_c_1956_n 0.0104892f $X=7.325 $Y=0.45 $X2=0
+ $Y2=0
cc_963 N_A_1354_413#_c_1425_n N_VGND_c_1956_n 0.0154767f $X=8.285 $Y=1.16 $X2=0
+ $Y2=0
cc_964 N_A_1354_413#_c_1427_n N_VGND_c_1956_n 0.00447237f $X=7.475 $Y=0.995
+ $X2=0 $Y2=0
cc_965 N_A_1354_413#_c_1422_n N_VGND_c_1957_n 0.00543148f $X=8.77 $Y=0.995 $X2=0
+ $Y2=0
cc_966 N_A_1354_413#_c_1422_n N_VGND_c_1958_n 0.00318378f $X=8.77 $Y=0.995 $X2=0
+ $Y2=0
cc_967 N_A_1354_413#_c_1437_n N_VGND_c_1966_n 0.0184388f $X=7.325 $Y=0.45 $X2=0
+ $Y2=0
cc_968 N_A_1354_413#_M1022_d N_VGND_c_1978_n 0.00333348f $X=6.9 $Y=0.235 $X2=0
+ $Y2=0
cc_969 N_A_1354_413#_c_1422_n N_VGND_c_1978_n 0.0109852f $X=8.77 $Y=0.995 $X2=0
+ $Y2=0
cc_970 N_A_1354_413#_c_1437_n N_VGND_c_1978_n 0.0182474f $X=7.325 $Y=0.45 $X2=0
+ $Y2=0
cc_971 N_A_1354_413#_c_1437_n A_1483_47# 0.00201232f $X=7.325 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_972 N_A_1354_413#_c_1427_n A_1483_47# 0.00127737f $X=7.475 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_973 N_A_2049_47#_c_1516_n N_VPWR_c_1586_n 0.0453751f $X=10.37 $Y=2 $X2=0
+ $Y2=0
cc_974 N_A_2049_47#_M1002_g N_VPWR_c_1587_n 0.0158665f $X=11.065 $Y=1.985 $X2=0
+ $Y2=0
cc_975 N_A_2049_47#_M1014_g N_VPWR_c_1587_n 0.00118467f $X=11.485 $Y=1.985 $X2=0
+ $Y2=0
cc_976 N_A_2049_47#_c_1516_n N_VPWR_c_1587_n 0.0691115f $X=10.37 $Y=2 $X2=0
+ $Y2=0
cc_977 N_A_2049_47#_c_1512_n N_VPWR_c_1587_n 0.0228967f $X=10.98 $Y=1.16 $X2=0
+ $Y2=0
cc_978 N_A_2049_47#_c_1513_n N_VPWR_c_1587_n 0.00320419f $X=11.485 $Y=1.16 $X2=0
+ $Y2=0
cc_979 N_A_2049_47#_M1014_g N_VPWR_c_1589_n 0.00505661f $X=11.485 $Y=1.985 $X2=0
+ $Y2=0
cc_980 N_A_2049_47#_c_1516_n N_VPWR_c_1598_n 0.016757f $X=10.37 $Y=2 $X2=0 $Y2=0
cc_981 N_A_2049_47#_M1002_g N_VPWR_c_1599_n 0.0046653f $X=11.065 $Y=1.985 $X2=0
+ $Y2=0
cc_982 N_A_2049_47#_M1014_g N_VPWR_c_1599_n 0.00546688f $X=11.485 $Y=1.985 $X2=0
+ $Y2=0
cc_983 N_A_2049_47#_M1038_s N_VPWR_c_1578_n 0.00211564f $X=10.245 $Y=1.845 $X2=0
+ $Y2=0
cc_984 N_A_2049_47#_M1002_g N_VPWR_c_1578_n 0.00796766f $X=11.065 $Y=1.985 $X2=0
+ $Y2=0
cc_985 N_A_2049_47#_M1014_g N_VPWR_c_1578_n 0.0105222f $X=11.485 $Y=1.985 $X2=0
+ $Y2=0
cc_986 N_A_2049_47#_c_1516_n N_VPWR_c_1578_n 0.0121755f $X=10.37 $Y=2 $X2=0
+ $Y2=0
cc_987 N_A_2049_47#_c_1516_n N_Q_c_1895_n 0.00251221f $X=10.37 $Y=2 $X2=0 $Y2=0
cc_988 N_A_2049_47#_c_1511_n N_Q_c_1892_n 0.00299495f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_989 N_A_2049_47#_c_1516_n N_Q_c_1892_n 0.00611401f $X=10.37 $Y=2 $X2=0 $Y2=0
cc_990 N_A_2049_47#_c_1532_n N_Q_c_1892_n 0.00896744f $X=10.37 $Y=1.16 $X2=0
+ $Y2=0
cc_991 N_A_2049_47#_c_1511_n N_Q_c_1893_n 0.00297195f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_992 N_A_2049_47#_c_1511_n N_Q_c_1911_n 0.00288832f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_993 N_A_2049_47#_c_1510_n N_Q_N_c_1933_n 0.00620145f $X=11.485 $Y=0.995 $X2=0
+ $Y2=0
cc_994 N_A_2049_47#_c_1510_n N_Q_N_c_1934_n 0.00137437f $X=11.485 $Y=0.995 $X2=0
+ $Y2=0
cc_995 N_A_2049_47#_c_1509_n Q_N 0.0043963f $X=11.065 $Y=0.995 $X2=0 $Y2=0
cc_996 N_A_2049_47#_M1002_g Q_N 0.00389879f $X=11.065 $Y=1.985 $X2=0 $Y2=0
cc_997 N_A_2049_47#_c_1510_n Q_N 0.00469373f $X=11.485 $Y=0.995 $X2=0 $Y2=0
cc_998 N_A_2049_47#_M1014_g Q_N 0.0159787f $X=11.485 $Y=1.985 $X2=0 $Y2=0
cc_999 N_A_2049_47#_c_1516_n Q_N 0.00120363f $X=10.37 $Y=2 $X2=0 $Y2=0
cc_1000 N_A_2049_47#_c_1512_n Q_N 0.0253118f $X=10.98 $Y=1.16 $X2=0 $Y2=0
cc_1001 N_A_2049_47#_c_1513_n Q_N 0.0276587f $X=11.485 $Y=1.16 $X2=0 $Y2=0
cc_1002 N_A_2049_47#_c_1511_n N_VGND_c_1959_n 0.0228544f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_1003 N_A_2049_47#_c_1509_n N_VGND_c_1960_n 0.0105018f $X=11.065 $Y=0.995
+ $X2=0 $Y2=0
cc_1004 N_A_2049_47#_c_1510_n N_VGND_c_1960_n 7.8737e-19 $X=11.485 $Y=0.995
+ $X2=0 $Y2=0
cc_1005 N_A_2049_47#_c_1511_n N_VGND_c_1960_n 0.00937628f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_1006 N_A_2049_47#_c_1512_n N_VGND_c_1960_n 0.0230938f $X=10.98 $Y=1.16 $X2=0
+ $Y2=0
cc_1007 N_A_2049_47#_c_1513_n N_VGND_c_1960_n 0.00315906f $X=11.485 $Y=1.16
+ $X2=0 $Y2=0
cc_1008 N_A_2049_47#_c_1510_n N_VGND_c_1962_n 0.00461523f $X=11.485 $Y=0.995
+ $X2=0 $Y2=0
cc_1009 N_A_2049_47#_c_1511_n N_VGND_c_1968_n 0.0109259f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_1010 N_A_2049_47#_c_1509_n N_VGND_c_1969_n 0.0046653f $X=11.065 $Y=0.995
+ $X2=0 $Y2=0
cc_1011 N_A_2049_47#_c_1510_n N_VGND_c_1969_n 0.00541763f $X=11.485 $Y=0.995
+ $X2=0 $Y2=0
cc_1012 N_A_2049_47#_M1025_s N_VGND_c_1978_n 0.00272276f $X=10.245 $Y=0.235
+ $X2=0 $Y2=0
cc_1013 N_A_2049_47#_c_1509_n N_VGND_c_1978_n 0.00796766f $X=11.065 $Y=0.995
+ $X2=0 $Y2=0
cc_1014 N_A_2049_47#_c_1510_n N_VGND_c_1978_n 0.0104998f $X=11.485 $Y=0.995
+ $X2=0 $Y2=0
cc_1015 N_A_2049_47#_c_1511_n N_VGND_c_1978_n 0.00910216f $X=10.37 $Y=0.51 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1578_n A_466_369# 0.00283439f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1017 N_VPWR_c_1578_n N_A_560_369#_M1010_d 0.00179277f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1578_n N_A_560_369#_M1015_s 0.0020818f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1580_n N_A_560_369#_c_1782_n 0.00569582f $X=2.045 $Y=2.33 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1581_n N_A_560_369#_c_1782_n 0.0133617f $X=3.845 $Y=2.33 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1596_n N_A_560_369#_c_1782_n 0.0382569f $X=3.76 $Y=2.72 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1578_n N_A_560_369#_c_1782_n 0.0141922f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1581_n N_A_560_369#_c_1806_n 0.00558244f $X=3.845 $Y=2.33 $X2=0
+ $Y2=0
cc_1024 N_VPWR_M1004_d N_A_560_369#_c_1778_n 0.00372198f $X=3.685 $Y=1.845 $X2=0
+ $Y2=0
cc_1025 N_VPWR_c_1581_n N_A_560_369#_c_1778_n 0.0119067f $X=3.845 $Y=2.33 $X2=0
+ $Y2=0
cc_1026 N_VPWR_c_1590_n N_A_560_369#_c_1778_n 0.00414556f $X=5.925 $Y=2.72 $X2=0
+ $Y2=0
cc_1027 N_VPWR_c_1596_n N_A_560_369#_c_1778_n 0.00196122f $X=3.76 $Y=2.72 $X2=0
+ $Y2=0
cc_1028 N_VPWR_c_1578_n N_A_560_369#_c_1778_n 0.00521764f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1029 N_VPWR_c_1581_n N_A_560_369#_c_1781_n 0.0150527f $X=3.845 $Y=2.33 $X2=0
+ $Y2=0
cc_1030 N_VPWR_c_1590_n N_A_560_369#_c_1781_n 0.0166939f $X=5.925 $Y=2.72 $X2=0
+ $Y2=0
cc_1031 N_VPWR_c_1578_n N_A_560_369#_c_1781_n 0.00499134f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1032 N_VPWR_c_1578_n A_644_369# 0.00210687f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1033 N_VPWR_c_1578_n A_1031_413# 0.00220519f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1034 N_VPWR_c_1578_n A_1438_413# 0.00377587f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1035 N_VPWR_c_1578_n N_Q_M1005_s 0.00217091f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1036 N_VPWR_c_1585_n N_Q_c_1895_n 0.0571095f $X=8.99 $Y=1.79 $X2=0 $Y2=0
cc_1037 N_VPWR_c_1586_n N_Q_c_1895_n 0.0575746f $X=9.85 $Y=1.78 $X2=0 $Y2=0
cc_1038 N_VPWR_c_1592_n N_Q_c_1895_n 0.0154695f $X=9.765 $Y=2.72 $X2=0 $Y2=0
cc_1039 N_VPWR_c_1578_n N_Q_c_1895_n 0.0120018f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1040 N_VPWR_c_1578_n N_Q_N_M1002_s 0.00409194f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1041 N_VPWR_c_1589_n Q_N 0.036666f $X=11.695 $Y=1.66 $X2=0 $Y2=0
cc_1042 N_VPWR_c_1599_n Q_N 0.00795791f $X=11.61 $Y=2.72 $X2=0 $Y2=0
cc_1043 N_VPWR_c_1578_n Q_N 0.00867074f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1044 N_VPWR_c_1589_n N_VGND_c_1962_n 0.00811802f $X=11.695 $Y=1.66 $X2=0
+ $Y2=0
cc_1045 N_A_560_369#_c_1782_n A_644_369# 0.00382565f $X=3.42 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_1046 N_A_560_369#_c_1806_n A_644_369# 0.00266005f $X=3.505 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_1047 N_A_560_369#_c_1779_n A_644_369# 9.25434e-19 $X=3.59 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_1048 N_A_560_369#_c_1794_n N_VGND_c_1952_n 9.32728e-19 $X=3.425 $Y=0.36 $X2=0
+ $Y2=0
cc_1049 N_A_560_369#_c_1794_n N_VGND_c_1953_n 0.0135146f $X=3.425 $Y=0.36 $X2=0
+ $Y2=0
cc_1050 N_A_560_369#_c_1771_n N_VGND_c_1953_n 0.00565411f $X=3.51 $Y=0.695 $X2=0
+ $Y2=0
cc_1051 N_A_560_369#_c_1772_n N_VGND_c_1953_n 0.0142693f $X=4.205 $Y=0.78 $X2=0
+ $Y2=0
cc_1052 N_A_560_369#_c_1776_n N_VGND_c_1953_n 0.00987265f $X=4.39 $Y=0.45 $X2=0
+ $Y2=0
cc_1053 N_A_560_369#_c_1772_n N_VGND_c_1954_n 0.00386218f $X=4.205 $Y=0.78 $X2=0
+ $Y2=0
cc_1054 N_A_560_369#_c_1776_n N_VGND_c_1954_n 0.012161f $X=4.39 $Y=0.45 $X2=0
+ $Y2=0
cc_1055 N_A_560_369#_c_1794_n N_VGND_c_1965_n 0.0381281f $X=3.425 $Y=0.36 $X2=0
+ $Y2=0
cc_1056 N_A_560_369#_c_1772_n N_VGND_c_1965_n 0.00256455f $X=4.205 $Y=0.78 $X2=0
+ $Y2=0
cc_1057 N_A_560_369#_M1017_d N_VGND_c_1978_n 0.00217379f $X=2.825 $Y=0.235 $X2=0
+ $Y2=0
cc_1058 N_A_560_369#_M1024_s N_VGND_c_1978_n 0.00195217f $X=4.265 $Y=0.235 $X2=0
+ $Y2=0
cc_1059 N_A_560_369#_c_1794_n N_VGND_c_1978_n 0.012717f $X=3.425 $Y=0.36 $X2=0
+ $Y2=0
cc_1060 N_A_560_369#_c_1772_n N_VGND_c_1978_n 0.00505516f $X=4.205 $Y=0.78 $X2=0
+ $Y2=0
cc_1061 N_A_560_369#_c_1776_n N_VGND_c_1978_n 0.00544577f $X=4.39 $Y=0.45 $X2=0
+ $Y2=0
cc_1062 N_A_560_369#_c_1794_n A_661_47# 0.00210886f $X=3.425 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1063 N_A_560_369#_c_1771_n A_661_47# 0.00222412f $X=3.51 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_1064 N_Q_c_1911_n N_VGND_c_1967_n 0.0188061f $X=9.42 $Y=0.36 $X2=0 $Y2=0
cc_1065 N_Q_M1028_s N_VGND_c_1978_n 0.00215201f $X=9.285 $Y=0.235 $X2=0 $Y2=0
cc_1066 N_Q_c_1893_n N_VGND_c_1978_n 9.95486e-19 $X=9.42 $Y=0.79 $X2=0 $Y2=0
cc_1067 N_Q_c_1911_n N_VGND_c_1978_n 0.0121925f $X=9.42 $Y=0.36 $X2=0 $Y2=0
cc_1068 Q_N N_VGND_c_1960_n 5.93491e-19 $X=11.235 $Y=1.445 $X2=0 $Y2=0
cc_1069 N_Q_N_c_1933_n N_VGND_c_1962_n 0.0271646f $X=11.315 $Y=0.67 $X2=0 $Y2=0
cc_1070 N_Q_N_c_1933_n N_VGND_c_1969_n 0.0142293f $X=11.315 $Y=0.67 $X2=0 $Y2=0
cc_1071 N_Q_N_M1006_s N_VGND_c_1978_n 0.0039413f $X=11.14 $Y=0.235 $X2=0 $Y2=0
cc_1072 N_Q_N_c_1933_n N_VGND_c_1978_n 0.00936105f $X=11.315 $Y=0.67 $X2=0 $Y2=0
cc_1073 N_VGND_c_1978_n A_487_47# 0.00171756f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1074 N_VGND_c_1978_n A_661_47# 0.00152414f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1075 N_VGND_c_1978_n A_1035_47# 0.00272292f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1076 N_VGND_c_1978_n A_1483_47# 0.0111093f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nor4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.240000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.075000 2.635000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.075000 3.535000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.805000 1.075000 5.435000 1.285000 ;
        RECT 5.185000 1.285000 5.435000 1.955000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 3.920000 0.905000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 2.750000 0.255000 3.080000 0.725000 ;
        RECT 3.590000 0.255000 3.920000 0.725000 ;
        RECT 3.630000 1.455000 4.035000 1.625000 ;
        RECT 3.630000 1.625000 3.880000 2.125000 ;
        RECT 3.715000 0.905000 3.920000 1.075000 ;
        RECT 3.715000 1.075000 4.035000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.085000  0.085000 0.345000 0.905000 ;
        RECT 1.015000  0.085000 1.185000 0.555000 ;
        RECT 1.855000  0.085000 2.580000 0.555000 ;
        RECT 3.250000  0.085000 3.420000 0.555000 ;
        RECT 4.090000  0.085000 4.295000 0.895000 ;
        RECT 4.990000  0.085000 5.240000 0.825000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.595000 1.795000 0.805000 2.635000 ;
        RECT 4.990000 2.135000 5.240000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.455000 2.105000 1.625000 ;
      RECT 0.085000 1.625000 0.425000 2.465000 ;
      RECT 0.975000 1.625000 1.225000 2.465000 ;
      RECT 1.395000 1.795000 1.605000 2.295000 ;
      RECT 1.395000 2.295000 3.040000 2.465000 ;
      RECT 1.775000 1.625000 2.105000 2.125000 ;
      RECT 2.275000 1.455000 3.460000 1.625000 ;
      RECT 2.275000 1.625000 2.660000 2.125000 ;
      RECT 2.830000 1.795000 3.040000 2.295000 ;
      RECT 3.210000 1.625000 3.460000 2.295000 ;
      RECT 3.210000 2.295000 4.295000 2.465000 ;
      RECT 4.050000 1.795000 4.295000 2.295000 ;
      RECT 4.320000 1.075000 4.635000 1.245000 ;
      RECT 4.465000 0.380000 4.820000 0.905000 ;
      RECT 4.465000 0.905000 4.635000 1.075000 ;
      RECT 4.465000 1.245000 4.635000 2.035000 ;
      RECT 4.465000 2.035000 4.820000 2.450000 ;
  END
END sky130_fd_sc_hd__nor4b_2
END LIBRARY

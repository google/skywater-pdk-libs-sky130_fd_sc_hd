* File: sky130_fd_sc_hd__a2111oi_1.spice
* Created: Thu Aug 27 13:58:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a2111oi_1  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_D1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.125125 AS=0.481 PD=1.035 PS=2.78 NRD=4.152 NRS=50.76 M=1 R=4.33333
+ SA=75000.7 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_C1_M1000_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.125125 PD=1.02 PS=1.035 NRD=0 NRS=15.228 M=1 R=4.33333
+ SA=75001.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19175 AS=0.12025 PD=1.24 PS=1.02 NRD=2.76 NRS=17.532 M=1 R=4.33333
+ SA=75001.7 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 A_568_47# N_A1_M1002_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.0845
+ AS=0.19175 PD=0.91 PS=1.24 NRD=13.836 NRS=54.456 M=1 R=4.33333 SA=75002.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g A_568_47# VNB NSHORT L=0.15 W=0.65 AD=0.19175
+ AS=0.0845 PD=1.89 PS=0.91 NRD=0.912 NRS=13.836 M=1 R=4.33333 SA=75002.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 A_217_297# N_D1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.1725
+ AS=0.755 PD=1.345 PS=3.51 NRD=23.1278 NRS=68.95 M=1 R=6.66667 SA=75000.7
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1001 A_316_297# N_C1_M1001_g A_217_297# VPB PHIGHVT L=0.15 W=1 AD=0.185
+ AS=0.1725 PD=1.37 PS=1.345 NRD=25.5903 NRS=23.1278 M=1 R=6.66667 SA=75001.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1008 N_A_420_297#_M1008_d N_B1_M1008_g A_316_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.29 AS=0.185 PD=1.58 PS=1.37 NRD=59.0803 NRS=25.5903 M=1 R=6.66667
+ SA=75001.7 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_420_297#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.29 PD=1.275 PS=1.58 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_420_297#_M1005_d N_A2_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.29 AS=0.1375 PD=2.58 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a2111oi_1.pxi.spice"
*
.ends
*
*

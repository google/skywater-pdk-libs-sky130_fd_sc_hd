* File: sky130_fd_sc_hd__o211ai_1.pex.spice
* Created: Tue Sep  1 19:20:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O211AI_1%A1 3 6 8 11 13
r26 11 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.16
+ $X2=0.362 $Y2=1.325
r27 11 13 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.16
+ $X2=0.362 $Y2=0.995
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.16 $X2=0.31 $Y2=1.16
r29 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r30 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%A2 3 7 12 13 15 18
c37 3 0 1.26957e-19 $X=0.835 $Y=1.985
r38 13 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.925 $Y2=1.325
r39 13 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.925 $Y2=0.995
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=1.16 $X2=0.895 $Y2=1.16
r41 9 15 14.7118 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.69 $Y=1.325
+ $X2=0.69 $Y2=1.53
r42 8 12 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.895 $Y2=1.16
r43 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.69
+ $Y2=1.325
r44 7 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.015 $Y=0.56
+ $X2=1.015 $Y2=0.995
r45 3 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.835 $Y=1.985
+ $X2=0.835 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%B1 3 7 8 9 13 15
c33 8 0 1.26957e-19 $X=1.61 $Y=1.19
r34 13 16 51.4573 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.465 $Y=1.16
+ $X2=1.465 $Y2=1.355
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.16
+ $X2=1.465 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.435
+ $Y=1.16 $X2=1.435 $Y2=1.16
r37 8 9 9.99518 $w=4.15e-07 $l=3.4e-07 $layer=LI1_cond $X=1.547 $Y=1.19
+ $X2=1.547 $Y2=1.53
r38 8 14 0.881928 $w=4.15e-07 $l=3e-08 $layer=LI1_cond $X=1.547 $Y=1.19
+ $X2=1.547 $Y2=1.16
r39 7 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.555 $Y=0.56
+ $X2=1.555 $Y2=0.995
r40 3 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.375 $Y=1.985
+ $X2=1.375 $Y2=1.355
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%C1 1 3 6 8 13 14
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.16 $X2=2.135 $Y2=1.16
r30 10 13 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.915 $Y=1.16
+ $X2=2.135 $Y2=1.16
r31 8 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.135 $Y=1.53
+ $X2=2.135 $Y2=1.16
r32 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.325
+ $X2=1.915 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.915 $Y=1.325
+ $X2=1.915 $Y2=1.985
r34 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%VPWR 1 2 7 9 15 17 19 26 27 33
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 27 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r42 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.61 $Y2=2.72
r43 24 26 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r45 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 20 30 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r47 20 22 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 19 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 17 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 17 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r52 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=2.635
+ $X2=1.61 $Y2=2.72
r53 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.61 $Y=2.635
+ $X2=1.61 $Y2=2.36
r54 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66 $X2=0.26
+ $Y2=2.34
r55 7 30 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r56 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r57 2 15 600 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.61 $Y2=2.36
r58 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r59 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%Y 1 2 3 15 17 21 24 25 27 34
r39 27 34 0.851446 $w=5.88e-07 $l=4.2e-08 $layer=LI1_cond $X=2.53 $Y=0.55
+ $X2=2.572 $Y2=0.55
r40 27 30 1.21635 $w=5.88e-07 $l=6e-08 $layer=LI1_cond $X=2.53 $Y=0.55 $X2=2.47
+ $Y2=0.55
r41 23 25 1.69291 $w=6.48e-07 $l=9.2e-08 $layer=LI1_cond $X=2.48 $Y=2.14
+ $X2=2.572 $Y2=2.14
r42 23 24 14.5837 $w=6.48e-07 $l=5.05e-07 $layer=LI1_cond $X=2.48 $Y=2.14
+ $X2=1.975 $Y2=2.14
r43 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.11 $Y=1.93 $X2=1.11
+ $Y2=2.02
r44 17 19 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.11 $Y=1.68
+ $X2=1.11 $Y2=1.93
r45 15 25 7.6405 $w=2.05e-07 $l=3.25e-07 $layer=LI1_cond $X=2.572 $Y=1.815
+ $X2=2.572 $Y2=2.14
r46 14 34 7.03101 $w=2.05e-07 $l=2.95e-07 $layer=LI1_cond $X=2.572 $Y=0.845
+ $X2=2.572 $Y2=0.55
r47 14 15 52.4789 $w=2.03e-07 $l=9.7e-07 $layer=LI1_cond $X=2.572 $Y=0.845
+ $X2=2.572 $Y2=1.815
r48 13 19 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=1.93
+ $X2=1.11 $Y2=1.93
r49 13 24 35.0744 $w=2.28e-07 $l=7e-07 $layer=LI1_cond $X=1.275 $Y=1.93
+ $X2=1.975 $Y2=1.93
r50 3 23 150 $w=1.7e-07 $l=7.40523e-07 $layer=licon1_PDIFF $count=4 $X=1.99
+ $Y=1.485 $X2=2.48 $Y2=2.02
r51 2 21 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=1.485 $X2=1.11 $Y2=2.02
r52 2 17 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.485 $X2=1.11 $Y2=1.68
r53 1 30 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=1.99
+ $Y=0.235 $X2=2.47 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%A_27_47# 1 2 9 11 12 13 15
r24 13 18 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.29 $Y=0.615
+ $X2=1.29 $Y2=0.72
r25 13 15 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.29 $Y=0.615
+ $X2=1.29 $Y2=0.38
r26 11 18 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=0.72
+ $X2=1.29 $Y2=0.72
r27 11 12 36.9697 $w=2.08e-07 $l=7e-07 $layer=LI1_cond $X=1.125 $Y=0.72
+ $X2=0.425 $Y2=0.72
r28 7 12 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.425 $Y2=0.72
r29 7 9 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.26 $Y2=0.38
r30 2 18 182 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.29 $Y2=0.72
r31 2 15 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.29 $Y2=0.38
r32 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211AI_1%VGND 1 6 8 10 20 21 24
r30 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r31 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r32 18 21 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r33 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r34 17 20 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r35 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r36 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.76
+ $Y2=0
r37 15 17 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r38 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.76
+ $Y2=0
r39 10 12 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r40 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r41 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r42 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r43 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.36
r44 1 6 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.76 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__a41oi_4.spice
* Created: Thu Aug 27 14:06:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a41oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a41oi_4  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_B1_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.4
+ A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_B1_M1024_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1024_d N_B1_M1025_g N_Y_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1036 N_VGND_M1036_d N_B1_M1036_g N_Y_M1025_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g N_A_493_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1003_d N_A1_M1004_g N_A_493_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1009_d N_A1_M1009_g N_A_493_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1009_d N_A1_M1012_g N_A_493_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1006 N_A_493_47#_M1012_s N_A2_M1006_g N_A_911_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1010 N_A_493_47#_M1010_d N_A2_M1010_g N_A_911_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1011 N_A_493_47#_M1010_d N_A2_M1011_g N_A_911_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1039 N_A_493_47#_M1039_d N_A2_M1039_g N_A_911_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_1269_47#_M1000_d N_A3_M1000_g N_A_911_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1029 N_A_1269_47#_M1029_d N_A3_M1029_g N_A_911_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1033 N_A_1269_47#_M1029_d N_A3_M1033_g N_A_911_47#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1034 N_A_1269_47#_M1034_d N_A3_M1034_g N_A_911_47#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A4_M1001_g N_A_1269_47#_M1034_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1001_d N_A4_M1008_g N_A_1269_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_A4_M1016_g N_A_1269_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1016_d N_A4_M1038_g N_A_1269_47#_M1038_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1885 PD=0.92 PS=1.88 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75009.4 A=0.15 P=2.3 MULT=1
MM1013 N_Y_M1005_d N_B1_M1013_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75008.9 A=0.15 P=2.3 MULT=1
MM1026 N_Y_M1026_d N_B1_M1026_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75008.5 A=0.15 P=2.3 MULT=1
MM1035 N_Y_M1026_d N_B1_M1035_g N_A_27_297#_M1035_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.29 PD=1.27 PS=1.58 NRD=0 NRS=60.0653 M=1 R=6.66667 SA=75001.4
+ SB=75008.1 A=0.15 P=2.3 MULT=1
MM1002 N_A_27_297#_M1035_s N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.29 AS=0.305 PD=1.58 PS=1.61 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.2
+ SB=75007.4 A=0.15 P=2.3 MULT=1
MM1018 N_A_27_297#_M1018_d N_A1_M1018_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.305 PD=1.27 PS=1.61 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1022 N_A_27_297#_M1018_d N_A1_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.4
+ SB=75006.2 A=0.15 P=2.3 MULT=1
MM1030 N_A_27_297#_M1030_d N_A1_M1030_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1825 AS=0.135 PD=1.365 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.8
+ SB=75005.8 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A2_M1014_g N_A_27_297#_M1030_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1825 PD=1.27 PS=1.365 NRD=0 NRS=17.73 M=1 R=6.66667 SA=75004.3
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1014_d N_A2_M1017_g N_A_27_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.7
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A2_M1019_g N_A_27_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3375 AS=0.135 PD=1.675 PS=1.27 NRD=5.8903 NRS=0 M=1 R=6.66667 SA=75005.1
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1019_d N_A2_M1028_g N_A_27_297#_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3375 AS=0.145 PD=1.675 PS=1.29 NRD=4.9053 NRS=2.9353 M=1 R=6.66667
+ SA=75006 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A3_M1007_g N_A_27_297#_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.4
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1027 N_VPWR_M1007_d N_A3_M1027_g N_A_27_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.8
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1031 N_VPWR_M1031_d N_A3_M1031_g N_A_27_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1037 N_VPWR_M1031_d N_A3_M1037_g N_A_27_297#_M1037_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.7
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 N_A_27_297#_M1037_s N_A4_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1020 N_A_27_297#_M1020_d N_A4_M1020_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1023 N_A_27_297#_M1020_d N_A4_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1032 N_A_27_297#_M1032_d N_A4_M1032_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.29 AS=0.135 PD=2.58 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75009.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.8525 P=24.21
*
.include "sky130_fd_sc_hd__a41oi_4.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 7.885000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965000 1.075000 6.295000 1.445000 ;
        RECT 5.965000 1.445000 8.265000 1.615000 ;
        RECT 8.095000 1.075000 9.575000 1.275000 ;
        RECT 8.095000 1.275000 8.265000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 0.995000 5.285000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415000 0.995000 3.765000 1.325000 ;
        RECT 3.595000 1.325000 3.765000 1.445000 ;
        RECT 3.595000 1.445000 5.795000 1.615000 ;
        RECT 5.465000 1.075000 5.795000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.335000 1.275000 ;
    END
  END C1
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.905000 ;
        RECT 0.575000 1.445000 1.705000 1.615000 ;
        RECT 0.575000 1.615000 0.825000 2.125000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 1.615000 1.665000 2.125000 ;
        RECT 1.505000 0.905000 1.705000 1.095000 ;
        RECT 1.505000 1.095000 3.245000 1.275000 ;
        RECT 1.505000 1.275000 1.705000 1.445000 ;
        RECT 3.075000 0.645000 5.680000 0.735000 ;
        RECT 3.075000 0.735000 7.765000 0.820000 ;
        RECT 3.075000 0.820000 3.245000 1.095000 ;
        RECT 5.510000 0.820000 6.460000 0.905000 ;
        RECT 6.290000 0.645000 7.765000 0.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  1.445000 0.405000 2.295000 ;
      RECT 0.090000  2.295000 2.125000 2.465000 ;
      RECT 0.115000  0.085000 0.365000 0.895000 ;
      RECT 0.995000  1.785000 1.245000 2.295000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.875000  0.085000 2.045000 0.645000 ;
      RECT 1.875000  0.645000 2.905000 0.925000 ;
      RECT 1.875000  1.445000 3.030000 1.615000 ;
      RECT 1.875000  1.615000 2.125000 2.295000 ;
      RECT 2.235000  0.255000 5.585000 0.425000 ;
      RECT 2.235000  0.425000 2.610000 0.475000 ;
      RECT 2.315000  1.795000 2.565000 2.215000 ;
      RECT 2.315000  2.215000 6.005000 2.465000 ;
      RECT 2.735000  0.595000 2.905000 0.645000 ;
      RECT 2.735000  1.615000 3.030000 1.835000 ;
      RECT 2.735000  1.835000 5.585000 2.045000 ;
      RECT 3.035000  0.425000 5.585000 0.475000 ;
      RECT 5.755000  1.785000 8.605000 2.045000 ;
      RECT 5.755000  2.045000 6.005000 2.215000 ;
      RECT 5.835000  0.085000 6.005000 0.555000 ;
      RECT 6.175000  0.255000 8.185000 0.475000 ;
      RECT 6.175000  2.215000 8.185000 2.635000 ;
      RECT 7.935000  0.475000 8.185000 0.725000 ;
      RECT 7.935000  0.725000 9.025000 0.905000 ;
      RECT 8.355000  0.085000 8.525000 0.555000 ;
      RECT 8.355000  2.045000 8.525000 2.465000 ;
      RECT 8.435000  1.445000 9.405000 1.615000 ;
      RECT 8.435000  1.615000 8.605000 1.785000 ;
      RECT 8.695000  0.255000 9.025000 0.725000 ;
      RECT 8.775000  1.795000 8.945000 2.635000 ;
      RECT 9.155000  1.615000 9.405000 2.465000 ;
      RECT 9.195000  0.085000 9.365000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_4
END LIBRARY

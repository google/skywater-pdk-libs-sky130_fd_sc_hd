* File: sky130_fd_sc_hd__a22oi_2.spice.pex
* Created: Thu Aug 27 14:02:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A22OI_2%B2 1 3 6 8 10 13 15 16 24
c40 16 0 1.52846e-19 $X=0.695 $Y=1.19
c41 8 0 8.29508e-20 $X=0.89 $Y=0.995
r42 23 24 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r43 20 23 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.41 $Y=1.16 $X2=0.47
+ $Y2=1.16
r44 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r45 16 21 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.41 $Y2=1.175
r46 15 21 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.41 $Y2=1.175
r47 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r48 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r49 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r50 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r51 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r52 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r53 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%B1 1 3 6 8 10 13 15 16 24
c46 24 0 1.52846e-19 $X=1.73 $Y=1.16
r47 22 24 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.4 $Y=1.16 $X2=1.73
+ $Y2=1.16
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=1.16 $X2=1.4 $Y2=1.16
r49 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.31 $Y=1.16 $X2=1.4
+ $Y2=1.16
r50 16 23 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.4 $Y2=1.175
r51 15 23 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.4 $Y2=1.175
r52 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r54 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r56 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%A1 1 3 6 8 10 13 15 16 24
r49 23 24 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=3.09 $Y2=1.16
r50 20 23 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.61 $Y=1.16 $X2=2.67
+ $Y2=1.16
r51 15 16 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=3.015 $Y2=1.175
r52 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.16 $X2=2.61 $Y2=1.16
r53 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.325
+ $X2=3.09 $Y2=1.16
r54 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.09 $Y=1.325
+ $X2=3.09 $Y2=1.985
r55 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=1.16
r56 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=0.56
r57 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.325
+ $X2=2.67 $Y2=1.16
r58 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.325 $X2=2.67
+ $Y2=1.985
r59 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=1.16
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995 $X2=2.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%A2 1 3 6 8 10 13 15 16 24
c39 1 0 8.29508e-20 $X=3.51 $Y=0.995
r40 22 24 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.6 $Y=1.16 $X2=3.93
+ $Y2=1.16
r41 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.16 $X2=3.6 $Y2=1.16
r42 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.51 $Y=1.16 $X2=3.6
+ $Y2=1.16
r43 16 23 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=3.6 $Y2=1.175
r44 15 23 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.6 $Y2=1.175
r45 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=1.325
+ $X2=3.93 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.93 $Y=1.325
+ $X2=3.93 $Y2=1.985
r47 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=0.56
r49 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=1.325
+ $X2=3.51 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.325 $X2=3.51
+ $Y2=1.985
r51 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995 $X2=3.51
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%Y 1 2 3 4 5 18 20 21 24 26 28 32 33 34 35 36
+ 47 54 60
c80 60 0 8.29508e-20 $X=2.88 $Y=0.76
c81 28 0 8.29508e-20 $X=1.87 $Y=0.76
r82 52 54 0.149668 $w=3.83e-07 $l=5e-09 $layer=LI1_cond $X=1.967 $Y=1.655
+ $X2=1.967 $Y2=1.66
r83 44 47 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=2.015 $Y=0.845
+ $X2=2.015 $Y2=0.85
r84 36 54 6.28605 $w=3.83e-07 $l=2.1e-07 $layer=LI1_cond $X=1.967 $Y=1.87
+ $X2=1.967 $Y2=1.66
r85 35 45 2.82881 $w=3.37e-07 $l=1.06325e-07 $layer=LI1_cond $X=1.967 $Y=1.57
+ $X2=2.015 $Y2=1.485
r86 35 52 2.82881 $w=3.37e-07 $l=8.5e-08 $layer=LI1_cond $X=1.967 $Y=1.57
+ $X2=1.967 $Y2=1.655
r87 35 45 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=2.015 $Y=1.465
+ $X2=2.015 $Y2=1.485
r88 34 35 10.9283 $w=2.88e-07 $l=2.75e-07 $layer=LI1_cond $X=2.015 $Y=1.19
+ $X2=2.015 $Y2=1.465
r89 33 44 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.76
+ $X2=2.015 $Y2=0.845
r90 33 60 34.3775 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=2.16 $Y=0.76
+ $X2=2.88 $Y2=0.76
r91 33 34 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=2.015 $Y=0.89
+ $X2=2.015 $Y2=1.19
r92 33 47 1.58958 $w=2.88e-07 $l=4e-08 $layer=LI1_cond $X=2.015 $Y=0.89
+ $X2=2.015 $Y2=0.85
r93 28 33 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.87 $Y=0.76
+ $X2=2.015 $Y2=0.76
r94 28 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.87 $Y=0.76
+ $X2=1.52 $Y2=0.76
r95 27 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=1.57
+ $X2=1.1 $Y2=1.57
r96 26 35 3.89502 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.775 $Y=1.57
+ $X2=1.967 $Y2=1.57
r97 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=1.57
+ $X2=1.265 $Y2=1.57
r98 22 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.655 $X2=1.1
+ $Y2=1.57
r99 22 24 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.1 $Y=1.655 $X2=1.1
+ $Y2=1.66
r100 20 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.57
+ $X2=1.1 $Y2=1.57
r101 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.935 $Y=1.57
+ $X2=0.345 $Y2=1.57
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=1.655
+ $X2=0.345 $Y2=1.57
r103 16 18 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.22 $Y=1.655
+ $X2=0.22 $Y2=1.8
r104 5 54 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.66
r105 4 24 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.66
r106 3 18 300 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.8
r107 2 60 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.76
r108 1 30 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%A_109_297# 1 2 3 4 5 18 20 21 24 26 29 31 32
+ 33 36 40 44 48 51
r72 44 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.14 $Y=1.66
+ $X2=4.14 $Y2=2.34
r73 42 44 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.14 $Y=1.655
+ $X2=4.14 $Y2=1.66
r74 41 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=1.57
+ $X2=3.3 $Y2=1.57
r75 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.975 $Y=1.57
+ $X2=4.14 $Y2=1.655
r76 40 41 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.975 $Y=1.57
+ $X2=3.465 $Y2=1.57
r77 36 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.3 $Y=1.66 $X2=3.3
+ $Y2=2.34
r78 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=1.655 $X2=3.3
+ $Y2=1.57
r79 34 36 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.3 $Y=1.655 $X2=3.3
+ $Y2=1.66
r80 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=1.57
+ $X2=3.3 $Y2=1.57
r81 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.135 $Y=1.57
+ $X2=2.625 $Y2=1.57
r82 29 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=2.295 $X2=2.5
+ $Y2=2.38
r83 29 31 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.5 $Y=2.295
+ $X2=2.5 $Y2=1.66
r84 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.5 $Y=1.655
+ $X2=2.625 $Y2=1.57
r85 28 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.5 $Y=1.655 $X2=2.5
+ $Y2=1.66
r86 27 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.38
+ $X2=1.52 $Y2=2.38
r87 26 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=2.5 $Y2=2.38
r88 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=1.605 $Y2=2.38
r89 22 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.295
+ $X2=1.52 $Y2=2.38
r90 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=2.295
+ $X2=1.52 $Y2=2
r91 20 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.38
+ $X2=1.52 $Y2=2.38
r92 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=2.38
+ $X2=0.765 $Y2=2.38
r93 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.64 $Y=2.295
+ $X2=0.765 $Y2=2.38
r94 16 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.64 $Y=2.295
+ $X2=0.64 $Y2=2
r95 5 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.34
r96 5 44 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=1.66
r97 4 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2.34
r98 4 36 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.66
r99 3 50 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=2.34
r100 3 31 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=1.66
r101 2 24 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
r102 1 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%VPWR 1 2 9 13 16 17 19 20 21 23 38 39
r57 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r58 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r59 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 23 33 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r63 23 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 21 32 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 21 26 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 19 35 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.72 $Y2=2.72
r68 18 38 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=4.37 $Y2=2.72
r69 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.72 $Y2=2.72
r70 16 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.88 $Y2=2.72
r72 15 35 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.88 $Y2=2.72
r74 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2.72
r75 11 13 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2
r76 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=2.635 $X2=2.88
+ $Y2=2.72
r77 7 9 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2
r78 2 13 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2
r79 1 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%A_27_47# 1 2 3 10 13 14 19 21
r37 19 21 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=1.185 $Y=0.38
+ $X2=1.94 $Y2=0.38
r38 16 18 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.1 $Y=0.68 $X2=1.1
+ $Y2=0.57
r39 15 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.1 $Y=0.505
+ $X2=1.185 $Y2=0.38
r40 15 18 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.1 $Y=0.505 $X2=1.1
+ $Y2=0.57
r41 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.015 $Y=0.765
+ $X2=1.1 $Y2=0.68
r42 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.765
+ $X2=0.345 $Y2=0.765
r43 10 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=0.68
+ $X2=0.345 $Y2=0.765
r44 10 12 5.368 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.22 $Y=0.68 $X2=0.22
+ $Y2=0.57
r45 3 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.42
r46 2 18 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.57
r47 1 12 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%VGND 1 2 9 12 13 14 17 19 32 33 41
r62 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r63 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r64 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r65 27 30 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r66 27 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r67 26 29 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r68 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r70 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r71 17 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r72 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 14 41 8.91899 $w=4.98e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r74 14 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r75 14 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0 $X2=0.515
+ $Y2=0
r76 14 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0 $X2=0.845
+ $Y2=0
r77 12 29 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.45
+ $Y2=0
r78 12 13 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.72
+ $Y2=0
r79 11 32 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=4.37
+ $Y2=0
r80 11 13 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.72
+ $Y2=0
r81 7 13 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085 $X2=3.72
+ $Y2=0
r82 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.4
r83 2 9 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.4
r84 1 41 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_2%A_467_47# 1 2 3 10 18 19 20
r27 20 22 4.19375 $w=3.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.215 $Y=0.68
+ $X2=4.215 $Y2=0.57
r28 18 20 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=4.055 $Y=0.765
+ $X2=4.215 $Y2=0.68
r29 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.055 $Y=0.765
+ $X2=3.385 $Y2=0.765
r30 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.3 $Y=0.68
+ $X2=3.385 $Y2=0.765
r31 15 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.3 $Y=0.68 $X2=3.3
+ $Y2=0.57
r32 14 17 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.3 $Y=0.505 $X2=3.3
+ $Y2=0.57
r33 10 14 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.215 $Y=0.38
+ $X2=3.3 $Y2=0.505
r34 10 12 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=3.215 $Y=0.38
+ $X2=2.46 $Y2=0.38
r35 3 22 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.57
r36 2 17 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.57
r37 1 12 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.42
.ends


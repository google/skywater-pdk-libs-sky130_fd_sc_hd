* File: sky130_fd_sc_hd__ha_2.spice
* Created: Tue Sep  1 19:09:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ha_2.pex.spice"
.subckt sky130_fd_sc_hd__ha_2  VNB VPB B A VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_79_21#_M1015_g N_SUM_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10075 PD=1.82 PS=0.96 NRD=0 NRS=6.456 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_A_79_21#_M1016_g N_SUM_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10075 PD=1.82 PS=0.96 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_389_47#_M1012_d N_A_342_199#_M1012_g N_A_79_21#_M1012_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_389_47#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_389_47#_M1017_d N_A_M1017_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 A_766_47# N_B_M1013_g N_A_342_199#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_M1014_g A_766_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.0441 PD=0.765421 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_COUT_M1002_d N_A_342_199#_M1002_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.65 AD=0.10075 AS=0.11785 PD=0.96 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_COUT_M1002_d N_A_342_199#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10075 AS=0.169 PD=0.96 PS=1.82 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_79_21#_M1004_g N_SUM_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.155 PD=2.52 PS=1.31 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75000.2
+ SB=75003.3 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_79_21#_M1010_g N_SUM_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.35561 AS=0.155 PD=2.15244 PS=1.31 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1005 N_A_79_21#_M1005_d N_A_342_199#_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.22759 PD=0.91 PS=1.37756 NRD=0 NRS=150.823 M=1 R=4.26667
+ SA=75001.6 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1003 A_468_369# N_B_M1003_g N_A_79_21#_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.128 AS=0.0864 PD=1.04 PS=0.91 NRD=44.6205 NRS=0 M=1 R=4.26667 SA=75002
+ SB=75003 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_468_369# VPB PHIGHVT L=0.15 W=0.64 AD=0.2272
+ AS=0.128 PD=1.35 PS=1.04 NRD=13.8491 NRS=44.6205 M=1 R=4.26667 SA=75002.5
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1009 N_A_342_199#_M1009_d N_B_M1009_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0928 AS=0.2272 PD=0.93 PS=1.35 NRD=1.5366 NRS=13.8491 M=1 R=4.26667
+ SA=75003.4 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_342_199#_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116293 AS=0.0928 PD=1.03415 PS=0.93 NRD=15.3857 NRS=1.5366 M=1 R=4.26667
+ SA=75003.8 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_COUT_M1000_d N_A_342_199#_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.181707 PD=1.31 PS=1.61585 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_COUT_M1000_d N_A_342_199#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.26 PD=1.31 PS=2.52 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__ha_2.pxi.spice"
*
.ends
*
*

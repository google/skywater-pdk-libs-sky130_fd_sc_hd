* File: sky130_fd_sc_hd__a21bo_2.pxi.spice
* Created: Tue Sep  1 18:51:27 2020
* 
x_PM_SKY130_FD_SC_HD__A21BO_2%A_79_21# N_A_79_21#_M1008_d N_A_79_21#_M1006_s
+ N_A_79_21#_M1009_g N_A_79_21#_M1001_g N_A_79_21#_M1010_g N_A_79_21#_M1007_g
+ N_A_79_21#_c_75_n N_A_79_21#_c_76_n N_A_79_21#_c_77_n N_A_79_21#_c_81_n
+ N_A_79_21#_c_94_p N_A_79_21#_c_144_p N_A_79_21#_c_125_p N_A_79_21#_c_82_n
+ N_A_79_21#_c_83_n N_A_79_21#_c_84_n N_A_79_21#_c_90_p N_A_79_21#_c_78_n
+ N_A_79_21#_c_86_n N_A_79_21#_c_102_p N_A_79_21#_c_103_p
+ PM_SKY130_FD_SC_HD__A21BO_2%A_79_21#
x_PM_SKY130_FD_SC_HD__A21BO_2%B1_N N_B1_N_M1003_g N_B1_N_M1002_g B1_N
+ N_B1_N_c_175_n N_B1_N_c_176_n PM_SKY130_FD_SC_HD__A21BO_2%B1_N
x_PM_SKY130_FD_SC_HD__A21BO_2%A_297_93# N_A_297_93#_M1003_d N_A_297_93#_M1002_d
+ N_A_297_93#_c_210_n N_A_297_93#_M1008_g N_A_297_93#_M1006_g
+ N_A_297_93#_c_211_n N_A_297_93#_c_216_n N_A_297_93#_c_212_n
+ N_A_297_93#_c_217_n N_A_297_93#_c_213_n PM_SKY130_FD_SC_HD__A21BO_2%A_297_93#
x_PM_SKY130_FD_SC_HD__A21BO_2%A1 N_A1_M1005_g N_A1_M1011_g A1 N_A1_c_266_n
+ N_A1_c_267_n N_A1_c_268_n PM_SKY130_FD_SC_HD__A21BO_2%A1
x_PM_SKY130_FD_SC_HD__A21BO_2%A2 N_A2_M1000_g N_A2_M1004_g A2 N_A2_c_305_n
+ N_A2_c_306_n A2 PM_SKY130_FD_SC_HD__A21BO_2%A2
x_PM_SKY130_FD_SC_HD__A21BO_2%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_M1005_d
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_336_n VPWR N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_330_n
+ N_VPWR_c_340_n PM_SKY130_FD_SC_HD__A21BO_2%VPWR
x_PM_SKY130_FD_SC_HD__A21BO_2%X N_X_M1009_d N_X_M1001_s N_X_c_397_n N_X_c_398_n
+ N_X_c_402_n N_X_c_404_n N_X_c_409_n X N_X_c_421_n
+ PM_SKY130_FD_SC_HD__A21BO_2%X
x_PM_SKY130_FD_SC_HD__A21BO_2%A_485_297# N_A_485_297#_M1006_d
+ N_A_485_297#_M1004_d N_A_485_297#_c_437_n N_A_485_297#_c_435_n
+ N_A_485_297#_c_432_n PM_SKY130_FD_SC_HD__A21BO_2%A_485_297#
x_PM_SKY130_FD_SC_HD__A21BO_2%VGND N_VGND_M1009_s N_VGND_M1010_s N_VGND_M1008_s
+ N_VGND_M1000_d N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n N_VGND_c_463_n
+ N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n VGND
+ N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n
+ PM_SKY130_FD_SC_HD__A21BO_2%VGND
cc_1 VNB N_A_79_21#_M1009_g 0.0208366f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_79_21#_M1001_g 4.87965e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_A_79_21#_M1010_g 0.0209558f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.56
cc_4 VNB N_A_79_21#_M1007_g 4.47996e-19 $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.985
cc_5 VNB N_A_79_21#_c_75_n 0.0108564f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_6 VNB N_A_79_21#_c_76_n 0.0131562f $X=-0.19 $Y=-0.24 $X2=0.825 $Y2=1.16
cc_7 VNB N_A_79_21#_c_77_n 0.0100782f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_8 VNB N_A_79_21#_c_78_n 0.00293881f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.505
cc_9 VNB B1_N 0.00733004f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_B1_N_c_175_n 0.0246054f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_11 VNB N_B1_N_c_176_n 0.019191f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_12 VNB N_A_297_93#_c_210_n 0.0533769f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_13 VNB N_A_297_93#_c_211_n 0.00393835f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.025
cc_14 VNB N_A_297_93#_c_212_n 0.00435252f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.985
cc_15 VNB N_A_297_93#_c_213_n 0.0064793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_266_n 0.020316f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_17 VNB N_A1_c_267_n 0.0107836f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_18 VNB N_A1_c_268_n 0.0164055f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_19 VNB A2 0.0120009f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_A2_c_305_n 0.0317419f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_21 VNB N_A2_c_306_n 0.0207298f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_22 VNB N_VPWR_c_330_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.14 $Y2=1.675
cc_23 VNB X 0.0205786f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_24 VNB N_VGND_c_460_n 0.00994884f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_25 VNB N_VGND_c_461_n 0.0180355f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.025
cc_26 VNB N_VGND_c_462_n 0.00435274f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.295
cc_27 VNB N_VGND_c_463_n 0.00899266f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_28 VNB N_VGND_c_464_n 0.010974f $X=-0.19 $Y=-0.24 $X2=0.825 $Y2=1.16
cc_29 VNB N_VGND_c_465_n 0.0258516f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=1.495
cc_30 VNB N_VGND_c_466_n 0.0179964f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=1.16
cc_31 VNB N_VGND_c_467_n 0.00384695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_468_n 0.0222114f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=2.105
cc_33 VNB N_VGND_c_469_n 0.0256823f $X=-0.19 $Y=-0.24 $X2=2.14 $Y2=1.895
cc_34 VNB N_VGND_c_470_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_471_n 0.213961f $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=0.73
cc_36 VPB N_A_79_21#_M1001_g 0.0221747f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A_79_21#_M1007_g 0.022489f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_38 VPB N_A_79_21#_c_81_n 0.00110605f $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.16
cc_39 VPB N_A_79_21#_c_82_n 0.0133751f $X=-0.19 $Y=1.305 $X2=1.975 $Y2=2
cc_40 VPB N_A_79_21#_c_83_n 2.08527e-19 $X=-0.19 $Y=1.305 $X2=1.285 $Y2=2
cc_41 VPB N_A_79_21#_c_84_n 0.00994564f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=2.105
cc_42 VPB N_A_79_21#_c_78_n 0.00108343f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.505
cc_43 VPB N_A_79_21#_c_86_n 7.80569e-19 $X=-0.19 $Y=1.305 $X2=2.1 $Y2=2
cc_44 VPB N_B1_N_M1002_g 0.0217604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB B1_N 0.00332064f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_46 VPB N_B1_N_c_175_n 0.00456326f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_47 VPB N_A_297_93#_c_210_n 0.0100666f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.025
cc_48 VPB N_A_297_93#_M1006_g 0.0220828f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_49 VPB N_A_297_93#_c_216_n 0.00520771f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_50 VPB N_A_297_93#_c_217_n 0.00338429f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_51 VPB N_A_297_93#_c_213_n 0.00205602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A1_M1005_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A1_c_266_n 0.0046406f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_54 VPB N_A1_c_267_n 0.00209405f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_55 VPB N_A2_M1004_g 0.0221372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB A2 0.0127749f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_57 VPB N_A2_c_305_n 0.00814369f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_58 VPB N_VPWR_c_331_n 0.0102396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_332_n 0.0133561f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_60 VPB N_VPWR_c_333_n 0.0050483f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_61 VPB N_VPWR_c_334_n 0.0046277f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_62 VPB N_VPWR_c_335_n 0.0393493f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_63 VPB N_VPWR_c_336_n 0.00323576f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_64 VPB N_VPWR_c_337_n 0.015606f $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.495
cc_65 VPB N_VPWR_c_338_n 0.0178228f $X=-0.19 $Y=1.305 $X2=2.14 $Y2=2.11
cc_66 VPB N_VPWR_c_330_n 0.051081f $X=-0.19 $Y=1.305 $X2=2.14 $Y2=1.675
cc_67 VPB N_VPWR_c_340_n 0.00631318f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=2
cc_68 VPB X 0.00900657f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_69 VPB N_A_485_297#_c_432_n 0.0251772f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_70 N_A_79_21#_M1007_g N_B1_N_M1002_g 0.0203057f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_81_n N_B1_N_M1002_g 8.68148e-19 $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_82_n N_B1_N_M1002_g 0.0127401f $X=1.975 $Y=2 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_90_p N_B1_N_M1002_g 0.00261208f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_74 N_A_79_21#_M1010_g B1_N 2.38958e-19 $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_77_n B1_N 0.00346303f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_81_n B1_N 0.0203601f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_94_p B1_N 0.0176891f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_82_n B1_N 0.00398434f $X=1.975 $Y=2 $X2=0 $Y2=0
cc_79 N_A_79_21#_M1010_g N_B1_N_c_175_n 0.0117365f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_80 N_A_79_21#_M1010_g N_B1_N_c_176_n 0.0112338f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_82_n N_A_297_93#_M1002_d 0.00217362f $X=1.975 $Y=2 $X2=0
+ $Y2=0
cc_82 N_A_79_21#_c_82_n N_A_297_93#_c_210_n 3.30674e-19 $X=1.975 $Y=2 $X2=0
+ $Y2=0
cc_83 N_A_79_21#_c_78_n N_A_297_93#_c_210_n 0.0130297f $X=2.43 $Y=1.505 $X2=0
+ $Y2=0
cc_84 N_A_79_21#_c_86_n N_A_297_93#_c_210_n 0.00140592f $X=2.1 $Y=2 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_102_p N_A_297_93#_c_210_n 0.00542686f $X=2.43 $Y=1.59 $X2=0
+ $Y2=0
cc_86 N_A_79_21#_c_103_p N_A_297_93#_c_210_n 0.00674728f $X=2.575 $Y=0.73 $X2=0
+ $Y2=0
cc_87 N_A_79_21#_c_78_n N_A_297_93#_M1006_g 0.00521756f $X=2.43 $Y=1.505 $X2=0
+ $Y2=0
cc_88 N_A_79_21#_c_102_p N_A_297_93#_M1006_g 0.0136386f $X=2.43 $Y=1.59 $X2=0
+ $Y2=0
cc_89 N_A_79_21#_c_78_n N_A_297_93#_c_211_n 0.00557939f $X=2.43 $Y=1.505 $X2=0
+ $Y2=0
cc_90 N_A_79_21#_c_78_n N_A_297_93#_c_216_n 0.00590914f $X=2.43 $Y=1.505 $X2=0
+ $Y2=0
cc_91 N_A_79_21#_c_102_p N_A_297_93#_c_216_n 0.00362224f $X=2.43 $Y=1.59 $X2=0
+ $Y2=0
cc_92 N_A_79_21#_c_103_p N_A_297_93#_c_212_n 0.00633165f $X=2.575 $Y=0.73 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_82_n N_A_297_93#_c_217_n 0.0261985f $X=1.975 $Y=2 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_90_p N_A_297_93#_c_217_n 0.003603f $X=2.14 $Y=1.77 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_102_p N_A_297_93#_c_217_n 0.00935054f $X=2.43 $Y=1.59 $X2=0
+ $Y2=0
cc_96 N_A_79_21#_c_82_n N_A_297_93#_c_213_n 0.00372524f $X=1.975 $Y=2 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_c_78_n N_A_297_93#_c_213_n 0.0242722f $X=2.43 $Y=1.505 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_86_n N_A_297_93#_c_213_n 0.00260016f $X=2.1 $Y=2 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_102_p N_A_297_93#_c_213_n 0.00847745f $X=2.43 $Y=1.59 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_78_n N_A1_M1005_g 5.50095e-19 $X=2.43 $Y=1.505 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_102_p N_A1_M1005_g 0.00185588f $X=2.43 $Y=1.59 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_78_n N_A1_c_266_n 0.00187393f $X=2.43 $Y=1.505 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_103_p N_A1_c_266_n 0.00222434f $X=2.575 $Y=0.73 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_78_n N_A1_c_267_n 0.0388417f $X=2.43 $Y=1.505 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_103_p N_A1_c_267_n 0.00268802f $X=2.575 $Y=0.73 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_78_n N_A1_c_268_n 0.00310267f $X=2.43 $Y=1.505 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_94_p N_VPWR_M1007_d 0.00591219f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_125_p N_VPWR_M1007_d 0.00293726f $X=1.2 $Y=1.895 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_83_n N_VPWR_M1007_d 0.00415349f $X=1.285 $Y=2 $X2=0 $Y2=0
cc_110 N_A_79_21#_M1001_g N_VPWR_c_332_n 0.00843941f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_79_21#_M1007_g N_VPWR_c_332_n 5.82214e-19 $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_79_21#_M1007_g N_VPWR_c_333_n 0.00812103f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_94_p N_VPWR_c_333_n 0.00224709f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_82_n N_VPWR_c_333_n 0.00652529f $X=1.975 $Y=2 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_83_n N_VPWR_c_333_n 0.0141627f $X=1.285 $Y=2 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_84_n N_VPWR_c_333_n 0.00608606f $X=2.1 $Y=2.105 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_82_n N_VPWR_c_335_n 0.0116969f $X=1.975 $Y=2 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_84_n N_VPWR_c_335_n 0.0172111f $X=2.1 $Y=2.105 $X2=0 $Y2=0
cc_119 N_A_79_21#_M1001_g N_VPWR_c_337_n 0.00348405f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_79_21#_M1007_g N_VPWR_c_337_n 0.00550269f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_79_21#_M1006_s N_VPWR_c_330_n 0.00387172f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_122 N_A_79_21#_M1001_g N_VPWR_c_330_n 0.00417296f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_M1007_g N_VPWR_c_330_n 0.0112454f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_82_n N_VPWR_c_330_n 0.0179781f $X=1.975 $Y=2 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_83_n N_VPWR_c_330_n 8.79686e-19 $X=1.285 $Y=2 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_84_n N_VPWR_c_330_n 0.00953699f $X=2.1 $Y=2.105 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_144_p N_X_M1001_s 0.00221225f $X=0.9 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_79_21#_M1001_g N_X_c_397_n 0.0156431f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_79_21#_M1009_g N_X_c_398_n 0.0154706f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_130 N_A_79_21#_M1010_g N_X_c_398_n 0.00241342f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_76_n N_X_c_398_n 0.0022528f $X=0.825 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_81_n N_X_c_398_n 0.0167974f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_79_21#_M1009_g N_X_c_402_n 0.0101786f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_79_21#_M1010_g N_X_c_402_n 0.00443252f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_135 N_A_79_21#_M1007_g N_X_c_404_n 0.00244371f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_76_n N_X_c_404_n 3.6121e-19 $X=0.825 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_144_p N_X_c_404_n 0.0166855f $X=0.9 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_125_p N_X_c_404_n 0.00332662f $X=1.2 $Y=1.895 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_83_n N_X_c_404_n 0.00683223f $X=1.285 $Y=2 $X2=0 $Y2=0
cc_140 N_A_79_21#_M1007_g N_X_c_409_n 0.0103519f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_83_n N_X_c_409_n 0.00574271f $X=1.285 $Y=2 $X2=0 $Y2=0
cc_142 N_A_79_21#_M1009_g X 0.0265638f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_81_n X 0.0297165f $X=0.735 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_78_n N_A_485_297#_M1006_d 2.62576e-19 $X=2.43 $Y=1.505
+ $X2=-0.19 $Y2=-0.24
cc_145 N_A_79_21#_c_102_p N_A_485_297#_M1006_d 0.00215305f $X=2.43 $Y=1.59
+ $X2=-0.19 $Y2=-0.24
cc_146 N_A_79_21#_c_102_p N_A_485_297#_c_435_n 0.00485487f $X=2.43 $Y=1.59 $X2=0
+ $Y2=0
cc_147 N_A_79_21#_M1009_g N_VGND_c_461_n 0.00322099f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A_79_21#_M1010_g N_VGND_c_462_n 0.00322196f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_94_p N_VGND_c_462_n 0.00115409f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_79_21#_M1009_g N_VGND_c_466_n 0.00425835f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_79_21#_M1010_g N_VGND_c_466_n 0.00549917f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_103_p N_VGND_c_469_n 0.00608897f $X=2.575 $Y=0.73 $X2=0
+ $Y2=0
cc_153 N_A_79_21#_M1008_d N_VGND_c_471_n 0.00431979f $X=2.425 $Y=0.235 $X2=0
+ $Y2=0
cc_154 N_A_79_21#_M1009_g N_VGND_c_471_n 0.00672289f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A_79_21#_M1010_g N_VGND_c_471_n 0.0109846f $X=0.9 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_103_p N_VGND_c_471_n 0.0108281f $X=2.575 $Y=0.73 $X2=0 $Y2=0
cc_157 B1_N N_A_297_93#_c_210_n 2.6446e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_158 N_B1_N_c_175_n N_A_297_93#_c_210_n 0.00909219f $X=1.44 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_B1_N_c_176_n N_A_297_93#_c_211_n 0.00407921f $X=1.44 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_B1_N_M1002_g N_A_297_93#_c_216_n 0.00566324f $X=1.41 $Y=1.695 $X2=0
+ $Y2=0
cc_161 B1_N N_A_297_93#_c_212_n 0.00362896f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_162 N_B1_N_c_175_n N_A_297_93#_c_212_n 0.00158354f $X=1.44 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_B1_N_c_176_n N_A_297_93#_c_212_n 0.00303643f $X=1.44 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_B1_N_M1002_g N_A_297_93#_c_217_n 0.00263532f $X=1.41 $Y=1.695 $X2=0
+ $Y2=0
cc_165 B1_N N_A_297_93#_c_217_n 0.00284653f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_166 N_B1_N_c_175_n N_A_297_93#_c_217_n 0.00148463f $X=1.44 $Y=1.16 $X2=0
+ $Y2=0
cc_167 B1_N N_A_297_93#_c_213_n 0.0274459f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_168 N_B1_N_c_175_n N_A_297_93#_c_213_n 0.00281016f $X=1.44 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_B1_N_M1002_g N_VPWR_c_333_n 2.15973e-19 $X=1.41 $Y=1.695 $X2=0 $Y2=0
cc_170 N_B1_N_M1002_g N_VPWR_c_335_n 4.03486e-19 $X=1.41 $Y=1.695 $X2=0 $Y2=0
cc_171 B1_N N_VGND_c_462_n 0.012858f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_172 N_B1_N_c_176_n N_VGND_c_462_n 0.00943349f $X=1.44 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B1_N_c_176_n N_VGND_c_463_n 0.0034467f $X=1.44 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B1_N_c_176_n N_VGND_c_468_n 0.00487013f $X=1.44 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B1_N_c_176_n N_VGND_c_471_n 0.00512902f $X=1.44 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_297_93#_M1006_g N_A1_M1005_g 0.0292483f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_297_93#_c_210_n N_A1_c_266_n 0.0202376f $X=2.35 $Y=0.99 $X2=0 $Y2=0
cc_178 N_A_297_93#_c_210_n N_A1_c_267_n 3.15782e-19 $X=2.35 $Y=0.99 $X2=0 $Y2=0
cc_179 N_A_297_93#_M1006_g N_A1_c_267_n 4.80424e-19 $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_297_93#_c_210_n N_A1_c_268_n 0.0209795f $X=2.35 $Y=0.99 $X2=0 $Y2=0
cc_181 N_A_297_93#_M1006_g N_VPWR_c_335_n 0.00541359f $X=2.35 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_297_93#_M1006_g N_VPWR_c_330_n 0.0111045f $X=2.35 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_297_93#_M1006_g N_A_485_297#_c_435_n 0.00745188f $X=2.35 $Y=1.985
+ $X2=0 $Y2=0
cc_184 N_A_297_93#_c_211_n N_VGND_c_462_n 0.00137223f $X=1.78 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_297_93#_c_212_n N_VGND_c_462_n 0.00998923f $X=1.78 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_297_93#_c_210_n N_VGND_c_463_n 0.0175576f $X=2.35 $Y=0.99 $X2=0 $Y2=0
cc_187 N_A_297_93#_c_213_n N_VGND_c_463_n 0.00672869f $X=2.09 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A_297_93#_c_212_n N_VGND_c_468_n 0.00649604f $X=1.78 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_297_93#_c_210_n N_VGND_c_469_n 0.00381042f $X=2.35 $Y=0.99 $X2=0
+ $Y2=0
cc_190 N_A_297_93#_c_210_n N_VGND_c_471_n 0.00549693f $X=2.35 $Y=0.99 $X2=0
+ $Y2=0
cc_191 N_A_297_93#_c_212_n N_VGND_c_471_n 0.0113942f $X=1.78 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_M1005_g N_A2_M1004_g 0.045132f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A1_c_266_n A2 2.30431e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A1_c_267_n A2 0.0398007f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A1_c_266_n N_A2_c_305_n 0.0378105f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A1_c_267_n N_A2_c_305_n 0.00455047f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A1_c_268_n N_A2_c_306_n 0.0378105f $X=2.77 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_267_n N_VPWR_M1005_d 0.00217416f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A1_M1005_g N_VPWR_c_334_n 0.00268723f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A1_M1005_g N_VPWR_c_335_n 0.00421138f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A1_M1005_g N_VPWR_c_330_n 0.00573126f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A1_M1005_g N_A_485_297#_c_437_n 0.00864432f $X=2.77 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A1_c_267_n N_A_485_297#_c_437_n 0.017153f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A1_M1005_g N_A_485_297#_c_435_n 0.00703925f $X=2.77 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A1_c_266_n N_A_485_297#_c_435_n 7.64552e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A1_c_267_n N_A_485_297#_c_435_n 0.00192944f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A1_M1005_g N_A_485_297#_c_432_n 5.37795e-19 $X=2.77 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A1_c_268_n N_VGND_c_463_n 0.00206618f $X=2.77 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_268_n N_VGND_c_465_n 0.00368972f $X=2.77 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_268_n N_VGND_c_469_n 0.00585385f $X=2.77 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A1_c_268_n N_VGND_c_471_n 0.0108513f $X=2.77 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A2_M1004_g N_VPWR_c_334_n 0.00268723f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A2_M1004_g N_VPWR_c_338_n 0.00421138f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A2_M1004_g N_VPWR_c_330_n 0.00667694f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_215 A2 N_A_485_297#_M1004_d 0.00379222f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A2_M1004_g N_A_485_297#_c_437_n 0.0120004f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A2_M1004_g N_A_485_297#_c_435_n 5.37795e-19 $X=3.19 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A2_M1004_g N_A_485_297#_c_432_n 0.00800369f $X=3.19 $Y=1.985 $X2=0
+ $Y2=0
cc_219 A2 N_A_485_297#_c_432_n 0.0169621f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_220 N_A2_c_305_n N_A_485_297#_c_432_n 8.30139e-19 $X=3.355 $Y=1.16 $X2=0
+ $Y2=0
cc_221 A2 N_VGND_c_465_n 0.0230961f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A2_c_305_n N_VGND_c_465_n 0.00506784f $X=3.355 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A2_c_306_n N_VGND_c_465_n 0.0239842f $X=3.302 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_306_n N_VGND_c_469_n 0.0046653f $X=3.302 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A2_c_306_n N_VGND_c_471_n 0.00783311f $X=3.302 $Y=0.995 $X2=0 $Y2=0
cc_226 N_VPWR_c_330_n N_X_M1001_s 0.00250132f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_c_332_n N_X_c_397_n 0.00143691f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_228 N_VPWR_c_337_n N_X_c_397_n 0.0020257f $X=1.04 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_330_n N_X_c_397_n 0.00413047f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_333_n N_X_c_409_n 0.0104876f $X=1.205 $Y=2.36 $X2=0 $Y2=0
cc_231 N_VPWR_c_337_n N_X_c_409_n 0.0122547f $X=1.04 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_330_n N_X_c_409_n 0.00938767f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_M1001_d X 0.0162128f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_234 N_VPWR_M1001_d N_X_c_421_n 0.0106914f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_235 N_VPWR_c_332_n N_X_c_421_n 0.0113976f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_236 N_VPWR_c_330_n N_X_c_421_n 0.00122621f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_330_n N_A_485_297#_M1006_d 0.00215201f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_238 N_VPWR_c_330_n N_A_485_297#_M1004_d 0.00209319f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_239 N_VPWR_M1005_d N_A_485_297#_c_437_n 0.0034719f $X=2.845 $Y=1.485 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_334_n N_A_485_297#_c_437_n 0.0121469f $X=2.98 $Y=2.36 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_335_n N_A_485_297#_c_437_n 0.00207171f $X=2.895 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_338_n N_A_485_297#_c_437_n 0.00207171f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_330_n N_A_485_297#_c_437_n 0.008494f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_335_n N_A_485_297#_c_435_n 0.0188044f $X=2.895 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_330_n N_A_485_297#_c_435_n 0.0121916f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_338_n N_A_485_297#_c_432_n 0.0209097f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_330_n N_A_485_297#_c_432_n 0.0123965f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_248 N_X_c_398_n N_VGND_M1009_s 0.0107097f $X=0.685 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_249 X N_VGND_M1009_s 5.52941e-19 $X=0.15 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_250 N_X_c_398_n N_VGND_c_461_n 0.0146773f $X=0.685 $Y=0.715 $X2=0 $Y2=0
cc_251 N_X_c_398_n N_VGND_c_466_n 0.00212719f $X=0.685 $Y=0.715 $X2=0 $Y2=0
cc_252 N_X_c_402_n N_VGND_c_466_n 0.0133207f $X=0.685 $Y=0.4 $X2=0 $Y2=0
cc_253 N_X_M1009_d N_VGND_c_471_n 0.00227848f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_254 N_X_c_398_n N_VGND_c_471_n 0.00479164f $X=0.685 $Y=0.715 $X2=0 $Y2=0
cc_255 N_X_c_402_n N_VGND_c_471_n 0.0116884f $X=0.685 $Y=0.4 $X2=0 $Y2=0
cc_256 N_VGND_c_471_n A_581_47# 0.00897657f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__and3b_4.spice
* Created: Tue Sep  1 18:57:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and3b_4.pex.spice"
.subckt sky130_fd_sc_hd__and3b_4  VNB VPB B C A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1010 A_152_47# N_A_98_199#_M1010_g N_A_56_297#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.121875 AS=0.19825 PD=1.025 PS=1.91 NRD=24.456 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1001 A_257_47# N_B_M1001_g A_152_47# VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.121875 PD=0.88 PS=1.025 NRD=11.076 NRS=24.456 M=1 R=4.33333 SA=75000.8
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_C_M1011_g A_257_47# VNB NSHORT L=0.15 W=0.65 AD=0.138125
+ AS=0.07475 PD=1.075 PS=0.88 NRD=25.836 NRS=11.076 M=1 R=4.33333 SA=75001.1
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1011_d N_A_56_297#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.138125 AS=0.091 PD=1.075 PS=0.93 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_56_297#_M1005_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1005_d N_A_56_297#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_56_297#_M1014_g N_X_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.131671 AS=0.091 PD=1.2271 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_98_199#_M1002_d N_A_N_M1002_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1491 AS=0.0850794 PD=1.55 PS=0.792897 NRD=19.992 NRS=42.156 M=1 R=2.8
+ SA=75003.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_98_199#_M1007_g N_A_56_297#_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.1875 AS=0.33 PD=1.375 PS=2.66 NRD=12.7853 NRS=8.8453 M=1 R=6.66667
+ SA=75000.3 SB=75003.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_56_297#_M1000_d N_B_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.1875 PD=1.3 PS=1.375 NRD=3.9203 NRS=5.8903 M=1 R=6.66667
+ SA=75000.8 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_A_56_297#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1775 AS=0.15 PD=1.355 PS=1.3 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_56_297#_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.1775 PD=1.29 PS=1.355 NRD=1.9503 NRS=7.8603 M=1 R=6.66667
+ SA=75001.7 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1003_d N_A_56_297#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.135 PD=1.29 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1013_d N_A_56_297#_M1013_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.6
+ SB=75000.9 A=0.15 P=2.3 MULT=1
MM1015 N_X_M1013_d N_A_56_297#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.222887 PD=1.28 PS=1.91549 NRD=0 NRS=0 M=1 R=6.66667 SA=75003
+ SB=75000.4 A=0.15 P=2.3 MULT=1
MM1009 N_A_98_199#_M1009_d N_A_N_M1009_g N_VPWR_M1015_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0936127 PD=1.41 PS=0.804507 NRD=0 NRS=78.7409 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__and3b_4.pxi.spice"
*
.ends
*
*

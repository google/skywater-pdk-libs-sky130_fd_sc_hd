# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o221ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965000 1.075000 6.295000 1.445000 ;
        RECT 5.965000 1.445000 8.420000 1.615000 ;
        RECT 8.155000 1.075000 9.575000 1.275000 ;
        RECT 8.155000 1.275000 8.420000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 7.885000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.360000 1.075000 4.505000 1.275000 ;
        RECT 4.335000 1.275000 4.505000 1.495000 ;
        RECT 4.335000 1.495000 5.795000 1.665000 ;
        RECT 5.465000 1.075000 5.795000 1.495000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 0.995000 5.285000 1.325000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.750000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 2.125000 0.865000 ;
        RECT 0.575000 1.445000 4.165000 1.615000 ;
        RECT 0.575000 1.615000 0.825000 2.465000 ;
        RECT 1.415000 1.615000 2.125000 1.955000 ;
        RECT 1.415000 1.955000 1.665000 2.465000 ;
        RECT 1.920000 0.865000 2.125000 1.445000 ;
        RECT 3.995000 1.615000 4.165000 1.835000 ;
        RECT 3.995000 1.835000 7.725000 1.955000 ;
        RECT 3.995000 1.955000 6.885000 2.005000 ;
        RECT 3.995000 2.005000 4.285000 2.125000 ;
        RECT 4.875000 2.005000 5.085000 2.125000 ;
        RECT 5.965000 1.785000 7.725000 1.835000 ;
        RECT 6.675000 2.005000 6.885000 2.125000 ;
        RECT 7.475000 1.955000 7.725000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 6.255000  0.085000 6.425000 0.555000 ;
        RECT 7.095000  0.085000 7.265000 0.555000 ;
        RECT 7.935000  0.085000 8.105000 0.555000 ;
        RECT 8.775000  0.085000 8.945000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.155000 1.485000 0.405000 2.635000 ;
        RECT 0.995000 1.825000 1.245000 2.635000 ;
        RECT 1.835000 2.125000 2.605000 2.635000 ;
        RECT 3.195000 2.125000 3.445000 2.635000 ;
        RECT 5.755000 2.175000 6.005000 2.635000 ;
        RECT 8.315000 2.125000 8.565000 2.635000 ;
        RECT 9.155000 1.445000 9.405000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.255000 5.585000 0.475000 ;
      RECT 0.115000 0.475000 0.365000 0.895000 ;
      RECT 2.315000 0.645000 6.085000 0.735000 ;
      RECT 2.315000 0.735000 9.445000 0.820000 ;
      RECT 2.775000 1.785000 3.825000 1.955000 ;
      RECT 2.775000 1.955000 3.025000 2.465000 ;
      RECT 3.615000 1.955000 3.825000 2.295000 ;
      RECT 3.615000 2.295000 5.585000 2.465000 ;
      RECT 4.455000 2.175000 4.705000 2.295000 ;
      RECT 5.255000 2.175000 5.585000 2.295000 ;
      RECT 5.465000 0.820000 9.445000 0.905000 ;
      RECT 5.755000 0.255000 6.085000 0.645000 ;
      RECT 6.175000 2.175000 6.505000 2.295000 ;
      RECT 6.175000 2.295000 8.145000 2.465000 ;
      RECT 6.595000 0.255000 6.925000 0.725000 ;
      RECT 6.595000 0.725000 7.765000 0.735000 ;
      RECT 7.055000 2.125000 7.305000 2.295000 ;
      RECT 7.435000 0.255000 7.765000 0.725000 ;
      RECT 7.895000 1.785000 8.985000 1.955000 ;
      RECT 7.895000 1.955000 8.145000 2.295000 ;
      RECT 8.275000 0.255000 8.605000 0.725000 ;
      RECT 8.275000 0.725000 9.445000 0.735000 ;
      RECT 8.735000 1.445000 8.985000 1.785000 ;
      RECT 8.735000 1.955000 8.985000 2.465000 ;
      RECT 9.115000 0.255000 9.445000 0.725000 ;
  END
END sky130_fd_sc_hd__o221ai_4

* File: sky130_fd_sc_hd__nand4_2.spice
* Created: Thu Aug 27 14:30:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4_2.pex.spice"
.subckt sky130_fd_sc_hd__nand4_2  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_A_27_47#_M1004_d N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1013 N_A_27_47#_M1013_d N_D_M1013_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 N_A_27_47#_M1013_d N_C_M1006_g N_A_277_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1007_d N_C_M1007_g N_A_277_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_471_47#_M1010_d N_B_M1010_g N_A_277_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1014 N_A_471_47#_M1014_d N_B_M1014_g N_A_277_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_A_471_47#_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1009_d N_A_M1015_g N_A_471_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.234 PD=0.92 PS=2.02 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75001.5
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_D_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75003.8
+ A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75003.4
+ A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75003 A=0.15
+ P=2.3 MULT=1
MM1011 N_Y_M1001_d N_C_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.215 PD=1.27 PS=1.43 NRD=0 NRS=14.7553 M=1 R=6.66667 SA=75001.4 SB=75002.6
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1011_s N_B_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.215
+ AS=0.135 PD=1.43 PS=1.27 NRD=14.7553 NRS=0 M=1 R=6.66667 SA=75002 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.335
+ AS=0.135 PD=1.67 PS=1.27 NRD=42.3353 NRS=0 M=1 R=6.66667 SA=75002.4 SB=75001.6
+ A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.335 PD=1.27 PS=1.67 NRD=0 NRS=34.4553 M=1 R=6.66667 SA=75003.3 SB=75000.8
+ A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1000_d N_A_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.42 PD=1.27 PS=2.84 NRD=0 NRS=14.775 M=1 R=6.66667 SA=75003.7 SB=75000.3
+ A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__nand4_2.pxi.spice"
*
.ends
*
*

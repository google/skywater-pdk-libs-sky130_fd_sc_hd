* File: sky130_fd_sc_hd__nand2_4.pxi.spice
* Created: Thu Aug 27 14:28:50 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2_4%B N_B_c_61_n N_B_M1004_g N_B_M1001_g N_B_c_62_n
+ N_B_M1005_g N_B_M1002_g N_B_c_63_n N_B_M1007_g N_B_M1008_g N_B_c_64_n
+ N_B_M1015_g N_B_M1013_g B B B B N_B_c_66_n PM_SKY130_FD_SC_HD__NAND2_4%B
x_PM_SKY130_FD_SC_HD__NAND2_4%A N_A_c_151_n N_A_M1006_g N_A_M1000_g N_A_c_152_n
+ N_A_M1009_g N_A_M1003_g N_A_c_153_n N_A_M1011_g N_A_M1010_g N_A_c_154_n
+ N_A_M1012_g N_A_M1014_g A A A N_A_c_156_n PM_SKY130_FD_SC_HD__NAND2_4%A
x_PM_SKY130_FD_SC_HD__NAND2_4%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1013_s
+ N_VPWR_M1003_s N_VPWR_M1014_s N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_226_n
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n
+ N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n
+ N_VPWR_c_237_n VPWR N_VPWR_c_238_n N_VPWR_c_223_n
+ PM_SKY130_FD_SC_HD__NAND2_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND2_4%Y N_Y_M1006_d N_Y_M1011_d N_Y_M1001_d N_Y_M1008_d
+ N_Y_M1000_d N_Y_M1010_d N_Y_c_291_n N_Y_c_295_n N_Y_c_298_n N_Y_c_302_n
+ N_Y_c_305_n N_Y_c_316_n N_Y_c_288_n N_Y_c_308_n N_Y_c_323_n N_Y_c_328_n
+ N_Y_c_289_n N_Y_c_336_n N_Y_c_340_n N_Y_c_311_n Y
+ PM_SKY130_FD_SC_HD__NAND2_4%Y
x_PM_SKY130_FD_SC_HD__NAND2_4%A_27_47# N_A_27_47#_M1004_d N_A_27_47#_M1005_d
+ N_A_27_47#_M1015_d N_A_27_47#_M1009_s N_A_27_47#_M1012_s N_A_27_47#_c_375_n
+ N_A_27_47#_c_376_n N_A_27_47#_c_377_n N_A_27_47#_c_392_n N_A_27_47#_c_378_n
+ N_A_27_47#_c_400_n N_A_27_47#_c_379_n N_A_27_47#_c_407_n N_A_27_47#_c_380_n
+ N_A_27_47#_c_381_n N_A_27_47#_c_382_n PM_SKY130_FD_SC_HD__NAND2_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND2_4%VGND N_VGND_M1004_s N_VGND_M1007_s N_VGND_c_450_n
+ N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n
+ VGND N_VGND_c_456_n N_VGND_c_457_n PM_SKY130_FD_SC_HD__NAND2_4%VGND
cc_1 VNB N_B_c_61_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B_c_62_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_B_c_63_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_B_c_64_n 0.016004f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB B 0.00932659f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_6 VNB N_B_c_66_n 0.0857113f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_7 VNB N_A_c_151_n 0.01577f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_A_c_152_n 0.0159731f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_9 VNB N_A_c_153_n 0.0160006f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_10 VNB N_A_c_154_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_11 VNB A 0.0255779f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_12 VNB N_A_c_156_n 0.0688989f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_13 VNB N_VPWR_c_223_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_288_n 0.00103672f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_15 VNB N_Y_c_289_n 0.00328583f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_16 VNB N_A_27_47#_c_375_n 0.0182049f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_17 VNB N_A_27_47#_c_376_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_18 VNB N_A_27_47#_c_377_n 0.0100781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_378_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_20 VNB N_A_27_47#_c_379_n 0.00290363f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_A_27_47#_c_380_n 0.00914706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_381_n 0.0180561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_382_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_24 VNB N_VGND_c_450_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_25 VNB N_VGND_c_451_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_26 VNB N_VGND_c_452_n 0.0171658f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_27 VNB N_VGND_c_453_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_28 VNB N_VGND_c_454_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_29 VNB N_VGND_c_455_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_30 VNB N_VGND_c_456_n 0.0626673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_457_n 0.229746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_B_M1001_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB N_B_M1002_g 0.0185065f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_34 VPB N_B_M1008_g 0.0185018f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_35 VPB N_B_M1013_g 0.0187899f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_36 VPB B 7.73822e-19 $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_37 VPB N_B_c_66_n 0.019304f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_38 VPB N_A_M1000_g 0.0172006f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB N_A_M1003_g 0.0184594f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_40 VPB N_A_M1010_g 0.0184995f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_41 VPB N_A_M1014_g 0.0259842f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_42 VPB A 0.0163038f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_43 VPB N_A_c_156_n 0.0107017f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_44 VPB N_VPWR_c_224_n 0.00994749f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_45 VPB N_VPWR_c_225_n 0.0423299f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_46 VPB N_VPWR_c_226_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_47 VPB N_VPWR_c_227_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_228_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_49 VPB N_VPWR_c_229_n 0.0294355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_230_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_51 VPB N_VPWR_c_231_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_232_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_53 VPB N_VPWR_c_233_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_54 VPB N_VPWR_c_234_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_55 VPB N_VPWR_c_235_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_56 VPB N_VPWR_c_236_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_237_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_58 VPB N_VPWR_c_238_n 0.0134401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_223_n 0.0537104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_Y_c_289_n 0.00347809f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_61 N_B_c_64_n N_A_c_151_n 0.0187942f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_62 N_B_M1013_g N_A_M1000_g 0.0187942f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_63 B N_A_c_156_n 2.09391e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_64 N_B_c_66_n N_A_c_156_n 0.0187942f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_65 N_B_M1001_g N_VPWR_c_225_n 0.00321527f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_66 B N_VPWR_c_225_n 0.0187309f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_67 N_B_c_66_n N_VPWR_c_225_n 0.0054329f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B_M1002_g N_VPWR_c_226_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_69 N_B_M1008_g N_VPWR_c_226_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_70 N_B_M1013_g N_VPWR_c_227_n 0.00146448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_71 N_B_M1001_g N_VPWR_c_230_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_72 N_B_M1002_g N_VPWR_c_230_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 N_B_M1008_g N_VPWR_c_232_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_74 N_B_M1013_g N_VPWR_c_232_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_75 N_B_M1001_g N_VPWR_c_223_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_76 N_B_M1002_g N_VPWR_c_223_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_77 N_B_M1008_g N_VPWR_c_223_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B_M1013_g N_VPWR_c_223_n 0.00952874f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B_M1001_g N_Y_c_291_n 0.00229676f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_80 N_B_M1002_g N_Y_c_291_n 8.84614e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_81 B N_Y_c_291_n 0.0213676f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_82 N_B_c_66_n N_Y_c_291_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B_M1001_g N_Y_c_295_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_84 N_B_M1002_g N_Y_c_295_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_85 N_B_M1008_g N_Y_c_295_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_86 N_B_M1002_g N_Y_c_298_n 0.0107189f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_87 N_B_M1008_g N_Y_c_298_n 0.0107189f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_88 B N_Y_c_298_n 0.0320704f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_89 N_B_c_66_n N_Y_c_298_n 0.00201785f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_M1002_g N_Y_c_302_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_91 N_B_M1008_g N_Y_c_302_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B_M1013_g N_Y_c_302_n 0.00975139f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_93 N_B_M1013_g N_Y_c_305_n 0.0116765f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_94 B N_Y_c_305_n 0.00310934f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B_c_64_n N_Y_c_288_n 9.48164e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B_M1013_g N_Y_c_308_n 6.1949e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_97 B N_Y_c_289_n 0.0207728f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B_c_66_n N_Y_c_289_n 0.00695919f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B_M1008_g N_Y_c_311_n 8.84614e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B_M1013_g N_Y_c_311_n 8.84614e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_101 B N_Y_c_311_n 0.0213676f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_102 N_B_c_66_n N_Y_c_311_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_c_61_n N_A_27_47#_c_375_n 0.00620543f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B_c_62_n N_A_27_47#_c_375_n 5.19198e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_c_61_n N_A_27_47#_c_376_n 0.00890471f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B_c_62_n N_A_27_47#_c_376_n 0.00890471f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_107 B N_A_27_47#_c_376_n 0.0368812f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B_c_66_n N_A_27_47#_c_376_n 0.00222429f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B_c_61_n N_A_27_47#_c_377_n 0.00132416f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_110 B N_A_27_47#_c_377_n 0.0258342f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B_c_66_n N_A_27_47#_c_377_n 0.00729406f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B_c_61_n N_A_27_47#_c_392_n 5.19281e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_62_n N_A_27_47#_c_392_n 0.00620543f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B_c_63_n N_A_27_47#_c_392_n 0.00620543f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_64_n N_A_27_47#_c_392_n 5.19281e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B_c_63_n N_A_27_47#_c_378_n 0.0088553f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_64_n N_A_27_47#_c_378_n 0.00949606f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_118 B N_A_27_47#_c_378_n 0.0337462f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B_c_66_n N_A_27_47#_c_378_n 0.00222429f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_c_64_n N_A_27_47#_c_400_n 0.00244813f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B_c_63_n N_A_27_47#_c_379_n 4.58193e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_64_n N_A_27_47#_c_379_n 0.00531461f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_62_n N_A_27_47#_c_382_n 0.00116017f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_63_n N_A_27_47#_c_382_n 0.00116017f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_125 B N_A_27_47#_c_382_n 0.0269421f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B_c_66_n N_A_27_47#_c_382_n 0.00230339f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B_c_61_n N_VGND_c_450_n 0.00268723f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B_c_62_n N_VGND_c_450_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B_c_63_n N_VGND_c_451_n 0.00146448f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B_c_64_n N_VGND_c_451_n 0.00268723f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B_c_61_n N_VGND_c_452_n 0.00422241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B_c_62_n N_VGND_c_454_n 0.00422241f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B_c_63_n N_VGND_c_454_n 0.00422241f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B_c_64_n N_VGND_c_456_n 0.00420723f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B_c_61_n N_VGND_c_457_n 0.00665076f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B_c_62_n N_VGND_c_457_n 0.00569656f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B_c_63_n N_VGND_c_457_n 0.00569656f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B_c_64_n N_VGND_c_457_n 0.00573284f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_VPWR_c_227_n 0.00146448f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1003_g N_VPWR_c_228_n 0.00146448f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1010_g N_VPWR_c_228_n 0.00146448f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1014_g N_VPWR_c_229_n 0.00321269f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_143 A N_VPWR_c_229_n 0.00950731f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_VPWR_c_234_n 0.00541359f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1003_g N_VPWR_c_234_n 0.00541359f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1010_g N_VPWR_c_236_n 0.00541359f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1014_g N_VPWR_c_236_n 0.00541359f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1000_g N_VPWR_c_223_n 0.00952874f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1003_g N_VPWR_c_223_n 0.00950154f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1010_g N_VPWR_c_223_n 0.00950154f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1014_g N_VPWR_c_223_n 0.0106288f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1000_g N_Y_c_302_n 6.1949e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_c_151_n N_Y_c_316_n 0.00219421f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_151_n N_Y_c_288_n 0.00358324f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_152_n N_Y_c_288_n 0.00280346f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_156_n N_Y_c_288_n 0.00860058f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_M1000_g N_Y_c_308_n 0.00975139f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_Y_c_308_n 0.00975139f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1010_g N_Y_c_308_n 6.1949e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_c_152_n N_Y_c_323_n 0.0121073f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_153_n N_Y_c_323_n 0.00893253f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_154_n N_Y_c_323_n 0.00275569f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_163 A N_Y_c_323_n 0.0315661f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A_c_156_n N_Y_c_323_n 0.00414123f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_M1003_g N_Y_c_328_n 0.0134371f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_M1010_g N_Y_c_328_n 0.0107189f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_167 A N_Y_c_328_n 0.0258179f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A_c_156_n N_Y_c_328_n 0.00201785f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_M1000_g N_Y_c_289_n 0.0154787f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_M1003_g N_Y_c_289_n 0.00672354f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_171 A N_Y_c_289_n 0.0206172f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A_c_156_n N_Y_c_289_n 0.0198408f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_M1010_g N_Y_c_336_n 8.84614e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_M1014_g N_Y_c_336_n 0.00849147f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_175 A N_Y_c_336_n 0.0213676f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A_c_156_n N_Y_c_336_n 0.00209661f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_M1003_g N_Y_c_340_n 6.1949e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_M1010_g N_Y_c_340_n 0.00975139f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_M1014_g N_Y_c_340_n 0.0145598f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_c_151_n N_A_27_47#_c_407_n 0.0103273f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_152_n N_A_27_47#_c_407_n 0.00866705f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_153_n N_A_27_47#_c_407_n 0.00866705f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_154_n N_A_27_47#_c_407_n 0.0103313f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_184 A N_A_27_47#_c_407_n 0.00376413f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_185 N_A_c_156_n N_A_27_47#_c_407_n 3.01257e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_186 A N_A_27_47#_c_381_n 0.0191425f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A_c_151_n N_VGND_c_456_n 0.00357877f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_152_n N_VGND_c_456_n 0.00357877f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_153_n N_VGND_c_456_n 0.00357877f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_154_n N_VGND_c_456_n 0.00357877f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_151_n N_VGND_c_457_n 0.00525237f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_152_n N_VGND_c_457_n 0.00522516f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_153_n N_VGND_c_457_n 0.00522516f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_154_n N_VGND_c_457_n 0.00635241f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_195 N_VPWR_c_223_n N_Y_M1001_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_223_n N_Y_M1008_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_197 N_VPWR_c_223_n N_Y_M1000_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_223_n N_Y_M1010_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_230_n N_Y_c_295_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_c_223_n N_Y_c_295_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_201 N_VPWR_M1002_s N_Y_c_298_n 0.00311483f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_202 N_VPWR_c_226_n N_Y_c_298_n 0.0126919f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_203 N_VPWR_c_232_n N_Y_c_302_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_c_223_n N_Y_c_302_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_M1013_s N_Y_c_305_n 0.00142612f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_206 N_VPWR_c_227_n N_Y_c_305_n 0.00386873f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_207 N_VPWR_c_234_n N_Y_c_308_n 0.0189039f $X=2.695 $Y=2.72 $X2=0 $Y2=0
cc_208 N_VPWR_c_223_n N_Y_c_308_n 0.0122165f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_209 N_VPWR_M1003_s N_Y_c_328_n 0.00311483f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_210 N_VPWR_c_228_n N_Y_c_328_n 0.0126919f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_211 N_VPWR_M1013_s N_Y_c_289_n 0.00131839f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_212 N_VPWR_c_227_n N_Y_c_289_n 0.00963603f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_213 N_VPWR_c_236_n N_Y_c_340_n 0.0189039f $X=3.535 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_223_n N_Y_c_340_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_c_225_n N_A_27_47#_c_377_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_216 N_Y_c_323_n N_A_27_47#_M1009_s 0.00337959f $X=3.2 $Y=0.72 $X2=0 $Y2=0
cc_217 N_Y_c_305_n N_A_27_47#_c_378_n 0.00108863f $X=1.91 $Y=1.58 $X2=0 $Y2=0
cc_218 N_Y_c_305_n N_A_27_47#_c_379_n 0.00353053f $X=1.91 $Y=1.58 $X2=0 $Y2=0
cc_219 N_Y_c_288_n N_A_27_47#_c_379_n 0.00446267f $X=2.32 $Y=1.075 $X2=0 $Y2=0
cc_220 N_Y_c_289_n N_A_27_47#_c_379_n 0.010625f $X=2.525 $Y=1.58 $X2=0 $Y2=0
cc_221 N_Y_M1006_d N_A_27_47#_c_407_n 0.00304479f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_222 N_Y_M1011_d N_A_27_47#_c_407_n 0.00304849f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_223 N_Y_c_316_n N_A_27_47#_c_407_n 0.0143215f $X=2.32 $Y=0.805 $X2=0 $Y2=0
cc_224 N_Y_c_323_n N_A_27_47#_c_407_n 0.0433054f $X=3.2 $Y=0.72 $X2=0 $Y2=0
cc_225 N_Y_c_289_n N_A_27_47#_c_407_n 0.0040954f $X=2.525 $Y=1.58 $X2=0 $Y2=0
cc_226 N_Y_M1006_d N_VGND_c_457_n 0.00216833f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_227 N_Y_M1011_d N_VGND_c_457_n 0.00216833f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_376_n N_VGND_M1004_s 0.00162148f $X=0.935 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_229 N_A_27_47#_c_378_n N_VGND_M1007_s 0.00162148f $X=1.775 $Y=0.81 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_376_n N_VGND_c_450_n 0.0122675f $X=0.935 $Y=0.81 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_378_n N_VGND_c_451_n 0.0122675f $X=1.775 $Y=0.81 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_375_n N_VGND_c_452_n 0.0213324f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_376_n N_VGND_c_452_n 0.00203746f $X=0.935 $Y=0.81 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_376_n N_VGND_c_454_n 0.00203746f $X=0.935 $Y=0.81 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_392_n N_VGND_c_454_n 0.0188551f $X=1.1 $Y=0.38 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_378_n N_VGND_c_454_n 0.00203746f $X=1.775 $Y=0.81 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_378_n N_VGND_c_456_n 0.00203746f $X=1.775 $Y=0.81 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_400_n N_VGND_c_456_n 0.0152108f $X=1.9 $Y=0.465 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_407_n N_VGND_c_456_n 0.0830015f $X=3.535 $Y=0.36 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_380_n N_VGND_c_456_n 0.0172955f $X=3.66 $Y=0.465 $X2=0 $Y2=0
cc_241 N_A_27_47#_M1004_d N_VGND_c_457_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1005_d N_VGND_c_457_n 0.00215201f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_M1015_d N_VGND_c_457_n 0.00215206f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1009_s N_VGND_c_457_n 0.00215227f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_M1012_s N_VGND_c_457_n 0.00209324f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_375_n N_VGND_c_457_n 0.0126042f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_376_n N_VGND_c_457_n 0.00845923f $X=0.935 $Y=0.81 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_392_n N_VGND_c_457_n 0.0122069f $X=1.1 $Y=0.38 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_378_n N_VGND_c_457_n 0.00845923f $X=1.775 $Y=0.81 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_400_n N_VGND_c_457_n 0.00940698f $X=1.9 $Y=0.465 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_407_n N_VGND_c_457_n 0.0534749f $X=3.535 $Y=0.36 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_380_n N_VGND_c_457_n 0.00960883f $X=3.66 $Y=0.465 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__inv_12.pxi.spice
* Created: Thu Aug 27 14:22:19 2020
* 
x_PM_SKY130_FD_SC_HD__INV_12%A N_A_c_88_n N_A_M1001_g N_A_M1000_g N_A_c_89_n
+ N_A_M1002_g N_A_M1003_g N_A_c_90_n N_A_M1004_g N_A_M1006_g N_A_c_91_n
+ N_A_M1005_g N_A_M1007_g N_A_c_92_n N_A_M1008_g N_A_M1012_g N_A_c_93_n
+ N_A_M1009_g N_A_M1015_g N_A_c_94_n N_A_M1010_g N_A_M1016_g N_A_c_95_n
+ N_A_M1011_g N_A_M1017_g N_A_c_96_n N_A_M1013_g N_A_M1018_g N_A_c_97_n
+ N_A_M1014_g N_A_M1019_g N_A_c_98_n N_A_M1020_g N_A_M1021_g N_A_c_99_n
+ N_A_M1022_g N_A_M1023_g A A A A A A A A A A N_A_c_100_n
+ PM_SKY130_FD_SC_HD__INV_12%A
x_PM_SKY130_FD_SC_HD__INV_12%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1007_s
+ N_VPWR_M1015_s N_VPWR_M1017_s N_VPWR_M1019_s N_VPWR_M1023_s N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ N_VPWR_c_341_n N_VPWR_c_342_n VPWR N_VPWR_c_343_n N_VPWR_c_344_n
+ N_VPWR_c_324_n PM_SKY130_FD_SC_HD__INV_12%VPWR
x_PM_SKY130_FD_SC_HD__INV_12%Y N_Y_M1001_d N_Y_M1004_d N_Y_M1008_d N_Y_M1010_d
+ N_Y_M1013_d N_Y_M1020_d N_Y_M1000_d N_Y_M1006_d N_Y_M1012_d N_Y_M1016_d
+ N_Y_M1018_d N_Y_M1021_d N_Y_c_435_n N_Y_c_438_n N_Y_c_417_n N_Y_c_418_n
+ N_Y_c_448_n N_Y_c_431_n N_Y_c_455_n N_Y_c_459_n N_Y_c_419_n N_Y_c_467_n
+ N_Y_c_471_n N_Y_c_475_n N_Y_c_420_n N_Y_c_483_n N_Y_c_487_n N_Y_c_491_n
+ N_Y_c_421_n N_Y_c_499_n N_Y_c_503_n N_Y_c_507_n N_Y_c_422_n N_Y_c_515_n
+ N_Y_c_519_n N_Y_c_522_n N_Y_c_423_n N_Y_c_432_n N_Y_c_424_n N_Y_c_533_n
+ N_Y_c_425_n N_Y_c_541_n N_Y_c_426_n N_Y_c_549_n N_Y_c_427_n N_Y_c_557_n
+ N_Y_c_428_n N_Y_c_565_n Y Y PM_SKY130_FD_SC_HD__INV_12%Y
x_PM_SKY130_FD_SC_HD__INV_12%VGND N_VGND_M1001_s N_VGND_M1002_s N_VGND_M1005_s
+ N_VGND_M1009_s N_VGND_M1011_s N_VGND_M1014_s N_VGND_M1022_s N_VGND_c_660_n
+ N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n
+ N_VGND_c_666_n N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n N_VGND_c_670_n
+ N_VGND_c_671_n N_VGND_c_672_n N_VGND_c_673_n N_VGND_c_674_n N_VGND_c_675_n
+ N_VGND_c_676_n N_VGND_c_677_n VGND N_VGND_c_678_n N_VGND_c_679_n
+ N_VGND_c_680_n PM_SKY130_FD_SC_HD__INV_12%VGND
cc_1 VNB N_A_c_88_n 0.0191475f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_2 VNB N_A_c_89_n 0.0157835f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_3 VNB N_A_c_90_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=0.995
cc_4 VNB N_A_c_91_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.995
cc_5 VNB N_A_c_92_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=0.995
cc_6 VNB N_A_c_93_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.995
cc_7 VNB N_A_c_94_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=0.995
cc_8 VNB N_A_c_95_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=0.995
cc_9 VNB N_A_c_96_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.995
cc_10 VNB N_A_c_97_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=4.415 $Y2=0.995
cc_11 VNB N_A_c_98_n 0.0157991f $X=-0.19 $Y=-0.24 $X2=4.835 $Y2=0.995
cc_12 VNB N_A_c_99_n 0.019292f $X=-0.19 $Y=-0.24 $X2=5.255 $Y2=0.995
cc_13 VNB N_A_c_100_n 0.196058f $X=-0.19 $Y=-0.24 $X2=5.255 $Y2=1.16
cc_14 VNB N_VPWR_c_324_n 0.250759f $X=-0.19 $Y=-0.24 $X2=3.745 $Y2=1.105
cc_15 VNB N_Y_c_417_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=0.56
cc_16 VNB N_Y_c_418_n 0.016096f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=1.325
cc_17 VNB N_Y_c_419_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.995
cc_18 VNB N_Y_c_420_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=4.415 $Y2=1.985
cc_19 VNB N_Y_c_421_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=5.255 $Y2=1.325
cc_20 VNB N_Y_c_422_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=4.585 $Y2=1.105
cc_21 VNB N_Y_c_423_n 0.0117589f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_22 VNB N_Y_c_424_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=4.415 $Y2=1.16
cc_23 VNB N_Y_c_425_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=5.045 $Y2=1.16
cc_24 VNB N_Y_c_426_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_427_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.2
cc_26 VNB N_Y_c_428_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB Y 0.0249933f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.2
cc_28 VNB Y 0.0236239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_660_n 0.0145634f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.995
cc_30 VNB N_VGND_c_661_n 0.0166345f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.56
cc_31 VNB N_VGND_c_662_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_663_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=0.56
cc_33 VNB N_VGND_c_664_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=1.985
cc_34 VNB N_VGND_c_665_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.56
cc_35 VNB N_VGND_c_666_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_667_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=1.325
cc_37 VNB N_VGND_c_668_n 0.0114236f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=1.985
cc_38 VNB N_VGND_c_669_n 0.018193f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=0.995
cc_39 VNB N_VGND_c_670_n 0.0166611f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=0.56
cc_40 VNB N_VGND_c_671_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=1.325
cc_41 VNB N_VGND_c_672_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=1.985
cc_42 VNB N_VGND_c_673_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_674_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.56
cc_44 VNB N_VGND_c_675_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.56
cc_45 VNB N_VGND_c_676_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=1.985
cc_46 VNB N_VGND_c_677_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=1.985
cc_47 VNB N_VGND_c_678_n 0.0215456f $X=-0.19 $Y=-0.24 $X2=5.255 $Y2=0.56
cc_48 VNB N_VGND_c_679_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=1.985 $Y2=1.105
cc_49 VNB N_VGND_c_680_n 0.295472f $X=-0.19 $Y=-0.24 $X2=3.745 $Y2=1.105
cc_50 VPB N_A_M1000_g 0.0218766f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.985
cc_51 VPB N_A_M1003_g 0.0184996f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.985
cc_52 VPB N_A_M1006_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=1.985
cc_53 VPB N_A_M1007_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=1.985
cc_54 VPB N_A_M1012_g 0.0185065f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.985
cc_55 VPB N_A_M1015_g 0.0185065f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=1.985
cc_56 VPB N_A_M1016_g 0.0185065f $X=-0.19 $Y=1.305 $X2=3.155 $Y2=1.985
cc_57 VPB N_A_M1017_g 0.0185065f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.985
cc_58 VPB N_A_M1018_g 0.0185065f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=1.985
cc_59 VPB N_A_M1019_g 0.0185065f $X=-0.19 $Y=1.305 $X2=4.415 $Y2=1.985
cc_60 VPB N_A_M1021_g 0.0185044f $X=-0.19 $Y=1.305 $X2=4.835 $Y2=1.985
cc_61 VPB N_A_M1023_g 0.0221422f $X=-0.19 $Y=1.305 $X2=5.255 $Y2=1.985
cc_62 VPB N_A_c_100_n 0.0350807f $X=-0.19 $Y=1.305 $X2=5.255 $Y2=1.16
cc_63 VPB N_VPWR_c_325_n 0.0152107f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=0.995
cc_64 VPB N_VPWR_c_326_n 0.0294655f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=0.56
cc_65 VPB N_VPWR_c_327_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_328_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=0.56
cc_67 VPB N_VPWR_c_329_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.985
cc_68 VPB N_VPWR_c_330_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=0.56
cc_69 VPB N_VPWR_c_331_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_332_n 0.00410835f $X=-0.19 $Y=1.305 $X2=3.155 $Y2=1.325
cc_71 VPB N_VPWR_c_333_n 0.0114263f $X=-0.19 $Y=1.305 $X2=3.155 $Y2=1.985
cc_72 VPB N_VPWR_c_334_n 0.0315275f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=0.995
cc_73 VPB N_VPWR_c_335_n 0.017949f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=0.56
cc_74 VPB N_VPWR_c_336_n 0.00323736f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.325
cc_75 VPB N_VPWR_c_337_n 0.017949f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.985
cc_76 VPB N_VPWR_c_338_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_339_n 0.017949f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=0.56
cc_78 VPB N_VPWR_c_340_n 0.00323736f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=0.56
cc_79 VPB N_VPWR_c_341_n 0.017949f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=1.985
cc_80 VPB N_VPWR_c_342_n 0.00323736f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=1.985
cc_81 VPB N_VPWR_c_343_n 0.0235145f $X=-0.19 $Y=1.305 $X2=5.255 $Y2=0.56
cc_82 VPB N_VPWR_c_344_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.985 $Y2=1.105
cc_83 VPB N_VPWR_c_324_n 0.0496249f $X=-0.19 $Y=1.305 $X2=3.745 $Y2=1.105
cc_84 VPB N_Y_c_431_n 0.0150327f $X=-0.19 $Y=1.305 $X2=3.155 $Y2=1.985
cc_85 VPB N_Y_c_432_n 0.00769728f $X=-0.19 $Y=1.305 $X2=0.845 $Y2=1.16
cc_86 VPB Y 0.0117253f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.2
cc_87 VPB Y 0.0113004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 N_A_M1000_g N_VPWR_c_326_n 0.00321527f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VPWR_c_327_n 0.00146448f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_M1006_g N_VPWR_c_327_n 0.00146448f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_M1006_g N_VPWR_c_328_n 0.00541359f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_VPWR_c_328_n 0.00541359f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_M1007_g N_VPWR_c_329_n 0.00146448f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_M1012_g N_VPWR_c_329_n 0.00146448f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_M1015_g N_VPWR_c_330_n 0.00146448f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_M1016_g N_VPWR_c_330_n 0.00146448f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_M1017_g N_VPWR_c_331_n 0.00146448f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_M1018_g N_VPWR_c_331_n 0.00146448f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_M1019_g N_VPWR_c_332_n 0.00146448f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_M1021_g N_VPWR_c_332_n 0.00268723f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_M1023_g N_VPWR_c_334_n 0.0167864f $X=5.255 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_M1000_g N_VPWR_c_335_n 0.00541359f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_M1003_g N_VPWR_c_335_n 0.00541359f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_M1012_g N_VPWR_c_337_n 0.00541359f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_M1015_g N_VPWR_c_337_n 0.00541359f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_M1016_g N_VPWR_c_339_n 0.00541359f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_M1017_g N_VPWR_c_339_n 0.00541359f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1018_g N_VPWR_c_341_n 0.00541359f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_M1019_g N_VPWR_c_341_n 0.00541359f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_M1021_g N_VPWR_c_343_n 0.00541359f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_M1023_g N_VPWR_c_343_n 0.00541359f $X=5.255 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_M1000_g N_VPWR_c_324_n 0.0105807f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_M1003_g N_VPWR_c_324_n 0.00950154f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_M1006_g N_VPWR_c_324_n 0.00950154f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_M1007_g N_VPWR_c_324_n 0.00950154f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_M1012_g N_VPWR_c_324_n 0.00950154f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_M1015_g N_VPWR_c_324_n 0.00950154f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_M1016_g N_VPWR_c_324_n 0.00950154f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1017_g N_VPWR_c_324_n 0.00950154f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_M1018_g N_VPWR_c_324_n 0.00950154f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_M1019_g N_VPWR_c_324_n 0.00950154f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_M1021_g N_VPWR_c_324_n 0.00950154f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_M1023_g N_VPWR_c_324_n 0.0108685f $X=5.255 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_c_88_n N_Y_c_435_n 0.0109535f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_89_n N_Y_c_435_n 0.00631111f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_90_n N_Y_c_435_n 5.2007e-19 $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_M1000_g N_Y_c_438_n 0.0146918f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_M1003_g N_Y_c_438_n 0.00985707f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1006_g N_Y_c_438_n 6.20279e-19 $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_c_89_n N_Y_c_417_n 0.00890471f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_90_n N_Y_c_417_n 0.00890471f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_100_n N_Y_c_417_n 0.00222429f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_c_88_n N_Y_c_418_n 0.0138243f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_89_n N_Y_c_418_n 0.0012996f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_135 A N_Y_c_418_n 0.0611532f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_c_100_n N_Y_c_418_n 0.00222429f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_M1003_g N_Y_c_448_n 0.0107189f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1006_g N_Y_c_448_n 0.0107189f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_c_100_n N_Y_c_448_n 0.00201785f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_Y_c_431_n 0.0151128f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_Y_c_431_n 9.43996e-19 $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_142 A N_Y_c_431_n 0.0515679f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_c_100_n N_Y_c_431_n 0.00201785f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_c_89_n N_Y_c_455_n 5.19281e-19 $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_90_n N_Y_c_455_n 0.00620543f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_91_n N_Y_c_455_n 0.00620543f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_92_n N_Y_c_455_n 5.19281e-19 $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_M1003_g N_Y_c_459_n 6.1949e-19 $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_Y_c_459_n 0.00975139f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_Y_c_459_n 0.00975139f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1012_g N_Y_c_459_n 6.1949e-19 $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_c_91_n N_Y_c_419_n 0.00890471f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_92_n N_Y_c_419_n 0.00890471f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_154 A N_Y_c_419_n 0.0368812f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_c_100_n N_Y_c_419_n 0.00222429f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_M1007_g N_Y_c_467_n 0.0107189f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1012_g N_Y_c_467_n 0.0107189f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_158 A N_Y_c_467_n 0.0320704f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A_c_100_n N_Y_c_467_n 0.00201785f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_91_n N_Y_c_471_n 5.19281e-19 $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_92_n N_Y_c_471_n 0.00620543f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_93_n N_Y_c_471_n 0.00620543f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_94_n N_Y_c_471_n 5.19281e-19 $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_M1007_g N_Y_c_475_n 6.1949e-19 $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_M1012_g N_Y_c_475_n 0.00975139f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_M1015_g N_Y_c_475_n 0.00975139f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_M1016_g N_Y_c_475_n 6.1949e-19 $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_c_93_n N_Y_c_420_n 0.00890471f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_94_n N_Y_c_420_n 0.00890471f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_170 A N_Y_c_420_n 0.0368812f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A_c_100_n N_Y_c_420_n 0.00222429f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_M1015_g N_Y_c_483_n 0.0107189f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_M1016_g N_Y_c_483_n 0.0107189f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_174 A N_Y_c_483_n 0.0320704f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A_c_100_n N_Y_c_483_n 0.00201785f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_c_93_n N_Y_c_487_n 5.19281e-19 $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_94_n N_Y_c_487_n 0.00620543f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_95_n N_Y_c_487_n 0.00620543f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_96_n N_Y_c_487_n 5.19281e-19 $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_M1015_g N_Y_c_491_n 6.1949e-19 $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_M1016_g N_Y_c_491_n 0.00975139f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1017_g N_Y_c_491_n 0.00975139f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1018_g N_Y_c_491_n 6.1949e-19 $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_c_95_n N_Y_c_421_n 0.00890471f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_96_n N_Y_c_421_n 0.00890471f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_186 A N_Y_c_421_n 0.0368812f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A_c_100_n N_Y_c_421_n 0.00222429f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_M1017_g N_Y_c_499_n 0.0107189f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_M1018_g N_Y_c_499_n 0.0107189f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_190 A N_Y_c_499_n 0.0320704f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A_c_100_n N_Y_c_499_n 0.00201785f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_c_95_n N_Y_c_503_n 5.19281e-19 $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_96_n N_Y_c_503_n 0.00620543f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_97_n N_Y_c_503_n 0.00620543f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_98_n N_Y_c_503_n 5.19281e-19 $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_M1017_g N_Y_c_507_n 6.1949e-19 $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_M1018_g N_Y_c_507_n 0.00975139f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_M1019_g N_Y_c_507_n 0.00975139f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_M1021_g N_Y_c_507_n 6.1949e-19 $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_c_97_n N_Y_c_422_n 0.00890471f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_98_n N_Y_c_422_n 0.00890471f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_202 A N_Y_c_422_n 0.0368812f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A_c_100_n N_Y_c_422_n 0.00222429f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_M1019_g N_Y_c_515_n 0.0107189f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_M1021_g N_Y_c_515_n 0.0107189f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_206 A N_Y_c_515_n 0.0320704f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_207 N_A_c_100_n N_Y_c_515_n 0.00201785f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_c_97_n N_Y_c_519_n 5.19281e-19 $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_c_98_n N_Y_c_519_n 0.00620543f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_c_99_n N_Y_c_519_n 0.0121304f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_M1019_g N_Y_c_522_n 6.1949e-19 $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_M1021_g N_Y_c_522_n 0.00975139f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_M1023_g N_Y_c_522_n 0.0174034f $X=5.255 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_c_99_n N_Y_c_423_n 0.0118214f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_215 A N_Y_c_423_n 0.00419161f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A_M1023_g N_Y_c_432_n 0.0134103f $X=5.255 $Y=1.985 $X2=0 $Y2=0
cc_217 A N_Y_c_432_n 0.00415709f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_218 N_A_c_90_n N_Y_c_424_n 0.00116017f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_91_n N_Y_c_424_n 0.00116017f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_220 A N_Y_c_424_n 0.0269421f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_221 N_A_c_100_n N_Y_c_424_n 0.00230339f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_M1006_g N_Y_c_533_n 8.84614e-19 $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_M1007_g N_Y_c_533_n 8.84614e-19 $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_224 A N_Y_c_533_n 0.0213676f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_225 N_A_c_100_n N_Y_c_533_n 0.00209661f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_c_92_n N_Y_c_425_n 0.00116017f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_93_n N_Y_c_425_n 0.00116017f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_228 A N_Y_c_425_n 0.0269421f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_229 N_A_c_100_n N_Y_c_425_n 0.00230339f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_M1012_g N_Y_c_541_n 8.84614e-19 $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A_M1015_g N_Y_c_541_n 8.84614e-19 $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_232 A N_Y_c_541_n 0.0213676f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A_c_100_n N_Y_c_541_n 0.00209661f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_c_94_n N_Y_c_426_n 0.00116017f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_c_95_n N_Y_c_426_n 0.00116017f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_236 A N_Y_c_426_n 0.0269421f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_237 N_A_c_100_n N_Y_c_426_n 0.00230339f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_M1016_g N_Y_c_549_n 8.84614e-19 $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A_M1017_g N_Y_c_549_n 8.84614e-19 $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_240 A N_Y_c_549_n 0.0213676f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_241 N_A_c_100_n N_Y_c_549_n 0.00209661f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_c_96_n N_Y_c_427_n 0.00116017f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_97_n N_Y_c_427_n 0.00116017f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_244 A N_Y_c_427_n 0.0269421f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_245 N_A_c_100_n N_Y_c_427_n 0.00230339f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_M1018_g N_Y_c_557_n 8.84614e-19 $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_M1019_g N_Y_c_557_n 8.84614e-19 $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_248 A N_Y_c_557_n 0.0213676f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_249 N_A_c_100_n N_Y_c_557_n 0.00209661f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_c_98_n N_Y_c_428_n 0.00116017f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_99_n N_Y_c_428_n 0.00116017f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_252 A N_Y_c_428_n 0.0269421f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A_c_100_n N_Y_c_428_n 0.00230339f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_M1021_g N_Y_c_565_n 8.84614e-19 $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_M1023_g N_Y_c_565_n 8.84614e-19 $X=5.255 $Y=1.985 $X2=0 $Y2=0
cc_256 A N_Y_c_565_n 0.0213676f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_257 N_A_c_100_n N_Y_c_565_n 0.00209661f $X=5.255 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_c_88_n Y 0.0229913f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_259 A Y 0.0212121f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_260 N_A_c_99_n Y 0.0192911f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_261 A Y 0.0145692f $X=5.005 $Y=1.105 $X2=0 $Y2=0
cc_262 N_A_c_88_n N_VGND_c_661_n 0.00321527f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_c_89_n N_VGND_c_662_n 0.00146448f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_c_90_n N_VGND_c_662_n 0.00146448f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_c_90_n N_VGND_c_663_n 0.00422241f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_c_91_n N_VGND_c_663_n 0.00422241f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_91_n N_VGND_c_664_n 0.00146448f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_c_92_n N_VGND_c_664_n 0.00146448f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_c_93_n N_VGND_c_665_n 0.00146448f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_c_94_n N_VGND_c_665_n 0.00146448f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_c_95_n N_VGND_c_666_n 0.00146448f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_c_96_n N_VGND_c_666_n 0.00146448f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_c_97_n N_VGND_c_667_n 0.00146448f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_c_98_n N_VGND_c_667_n 0.00268723f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A_c_99_n N_VGND_c_669_n 0.00988424f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A_c_88_n N_VGND_c_670_n 0.00421248f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A_c_89_n N_VGND_c_670_n 0.00421248f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_c_92_n N_VGND_c_672_n 0.00422241f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_c_93_n N_VGND_c_672_n 0.00422241f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A_c_94_n N_VGND_c_674_n 0.00422241f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A_c_95_n N_VGND_c_674_n 0.00422241f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_c_96_n N_VGND_c_676_n 0.00422241f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A_c_97_n N_VGND_c_676_n 0.00422241f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A_c_98_n N_VGND_c_678_n 0.00422241f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A_c_99_n N_VGND_c_678_n 0.00422241f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_c_88_n N_VGND_c_680_n 0.0067902f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A_c_89_n N_VGND_c_680_n 0.00571103f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_c_90_n N_VGND_c_680_n 0.00569656f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_c_91_n N_VGND_c_680_n 0.00569656f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A_c_92_n N_VGND_c_680_n 0.00569656f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A_c_93_n N_VGND_c_680_n 0.00569656f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_292 N_A_c_94_n N_VGND_c_680_n 0.00569656f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_c_95_n N_VGND_c_680_n 0.00569656f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_c_96_n N_VGND_c_680_n 0.00569656f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_c_97_n N_VGND_c_680_n 0.00569656f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_c_98_n N_VGND_c_680_n 0.00569656f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A_c_99_n N_VGND_c_680_n 0.00703192f $X=5.255 $Y=0.995 $X2=0 $Y2=0
cc_298 N_VPWR_c_324_n N_Y_M1000_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_c_324_n N_Y_M1006_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_324_n N_Y_M1012_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_324_n N_Y_M1016_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_324_n N_Y_M1018_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_303 N_VPWR_c_324_n N_Y_M1021_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_304 N_VPWR_c_335_n N_Y_c_438_n 0.0189039f $X=1.18 $Y=2.72 $X2=0 $Y2=0
cc_305 N_VPWR_c_324_n N_Y_c_438_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_306 N_VPWR_M1003_s N_Y_c_448_n 0.00311483f $X=1.13 $Y=1.485 $X2=0 $Y2=0
cc_307 N_VPWR_c_327_n N_Y_c_448_n 0.0126919f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_308 N_VPWR_M1000_s N_Y_c_431_n 0.00350209f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_309 N_VPWR_c_326_n N_Y_c_431_n 0.020232f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_310 N_VPWR_c_328_n N_Y_c_459_n 0.0189039f $X=2.02 $Y=2.72 $X2=0 $Y2=0
cc_311 N_VPWR_c_324_n N_Y_c_459_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_312 N_VPWR_M1007_s N_Y_c_467_n 0.00311483f $X=1.97 $Y=1.485 $X2=0 $Y2=0
cc_313 N_VPWR_c_329_n N_Y_c_467_n 0.0126919f $X=2.105 $Y=2 $X2=0 $Y2=0
cc_314 N_VPWR_c_337_n N_Y_c_475_n 0.0189039f $X=2.86 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_324_n N_Y_c_475_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_M1015_s N_Y_c_483_n 0.00311483f $X=2.81 $Y=1.485 $X2=0 $Y2=0
cc_317 N_VPWR_c_330_n N_Y_c_483_n 0.0126919f $X=2.945 $Y=2 $X2=0 $Y2=0
cc_318 N_VPWR_c_339_n N_Y_c_491_n 0.0189039f $X=3.7 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_c_324_n N_Y_c_491_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_M1017_s N_Y_c_499_n 0.00311483f $X=3.65 $Y=1.485 $X2=0 $Y2=0
cc_321 N_VPWR_c_331_n N_Y_c_499_n 0.0126919f $X=3.785 $Y=2 $X2=0 $Y2=0
cc_322 N_VPWR_c_341_n N_Y_c_507_n 0.0189039f $X=4.54 $Y=2.72 $X2=0 $Y2=0
cc_323 N_VPWR_c_324_n N_Y_c_507_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_M1019_s N_Y_c_515_n 0.00311483f $X=4.49 $Y=1.485 $X2=0 $Y2=0
cc_325 N_VPWR_c_332_n N_Y_c_515_n 0.0126919f $X=4.625 $Y=2 $X2=0 $Y2=0
cc_326 N_VPWR_c_334_n N_Y_c_522_n 0.02848f $X=5.72 $Y=2 $X2=0 $Y2=0
cc_327 N_VPWR_c_343_n N_Y_c_522_n 0.0189039f $X=5.555 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_c_324_n N_Y_c_522_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_329 N_VPWR_M1023_s N_Y_c_432_n 0.015685f $X=5.33 $Y=1.485 $X2=0 $Y2=0
cc_330 N_VPWR_c_334_n N_Y_c_432_n 0.0306479f $X=5.72 $Y=2 $X2=0 $Y2=0
cc_331 N_VPWR_M1000_s Y 6.44532e-19 $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_332 N_VPWR_M1023_s Y 2.66588e-19 $X=5.33 $Y=1.485 $X2=0 $Y2=0
cc_333 N_Y_c_418_n N_VGND_M1001_s 0.00285834f $X=1.01 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_334 N_Y_c_417_n N_VGND_M1002_s 0.00162148f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_335 N_Y_c_419_n N_VGND_M1005_s 0.00162148f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_336 N_Y_c_420_n N_VGND_M1009_s 0.00162148f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_337 N_Y_c_421_n N_VGND_M1011_s 0.00162148f $X=4.04 $Y=0.81 $X2=0 $Y2=0
cc_338 N_Y_c_422_n N_VGND_M1014_s 0.00162148f $X=4.88 $Y=0.81 $X2=0 $Y2=0
cc_339 N_Y_c_423_n N_VGND_M1022_s 0.009453f $X=5.545 $Y=0.81 $X2=0 $Y2=0
cc_340 N_Y_c_418_n N_VGND_c_660_n 0.00267039f $X=1.01 $Y=0.81 $X2=0 $Y2=0
cc_341 N_Y_c_418_n N_VGND_c_661_n 0.0195556f $X=1.01 $Y=0.81 $X2=0 $Y2=0
cc_342 N_Y_c_417_n N_VGND_c_662_n 0.0122675f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_343 N_Y_c_417_n N_VGND_c_663_n 0.00203746f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_344 N_Y_c_455_n N_VGND_c_663_n 0.0188551f $X=1.685 $Y=0.38 $X2=0 $Y2=0
cc_345 N_Y_c_419_n N_VGND_c_663_n 0.00203746f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_346 N_Y_c_419_n N_VGND_c_664_n 0.0122675f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_347 N_Y_c_420_n N_VGND_c_665_n 0.0122675f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_348 N_Y_c_421_n N_VGND_c_666_n 0.0122675f $X=4.04 $Y=0.81 $X2=0 $Y2=0
cc_349 N_Y_c_422_n N_VGND_c_667_n 0.0122675f $X=4.88 $Y=0.81 $X2=0 $Y2=0
cc_350 N_Y_c_519_n N_VGND_c_669_n 0.0131099f $X=5.045 $Y=0.38 $X2=0 $Y2=0
cc_351 N_Y_c_423_n N_VGND_c_669_n 0.0293195f $X=5.545 $Y=0.81 $X2=0 $Y2=0
cc_352 N_Y_c_435_n N_VGND_c_670_n 0.0184921f $X=0.845 $Y=0.38 $X2=0 $Y2=0
cc_353 N_Y_c_418_n N_VGND_c_670_n 0.0041083f $X=1.01 $Y=0.81 $X2=0 $Y2=0
cc_354 N_Y_c_419_n N_VGND_c_672_n 0.00203746f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_355 N_Y_c_471_n N_VGND_c_672_n 0.0188551f $X=2.525 $Y=0.38 $X2=0 $Y2=0
cc_356 N_Y_c_420_n N_VGND_c_672_n 0.00203746f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_357 N_Y_c_420_n N_VGND_c_674_n 0.00203746f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_358 N_Y_c_487_n N_VGND_c_674_n 0.0188551f $X=3.365 $Y=0.38 $X2=0 $Y2=0
cc_359 N_Y_c_421_n N_VGND_c_674_n 0.00203746f $X=4.04 $Y=0.81 $X2=0 $Y2=0
cc_360 N_Y_c_421_n N_VGND_c_676_n 0.00203746f $X=4.04 $Y=0.81 $X2=0 $Y2=0
cc_361 N_Y_c_503_n N_VGND_c_676_n 0.0188551f $X=4.205 $Y=0.38 $X2=0 $Y2=0
cc_362 N_Y_c_422_n N_VGND_c_676_n 0.00203746f $X=4.88 $Y=0.81 $X2=0 $Y2=0
cc_363 N_Y_c_422_n N_VGND_c_678_n 0.00203746f $X=4.88 $Y=0.81 $X2=0 $Y2=0
cc_364 N_Y_c_519_n N_VGND_c_678_n 0.0188551f $X=5.045 $Y=0.38 $X2=0 $Y2=0
cc_365 N_Y_c_423_n N_VGND_c_678_n 0.00460273f $X=5.545 $Y=0.81 $X2=0 $Y2=0
cc_366 N_Y_M1001_d N_VGND_c_680_n 0.00215201f $X=0.71 $Y=0.235 $X2=0 $Y2=0
cc_367 N_Y_M1004_d N_VGND_c_680_n 0.00215201f $X=1.55 $Y=0.235 $X2=0 $Y2=0
cc_368 N_Y_M1008_d N_VGND_c_680_n 0.00215201f $X=2.39 $Y=0.235 $X2=0 $Y2=0
cc_369 N_Y_M1010_d N_VGND_c_680_n 0.00215201f $X=3.23 $Y=0.235 $X2=0 $Y2=0
cc_370 N_Y_M1013_d N_VGND_c_680_n 0.00215201f $X=4.07 $Y=0.235 $X2=0 $Y2=0
cc_371 N_Y_M1020_d N_VGND_c_680_n 0.00215201f $X=4.91 $Y=0.235 $X2=0 $Y2=0
cc_372 N_Y_c_435_n N_VGND_c_680_n 0.012098f $X=0.845 $Y=0.38 $X2=0 $Y2=0
cc_373 N_Y_c_417_n N_VGND_c_680_n 0.00455756f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_374 N_Y_c_418_n N_VGND_c_680_n 0.0134275f $X=1.01 $Y=0.81 $X2=0 $Y2=0
cc_375 N_Y_c_455_n N_VGND_c_680_n 0.0122069f $X=1.685 $Y=0.38 $X2=0 $Y2=0
cc_376 N_Y_c_419_n N_VGND_c_680_n 0.00845923f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_377 N_Y_c_471_n N_VGND_c_680_n 0.0122069f $X=2.525 $Y=0.38 $X2=0 $Y2=0
cc_378 N_Y_c_420_n N_VGND_c_680_n 0.00845923f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_379 N_Y_c_487_n N_VGND_c_680_n 0.0122069f $X=3.365 $Y=0.38 $X2=0 $Y2=0
cc_380 N_Y_c_421_n N_VGND_c_680_n 0.00845923f $X=4.04 $Y=0.81 $X2=0 $Y2=0
cc_381 N_Y_c_503_n N_VGND_c_680_n 0.0122069f $X=4.205 $Y=0.38 $X2=0 $Y2=0
cc_382 N_Y_c_422_n N_VGND_c_680_n 0.00845923f $X=4.88 $Y=0.81 $X2=0 $Y2=0
cc_383 N_Y_c_519_n N_VGND_c_680_n 0.0122069f $X=5.045 $Y=0.38 $X2=0 $Y2=0
cc_384 N_Y_c_423_n N_VGND_c_680_n 0.0101637f $X=5.545 $Y=0.81 $X2=0 $Y2=0

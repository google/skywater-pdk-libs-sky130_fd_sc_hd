* File: sky130_fd_sc_hd__lpflow_decapkapwr_8.pxi.spice
* Created: Tue Sep  1 19:11:56 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%VGND N_VGND_M1001_s N_VGND_M1000_g
+ N_VGND_c_18_n N_VGND_c_19_n VGND N_VGND_c_20_n N_VGND_c_21_n N_VGND_c_22_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%KAPWR N_KAPWR_M1000_s N_KAPWR_M1001_g
+ KAPWR N_KAPWR_c_40_n N_KAPWR_c_41_n N_KAPWR_c_43_n N_KAPWR_c_42_n
+ N_KAPWR_c_45_n N_KAPWR_c_46_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%VPWR VPWR N_VPWR_c_66_n N_VPWR_c_65_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%VPWR
cc_1 VNB N_VGND_c_18_n 0.0184325f $X=-0.19 $Y=-0.24 $X2=3.125 $Y2=0.385
cc_2 VNB N_VGND_c_19_n 0.0803762f $X=-0.19 $Y=-0.24 $X2=1.735 $Y2=0.385
cc_3 VNB N_VGND_c_20_n 0.0461317f $X=-0.19 $Y=-0.24 $X2=1.715 $Y2=1.87
cc_4 VNB N_VGND_c_21_n 0.0439808f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.475
cc_5 VNB N_VGND_c_22_n 0.19806f $X=-0.19 $Y=-0.24 $X2=3.45 $Y2=0
cc_6 VNB N_KAPWR_c_40_n 0.112251f $X=-0.19 $Y=-0.24 $X2=1.55 $Y2=1.87
cc_7 VNB N_KAPWR_c_41_n 0.171284f $X=-0.19 $Y=-0.24 $X2=1.55 $Y2=1.29
cc_8 VNB N_KAPWR_c_42_n 0.017777f $X=-0.19 $Y=-0.24 $X2=3.45 $Y2=0
cc_9 VNB N_VPWR_c_65_n 0.155873f $X=-0.19 $Y=-0.24 $X2=1.84 $Y2=2.05
cc_10 VPB N_VGND_c_19_n 0.00687456f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=0.385
cc_11 VPB N_VGND_c_20_n 0.253553f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=1.87
cc_12 VPB N_KAPWR_c_43_n 0.0353425f $X=-0.19 $Y=1.305 $X2=1.55 $Y2=0.645
cc_13 VPB N_KAPWR_c_42_n 0.045107f $X=-0.19 $Y=1.305 $X2=3.45 $Y2=0
cc_14 VPB N_KAPWR_c_45_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0
cc_15 VPB N_KAPWR_c_46_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_16 VPB N_VPWR_c_66_n 0.0875376f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=2.05
cc_17 VPB N_VPWR_c_65_n 0.0421982f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=2.05
cc_18 N_VGND_c_18_n N_KAPWR_c_40_n 0.0203072f $X=3.125 $Y=0.385 $X2=0 $Y2=0
cc_19 N_VGND_c_19_n N_KAPWR_c_40_n 0.150639f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_20 N_VGND_c_20_n N_KAPWR_c_40_n 0.0905514f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_21 N_VGND_c_18_n N_KAPWR_c_41_n 0.123274f $X=3.125 $Y=0.385 $X2=0 $Y2=0
cc_22 N_VGND_c_19_n N_KAPWR_c_41_n 0.00652589f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_23 N_VGND_c_20_n N_KAPWR_c_41_n 0.0987678f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_24 N_VGND_c_21_n N_KAPWR_c_41_n 0.0237254f $X=3.42 $Y=0.475 $X2=0 $Y2=0
cc_25 N_VGND_c_19_n N_KAPWR_c_43_n 0.141865f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_26 N_VGND_c_20_n N_KAPWR_c_43_n 0.169718f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_27 N_VGND_c_18_n N_KAPWR_c_42_n 0.102303f $X=3.125 $Y=0.385 $X2=0 $Y2=0
cc_28 N_VGND_c_19_n N_KAPWR_c_42_n 0.0326918f $X=1.735 $Y=0.385 $X2=0 $Y2=0
cc_29 N_VGND_c_20_n N_KAPWR_c_42_n 0.166937f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_30 N_VGND_c_21_n N_KAPWR_c_42_n 0.0424044f $X=3.42 $Y=0.475 $X2=0 $Y2=0
cc_31 N_VGND_c_20_n N_VPWR_c_66_n 0.0689298f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_32 N_VGND_c_20_n N_VPWR_c_65_n 0.0625156f $X=1.715 $Y=1.87 $X2=0 $Y2=0
cc_33 N_KAPWR_c_43_n N_VPWR_c_66_n 0.23514f $X=1.905 $Y=1.745 $X2=0 $Y2=0
cc_34 N_KAPWR_c_46_n N_VPWR_c_66_n 0.00247149f $X=0.215 $Y=2.21 $X2=0 $Y2=0
cc_35 N_KAPWR_M1000_s N_VPWR_c_65_n 0.00214099f $X=0.135 $Y=1.615 $X2=0 $Y2=0
cc_36 N_KAPWR_c_43_n N_VPWR_c_65_n 0.0294489f $X=1.905 $Y=1.745 $X2=0 $Y2=0
cc_37 N_KAPWR_c_46_n N_VPWR_c_65_n 0.361635f $X=0.215 $Y=2.21 $X2=0 $Y2=0

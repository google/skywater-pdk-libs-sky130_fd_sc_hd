* File: sky130_fd_sc_hd__nor4bb_1.pex.spice
* Created: Tue Sep  1 19:19:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%C_N 3 7 8 9 13 14 15
r33 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r34 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r36 8 9 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.53
r37 8 14 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.16
r38 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.51 $Y=0.675
+ $X2=0.51 $Y2=0.995
r39 3 16 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.47 $Y=2.26
+ $X2=0.47 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%D_N 3 6 8 11 13
r33 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.16
+ $X2=1.035 $Y2=1.325
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.16
+ $X2=1.035 $Y2=0.995
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r36 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.035 $Y2=1.16
r37 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.955 $Y=1.695
+ $X2=0.955 $Y2=1.325
r38 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.95 $Y=0.675
+ $X2=0.95 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%A_205_93# 1 2 7 9 12 14 15 16 23 25 28 30
r65 28 31 8.28933 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.547 $Y=1.16
+ $X2=1.547 $Y2=1.325
r66 28 30 8.28933 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.547 $Y=1.16
+ $X2=1.547 $Y2=0.995
r67 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r68 25 26 17.5021 $w=2.37e-07 $l=3.4e-07 $layer=LI1_cond $X=1.16 $Y=0.655
+ $X2=1.5 $Y2=0.655
r69 23 31 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=1.5 $Y=1.525 $X2=1.5
+ $Y2=1.325
r70 20 26 2.35055 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=1.5 $Y=0.825 $X2=1.5
+ $Y2=0.655
r71 20 30 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.5 $Y=0.825 $X2=1.5
+ $Y2=0.995
r72 16 23 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=1.41 $Y=1.62
+ $X2=1.5 $Y2=1.525
r73 16 18 14.3014 $w=1.88e-07 $l=2.45e-07 $layer=LI1_cond $X=1.41 $Y=1.62
+ $X2=1.165 $Y2=1.62
r74 14 29 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=1.6 $Y2=1.16
r75 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=1.89 $Y2=1.16
r76 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=1.89 $Y2=1.16
r77 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=1.89 $Y2=1.985
r78 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=0.995
+ $X2=1.89 $Y2=1.16
r79 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.89 $Y=0.995 $X2=1.89
+ $Y2=0.56
r80 2 18 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.63
r81 1 25 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.465 $X2=1.16 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%A_27_410# 1 2 7 9 12 15 18 20 23 24 25 28
+ 29 34 36
c81 28 0 1.59638e-19 $X=2.31 $Y=1.16
r82 31 34 3.93367 $w=3.73e-07 $l=1.28e-07 $layer=LI1_cond $X=0.172 $Y=0.637
+ $X2=0.3 $Y2=0.637
r83 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.16 $X2=2.31 $Y2=1.16
r84 26 28 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.31 $Y=2.295
+ $X2=2.31 $Y2=1.16
r85 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.225 $Y=2.38
+ $X2=2.31 $Y2=2.295
r86 24 25 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.225 $Y=2.38
+ $X2=1.205 $Y2=2.38
r87 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=2.295
+ $X2=1.205 $Y2=2.38
r88 22 23 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.12 $Y=2.07
+ $X2=1.12 $Y2=2.295
r89 21 36 1.93133 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.977
+ $X2=0.215 $Y2=1.977
r90 20 22 6.83233 $w=1.85e-07 $l=1.28662e-07 $layer=LI1_cond $X=1.035 $Y=1.977
+ $X2=1.12 $Y2=2.07
r91 20 21 41.3661 $w=1.83e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.977
+ $X2=0.345 $Y2=1.977
r92 16 36 4.5059 $w=2.17e-07 $l=9.3e-08 $layer=LI1_cond $X=0.215 $Y=2.07
+ $X2=0.215 $Y2=1.977
r93 16 18 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.215 $Y=2.07
+ $X2=0.215 $Y2=2.29
r94 15 36 4.5059 $w=2.17e-07 $l=1.11445e-07 $layer=LI1_cond $X=0.172 $Y=1.885
+ $X2=0.215 $Y2=1.977
r95 14 31 5.2298 $w=1.75e-07 $l=1.88e-07 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=0.637
r96 14 15 67.1792 $w=1.73e-07 $l=1.06e-06 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=1.885
r97 10 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.325
+ $X2=2.31 $Y2=1.16
r98 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.31 $Y=1.325
+ $X2=2.31 $Y2=1.985
r99 7 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=0.995
+ $X2=2.31 $Y2=1.16
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.31 $Y=0.995
+ $X2=2.31 $Y2=0.56
r101 2 18 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r102 1 34 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.465 $X2=0.3 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%B 1 3 6 10 14 15
c40 14 0 4.81382e-20 $X=2.79 $Y=1.16
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.16 $X2=2.79 $Y2=1.16
r42 10 15 9.03851 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.78 $Y=1.445
+ $X2=2.78 $Y2=1.16
r43 4 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.325
+ $X2=2.79 $Y2=1.16
r44 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.79 $Y=1.325 $X2=2.79
+ $Y2=1.985
r45 1 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.995
+ $X2=2.79 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.79 $Y=0.995 $X2=2.79
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%A 3 6 8 12 14 19
c28 19 0 4.81382e-20 $X=3.45 $Y=1.49
r29 17 23 0.291325 $w=3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.445 $Y=1.275
+ $X2=3.445 $Y2=1.135
r30 16 19 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=3.445 $Y=1.49
+ $X2=3.45 $Y2=1.49
r31 16 17 2.84566 $w=3e-07 $l=2.15e-07 $layer=LI1_cond $X=3.445 $Y=1.49
+ $X2=3.445 $Y2=1.275
r32 13 23 5.96801 $w=2.78e-07 $l=1.45e-07 $layer=LI1_cond $X=3.3 $Y=1.135
+ $X2=3.445 $Y2=1.135
r33 12 15 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.302 $Y=1.16
+ $X2=3.302 $Y2=1.325
r34 12 14 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.302 $Y=1.16
+ $X2=3.302 $Y2=0.995
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.3
+ $Y=1.16 $X2=3.3 $Y2=1.16
r36 8 23 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.135
+ $X2=3.445 $Y2=1.135
r37 8 19 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.45 $Y=1.275
+ $X2=3.45 $Y2=1.49
r38 6 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.985
+ $X2=3.21 $Y2=1.325
r39 3 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.56 $X2=3.21
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%VPWR 1 2 9 11 13 15 17 22 31 35
r46 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r49 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r55 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 22 34 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=3.467 $Y2=2.72
r57 22 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r59 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 11 34 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.42 $Y=2.635
+ $X2=3.467 $Y2=2.72
r63 11 13 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.42 $Y=2.635
+ $X2=3.42 $Y2=2
r64 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r65 7 9 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.325
r66 2 13 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=2
r67 1 9 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.05 $X2=0.68 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%Y 1 2 3 10 15 18 20 21 26
r52 25 26 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.985 $Y=0.655
+ $X2=2.985 $Y2=0.495
r53 20 25 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.885 $Y=0.74
+ $X2=2.985 $Y2=0.655
r54 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.885 $Y=0.74
+ $X2=2.215 $Y2=0.74
r55 16 21 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.115 $Y=0.74
+ $X2=2.215 $Y2=0.74
r56 16 18 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.115 $Y=0.655
+ $X2=2.115 $Y2=0.495
r57 14 16 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=2.115 $Y2=0.74
r58 14 15 62.6636 $w=1.98e-07 $l=1.13e-06 $layer=LI1_cond $X=1.955 $Y=0.825
+ $X2=1.955 $Y2=1.955
r59 10 15 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.855 $Y=2.04
+ $X2=1.955 $Y2=1.955
r60 10 12 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=2.04
+ $X2=1.68 $Y2=2.04
r61 3 12 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.895 $X2=1.68 $Y2=2.04
r62 2 26 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3 $Y2=0.495
r63 1 18 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.235 $X2=2.1 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_1%VGND 1 2 3 4 17 21 25 27 29 31 33 38 43 49
+ 52 55 59 61
r59 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r60 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r61 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r62 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r63 47 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r64 47 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r65 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r66 44 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.55
+ $Y2=0
r67 44 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.99
+ $Y2=0
r68 43 58 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r69 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r70 42 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r71 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r72 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 39 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.68
+ $Y2=0
r74 39 41 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=2.07
+ $Y2=0
r75 38 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.55
+ $Y2=0
r76 38 41 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.07
+ $Y2=0
r77 37 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r78 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r79 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r80 34 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.74
+ $Y2=0
r81 34 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=1.15
+ $Y2=0
r82 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.68
+ $Y2=0
r83 33 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.15
+ $Y2=0
r84 31 50 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r85 31 61 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r86 27 58 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.467 $Y2=0
r87 27 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.39
r88 23 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=0.085
+ $X2=2.55 $Y2=0
r89 23 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.55 $Y=0.085
+ $X2=2.55 $Y2=0.39
r90 19 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0
r91 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0.38
r92 15 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r93 15 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.66
r94 4 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.39
r95 3 25 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.235 $X2=2.55 $Y2=0.39
r96 2 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.68 $Y2=0.38
r97 1 17 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.465 $X2=0.74 $Y2=0.66
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
M1000 Y B a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.08e+12p pd=1.016e+07u as=2.44e+12p ps=2.288e+07u
M1001 a_27_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.08e+12p ps=1.016e+07u
M1002 a_27_297# B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.404e+12p pd=1.472e+07u as=1.5795e+12p ps=1.656e+07u
M1005 Y B a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_297# B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_297# B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y B a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND B Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_27_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y B a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__mux4_1.pxi.spice
* Created: Tue Sep  1 19:15:00 2020
* 
x_PM_SKY130_FD_SC_HD__MUX4_1%A1 N_A1_M1021_g N_A1_M1010_g A1 A1 N_A1_c_191_n
+ N_A1_c_192_n PM_SKY130_FD_SC_HD__MUX4_1%A1
x_PM_SKY130_FD_SC_HD__MUX4_1%A0 N_A0_M1013_g N_A0_M1025_g A0 A0 N_A0_c_221_n
+ N_A0_c_222_n PM_SKY130_FD_SC_HD__MUX4_1%A0
x_PM_SKY130_FD_SC_HD__MUX4_1%A_247_21# N_A_247_21#_M1006_s N_A_247_21#_M1002_s
+ N_A_247_21#_M1017_g N_A_247_21#_c_259_n N_A_247_21#_c_260_n
+ N_A_247_21#_M1014_g N_A_247_21#_c_261_n N_A_247_21#_M1022_g
+ N_A_247_21#_M1008_g N_A_247_21#_c_262_n N_A_247_21#_c_263_n
+ N_A_247_21#_c_277_n N_A_247_21#_c_264_n N_A_247_21#_c_265_n
+ N_A_247_21#_c_266_n N_A_247_21#_c_267_n N_A_247_21#_c_268_n
+ N_A_247_21#_c_269_n N_A_247_21#_c_270_n N_A_247_21#_c_271_n
+ PM_SKY130_FD_SC_HD__MUX4_1%A_247_21#
x_PM_SKY130_FD_SC_HD__MUX4_1%S0 N_S0_M1011_g N_S0_c_421_n N_S0_c_422_n
+ N_S0_c_428_n N_S0_M1012_g N_S0_c_429_n N_S0_c_430_n N_S0_M1006_g N_S0_c_424_n
+ N_S0_M1002_g N_S0_c_433_n N_S0_c_425_n N_S0_M1018_g N_S0_c_434_n N_S0_M1000_g
+ N_S0_c_426_n S0 S0 N_S0_c_427_n PM_SKY130_FD_SC_HD__MUX4_1%S0
x_PM_SKY130_FD_SC_HD__MUX4_1%A3 N_A3_M1004_g N_A3_M1023_g A3 A3 N_A3_c_529_n
+ PM_SKY130_FD_SC_HD__MUX4_1%A3
x_PM_SKY130_FD_SC_HD__MUX4_1%A2 N_A2_M1019_g N_A2_M1024_g A2 N_A2_c_576_n
+ N_A2_c_577_n PM_SKY130_FD_SC_HD__MUX4_1%A2
x_PM_SKY130_FD_SC_HD__MUX4_1%S1 N_S1_M1009_g N_S1_M1015_g N_S1_c_618_n
+ N_S1_M1001_g N_S1_M1005_g N_S1_c_620_n S1 N_S1_c_621_n
+ PM_SKY130_FD_SC_HD__MUX4_1%S1
x_PM_SKY130_FD_SC_HD__MUX4_1%A_1290_413# N_A_1290_413#_M1015_d
+ N_A_1290_413#_M1009_d N_A_1290_413#_M1003_g N_A_1290_413#_c_697_n
+ N_A_1290_413#_M1007_g N_A_1290_413#_c_698_n N_A_1290_413#_c_699_n
+ N_A_1290_413#_c_747_p N_A_1290_413#_c_706_n N_A_1290_413#_c_718_n
+ N_A_1290_413#_c_700_n N_A_1290_413#_c_721_n N_A_1290_413#_c_723_n
+ N_A_1290_413#_c_701_n N_A_1290_413#_c_702_n N_A_1290_413#_c_703_n
+ PM_SKY130_FD_SC_HD__MUX4_1%A_1290_413#
x_PM_SKY130_FD_SC_HD__MUX4_1%A_1478_413# N_A_1478_413#_M1005_d
+ N_A_1478_413#_M1001_d N_A_1478_413#_M1020_g N_A_1478_413#_M1016_g
+ N_A_1478_413#_c_805_n N_A_1478_413#_c_797_n N_A_1478_413#_c_806_n
+ N_A_1478_413#_c_798_n N_A_1478_413#_c_807_n N_A_1478_413#_c_808_n
+ N_A_1478_413#_c_799_n N_A_1478_413#_c_800_n N_A_1478_413#_c_801_n
+ N_A_1478_413#_c_802_n N_A_1478_413#_c_811_n N_A_1478_413#_c_813_n
+ N_A_1478_413#_c_803_n PM_SKY130_FD_SC_HD__MUX4_1%A_1478_413#
x_PM_SKY130_FD_SC_HD__MUX4_1%A_27_413# N_A_27_413#_M1010_s N_A_27_413#_M1014_s
+ N_A_27_413#_c_892_n N_A_27_413#_c_893_n N_A_27_413#_c_894_n
+ N_A_27_413#_c_895_n PM_SKY130_FD_SC_HD__MUX4_1%A_27_413#
x_PM_SKY130_FD_SC_HD__MUX4_1%VPWR N_VPWR_M1010_d N_VPWR_M1002_d N_VPWR_M1004_d
+ N_VPWR_M1009_s N_VPWR_M1016_s N_VPWR_c_924_n N_VPWR_c_925_n N_VPWR_c_926_n
+ N_VPWR_c_927_n N_VPWR_c_928_n VPWR N_VPWR_c_929_n N_VPWR_c_930_n
+ N_VPWR_c_931_n N_VPWR_c_932_n N_VPWR_c_933_n N_VPWR_c_934_n N_VPWR_c_923_n
+ N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_940_n
+ PM_SKY130_FD_SC_HD__MUX4_1%VPWR
x_PM_SKY130_FD_SC_HD__MUX4_1%A_193_413# N_A_193_413#_M1025_d
+ N_A_193_413#_M1012_d N_A_193_413#_c_1038_n N_A_193_413#_c_1039_n
+ N_A_193_413#_c_1046_n PM_SKY130_FD_SC_HD__MUX4_1%A_193_413#
x_PM_SKY130_FD_SC_HD__MUX4_1%A_277_47# N_A_277_47#_M1017_d N_A_277_47#_M1007_d
+ N_A_277_47#_M1014_d N_A_277_47#_M1001_s N_A_277_47#_c_1061_n
+ N_A_277_47#_c_1062_n N_A_277_47#_c_1072_n N_A_277_47#_c_1073_n
+ N_A_277_47#_c_1074_n N_A_277_47#_c_1094_n N_A_277_47#_c_1142_n
+ N_A_277_47#_c_1063_n N_A_277_47#_c_1064_n N_A_277_47#_c_1065_n
+ N_A_277_47#_c_1066_n N_A_277_47#_c_1067_n N_A_277_47#_c_1068_n
+ N_A_277_47#_c_1069_n N_A_277_47#_c_1070_n PM_SKY130_FD_SC_HD__MUX4_1%A_277_47#
x_PM_SKY130_FD_SC_HD__MUX4_1%A_757_363# N_A_757_363#_M1000_s
+ N_A_757_363#_M1019_d N_A_757_363#_c_1227_n N_A_757_363#_c_1228_n
+ N_A_757_363#_c_1229_n N_A_757_363#_c_1230_n N_A_757_363#_c_1231_n
+ N_A_757_363#_c_1235_n N_A_757_363#_c_1251_n
+ PM_SKY130_FD_SC_HD__MUX4_1%A_757_363#
x_PM_SKY130_FD_SC_HD__MUX4_1%A_750_97# N_A_750_97#_M1018_d N_A_750_97#_M1005_s
+ N_A_750_97#_M1000_d N_A_750_97#_M1003_d N_A_750_97#_c_1284_n
+ N_A_750_97#_c_1285_n N_A_750_97#_c_1288_n N_A_750_97#_c_1289_n
+ N_A_750_97#_c_1334_n N_A_750_97#_c_1286_n N_A_750_97#_c_1338_n
+ N_A_750_97#_c_1291_n N_A_750_97#_c_1292_n N_A_750_97#_c_1293_n
+ N_A_750_97#_c_1294_n N_A_750_97#_c_1309_n N_A_750_97#_c_1312_n
+ N_A_750_97#_c_1295_n PM_SKY130_FD_SC_HD__MUX4_1%A_750_97#
x_PM_SKY130_FD_SC_HD__MUX4_1%X N_X_M1020_d N_X_M1016_d X X X X N_X_c_1428_n
+ PM_SKY130_FD_SC_HD__MUX4_1%X
x_PM_SKY130_FD_SC_HD__MUX4_1%A_27_47# N_A_27_47#_M1021_s N_A_27_47#_M1011_d
+ N_A_27_47#_c_1470_p N_A_27_47#_c_1438_n N_A_27_47#_c_1439_n
+ N_A_27_47#_c_1440_n N_A_27_47#_c_1474_p N_A_27_47#_c_1452_n
+ PM_SKY130_FD_SC_HD__MUX4_1%A_27_47#
x_PM_SKY130_FD_SC_HD__MUX4_1%VGND N_VGND_M1021_d N_VGND_M1006_d N_VGND_M1023_d
+ N_VGND_M1015_s N_VGND_M1020_s N_VGND_c_1481_n N_VGND_c_1482_n N_VGND_c_1483_n
+ N_VGND_c_1484_n N_VGND_c_1485_n N_VGND_c_1486_n N_VGND_c_1487_n VGND
+ N_VGND_c_1488_n N_VGND_c_1489_n N_VGND_c_1490_n N_VGND_c_1491_n
+ N_VGND_c_1492_n N_VGND_c_1493_n N_VGND_c_1494_n N_VGND_c_1495_n
+ N_VGND_c_1496_n N_VGND_c_1497_n VGND PM_SKY130_FD_SC_HD__MUX4_1%VGND
x_PM_SKY130_FD_SC_HD__MUX4_1%A_668_97# N_A_668_97#_M1018_s N_A_668_97#_M1023_s
+ N_A_668_97#_c_1607_n N_A_668_97#_c_1608_n N_A_668_97#_c_1609_n
+ N_A_668_97#_c_1610_n PM_SKY130_FD_SC_HD__MUX4_1%A_668_97#
x_PM_SKY130_FD_SC_HD__MUX4_1%A_834_97# N_A_834_97#_M1022_d N_A_834_97#_M1024_d
+ N_A_834_97#_c_1638_n N_A_834_97#_c_1639_n N_A_834_97#_c_1640_n
+ PM_SKY130_FD_SC_HD__MUX4_1%A_834_97#
cc_1 VNB N_A1_M1021_g 0.0370886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_A1_c_191_n 0.0263062f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_3 VNB N_A1_c_192_n 0.0147234f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_4 VNB N_A0_M1013_g 0.0267303f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB N_A0_c_221_n 0.0203849f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_6 VNB N_A0_c_222_n 0.00302416f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_7 VNB N_A_247_21#_M1017_g 0.039604f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_247_21#_c_259_n 0.0145372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_247_21#_c_260_n 0.00312847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_247_21#_c_261_n 0.0396449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_247_21#_c_262_n 0.00536329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_247_21#_c_263_n 0.0155941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_247_21#_c_264_n 0.00124855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_247_21#_c_265_n 3.18678e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_247_21#_c_266_n 0.00292092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_247_21#_c_267_n 0.00128471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_247_21#_c_268_n 0.0249485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_247_21#_c_269_n 0.00693159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_247_21#_c_270_n 0.0346971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_247_21#_c_271_n 7.28774e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_S0_M1011_g 0.0195856f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_22 VNB N_S0_c_421_n 0.0675826f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_23 VNB N_S0_c_422_n 0.00996749f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_24 VNB N_S0_M1006_g 0.0219522f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_25 VNB N_S0_c_424_n 0.0336865f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_26 VNB N_S0_c_425_n 0.0341692f $X=-0.19 $Y=-0.24 $X2=0.322 $Y2=1.53
cc_27 VNB N_S0_c_426_n 0.0296253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_S0_c_427_n 0.0023899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A3_M1023_g 0.0398286f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_30 VNB A3 0.0027769f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_31 VNB N_A3_c_529_n 0.0210206f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_32 VNB N_A2_M1024_g 0.0387257f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_33 VNB N_A2_c_576_n 0.0183248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_c_577_n 0.00238465f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_35 VNB N_S1_M1015_g 0.0413384f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_36 VNB N_S1_c_618_n 0.0446949f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_37 VNB N_S1_M1005_g 0.0386981f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.325
cc_38 VNB N_S1_c_620_n 0.0110613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_S1_c_621_n 0.0321546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_1290_413#_c_697_n 0.0443346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_1290_413#_c_698_n 0.023361f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_42 VNB N_A_1290_413#_c_699_n 0.0073821f $X=-0.19 $Y=-0.24 $X2=0.322 $Y2=1.16
cc_43 VNB N_A_1290_413#_c_700_n 0.00420902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_1290_413#_c_701_n 0.00433766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_1290_413#_c_702_n 0.00262343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1290_413#_c_703_n 0.0232052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1478_413#_c_797_n 0.01374f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_48 VNB N_A_1478_413#_c_798_n 0.00693865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1478_413#_c_799_n 0.00685641f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1478_413#_c_800_n 0.00446709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1478_413#_c_801_n 0.00281946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1478_413#_c_802_n 0.0341616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1478_413#_c_803_n 0.0231009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_923_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_277_47#_c_1061_n 0.00488695f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_56 VNB N_A_277_47#_c_1062_n 0.00720023f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_57 VNB N_A_277_47#_c_1063_n 8.87589e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_277_47#_c_1064_n 0.0594603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_277_47#_c_1065_n 0.00202786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_277_47#_c_1066_n 0.00531848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_277_47#_c_1067_n 0.00261641f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_277_47#_c_1068_n 0.0043336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_277_47#_c_1069_n 0.00235731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_277_47#_c_1070_n 0.00253606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_750_97#_c_1284_n 9.2887e-19 $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_66 VNB N_A_750_97#_c_1285_n 0.0022651f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_67 VNB N_A_750_97#_c_1286_n 0.00616232f $X=-0.19 $Y=-0.24 $X2=0.322 $Y2=1.19
cc_68 VNB N_X_c_1428_n 0.0459692f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_69 VNB N_A_27_47#_c_1438_n 0.0111123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_27_47#_c_1439_n 0.00773178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_27_47#_c_1440_n 0.0058115f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_72 VNB N_VGND_c_1481_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.322 $Y2=1.16
cc_73 VNB N_VGND_c_1482_n 0.00900064f $X=-0.19 $Y=-0.24 $X2=0.322 $Y2=1.53
cc_74 VNB N_VGND_c_1483_n 0.00465285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1484_n 0.00563081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1485_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1486_n 0.049433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1487_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1488_n 0.015156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1489_n 0.0465196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1490_n 0.0191075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1491_n 0.0645756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1492_n 0.0184263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1493_n 0.472375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1494_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1495_n 0.00445369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1496_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1497_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_668_97#_c_1607_n 0.00113673f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_90 VNB N_A_668_97#_c_1608_n 0.00302147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_668_97#_c_1609_n 0.00208227f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_92 VNB N_A_668_97#_c_1610_n 0.013963f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_93 VNB N_A_834_97#_c_1638_n 0.0221352f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_94 VNB N_A_834_97#_c_1639_n 9.27166e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_834_97#_c_1640_n 0.00120445f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_96 VPB N_A1_M1010_g 0.06139f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_97 VPB N_A1_c_191_n 0.0049065f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_98 VPB N_A1_c_192_n 0.0149434f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_99 VPB N_A0_M1025_g 0.0602517f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_100 VPB N_A0_c_221_n 0.00460787f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_101 VPB N_A0_c_222_n 0.00737362f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_102 VPB N_A_247_21#_c_259_n 0.0104228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_247_21#_c_260_n 0.005512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_247_21#_M1014_g 0.0618159f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_105 VPB N_A_247_21#_M1008_g 0.0506501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_247_21#_c_262_n 4.7758e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_247_21#_c_277_n 0.0124205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_247_21#_c_265_n 2.6814e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_247_21#_c_266_n 0.00380445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_247_21#_c_268_n 0.00790865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_247_21#_c_269_n 0.00461028f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_247_21#_c_270_n 0.0114912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_S0_c_428_n 0.0323478f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_114 VPB N_S0_c_429_n 0.0216189f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_115 VPB N_S0_c_430_n 0.00769376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_S0_c_424_n 0.0453787f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_117 VPB N_S0_M1002_g 0.0345364f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.16
cc_118 VPB N_S0_c_433_n 0.0536074f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.19
cc_119 VPB N_S0_c_434_n 0.0317412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_S0_c_426_n 0.0111026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_S0_c_427_n 0.0119741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A3_M1004_g 0.0437263f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_123 VPB A3 0.00428172f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_124 VPB N_A3_c_529_n 0.0100844f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_125 VPB N_A2_M1019_g 0.0557383f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_126 VPB N_A2_c_576_n 0.00897023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A2_c_577_n 0.00798755f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_128 VPB N_S1_M1009_g 0.0683492f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_129 VPB N_S1_c_618_n 0.0218761f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_130 VPB N_S1_M1001_g 0.0571198f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_131 VPB N_S1_c_620_n 8.97301e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB S1 0.00700498f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.19
cc_133 VPB N_S1_c_621_n 0.0103462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_1290_413#_M1003_g 0.0672785f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_135 VPB N_A_1290_413#_c_698_n 0.00984038f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_136 VPB N_A_1290_413#_c_706_n 0.0155675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_1290_413#_c_701_n 0.00168011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_1290_413#_c_703_n 0.0176975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_1478_413#_M1016_g 0.0254972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_1478_413#_c_805_n 0.0240254f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_141 VPB N_A_1478_413#_c_806_n 0.00811431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_1478_413#_c_807_n 0.0136122f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.53
cc_143 VPB N_A_1478_413#_c_808_n 0.00499843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_1478_413#_c_801_n 0.00549657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_1478_413#_c_802_n 0.00789238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_1478_413#_c_811_n 0.00103517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_413#_c_892_n 0.00443274f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_148 VPB N_A_27_413#_c_893_n 0.0250146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_413#_c_894_n 0.00862673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_27_413#_c_895_n 0.00141558f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_151 VPB N_VPWR_c_924_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.16
cc_152 VPB N_VPWR_c_925_n 0.00547095f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.53
cc_153 VPB N_VPWR_c_926_n 4.09336e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_927_n 0.00558492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_928_n 0.00625317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_929_n 0.0153006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_930_n 0.0553846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_931_n 0.0357036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_932_n 0.0153204f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_933_n 0.0619547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_934_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_923_n 0.0967259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_936_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_937_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_938_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_939_n 0.00545594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_940_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_193_413#_c_1038_n 0.0203731f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_169 VPB N_A_193_413#_c_1039_n 0.00237213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_277_47#_c_1062_n 0.00197524f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_171 VPB N_A_277_47#_c_1072_n 0.00524683f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_172 VPB N_A_277_47#_c_1073_n 0.00353869f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_173 VPB N_A_277_47#_c_1074_n 0.00179107f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.16
cc_174 VPB N_A_277_47#_c_1063_n 0.014198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_757_363#_c_1227_n 0.00275204f $X=-0.19 $Y=1.305 $X2=0.15
+ $Y2=1.105
cc_176 VPB N_A_757_363#_c_1228_n 0.00738038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_757_363#_c_1229_n 0.00295611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_757_363#_c_1230_n 4.98462e-19 $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_179 VPB N_A_757_363#_c_1231_n 0.00770732f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_180 VPB N_A_750_97#_c_1285_n 0.00252139f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_181 VPB N_A_750_97#_c_1288_n 0.00326526f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_182 VPB N_A_750_97#_c_1289_n 0.00127018f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_183 VPB N_A_750_97#_c_1286_n 0.00850746f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=1.19
cc_184 VPB N_A_750_97#_c_1291_n 0.00162979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_750_97#_c_1292_n 0.00300209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_750_97#_c_1293_n 0.00210497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_750_97#_c_1294_n 0.0473489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_750_97#_c_1295_n 0.00198097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_X_c_1428_n 0.0469154f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_190 N_A1_M1021_g N_A0_M1013_g 0.0266891f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A1_M1010_g N_A0_M1025_g 0.0447338f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_192 N_A1_c_192_n N_A0_M1025_g 3.41851e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A1_c_191_n N_A0_c_221_n 0.0198624f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A1_c_192_n N_A0_c_221_n 0.00106441f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A1_M1010_g N_A0_c_222_n 0.00193042f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_196 N_A1_c_191_n N_A0_c_222_n 0.00106296f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A1_c_192_n N_A0_c_222_n 0.03074f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A1_M1010_g N_A_27_413#_c_892_n 0.0046335f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_199 N_A1_M1010_g N_A_27_413#_c_893_n 0.0147274f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_200 N_A1_c_192_n N_A_27_413#_c_893_n 0.0111339f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A1_c_191_n N_A_27_413#_c_894_n 2.94677e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A1_c_192_n N_A_27_413#_c_894_n 0.0151696f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A1_M1010_g N_VPWR_c_924_n 0.00844918f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_204 N_A1_M1010_g N_VPWR_c_929_n 0.0035268f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_205 N_A1_M1010_g N_VPWR_c_923_n 0.00513527f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_206 N_A1_M1021_g N_A_27_47#_c_1438_n 0.0142497f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A1_c_191_n N_A_27_47#_c_1438_n 3.41787e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A1_c_192_n N_A_27_47#_c_1438_n 0.010452f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A1_c_191_n N_A_27_47#_c_1439_n 5.32462e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A1_c_192_n N_A_27_47#_c_1439_n 0.0140568f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A1_M1021_g N_VGND_c_1481_n 0.00847734f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_212 N_A1_M1021_g N_VGND_c_1488_n 0.00339367f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A1_M1021_g N_VGND_c_1493_n 0.00489827f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A0_M1013_g N_A_247_21#_M1017_g 0.0388251f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A0_c_221_n N_A_247_21#_M1017_g 0.0213451f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A0_c_222_n N_A_247_21#_M1017_g 0.0034624f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A0_M1025_g N_A_247_21#_c_260_n 4.51557e-19 $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_218 N_A0_c_222_n N_A_247_21#_c_260_n 0.00359631f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A0_c_222_n N_A_247_21#_M1014_g 7.74559e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A0_M1025_g N_A_27_413#_c_893_n 0.0139122f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_221 N_A0_c_221_n N_A_27_413#_c_893_n 0.00165433f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A0_c_222_n N_A_27_413#_c_893_n 0.033605f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A0_M1025_g N_A_27_413#_c_895_n 0.00375953f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_224 N_A0_M1025_g N_VPWR_c_924_n 0.00844082f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_225 N_A0_M1025_g N_VPWR_c_930_n 0.0035268f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_226 N_A0_M1025_g N_VPWR_c_923_n 0.00550713f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_227 N_A0_M1025_g N_A_277_47#_c_1062_n 4.70277e-19 $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_228 N_A0_c_222_n N_A_277_47#_c_1062_n 0.0351905f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A0_M1025_g N_A_277_47#_c_1073_n 9.97182e-19 $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_230 N_A0_c_222_n N_A_277_47#_c_1073_n 0.0143623f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A0_M1013_g N_A_27_47#_c_1438_n 0.0110469f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A0_c_221_n N_A_27_47#_c_1438_n 0.00235482f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A0_c_222_n N_A_27_47#_c_1438_n 0.0289705f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A0_c_222_n N_A_27_47#_c_1440_n 0.0011019f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A0_M1013_g N_VGND_c_1481_n 0.00779668f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A0_M1013_g N_VGND_c_1489_n 0.00339367f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A0_M1013_g N_VGND_c_1493_n 0.00401529f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_238 N_A_247_21#_c_259_n N_S0_M1011_g 0.0101534f $X=1.755 $Y=1.26 $X2=0 $Y2=0
cc_239 N_A_247_21#_c_263_n N_S0_M1011_g 0.00351379f $X=2.525 $Y=0.595 $X2=0
+ $Y2=0
cc_240 N_A_247_21#_c_263_n N_S0_c_421_n 0.00696405f $X=2.525 $Y=0.595 $X2=0
+ $Y2=0
cc_241 N_A_247_21#_M1017_g N_S0_c_422_n 0.0238872f $X=1.31 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_247_21#_c_277_n N_S0_c_428_n 0.00267135f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_243 N_A_247_21#_c_266_n N_S0_c_429_n 0.0158556f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_244 N_A_247_21#_M1014_g N_S0_c_430_n 0.0302898f $X=1.83 $Y=2.025 $X2=0 $Y2=0
cc_245 N_A_247_21#_c_266_n N_S0_c_430_n 0.00372075f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_246 N_A_247_21#_c_268_n N_S0_c_430_n 0.0124712f $X=2.245 $Y=1.2 $X2=0 $Y2=0
cc_247 N_A_247_21#_c_263_n N_S0_M1006_g 0.0106695f $X=2.525 $Y=0.595 $X2=0 $Y2=0
cc_248 N_A_247_21#_c_277_n N_S0_c_424_n 0.0162487f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_249 N_A_247_21#_c_264_n N_S0_c_424_n 0.0167386f $X=4.23 $Y=1.19 $X2=0 $Y2=0
cc_250 N_A_247_21#_c_265_n N_S0_c_424_n 0.00308163f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_251 N_A_247_21#_c_266_n N_S0_c_424_n 0.0302191f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_252 N_A_247_21#_c_268_n N_S0_c_424_n 0.0150137f $X=2.245 $Y=1.2 $X2=0 $Y2=0
cc_253 N_A_247_21#_c_277_n N_S0_M1002_g 0.00960136f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_254 N_A_247_21#_M1008_g N_S0_c_433_n 0.0302956f $X=4.54 $Y=2.025 $X2=0 $Y2=0
cc_255 N_A_247_21#_c_270_n N_S0_c_433_n 0.00844233f $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_256 N_A_247_21#_c_261_n N_S0_c_425_n 0.0210934f $X=4.095 $Y=1.045 $X2=0 $Y2=0
cc_257 N_A_247_21#_M1008_g N_S0_c_426_n 4.03439e-19 $X=4.54 $Y=2.025 $X2=0 $Y2=0
cc_258 N_A_247_21#_c_264_n N_S0_c_426_n 0.00527604f $X=4.23 $Y=1.19 $X2=0 $Y2=0
cc_259 N_A_247_21#_c_270_n N_S0_c_426_n 0.0210934f $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_260 N_A_247_21#_c_271_n N_S0_c_426_n 2.26862e-19 $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_261 N_A_247_21#_c_263_n N_S0_c_427_n 0.00270649f $X=2.525 $Y=0.595 $X2=0
+ $Y2=0
cc_262 N_A_247_21#_c_277_n N_S0_c_427_n 0.0263973f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_263 N_A_247_21#_c_264_n N_S0_c_427_n 0.0202263f $X=4.23 $Y=1.19 $X2=0 $Y2=0
cc_264 N_A_247_21#_c_265_n N_S0_c_427_n 0.00161848f $X=2.68 $Y=1.19 $X2=0 $Y2=0
cc_265 N_A_247_21#_c_266_n N_S0_c_427_n 0.022126f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_266 N_A_247_21#_M1008_g N_A3_M1004_g 0.0427779f $X=4.54 $Y=2.025 $X2=0 $Y2=0
cc_267 N_A_247_21#_c_270_n N_A3_M1023_g 2.83612e-19 $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_268 N_A_247_21#_c_267_n A3 0.00734503f $X=4.375 $Y=1.19 $X2=0 $Y2=0
cc_269 N_A_247_21#_c_270_n A3 0.00723458f $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_270 N_A_247_21#_c_271_n A3 0.00556885f $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_271 N_A_247_21#_c_270_n N_A3_c_529_n 0.0165262f $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_272 N_A_247_21#_c_271_n N_A3_c_529_n 3.96659e-19 $X=4.24 $Y=1.18 $X2=0 $Y2=0
cc_273 N_A_247_21#_c_259_n N_A_27_413#_c_893_n 4.67198e-19 $X=1.755 $Y=1.26
+ $X2=0 $Y2=0
cc_274 N_A_247_21#_c_260_n N_A_27_413#_c_893_n 0.00509772f $X=1.385 $Y=1.26
+ $X2=0 $Y2=0
cc_275 N_A_247_21#_c_259_n N_A_27_413#_c_895_n 3.6921e-19 $X=1.755 $Y=1.26 $X2=0
+ $Y2=0
cc_276 N_A_247_21#_M1014_g N_A_27_413#_c_895_n 4.38572e-19 $X=1.83 $Y=2.025
+ $X2=0 $Y2=0
cc_277 N_A_247_21#_M1008_g N_VPWR_c_926_n 0.00117811f $X=4.54 $Y=2.025 $X2=0
+ $Y2=0
cc_278 N_A_247_21#_M1014_g N_VPWR_c_930_n 0.00357877f $X=1.83 $Y=2.025 $X2=0
+ $Y2=0
cc_279 N_A_247_21#_c_277_n N_VPWR_c_930_n 0.0244536f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_280 N_A_247_21#_M1008_g N_VPWR_c_931_n 0.00354535f $X=4.54 $Y=2.025 $X2=0
+ $Y2=0
cc_281 N_A_247_21#_M1002_s N_VPWR_c_923_n 0.00382897f $X=2.855 $Y=2.155 $X2=0
+ $Y2=0
cc_282 N_A_247_21#_M1014_g N_VPWR_c_923_n 0.00666029f $X=1.83 $Y=2.025 $X2=0
+ $Y2=0
cc_283 N_A_247_21#_M1008_g N_VPWR_c_923_n 0.00531323f $X=4.54 $Y=2.025 $X2=0
+ $Y2=0
cc_284 N_A_247_21#_c_277_n N_VPWR_c_923_n 0.0134021f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_285 N_A_247_21#_M1014_g N_A_193_413#_c_1038_n 0.0133031f $X=1.83 $Y=2.025
+ $X2=0 $Y2=0
cc_286 N_A_247_21#_c_277_n N_A_193_413#_c_1038_n 0.0151015f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_287 N_A_247_21#_c_266_n N_A_193_413#_c_1038_n 0.00293046f $X=2.535 $Y=1.19
+ $X2=0 $Y2=0
cc_288 N_A_247_21#_c_277_n N_A_193_413#_c_1039_n 0.0392297f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_289 N_A_247_21#_c_265_n N_A_193_413#_c_1039_n 6.76379e-19 $X=2.68 $Y=1.19
+ $X2=0 $Y2=0
cc_290 N_A_247_21#_c_266_n N_A_193_413#_c_1039_n 0.0144458f $X=2.535 $Y=1.19
+ $X2=0 $Y2=0
cc_291 N_A_247_21#_M1014_g N_A_193_413#_c_1046_n 0.00375953f $X=1.83 $Y=2.025
+ $X2=0 $Y2=0
cc_292 N_A_247_21#_M1017_g N_A_277_47#_c_1061_n 0.00543554f $X=1.31 $Y=0.445
+ $X2=0 $Y2=0
cc_293 N_A_247_21#_c_259_n N_A_277_47#_c_1061_n 0.00293494f $X=1.755 $Y=1.26
+ $X2=0 $Y2=0
cc_294 N_A_247_21#_c_263_n N_A_277_47#_c_1061_n 0.00312887f $X=2.525 $Y=0.595
+ $X2=0 $Y2=0
cc_295 N_A_247_21#_M1017_g N_A_277_47#_c_1062_n 0.00515412f $X=1.31 $Y=0.445
+ $X2=0 $Y2=0
cc_296 N_A_247_21#_c_259_n N_A_277_47#_c_1062_n 0.0162054f $X=1.755 $Y=1.26
+ $X2=0 $Y2=0
cc_297 N_A_247_21#_M1014_g N_A_277_47#_c_1062_n 0.00405222f $X=1.83 $Y=2.025
+ $X2=0 $Y2=0
cc_298 N_A_247_21#_c_266_n N_A_277_47#_c_1062_n 0.00586601f $X=2.535 $Y=1.19
+ $X2=0 $Y2=0
cc_299 N_A_247_21#_c_268_n N_A_277_47#_c_1062_n 9.99087e-19 $X=2.245 $Y=1.2
+ $X2=0 $Y2=0
cc_300 N_A_247_21#_c_259_n N_A_277_47#_c_1072_n 0.00487332f $X=1.755 $Y=1.26
+ $X2=0 $Y2=0
cc_301 N_A_247_21#_M1014_g N_A_277_47#_c_1072_n 0.0135239f $X=1.83 $Y=2.025
+ $X2=0 $Y2=0
cc_302 N_A_247_21#_c_266_n N_A_277_47#_c_1072_n 0.0132538f $X=2.535 $Y=1.19
+ $X2=0 $Y2=0
cc_303 N_A_247_21#_c_269_n N_A_277_47#_c_1072_n 0.00577479f $X=2.08 $Y=1.2 $X2=0
+ $Y2=0
cc_304 N_A_247_21#_M1014_g N_A_277_47#_c_1074_n 0.01033f $X=1.83 $Y=2.025 $X2=0
+ $Y2=0
cc_305 N_A_247_21#_c_277_n N_A_277_47#_c_1074_n 0.00464826f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_306 N_A_247_21#_M1014_g N_A_277_47#_c_1094_n 0.00233366f $X=1.83 $Y=2.025
+ $X2=0 $Y2=0
cc_307 N_A_247_21#_c_266_n N_A_277_47#_c_1094_n 0.00216555f $X=2.535 $Y=1.19
+ $X2=0 $Y2=0
cc_308 N_A_247_21#_c_269_n N_A_277_47#_c_1094_n 0.0020311f $X=2.08 $Y=1.2 $X2=0
+ $Y2=0
cc_309 N_A_247_21#_M1006_s N_A_277_47#_c_1064_n 5.39371e-19 $X=2.4 $Y=0.45 $X2=0
+ $Y2=0
cc_310 N_A_247_21#_c_261_n N_A_277_47#_c_1064_n 0.00252647f $X=4.095 $Y=1.045
+ $X2=0 $Y2=0
cc_311 N_A_247_21#_c_262_n N_A_277_47#_c_1064_n 0.00504867f $X=1.83 $Y=1.26
+ $X2=0 $Y2=0
cc_312 N_A_247_21#_c_263_n N_A_277_47#_c_1064_n 0.028474f $X=2.525 $Y=0.595
+ $X2=0 $Y2=0
cc_313 N_A_247_21#_c_264_n N_A_277_47#_c_1064_n 0.12321f $X=4.23 $Y=1.19 $X2=0
+ $Y2=0
cc_314 N_A_247_21#_c_265_n N_A_277_47#_c_1064_n 0.0255397f $X=2.68 $Y=1.19 $X2=0
+ $Y2=0
cc_315 N_A_247_21#_c_266_n N_A_277_47#_c_1064_n 0.00730746f $X=2.535 $Y=1.19
+ $X2=0 $Y2=0
cc_316 N_A_247_21#_c_267_n N_A_277_47#_c_1064_n 0.0269008f $X=4.375 $Y=1.19
+ $X2=0 $Y2=0
cc_317 N_A_247_21#_c_268_n N_A_277_47#_c_1064_n 0.00428297f $X=2.245 $Y=1.2
+ $X2=0 $Y2=0
cc_318 N_A_247_21#_c_270_n N_A_277_47#_c_1064_n 0.00380009f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_319 N_A_247_21#_c_271_n N_A_277_47#_c_1064_n 0.00218034f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_320 N_A_247_21#_c_259_n N_A_277_47#_c_1065_n 0.00368177f $X=1.755 $Y=1.26
+ $X2=0 $Y2=0
cc_321 N_A_247_21#_c_263_n N_A_277_47#_c_1065_n 0.00184116f $X=2.525 $Y=0.595
+ $X2=0 $Y2=0
cc_322 N_A_247_21#_c_264_n N_A_757_363#_c_1227_n 5.3144e-19 $X=4.23 $Y=1.19
+ $X2=0 $Y2=0
cc_323 N_A_247_21#_M1008_g N_A_757_363#_c_1228_n 0.00986166f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_324 N_A_247_21#_M1008_g N_A_757_363#_c_1230_n 0.00153332f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_325 N_A_247_21#_M1008_g N_A_757_363#_c_1235_n 8.44061e-19 $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_326 N_A_247_21#_c_261_n N_A_750_97#_c_1284_n 0.00410949f $X=4.095 $Y=1.045
+ $X2=0 $Y2=0
cc_327 N_A_247_21#_c_264_n N_A_750_97#_c_1284_n 9.16332e-19 $X=4.23 $Y=1.19
+ $X2=0 $Y2=0
cc_328 N_A_247_21#_c_261_n N_A_750_97#_c_1285_n 0.00605631f $X=4.095 $Y=1.045
+ $X2=0 $Y2=0
cc_329 N_A_247_21#_M1008_g N_A_750_97#_c_1285_n 0.00242124f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_330 N_A_247_21#_c_264_n N_A_750_97#_c_1285_n 0.0115317f $X=4.23 $Y=1.19 $X2=0
+ $Y2=0
cc_331 N_A_247_21#_c_267_n N_A_750_97#_c_1285_n 0.00228911f $X=4.375 $Y=1.19
+ $X2=0 $Y2=0
cc_332 N_A_247_21#_c_271_n N_A_750_97#_c_1285_n 0.0119604f $X=4.24 $Y=1.18 $X2=0
+ $Y2=0
cc_333 N_A_247_21#_M1008_g N_A_750_97#_c_1288_n 0.00665247f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_334 N_A_247_21#_c_264_n N_A_750_97#_c_1288_n 0.00643575f $X=4.23 $Y=1.19
+ $X2=0 $Y2=0
cc_335 N_A_247_21#_c_267_n N_A_750_97#_c_1288_n 0.00356155f $X=4.375 $Y=1.19
+ $X2=0 $Y2=0
cc_336 N_A_247_21#_c_270_n N_A_750_97#_c_1288_n 0.00817365f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_337 N_A_247_21#_c_271_n N_A_750_97#_c_1288_n 0.0259392f $X=4.24 $Y=1.18 $X2=0
+ $Y2=0
cc_338 N_A_247_21#_M1008_g N_A_750_97#_c_1294_n 0.00406871f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_339 N_A_247_21#_M1008_g N_A_750_97#_c_1309_n 0.00363402f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_340 N_A_247_21#_c_267_n N_A_750_97#_c_1309_n 0.0130653f $X=4.375 $Y=1.19
+ $X2=0 $Y2=0
cc_341 N_A_247_21#_c_271_n N_A_750_97#_c_1309_n 2.59353e-19 $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_342 N_A_247_21#_M1008_g N_A_750_97#_c_1312_n 0.0108127f $X=4.54 $Y=2.025
+ $X2=0 $Y2=0
cc_343 N_A_247_21#_M1017_g N_A_27_47#_c_1438_n 0.00144871f $X=1.31 $Y=0.445
+ $X2=0 $Y2=0
cc_344 N_A_247_21#_M1017_g N_A_27_47#_c_1440_n 0.0138537f $X=1.31 $Y=0.445 $X2=0
+ $Y2=0
cc_345 N_A_247_21#_c_263_n N_A_27_47#_c_1452_n 0.0258306f $X=2.525 $Y=0.595
+ $X2=0 $Y2=0
cc_346 N_A_247_21#_c_266_n N_A_27_47#_c_1452_n 2.2046e-19 $X=2.535 $Y=1.19 $X2=0
+ $Y2=0
cc_347 N_A_247_21#_c_269_n N_A_27_47#_c_1452_n 0.00464914f $X=2.08 $Y=1.2 $X2=0
+ $Y2=0
cc_348 N_A_247_21#_M1017_g N_VGND_c_1481_n 0.00128204f $X=1.31 $Y=0.445 $X2=0
+ $Y2=0
cc_349 N_A_247_21#_c_263_n N_VGND_c_1482_n 0.0142589f $X=2.525 $Y=0.595 $X2=0
+ $Y2=0
cc_350 N_A_247_21#_c_264_n N_VGND_c_1482_n 9.35884e-19 $X=4.23 $Y=1.19 $X2=0
+ $Y2=0
cc_351 N_A_247_21#_c_266_n N_VGND_c_1482_n 0.00332889f $X=2.535 $Y=1.19 $X2=0
+ $Y2=0
cc_352 N_A_247_21#_c_261_n N_VGND_c_1486_n 0.00357877f $X=4.095 $Y=1.045 $X2=0
+ $Y2=0
cc_353 N_A_247_21#_M1017_g N_VGND_c_1489_n 0.00357877f $X=1.31 $Y=0.445 $X2=0
+ $Y2=0
cc_354 N_A_247_21#_c_263_n N_VGND_c_1489_n 0.0120781f $X=2.525 $Y=0.595 $X2=0
+ $Y2=0
cc_355 N_A_247_21#_M1017_g N_VGND_c_1493_n 0.00547802f $X=1.31 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_247_21#_c_261_n N_VGND_c_1493_n 0.00661646f $X=4.095 $Y=1.045 $X2=0
+ $Y2=0
cc_357 N_A_247_21#_c_263_n N_VGND_c_1493_n 0.00540324f $X=2.525 $Y=0.595 $X2=0
+ $Y2=0
cc_358 N_A_247_21#_c_261_n N_A_668_97#_c_1609_n 0.00108334f $X=4.095 $Y=1.045
+ $X2=0 $Y2=0
cc_359 N_A_247_21#_c_261_n N_A_668_97#_c_1610_n 0.0130507f $X=4.095 $Y=1.045
+ $X2=0 $Y2=0
cc_360 N_A_247_21#_c_270_n N_A_668_97#_c_1610_n 9.96285e-19 $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_361 N_A_247_21#_c_271_n N_A_668_97#_c_1610_n 0.00131554f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_362 N_A_247_21#_c_267_n N_A_834_97#_c_1638_n 5.63717e-19 $X=4.375 $Y=1.19
+ $X2=0 $Y2=0
cc_363 N_A_247_21#_c_270_n N_A_834_97#_c_1638_n 0.00486156f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_364 N_A_247_21#_c_271_n N_A_834_97#_c_1638_n 0.00380593f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_365 N_A_247_21#_c_261_n N_A_834_97#_c_1640_n 5.53411e-19 $X=4.095 $Y=1.045
+ $X2=0 $Y2=0
cc_366 N_A_247_21#_c_267_n N_A_834_97#_c_1640_n 9.41603e-19 $X=4.375 $Y=1.19
+ $X2=0 $Y2=0
cc_367 N_A_247_21#_c_270_n N_A_834_97#_c_1640_n 0.00393073f $X=4.24 $Y=1.18
+ $X2=0 $Y2=0
cc_368 N_A_247_21#_c_271_n N_A_834_97#_c_1640_n 0.0111811f $X=4.24 $Y=1.18 $X2=0
+ $Y2=0
cc_369 N_S0_M1002_g N_VPWR_c_925_n 0.0104129f $X=3.19 $Y=2.275 $X2=0 $Y2=0
cc_370 N_S0_c_433_n N_VPWR_c_925_n 9.44261e-19 $X=4.045 $Y=1.665 $X2=0 $Y2=0
cc_371 N_S0_c_434_n N_VPWR_c_925_n 0.00348769f $X=4.12 $Y=1.74 $X2=0 $Y2=0
cc_372 N_S0_c_427_n N_VPWR_c_925_n 0.0162672f $X=3.415 $Y=1.18 $X2=0 $Y2=0
cc_373 N_S0_c_428_n N_VPWR_c_930_n 0.00357877f $X=2.25 $Y=1.74 $X2=0 $Y2=0
cc_374 N_S0_M1002_g N_VPWR_c_930_n 0.0046653f $X=3.19 $Y=2.275 $X2=0 $Y2=0
cc_375 N_S0_c_434_n N_VPWR_c_931_n 0.00357877f $X=4.12 $Y=1.74 $X2=0 $Y2=0
cc_376 N_S0_c_428_n N_VPWR_c_923_n 0.00666937f $X=2.25 $Y=1.74 $X2=0 $Y2=0
cc_377 N_S0_M1002_g N_VPWR_c_923_n 0.00921786f $X=3.19 $Y=2.275 $X2=0 $Y2=0
cc_378 N_S0_c_434_n N_VPWR_c_923_n 0.00671933f $X=4.12 $Y=1.74 $X2=0 $Y2=0
cc_379 N_S0_c_427_n N_VPWR_c_923_n 0.00160573f $X=3.415 $Y=1.18 $X2=0 $Y2=0
cc_380 N_S0_c_428_n N_A_193_413#_c_1038_n 0.013436f $X=2.25 $Y=1.74 $X2=0 $Y2=0
cc_381 N_S0_c_428_n N_A_193_413#_c_1039_n 0.00432427f $X=2.25 $Y=1.74 $X2=0
+ $Y2=0
cc_382 N_S0_c_429_n N_A_193_413#_c_1039_n 0.00296089f $X=2.66 $Y=1.665 $X2=0
+ $Y2=0
cc_383 N_S0_M1011_g N_A_277_47#_c_1061_n 0.00435613f $X=1.795 $Y=0.615 $X2=0
+ $Y2=0
cc_384 N_S0_M1011_g N_A_277_47#_c_1062_n 3.40765e-19 $X=1.795 $Y=0.615 $X2=0
+ $Y2=0
cc_385 N_S0_M1011_g N_A_277_47#_c_1072_n 5.12805e-19 $X=1.795 $Y=0.615 $X2=0
+ $Y2=0
cc_386 N_S0_c_430_n N_A_277_47#_c_1072_n 3.14271e-19 $X=2.325 $Y=1.665 $X2=0
+ $Y2=0
cc_387 N_S0_c_430_n N_A_277_47#_c_1074_n 0.00292337f $X=2.325 $Y=1.665 $X2=0
+ $Y2=0
cc_388 N_S0_c_428_n N_A_277_47#_c_1094_n 0.00289673f $X=2.25 $Y=1.74 $X2=0 $Y2=0
cc_389 N_S0_M1011_g N_A_277_47#_c_1064_n 0.0049719f $X=1.795 $Y=0.615 $X2=0
+ $Y2=0
cc_390 N_S0_c_421_n N_A_277_47#_c_1064_n 0.00188296f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_391 N_S0_M1006_g N_A_277_47#_c_1064_n 0.00696464f $X=2.735 $Y=0.66 $X2=0
+ $Y2=0
cc_392 N_S0_c_424_n N_A_277_47#_c_1064_n 0.00721948f $X=3.19 $Y=1.74 $X2=0 $Y2=0
cc_393 N_S0_c_425_n N_A_277_47#_c_1064_n 0.00418482f $X=3.675 $Y=0.995 $X2=0
+ $Y2=0
cc_394 N_S0_c_427_n N_A_277_47#_c_1064_n 0.00552765f $X=3.415 $Y=1.18 $X2=0
+ $Y2=0
cc_395 N_S0_M1011_g N_A_277_47#_c_1065_n 0.00144514f $X=1.795 $Y=0.615 $X2=0
+ $Y2=0
cc_396 N_S0_M1002_g N_A_757_363#_c_1227_n 0.00502654f $X=3.19 $Y=2.275 $X2=0
+ $Y2=0
cc_397 N_S0_c_433_n N_A_757_363#_c_1227_n 0.0030015f $X=4.045 $Y=1.665 $X2=0
+ $Y2=0
cc_398 N_S0_c_434_n N_A_757_363#_c_1227_n 0.0038722f $X=4.12 $Y=1.74 $X2=0 $Y2=0
cc_399 N_S0_c_427_n N_A_757_363#_c_1227_n 0.0120326f $X=3.415 $Y=1.18 $X2=0
+ $Y2=0
cc_400 N_S0_c_434_n N_A_757_363#_c_1228_n 0.0144646f $X=4.12 $Y=1.74 $X2=0 $Y2=0
cc_401 N_S0_c_433_n N_A_750_97#_c_1284_n 4.13482e-19 $X=4.045 $Y=1.665 $X2=0
+ $Y2=0
cc_402 N_S0_c_425_n N_A_750_97#_c_1284_n 0.00564278f $X=3.675 $Y=0.995 $X2=0
+ $Y2=0
cc_403 N_S0_c_425_n N_A_750_97#_c_1285_n 0.00338926f $X=3.675 $Y=0.995 $X2=0
+ $Y2=0
cc_404 N_S0_c_426_n N_A_750_97#_c_1285_n 0.00780516f $X=3.6 $Y=1.18 $X2=0 $Y2=0
cc_405 N_S0_c_427_n N_A_750_97#_c_1285_n 0.0316639f $X=3.415 $Y=1.18 $X2=0 $Y2=0
cc_406 N_S0_c_433_n N_A_750_97#_c_1288_n 0.0125249f $X=4.045 $Y=1.665 $X2=0
+ $Y2=0
cc_407 N_S0_c_433_n N_A_750_97#_c_1289_n 0.00938569f $X=4.045 $Y=1.665 $X2=0
+ $Y2=0
cc_408 N_S0_c_427_n N_A_750_97#_c_1289_n 0.0147221f $X=3.415 $Y=1.18 $X2=0 $Y2=0
cc_409 N_S0_c_433_n N_A_750_97#_c_1312_n 0.00526604f $X=4.045 $Y=1.665 $X2=0
+ $Y2=0
cc_410 N_S0_c_434_n N_A_750_97#_c_1312_n 0.00626168f $X=4.12 $Y=1.74 $X2=0 $Y2=0
cc_411 N_S0_c_427_n N_A_750_97#_c_1312_n 0.00461702f $X=3.415 $Y=1.18 $X2=0
+ $Y2=0
cc_412 N_S0_M1011_g N_A_27_47#_c_1440_n 0.0112486f $X=1.795 $Y=0.615 $X2=0 $Y2=0
cc_413 N_S0_c_421_n N_A_27_47#_c_1440_n 0.00435006f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_414 N_S0_M1006_g N_A_27_47#_c_1440_n 0.00216821f $X=2.735 $Y=0.66 $X2=0 $Y2=0
cc_415 N_S0_M1006_g N_A_27_47#_c_1452_n 4.51098e-19 $X=2.735 $Y=0.66 $X2=0 $Y2=0
cc_416 N_S0_c_421_n N_VGND_c_1482_n 0.00720059f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_417 N_S0_M1006_g N_VGND_c_1482_n 0.0153813f $X=2.735 $Y=0.66 $X2=0 $Y2=0
cc_418 N_S0_c_424_n N_VGND_c_1482_n 0.00580626f $X=3.19 $Y=1.74 $X2=0 $Y2=0
cc_419 N_S0_c_425_n N_VGND_c_1482_n 0.00405432f $X=3.675 $Y=0.995 $X2=0 $Y2=0
cc_420 N_S0_c_425_n N_VGND_c_1486_n 0.00357877f $X=3.675 $Y=0.995 $X2=0 $Y2=0
cc_421 N_S0_c_422_n N_VGND_c_1489_n 0.0295744f $X=1.87 $Y=0.18 $X2=0 $Y2=0
cc_422 N_S0_c_421_n N_VGND_c_1493_n 0.0223142f $X=2.66 $Y=0.18 $X2=0 $Y2=0
cc_423 N_S0_c_422_n N_VGND_c_1493_n 0.0046026f $X=1.87 $Y=0.18 $X2=0 $Y2=0
cc_424 N_S0_c_425_n N_VGND_c_1493_n 0.00661646f $X=3.675 $Y=0.995 $X2=0 $Y2=0
cc_425 N_S0_M1006_g N_A_668_97#_c_1607_n 6.83003e-19 $X=2.735 $Y=0.66 $X2=0
+ $Y2=0
cc_426 N_S0_c_425_n N_A_668_97#_c_1607_n 0.0023199f $X=3.675 $Y=0.995 $X2=0
+ $Y2=0
cc_427 N_S0_c_426_n N_A_668_97#_c_1607_n 8.43873e-19 $X=3.6 $Y=1.18 $X2=0 $Y2=0
cc_428 N_S0_c_427_n N_A_668_97#_c_1607_n 0.00951121f $X=3.415 $Y=1.18 $X2=0
+ $Y2=0
cc_429 N_S0_M1006_g N_A_668_97#_c_1608_n 7.54046e-19 $X=2.735 $Y=0.66 $X2=0
+ $Y2=0
cc_430 N_S0_c_425_n N_A_668_97#_c_1610_n 0.0114064f $X=3.675 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_A3_M1004_g N_A2_M1019_g 0.0416743f $X=5.015 $Y=2.275 $X2=0 $Y2=0
cc_432 N_A3_M1023_g N_A2_M1024_g 0.0303284f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_433 A3 N_A2_c_576_n 5.79079e-19 $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_434 N_A3_c_529_n N_A2_c_576_n 0.020411f $X=4.96 $Y=1.22 $X2=0 $Y2=0
cc_435 N_A3_M1004_g N_A2_c_577_n 0.00184497f $X=5.015 $Y=2.275 $X2=0 $Y2=0
cc_436 A3 N_A2_c_577_n 0.041759f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_437 N_A3_c_529_n N_A2_c_577_n 0.00231347f $X=4.96 $Y=1.22 $X2=0 $Y2=0
cc_438 N_A3_M1004_g N_VPWR_c_926_n 0.00808692f $X=5.015 $Y=2.275 $X2=0 $Y2=0
cc_439 N_A3_M1004_g N_VPWR_c_931_n 0.00339367f $X=5.015 $Y=2.275 $X2=0 $Y2=0
cc_440 N_A3_M1004_g N_VPWR_c_923_n 0.00397532f $X=5.015 $Y=2.275 $X2=0 $Y2=0
cc_441 N_A3_M1023_g N_A_277_47#_c_1064_n 0.00387417f $X=5.025 $Y=0.445 $X2=0
+ $Y2=0
cc_442 A3 N_A_277_47#_c_1064_n 0.0061336f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_443 N_A3_c_529_n N_A_277_47#_c_1064_n 0.00123205f $X=4.96 $Y=1.22 $X2=0 $Y2=0
cc_444 N_A3_M1004_g N_A_757_363#_c_1228_n 0.00150156f $X=5.015 $Y=2.275 $X2=0
+ $Y2=0
cc_445 N_A3_M1004_g N_A_757_363#_c_1230_n 0.00418034f $X=5.015 $Y=2.275 $X2=0
+ $Y2=0
cc_446 N_A3_M1004_g N_A_757_363#_c_1231_n 0.0114586f $X=5.015 $Y=2.275 $X2=0
+ $Y2=0
cc_447 A3 N_A_757_363#_c_1231_n 0.00969037f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_448 N_A3_c_529_n N_A_757_363#_c_1231_n 0.00161983f $X=4.96 $Y=1.22 $X2=0
+ $Y2=0
cc_449 A3 N_A_757_363#_c_1235_n 0.00168148f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_450 A3 N_A_750_97#_c_1288_n 0.00899167f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_451 N_A3_M1004_g N_A_750_97#_c_1294_n 0.00442447f $X=5.015 $Y=2.275 $X2=0
+ $Y2=0
cc_452 A3 N_A_750_97#_c_1294_n 0.00658083f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_453 N_A3_c_529_n N_A_750_97#_c_1294_n 0.00128625f $X=4.96 $Y=1.22 $X2=0 $Y2=0
cc_454 N_A3_M1004_g N_A_750_97#_c_1309_n 2.19299e-19 $X=5.015 $Y=2.275 $X2=0
+ $Y2=0
cc_455 N_A3_M1004_g N_A_750_97#_c_1312_n 0.00180779f $X=5.015 $Y=2.275 $X2=0
+ $Y2=0
cc_456 A3 N_A_750_97#_c_1312_n 0.00297673f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_457 N_A3_M1023_g N_VGND_c_1483_n 0.00268723f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_458 N_A3_M1023_g N_VGND_c_1486_n 0.00420765f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_459 N_A3_M1023_g N_VGND_c_1493_n 0.00676015f $X=5.025 $Y=0.445 $X2=0 $Y2=0
cc_460 N_A3_M1023_g N_A_668_97#_c_1609_n 0.00290799f $X=5.025 $Y=0.445 $X2=0
+ $Y2=0
cc_461 N_A3_M1023_g N_A_834_97#_c_1638_n 0.0136885f $X=5.025 $Y=0.445 $X2=0
+ $Y2=0
cc_462 A3 N_A_834_97#_c_1638_n 0.0165172f $X=4.8 $Y=1.105 $X2=0 $Y2=0
cc_463 N_A3_c_529_n N_A_834_97#_c_1638_n 0.00251569f $X=4.96 $Y=1.22 $X2=0 $Y2=0
cc_464 N_A3_M1023_g N_A_834_97#_c_1639_n 8.44629e-19 $X=5.025 $Y=0.445 $X2=0
+ $Y2=0
cc_465 N_A3_M1023_g N_A_834_97#_c_1640_n 0.00371709f $X=5.025 $Y=0.445 $X2=0
+ $Y2=0
cc_466 N_A2_c_576_n N_S1_M1009_g 6.8064e-19 $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_467 N_A2_M1019_g S1 0.00154017f $X=5.435 $Y=2.275 $X2=0 $Y2=0
cc_468 N_A2_M1024_g S1 2.91523e-19 $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_469 N_A2_c_576_n S1 0.00156318f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_470 N_A2_c_577_n S1 0.0226551f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_471 N_A2_M1024_g N_S1_c_621_n 0.00176601f $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_472 N_A2_c_576_n N_S1_c_621_n 0.00874089f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_473 N_A2_c_577_n N_S1_c_621_n 0.00122824f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_474 N_A2_M1019_g N_VPWR_c_926_n 0.00694328f $X=5.435 $Y=2.275 $X2=0 $Y2=0
cc_475 N_A2_M1019_g N_VPWR_c_927_n 0.00190345f $X=5.435 $Y=2.275 $X2=0 $Y2=0
cc_476 N_A2_M1019_g N_VPWR_c_932_n 0.00339367f $X=5.435 $Y=2.275 $X2=0 $Y2=0
cc_477 N_A2_M1019_g N_VPWR_c_923_n 0.00505257f $X=5.435 $Y=2.275 $X2=0 $Y2=0
cc_478 N_A2_M1024_g N_A_277_47#_c_1064_n 0.00207269f $X=5.445 $Y=0.445 $X2=0
+ $Y2=0
cc_479 N_A2_c_576_n N_A_277_47#_c_1064_n 0.0029949f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_480 N_A2_c_577_n N_A_277_47#_c_1064_n 0.00828149f $X=5.495 $Y=1.22 $X2=0
+ $Y2=0
cc_481 N_A2_M1019_g N_A_757_363#_c_1231_n 0.0121453f $X=5.435 $Y=2.275 $X2=0
+ $Y2=0
cc_482 N_A2_c_576_n N_A_757_363#_c_1231_n 0.00133384f $X=5.495 $Y=1.22 $X2=0
+ $Y2=0
cc_483 N_A2_c_577_n N_A_757_363#_c_1231_n 0.0154002f $X=5.495 $Y=1.22 $X2=0
+ $Y2=0
cc_484 N_A2_M1019_g N_A_750_97#_c_1294_n 0.00397048f $X=5.435 $Y=2.275 $X2=0
+ $Y2=0
cc_485 N_A2_c_576_n N_A_750_97#_c_1294_n 0.00104503f $X=5.495 $Y=1.22 $X2=0
+ $Y2=0
cc_486 N_A2_c_577_n N_A_750_97#_c_1294_n 0.0088926f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_487 N_A2_M1024_g N_VGND_c_1483_n 0.00268723f $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_488 N_A2_M1024_g N_VGND_c_1484_n 0.00326758f $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_489 N_A2_M1024_g N_VGND_c_1490_n 0.00426187f $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_490 N_A2_M1024_g N_VGND_c_1493_n 0.00685926f $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_491 N_A2_M1024_g N_A_834_97#_c_1638_n 0.011679f $X=5.445 $Y=0.445 $X2=0 $Y2=0
cc_492 N_A2_c_576_n N_A_834_97#_c_1638_n 0.00340435f $X=5.495 $Y=1.22 $X2=0
+ $Y2=0
cc_493 N_A2_c_577_n N_A_834_97#_c_1638_n 0.022595f $X=5.495 $Y=1.22 $X2=0 $Y2=0
cc_494 N_A2_M1024_g N_A_834_97#_c_1639_n 0.00685241f $X=5.445 $Y=0.445 $X2=0
+ $Y2=0
cc_495 N_S1_M1001_g N_A_1290_413#_M1003_g 0.0366051f $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_496 N_S1_M1005_g N_A_1290_413#_c_697_n 0.00746374f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_497 N_S1_c_620_n N_A_1290_413#_c_698_n 0.0133929f $X=7.32 $Y=1.162 $X2=0
+ $Y2=0
cc_498 N_S1_M1015_g N_A_1290_413#_c_699_n 0.0125239f $X=6.385 $Y=0.445 $X2=0
+ $Y2=0
cc_499 N_S1_c_618_n N_A_1290_413#_c_699_n 0.00821217f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_500 S1 N_A_1290_413#_c_699_n 0.00757716f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_501 N_S1_M1009_g N_A_1290_413#_c_706_n 0.023837f $X=6.375 $Y=2.275 $X2=0
+ $Y2=0
cc_502 N_S1_c_618_n N_A_1290_413#_c_706_n 0.00595074f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_503 S1 N_A_1290_413#_c_706_n 0.0294324f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_504 N_S1_M1005_g N_A_1290_413#_c_718_n 0.00392615f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_505 N_S1_c_618_n N_A_1290_413#_c_700_n 0.00376716f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_506 N_S1_c_620_n N_A_1290_413#_c_700_n 0.0038942f $X=7.32 $Y=1.162 $X2=0
+ $Y2=0
cc_507 N_S1_c_618_n N_A_1290_413#_c_721_n 0.00319316f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_508 S1 N_A_1290_413#_c_721_n 0.00139444f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_509 N_S1_c_618_n N_A_1290_413#_c_723_n 0.0130333f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_510 S1 N_A_1290_413#_c_723_n 0.0114761f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_511 N_S1_M1001_g N_A_1478_413#_c_811_n 0.00308722f $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_512 N_S1_M1005_g N_A_1478_413#_c_813_n 0.00195037f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_513 N_S1_M1009_g N_VPWR_c_927_n 0.00983056f $X=6.375 $Y=2.275 $X2=0 $Y2=0
cc_514 S1 N_VPWR_c_927_n 0.00364539f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_515 N_S1_M1009_g N_VPWR_c_933_n 0.0046653f $X=6.375 $Y=2.275 $X2=0 $Y2=0
cc_516 N_S1_M1001_g N_VPWR_c_933_n 0.00539883f $X=7.315 $Y=2.275 $X2=0 $Y2=0
cc_517 N_S1_M1009_g N_VPWR_c_923_n 0.00571875f $X=6.375 $Y=2.275 $X2=0 $Y2=0
cc_518 N_S1_M1001_g N_VPWR_c_923_n 0.00761208f $X=7.315 $Y=2.275 $X2=0 $Y2=0
cc_519 N_S1_c_618_n N_A_277_47#_c_1063_n 0.0211849f $X=7.24 $Y=1.162 $X2=0 $Y2=0
cc_520 N_S1_M1001_g N_A_277_47#_c_1063_n 0.0190088f $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_521 N_S1_M1005_g N_A_277_47#_c_1063_n 0.0012803f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_522 N_S1_M1015_g N_A_277_47#_c_1064_n 0.012491f $X=6.385 $Y=0.445 $X2=0 $Y2=0
cc_523 N_S1_c_618_n N_A_277_47#_c_1064_n 0.00471169f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_524 S1 N_A_277_47#_c_1064_n 0.0102478f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_525 N_S1_c_621_n N_A_277_47#_c_1064_n 0.00782676f $X=6.46 $Y=1.16 $X2=0 $Y2=0
cc_526 N_S1_M1005_g N_A_277_47#_c_1066_n 0.00211374f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_527 N_S1_c_618_n N_A_277_47#_c_1067_n 2.22056e-19 $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_528 N_S1_M1005_g N_A_277_47#_c_1067_n 0.0045786f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_529 N_S1_c_618_n N_A_277_47#_c_1068_n 4.35966e-19 $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_530 N_S1_M1005_g N_A_277_47#_c_1068_n 0.00337688f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_531 N_S1_M1005_g N_A_277_47#_c_1070_n 2.5916e-19 $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_532 N_S1_M1009_g N_A_757_363#_c_1231_n 0.00429839f $X=6.375 $Y=2.275 $X2=0
+ $Y2=0
cc_533 N_S1_M1009_g N_A_757_363#_c_1251_n 0.00260065f $X=6.375 $Y=2.275 $X2=0
+ $Y2=0
cc_534 N_S1_M1005_g N_A_750_97#_c_1334_n 0.00907316f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_535 N_S1_M1001_g N_A_750_97#_c_1286_n 0.00419445f $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_536 N_S1_M1005_g N_A_750_97#_c_1286_n 0.0135832f $X=7.325 $Y=0.445 $X2=0
+ $Y2=0
cc_537 N_S1_c_620_n N_A_750_97#_c_1286_n 0.00862266f $X=7.32 $Y=1.162 $X2=0
+ $Y2=0
cc_538 N_S1_M1015_g N_A_750_97#_c_1338_n 0.00177555f $X=6.385 $Y=0.445 $X2=0
+ $Y2=0
cc_539 N_S1_c_618_n N_A_750_97#_c_1338_n 5.48304e-19 $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_540 N_S1_M1001_g N_A_750_97#_c_1291_n 0.00234697f $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_541 N_S1_M1001_g N_A_750_97#_c_1292_n 7.85391e-19 $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_542 N_S1_M1009_g N_A_750_97#_c_1294_n 0.012239f $X=6.375 $Y=2.275 $X2=0 $Y2=0
cc_543 N_S1_c_618_n N_A_750_97#_c_1294_n 0.00408442f $X=7.24 $Y=1.162 $X2=0
+ $Y2=0
cc_544 N_S1_M1001_g N_A_750_97#_c_1294_n 0.00728345f $X=7.315 $Y=2.275 $X2=0
+ $Y2=0
cc_545 S1 N_A_750_97#_c_1294_n 0.0103038f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_546 N_S1_c_621_n N_A_750_97#_c_1294_n 0.00100909f $X=6.46 $Y=1.16 $X2=0 $Y2=0
cc_547 N_S1_M1015_g N_VGND_c_1484_n 0.0120496f $X=6.385 $Y=0.445 $X2=0 $Y2=0
cc_548 S1 N_VGND_c_1484_n 0.00382302f $X=6.175 $Y=1.105 $X2=0 $Y2=0
cc_549 N_S1_c_621_n N_VGND_c_1484_n 0.0056914f $X=6.46 $Y=1.16 $X2=0 $Y2=0
cc_550 N_S1_M1015_g N_VGND_c_1491_n 0.0046653f $X=6.385 $Y=0.445 $X2=0 $Y2=0
cc_551 N_S1_M1005_g N_VGND_c_1491_n 0.00389055f $X=7.325 $Y=0.445 $X2=0 $Y2=0
cc_552 N_S1_M1015_g N_VGND_c_1493_n 0.00581646f $X=6.385 $Y=0.445 $X2=0 $Y2=0
cc_553 N_S1_M1005_g N_VGND_c_1493_n 0.00728031f $X=7.325 $Y=0.445 $X2=0 $Y2=0
cc_554 N_S1_M1015_g N_A_834_97#_c_1638_n 0.0033094f $X=6.385 $Y=0.445 $X2=0
+ $Y2=0
cc_555 N_S1_M1015_g N_A_834_97#_c_1639_n 0.00465666f $X=6.385 $Y=0.445 $X2=0
+ $Y2=0
cc_556 N_A_1290_413#_M1003_g N_A_1478_413#_c_805_n 0.0126095f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_557 N_A_1290_413#_c_697_n N_A_1478_413#_c_797_n 0.0124643f $X=8.09 $Y=1.055
+ $X2=0 $Y2=0
cc_558 N_A_1290_413#_c_703_n N_A_1478_413#_c_797_n 0.00332368f $X=8.355 $Y=1.19
+ $X2=0 $Y2=0
cc_559 N_A_1290_413#_M1003_g N_A_1478_413#_c_806_n 0.00303767f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_560 N_A_1290_413#_c_697_n N_A_1478_413#_c_798_n 0.00293873f $X=8.09 $Y=1.055
+ $X2=0 $Y2=0
cc_561 N_A_1290_413#_c_701_n N_A_1478_413#_c_807_n 0.00235591f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_562 N_A_1290_413#_M1003_g N_A_1478_413#_c_808_n 0.00267877f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_563 N_A_1290_413#_c_701_n N_A_1478_413#_c_808_n 0.00428389f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_564 N_A_1290_413#_c_702_n N_A_1478_413#_c_808_n 0.00517385f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_565 N_A_1290_413#_c_703_n N_A_1478_413#_c_808_n 9.37022e-19 $X=8.355 $Y=1.19
+ $X2=0 $Y2=0
cc_566 N_A_1290_413#_c_701_n N_A_1478_413#_c_800_n 0.00578808f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_567 N_A_1290_413#_c_702_n N_A_1478_413#_c_800_n 0.00501793f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_568 N_A_1290_413#_c_701_n N_A_1478_413#_c_801_n 0.00775382f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_569 N_A_1290_413#_c_702_n N_A_1478_413#_c_801_n 0.00565031f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_570 N_A_1290_413#_c_703_n N_A_1478_413#_c_801_n 7.08169e-19 $X=8.355 $Y=1.19
+ $X2=0 $Y2=0
cc_571 N_A_1290_413#_c_701_n N_A_1478_413#_c_802_n 0.00437988f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_572 N_A_1290_413#_c_702_n N_A_1478_413#_c_802_n 0.00122539f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_573 N_A_1290_413#_c_703_n N_A_1478_413#_c_802_n 0.00886286f $X=8.355 $Y=1.19
+ $X2=0 $Y2=0
cc_574 N_A_1290_413#_M1003_g N_A_1478_413#_c_811_n 0.00111553f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_575 N_A_1290_413#_c_697_n N_A_1478_413#_c_813_n 0.00283078f $X=8.09 $Y=1.055
+ $X2=0 $Y2=0
cc_576 N_A_1290_413#_c_698_n N_A_1478_413#_c_813_n 0.00347588f $X=8.165 $Y=1.19
+ $X2=0 $Y2=0
cc_577 N_A_1290_413#_M1003_g N_VPWR_c_933_n 0.00357877f $X=7.8 $Y=2.04 $X2=0
+ $Y2=0
cc_578 N_A_1290_413#_c_747_p N_VPWR_c_933_n 0.0126313f $X=6.585 $Y=2.3 $X2=0
+ $Y2=0
cc_579 N_A_1290_413#_M1009_d N_VPWR_c_923_n 0.00231546f $X=6.45 $Y=2.065 $X2=0
+ $Y2=0
cc_580 N_A_1290_413#_M1003_g N_VPWR_c_923_n 0.00677725f $X=7.8 $Y=2.04 $X2=0
+ $Y2=0
cc_581 N_A_1290_413#_c_747_p N_VPWR_c_923_n 0.00334754f $X=6.585 $Y=2.3 $X2=0
+ $Y2=0
cc_582 N_A_1290_413#_c_747_p N_A_277_47#_c_1142_n 0.0290155f $X=6.585 $Y=2.3
+ $X2=0 $Y2=0
cc_583 N_A_1290_413#_c_706_n N_A_277_47#_c_1063_n 0.0290155f $X=6.592 $Y=2.135
+ $X2=0 $Y2=0
cc_584 N_A_1290_413#_c_700_n N_A_277_47#_c_1063_n 0.0127356f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_585 N_A_1290_413#_c_721_n N_A_277_47#_c_1063_n 0.00246125f $X=6.865 $Y=1.19
+ $X2=0 $Y2=0
cc_586 N_A_1290_413#_c_723_n N_A_277_47#_c_1063_n 0.0104926f $X=6.72 $Y=1.19
+ $X2=0 $Y2=0
cc_587 N_A_1290_413#_c_699_n N_A_277_47#_c_1064_n 0.0161147f $X=6.6 $Y=1.105
+ $X2=0 $Y2=0
cc_588 N_A_1290_413#_c_700_n N_A_277_47#_c_1064_n 0.0101537f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_589 N_A_1290_413#_c_721_n N_A_277_47#_c_1064_n 0.0265663f $X=6.865 $Y=1.19
+ $X2=0 $Y2=0
cc_590 N_A_1290_413#_c_723_n N_A_277_47#_c_1064_n 0.0020644f $X=6.72 $Y=1.19
+ $X2=0 $Y2=0
cc_591 N_A_1290_413#_c_698_n N_A_277_47#_c_1066_n 9.26818e-19 $X=8.165 $Y=1.19
+ $X2=0 $Y2=0
cc_592 N_A_1290_413#_c_700_n N_A_277_47#_c_1066_n 0.0507053f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_593 N_A_1290_413#_c_699_n N_A_277_47#_c_1067_n 0.00169288f $X=6.6 $Y=1.105
+ $X2=0 $Y2=0
cc_594 N_A_1290_413#_c_700_n N_A_277_47#_c_1067_n 0.0260895f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_595 N_A_1290_413#_c_699_n N_A_277_47#_c_1068_n 0.0143668f $X=6.6 $Y=1.105
+ $X2=0 $Y2=0
cc_596 N_A_1290_413#_c_700_n N_A_277_47#_c_1068_n 4.61094e-19 $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_597 N_A_1290_413#_c_697_n N_A_277_47#_c_1069_n 0.00339231f $X=8.09 $Y=1.055
+ $X2=0 $Y2=0
cc_598 N_A_1290_413#_c_698_n N_A_277_47#_c_1069_n 5.16123e-19 $X=8.165 $Y=1.19
+ $X2=0 $Y2=0
cc_599 N_A_1290_413#_c_700_n N_A_277_47#_c_1069_n 0.0274791f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_600 N_A_1290_413#_c_703_n N_A_277_47#_c_1069_n 5.13169e-19 $X=8.355 $Y=1.19
+ $X2=0 $Y2=0
cc_601 N_A_1290_413#_c_697_n N_A_277_47#_c_1070_n 0.01007f $X=8.09 $Y=1.055
+ $X2=0 $Y2=0
cc_602 N_A_1290_413#_c_698_n N_A_277_47#_c_1070_n 0.00108071f $X=8.165 $Y=1.19
+ $X2=0 $Y2=0
cc_603 N_A_1290_413#_c_700_n N_A_277_47#_c_1070_n 0.00404564f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_604 N_A_1290_413#_c_702_n N_A_277_47#_c_1070_n 0.0132318f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_605 N_A_1290_413#_c_703_n N_A_277_47#_c_1070_n 0.0053863f $X=8.355 $Y=1.19
+ $X2=0 $Y2=0
cc_606 N_A_1290_413#_c_697_n N_A_750_97#_c_1286_n 0.00531349f $X=8.09 $Y=1.055
+ $X2=0 $Y2=0
cc_607 N_A_1290_413#_c_698_n N_A_750_97#_c_1286_n 0.0112934f $X=8.165 $Y=1.19
+ $X2=0 $Y2=0
cc_608 N_A_1290_413#_c_700_n N_A_750_97#_c_1286_n 0.0151935f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_609 N_A_1290_413#_c_702_n N_A_750_97#_c_1286_n 0.00258915f $X=8.56 $Y=1.19
+ $X2=0 $Y2=0
cc_610 N_A_1290_413#_c_718_n N_A_750_97#_c_1338_n 0.0112497f $X=6.595 $Y=0.49
+ $X2=0 $Y2=0
cc_611 N_A_1290_413#_M1003_g N_A_750_97#_c_1292_n 0.00687788f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_612 N_A_1290_413#_c_698_n N_A_750_97#_c_1292_n 0.00939747f $X=8.165 $Y=1.19
+ $X2=0 $Y2=0
cc_613 N_A_1290_413#_c_700_n N_A_750_97#_c_1292_n 0.0106042f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_614 N_A_1290_413#_M1003_g N_A_750_97#_c_1293_n 0.0109887f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_615 N_A_1290_413#_c_700_n N_A_750_97#_c_1293_n 0.00338754f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_616 N_A_1290_413#_c_747_p N_A_750_97#_c_1294_n 4.63669e-19 $X=6.585 $Y=2.3
+ $X2=0 $Y2=0
cc_617 N_A_1290_413#_c_706_n N_A_750_97#_c_1294_n 0.0181776f $X=6.592 $Y=2.135
+ $X2=0 $Y2=0
cc_618 N_A_1290_413#_c_700_n N_A_750_97#_c_1294_n 0.0270737f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_619 N_A_1290_413#_c_721_n N_A_750_97#_c_1294_n 0.0140097f $X=6.865 $Y=1.19
+ $X2=0 $Y2=0
cc_620 N_A_1290_413#_c_723_n N_A_750_97#_c_1294_n 0.00159146f $X=6.72 $Y=1.19
+ $X2=0 $Y2=0
cc_621 N_A_1290_413#_M1003_g N_A_750_97#_c_1295_n 0.00155484f $X=7.8 $Y=2.04
+ $X2=0 $Y2=0
cc_622 N_A_1290_413#_c_700_n N_A_750_97#_c_1295_n 0.0146458f $X=8.415 $Y=1.19
+ $X2=0 $Y2=0
cc_623 N_A_1290_413#_c_697_n N_VGND_c_1491_n 0.00357877f $X=8.09 $Y=1.055 $X2=0
+ $Y2=0
cc_624 N_A_1290_413#_c_718_n N_VGND_c_1491_n 0.00823101f $X=6.595 $Y=0.49 $X2=0
+ $Y2=0
cc_625 N_A_1290_413#_M1015_d N_VGND_c_1493_n 0.00243204f $X=6.46 $Y=0.235 $X2=0
+ $Y2=0
cc_626 N_A_1290_413#_c_697_n N_VGND_c_1493_n 0.00722627f $X=8.09 $Y=1.055 $X2=0
+ $Y2=0
cc_627 N_A_1290_413#_c_718_n N_VGND_c_1493_n 0.00305688f $X=6.595 $Y=0.49 $X2=0
+ $Y2=0
cc_628 N_A_1478_413#_c_807_n N_VPWR_M1016_s 0.00643848f $X=8.955 $Y=1.75 $X2=0
+ $Y2=0
cc_629 N_A_1478_413#_c_801_n N_VPWR_M1016_s 0.00682984f $X=9.04 $Y=1.16 $X2=0
+ $Y2=0
cc_630 N_A_1478_413#_M1016_g N_VPWR_c_928_n 0.0101988f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_631 N_A_1478_413#_c_805_n N_VPWR_c_928_n 0.0150383f $X=8.475 $Y=2.38 $X2=0
+ $Y2=0
cc_632 N_A_1478_413#_c_806_n N_VPWR_c_928_n 0.00313373f $X=8.56 $Y=2.295 $X2=0
+ $Y2=0
cc_633 N_A_1478_413#_c_807_n N_VPWR_c_928_n 0.0108139f $X=8.955 $Y=1.75 $X2=0
+ $Y2=0
cc_634 N_A_1478_413#_c_805_n N_VPWR_c_933_n 0.0121882f $X=8.475 $Y=2.38 $X2=0
+ $Y2=0
cc_635 N_A_1478_413#_c_811_n N_VPWR_c_933_n 0.0696014f $X=7.69 $Y=2.36 $X2=0
+ $Y2=0
cc_636 N_A_1478_413#_M1016_g N_VPWR_c_934_n 0.0046653f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_637 N_A_1478_413#_M1001_d N_VPWR_c_923_n 0.00167498f $X=7.39 $Y=2.065 $X2=0
+ $Y2=0
cc_638 N_A_1478_413#_M1016_g N_VPWR_c_923_n 0.008846f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_639 N_A_1478_413#_c_805_n N_VPWR_c_923_n 0.006547f $X=8.475 $Y=2.38 $X2=0
+ $Y2=0
cc_640 N_A_1478_413#_c_811_n N_VPWR_c_923_n 0.0321333f $X=7.69 $Y=2.36 $X2=0
+ $Y2=0
cc_641 N_A_1478_413#_M1005_d N_A_277_47#_c_1066_n 0.00148146f $X=7.4 $Y=0.235
+ $X2=0 $Y2=0
cc_642 N_A_1478_413#_c_797_n N_A_277_47#_c_1066_n 2.43387e-19 $X=8.555 $Y=0.34
+ $X2=0 $Y2=0
cc_643 N_A_1478_413#_c_813_n N_A_277_47#_c_1066_n 0.00556402f $X=7.815 $Y=0.42
+ $X2=0 $Y2=0
cc_644 N_A_1478_413#_M1005_d N_A_277_47#_c_1069_n 0.00128971f $X=7.4 $Y=0.235
+ $X2=0 $Y2=0
cc_645 N_A_1478_413#_c_797_n N_A_277_47#_c_1069_n 0.00369139f $X=8.555 $Y=0.34
+ $X2=0 $Y2=0
cc_646 N_A_1478_413#_c_800_n N_A_277_47#_c_1069_n 6.35163e-19 $X=8.725 $Y=0.8
+ $X2=0 $Y2=0
cc_647 N_A_1478_413#_c_797_n N_A_277_47#_c_1070_n 0.0186252f $X=8.555 $Y=0.34
+ $X2=0 $Y2=0
cc_648 N_A_1478_413#_c_798_n N_A_277_47#_c_1070_n 0.00890264f $X=8.64 $Y=0.715
+ $X2=0 $Y2=0
cc_649 N_A_1478_413#_c_800_n N_A_277_47#_c_1070_n 0.0138488f $X=8.725 $Y=0.8
+ $X2=0 $Y2=0
cc_650 N_A_1478_413#_c_801_n N_A_277_47#_c_1070_n 0.00169236f $X=9.04 $Y=1.16
+ $X2=0 $Y2=0
cc_651 N_A_1478_413#_c_806_n N_A_750_97#_M1003_d 0.00658385f $X=8.56 $Y=2.295
+ $X2=0 $Y2=0
cc_652 N_A_1478_413#_M1005_d N_A_750_97#_c_1334_n 0.0029748f $X=7.4 $Y=0.235
+ $X2=0 $Y2=0
cc_653 N_A_1478_413#_c_813_n N_A_750_97#_c_1334_n 0.0131522f $X=7.815 $Y=0.42
+ $X2=0 $Y2=0
cc_654 N_A_1478_413#_M1005_d N_A_750_97#_c_1286_n 0.00113817f $X=7.4 $Y=0.235
+ $X2=0 $Y2=0
cc_655 N_A_1478_413#_M1001_d N_A_750_97#_c_1291_n 0.00155728f $X=7.39 $Y=2.065
+ $X2=0 $Y2=0
cc_656 N_A_1478_413#_c_811_n N_A_750_97#_c_1291_n 0.00640458f $X=7.69 $Y=2.36
+ $X2=0 $Y2=0
cc_657 N_A_1478_413#_c_805_n N_A_750_97#_c_1292_n 0.0220258f $X=8.475 $Y=2.38
+ $X2=0 $Y2=0
cc_658 N_A_1478_413#_c_806_n N_A_750_97#_c_1292_n 0.0145729f $X=8.56 $Y=2.295
+ $X2=0 $Y2=0
cc_659 N_A_1478_413#_c_808_n N_A_750_97#_c_1292_n 0.00472949f $X=8.645 $Y=1.75
+ $X2=0 $Y2=0
cc_660 N_A_1478_413#_M1001_d N_A_750_97#_c_1293_n 7.77934e-19 $X=7.39 $Y=2.065
+ $X2=0 $Y2=0
cc_661 N_A_1478_413#_c_805_n N_A_750_97#_c_1293_n 0.00499274f $X=8.475 $Y=2.38
+ $X2=0 $Y2=0
cc_662 N_A_1478_413#_c_811_n N_A_750_97#_c_1293_n 0.00501044f $X=7.69 $Y=2.36
+ $X2=0 $Y2=0
cc_663 N_A_1478_413#_c_811_n N_A_750_97#_c_1294_n 0.00111916f $X=7.69 $Y=2.36
+ $X2=0 $Y2=0
cc_664 N_A_1478_413#_M1001_d N_A_750_97#_c_1295_n 0.00129512f $X=7.39 $Y=2.065
+ $X2=0 $Y2=0
cc_665 N_A_1478_413#_c_805_n N_A_750_97#_c_1295_n 8.49371e-19 $X=8.475 $Y=2.38
+ $X2=0 $Y2=0
cc_666 N_A_1478_413#_c_811_n N_A_750_97#_c_1295_n 0.0016832f $X=7.69 $Y=2.36
+ $X2=0 $Y2=0
cc_667 N_A_1478_413#_c_801_n N_X_c_1428_n 0.0456935f $X=9.04 $Y=1.16 $X2=0 $Y2=0
cc_668 N_A_1478_413#_c_803_n N_X_c_1428_n 0.0321632f $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_669 N_A_1478_413#_c_799_n N_VGND_M1020_s 0.00508641f $X=8.955 $Y=0.8 $X2=0
+ $Y2=0
cc_670 N_A_1478_413#_c_797_n N_VGND_c_1485_n 0.0141315f $X=8.555 $Y=0.34 $X2=0
+ $Y2=0
cc_671 N_A_1478_413#_c_798_n N_VGND_c_1485_n 0.00883814f $X=8.64 $Y=0.715 $X2=0
+ $Y2=0
cc_672 N_A_1478_413#_c_799_n N_VGND_c_1485_n 0.0134567f $X=8.955 $Y=0.8 $X2=0
+ $Y2=0
cc_673 N_A_1478_413#_c_802_n N_VGND_c_1485_n 5.67641e-19 $X=9.04 $Y=1.16 $X2=0
+ $Y2=0
cc_674 N_A_1478_413#_c_803_n N_VGND_c_1485_n 0.00438629f $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_675 N_A_1478_413#_c_797_n N_VGND_c_1491_n 0.0538095f $X=8.555 $Y=0.34 $X2=0
+ $Y2=0
cc_676 N_A_1478_413#_c_799_n N_VGND_c_1491_n 0.00259545f $X=8.955 $Y=0.8 $X2=0
+ $Y2=0
cc_677 N_A_1478_413#_c_813_n N_VGND_c_1491_n 0.0112187f $X=7.815 $Y=0.42 $X2=0
+ $Y2=0
cc_678 N_A_1478_413#_c_799_n N_VGND_c_1492_n 5.41497e-19 $X=8.955 $Y=0.8 $X2=0
+ $Y2=0
cc_679 N_A_1478_413#_c_803_n N_VGND_c_1492_n 0.00575449f $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_680 N_A_1478_413#_M1005_d N_VGND_c_1493_n 0.00501753f $X=7.4 $Y=0.235 $X2=0
+ $Y2=0
cc_681 N_A_1478_413#_c_797_n N_VGND_c_1493_n 0.0243252f $X=8.555 $Y=0.34 $X2=0
+ $Y2=0
cc_682 N_A_1478_413#_c_799_n N_VGND_c_1493_n 0.0068784f $X=8.955 $Y=0.8 $X2=0
+ $Y2=0
cc_683 N_A_1478_413#_c_813_n N_VGND_c_1493_n 0.00296679f $X=7.815 $Y=0.42 $X2=0
+ $Y2=0
cc_684 N_A_1478_413#_c_803_n N_VGND_c_1493_n 0.012533f $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_685 N_A_27_413#_c_893_n N_VPWR_c_924_n 0.0126961f $X=1.535 $Y=1.88 $X2=0
+ $Y2=0
cc_686 N_A_27_413#_c_892_n N_VPWR_c_929_n 0.0115924f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_687 N_A_27_413#_c_893_n N_VPWR_c_929_n 0.00221328f $X=1.535 $Y=1.88 $X2=0
+ $Y2=0
cc_688 N_A_27_413#_c_893_n N_VPWR_c_930_n 0.00224929f $X=1.535 $Y=1.88 $X2=0
+ $Y2=0
cc_689 N_A_27_413#_M1010_s N_VPWR_c_923_n 0.00377405f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_690 N_A_27_413#_c_892_n N_VPWR_c_923_n 0.00646745f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_691 N_A_27_413#_c_893_n N_VPWR_c_923_n 0.0104103f $X=1.535 $Y=1.88 $X2=0
+ $Y2=0
cc_692 N_A_27_413#_c_893_n N_A_193_413#_c_1038_n 0.0144965f $X=1.535 $Y=1.88
+ $X2=0 $Y2=0
cc_693 N_A_27_413#_c_895_n N_A_193_413#_c_1038_n 0.0121319f $X=1.62 $Y=1.96
+ $X2=0 $Y2=0
cc_694 N_A_27_413#_c_893_n N_A_193_413#_c_1046_n 0.0124642f $X=1.535 $Y=1.88
+ $X2=0 $Y2=0
cc_695 N_A_27_413#_c_895_n N_A_277_47#_c_1072_n 0.00983927f $X=1.62 $Y=1.96
+ $X2=0 $Y2=0
cc_696 N_A_27_413#_c_893_n N_A_277_47#_c_1073_n 0.0105574f $X=1.535 $Y=1.88
+ $X2=0 $Y2=0
cc_697 N_A_27_413#_c_895_n N_A_277_47#_c_1073_n 0.00391032f $X=1.62 $Y=1.96
+ $X2=0 $Y2=0
cc_698 N_A_27_413#_c_895_n N_A_277_47#_c_1074_n 0.00613728f $X=1.62 $Y=1.96
+ $X2=0 $Y2=0
cc_699 N_VPWR_c_923_n N_A_193_413#_M1025_d 0.00235617f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_700 N_VPWR_c_930_n N_A_193_413#_c_1038_n 0.0878972f $X=3.235 $Y=2.72 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_923_n N_A_193_413#_c_1038_n 0.0494983f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_930_n N_A_193_413#_c_1046_n 0.0110309f $X=3.235 $Y=2.72 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_923_n N_A_193_413#_c_1046_n 0.0063548f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_923_n N_A_277_47#_M1001_s 0.00210659f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_705 N_VPWR_c_933_n N_A_277_47#_c_1142_n 0.0143008f $X=8.815 $Y=2.72 $X2=0
+ $Y2=0
cc_706 N_VPWR_c_923_n N_A_277_47#_c_1142_n 0.00378903f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_707 N_VPWR_c_923_n N_A_757_363#_M1019_d 0.00214318f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_925_n N_A_757_363#_c_1227_n 0.00233153f $X=3.4 $Y=2.34 $X2=0
+ $Y2=0
cc_709 N_VPWR_c_926_n N_A_757_363#_c_1228_n 0.0113113f $X=5.225 $Y=2.34 $X2=0
+ $Y2=0
cc_710 N_VPWR_c_931_n N_A_757_363#_c_1228_n 0.0540373f $X=5.06 $Y=2.72 $X2=0
+ $Y2=0
cc_711 N_VPWR_c_923_n N_A_757_363#_c_1228_n 0.0187248f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_712 N_VPWR_c_925_n N_A_757_363#_c_1229_n 0.0111717f $X=3.4 $Y=2.34 $X2=0
+ $Y2=0
cc_713 N_VPWR_c_931_n N_A_757_363#_c_1229_n 0.0121882f $X=5.06 $Y=2.72 $X2=0
+ $Y2=0
cc_714 N_VPWR_c_923_n N_A_757_363#_c_1229_n 0.006547f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_715 N_VPWR_c_926_n N_A_757_363#_c_1230_n 0.00235085f $X=5.225 $Y=2.34 $X2=0
+ $Y2=0
cc_716 N_VPWR_M1004_d N_A_757_363#_c_1231_n 0.00159539f $X=5.09 $Y=2.065 $X2=0
+ $Y2=0
cc_717 N_VPWR_c_926_n N_A_757_363#_c_1231_n 0.0147822f $X=5.225 $Y=2.34 $X2=0
+ $Y2=0
cc_718 N_VPWR_c_931_n N_A_757_363#_c_1231_n 0.00334403f $X=5.06 $Y=2.72 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_932_n N_A_757_363#_c_1231_n 0.00244309f $X=5.98 $Y=2.72 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_923_n N_A_757_363#_c_1231_n 0.00518035f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_721 N_VPWR_c_927_n N_A_757_363#_c_1251_n 0.0124821f $X=6.165 $Y=2.34 $X2=0
+ $Y2=0
cc_722 N_VPWR_c_932_n N_A_757_363#_c_1251_n 0.01143f $X=5.98 $Y=2.72 $X2=0 $Y2=0
cc_723 N_VPWR_c_923_n N_A_757_363#_c_1251_n 0.00304647f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_724 N_VPWR_c_926_n N_A_750_97#_c_1294_n 0.00121475f $X=5.225 $Y=2.34 $X2=0
+ $Y2=0
cc_725 N_VPWR_c_927_n N_A_750_97#_c_1294_n 0.0061602f $X=6.165 $Y=2.34 $X2=0
+ $Y2=0
cc_726 N_VPWR_c_923_n N_A_750_97#_c_1294_n 0.139329f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_727 N_VPWR_c_923_n N_A_750_97#_c_1309_n 0.0148176f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_728 N_VPWR_c_923_n N_A_750_97#_c_1295_n 0.0156335f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_729 N_VPWR_c_923_n A_923_363# 0.00187976f $X=9.43 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_730 N_VPWR_c_923_n N_X_M1016_d 0.00382897f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_731 N_VPWR_c_934_n N_X_c_1428_n 0.018001f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_732 N_VPWR_c_923_n N_X_c_1428_n 0.00993603f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_733 N_A_193_413#_c_1038_n N_A_277_47#_c_1072_n 0.00404715f $X=2.375 $Y=2.38
+ $X2=0 $Y2=0
cc_734 N_A_193_413#_c_1039_n N_A_277_47#_c_1074_n 0.00404507f $X=2.46 $Y=1.96
+ $X2=0 $Y2=0
cc_735 N_A_193_413#_c_1038_n N_A_277_47#_c_1094_n 0.0189439f $X=2.375 $Y=2.38
+ $X2=0 $Y2=0
cc_736 N_A_277_47#_c_1064_n N_A_750_97#_c_1284_n 0.0190611f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_737 N_A_277_47#_c_1066_n N_A_750_97#_c_1334_n 0.00271972f $X=7.91 $Y=0.85
+ $X2=0 $Y2=0
cc_738 N_A_277_47#_c_1067_n N_A_750_97#_c_1334_n 0.0019625f $X=7.28 $Y=0.85
+ $X2=0 $Y2=0
cc_739 N_A_277_47#_c_1063_n N_A_750_97#_c_1286_n 0.0439132f $X=7.085 $Y=2.135
+ $X2=0 $Y2=0
cc_740 N_A_277_47#_c_1066_n N_A_750_97#_c_1286_n 0.0135132f $X=7.91 $Y=0.85
+ $X2=0 $Y2=0
cc_741 N_A_277_47#_c_1067_n N_A_750_97#_c_1286_n 0.00292803f $X=7.28 $Y=0.85
+ $X2=0 $Y2=0
cc_742 N_A_277_47#_c_1068_n N_A_750_97#_c_1286_n 0.0114082f $X=7.135 $Y=0.85
+ $X2=0 $Y2=0
cc_743 N_A_277_47#_c_1069_n N_A_750_97#_c_1286_n 0.00286468f $X=8.055 $Y=0.85
+ $X2=0 $Y2=0
cc_744 N_A_277_47#_c_1070_n N_A_750_97#_c_1286_n 0.00385068f $X=8.055 $Y=0.85
+ $X2=0 $Y2=0
cc_745 N_A_277_47#_c_1067_n N_A_750_97#_c_1338_n 0.00199109f $X=7.28 $Y=0.85
+ $X2=0 $Y2=0
cc_746 N_A_277_47#_c_1068_n N_A_750_97#_c_1338_n 0.0107937f $X=7.135 $Y=0.85
+ $X2=0 $Y2=0
cc_747 N_A_277_47#_c_1063_n N_A_750_97#_c_1291_n 0.0114554f $X=7.085 $Y=2.135
+ $X2=0 $Y2=0
cc_748 N_A_277_47#_c_1142_n N_A_750_97#_c_1294_n 0.00129165f $X=7.105 $Y=2.3
+ $X2=0 $Y2=0
cc_749 N_A_277_47#_c_1063_n N_A_750_97#_c_1294_n 0.0161103f $X=7.085 $Y=2.135
+ $X2=0 $Y2=0
cc_750 N_A_277_47#_c_1063_n N_A_750_97#_c_1295_n 5.19965e-19 $X=7.085 $Y=2.135
+ $X2=0 $Y2=0
cc_751 N_A_277_47#_c_1064_n N_A_27_47#_M1011_d 0.00212372f $X=6.99 $Y=0.85 $X2=0
+ $Y2=0
cc_752 N_A_277_47#_c_1061_n N_A_27_47#_c_1438_n 0.0102283f $X=1.495 $Y=0.935
+ $X2=0 $Y2=0
cc_753 N_A_277_47#_c_1065_n N_A_27_47#_c_1438_n 5.05319e-19 $X=1.76 $Y=0.85
+ $X2=0 $Y2=0
cc_754 N_A_277_47#_M1017_d N_A_27_47#_c_1440_n 0.00404773f $X=1.385 $Y=0.235
+ $X2=0 $Y2=0
cc_755 N_A_277_47#_c_1061_n N_A_27_47#_c_1440_n 0.0173523f $X=1.495 $Y=0.935
+ $X2=0 $Y2=0
cc_756 N_A_277_47#_c_1064_n N_A_27_47#_c_1440_n 0.00341193f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_757 N_A_277_47#_c_1065_n N_A_27_47#_c_1440_n 0.00108867f $X=1.76 $Y=0.85
+ $X2=0 $Y2=0
cc_758 N_A_277_47#_c_1064_n N_A_27_47#_c_1452_n 0.00711651f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_759 N_A_277_47#_c_1065_n N_A_27_47#_c_1452_n 6.25841e-19 $X=1.76 $Y=0.85
+ $X2=0 $Y2=0
cc_760 N_A_277_47#_c_1064_n N_VGND_c_1482_n 0.0136774f $X=6.99 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_A_277_47#_c_1064_n N_VGND_c_1483_n 7.79929e-19 $X=6.99 $Y=0.85 $X2=0
+ $Y2=0
cc_762 N_A_277_47#_c_1064_n N_VGND_c_1484_n 0.00520094f $X=6.99 $Y=0.85 $X2=0
+ $Y2=0
cc_763 N_A_277_47#_M1017_d N_VGND_c_1493_n 0.00173431f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_764 N_A_277_47#_c_1064_n N_VGND_c_1493_n 0.247886f $X=6.99 $Y=0.85 $X2=0
+ $Y2=0
cc_765 N_A_277_47#_c_1065_n N_VGND_c_1493_n 0.0146066f $X=1.76 $Y=0.85 $X2=0
+ $Y2=0
cc_766 N_A_277_47#_c_1066_n N_VGND_c_1493_n 0.0311099f $X=7.91 $Y=0.85 $X2=0
+ $Y2=0
cc_767 N_A_277_47#_c_1067_n N_VGND_c_1493_n 0.0160105f $X=7.28 $Y=0.85 $X2=0
+ $Y2=0
cc_768 N_A_277_47#_c_1068_n N_VGND_c_1493_n 5.77745e-19 $X=7.135 $Y=0.85 $X2=0
+ $Y2=0
cc_769 N_A_277_47#_c_1069_n N_VGND_c_1493_n 0.0157283f $X=8.055 $Y=0.85 $X2=0
+ $Y2=0
cc_770 N_A_277_47#_c_1064_n N_A_668_97#_M1018_s 0.00101014f $X=6.99 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_771 N_A_277_47#_c_1064_n N_A_668_97#_c_1607_n 0.00654267f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_772 N_A_277_47#_c_1064_n N_A_668_97#_c_1609_n 0.0015134f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_773 N_A_277_47#_c_1064_n N_A_668_97#_c_1610_n 0.00802406f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_774 N_A_277_47#_c_1064_n N_A_834_97#_M1022_d 4.01287e-19 $X=6.99 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_775 N_A_277_47#_c_1064_n N_A_834_97#_c_1638_n 0.059044f $X=6.99 $Y=0.85 $X2=0
+ $Y2=0
cc_776 N_A_277_47#_c_1064_n N_A_834_97#_c_1640_n 0.00901372f $X=6.99 $Y=0.85
+ $X2=0 $Y2=0
cc_777 N_A_757_363#_c_1227_n N_A_750_97#_c_1288_n 0.00688205f $X=3.91 $Y=1.96
+ $X2=0 $Y2=0
cc_778 N_A_757_363#_c_1227_n N_A_750_97#_c_1289_n 0.00680993f $X=3.91 $Y=1.96
+ $X2=0 $Y2=0
cc_779 N_A_757_363#_c_1228_n N_A_750_97#_c_1294_n 0.00242959f $X=4.665 $Y=2.38
+ $X2=0 $Y2=0
cc_780 N_A_757_363#_c_1231_n N_A_750_97#_c_1294_n 0.0338788f $X=5.56 $Y=2 $X2=0
+ $Y2=0
cc_781 N_A_757_363#_c_1235_n N_A_750_97#_c_1294_n 0.00899014f $X=4.835 $Y=2
+ $X2=0 $Y2=0
cc_782 N_A_757_363#_c_1227_n N_A_750_97#_c_1309_n 0.00114113f $X=3.91 $Y=1.96
+ $X2=0 $Y2=0
cc_783 N_A_757_363#_c_1228_n N_A_750_97#_c_1309_n 0.0020302f $X=4.665 $Y=2.38
+ $X2=0 $Y2=0
cc_784 N_A_757_363#_c_1235_n N_A_750_97#_c_1309_n 0.00124814f $X=4.835 $Y=2
+ $X2=0 $Y2=0
cc_785 N_A_757_363#_c_1227_n N_A_750_97#_c_1312_n 0.0136858f $X=3.91 $Y=1.96
+ $X2=0 $Y2=0
cc_786 N_A_757_363#_c_1228_n N_A_750_97#_c_1312_n 0.0193407f $X=4.665 $Y=2.38
+ $X2=0 $Y2=0
cc_787 N_A_757_363#_c_1235_n N_A_750_97#_c_1312_n 0.00653226f $X=4.835 $Y=2
+ $X2=0 $Y2=0
cc_788 N_A_757_363#_c_1228_n A_923_363# 0.00340842f $X=4.665 $Y=2.38 $X2=-0.19
+ $Y2=1.305
cc_789 N_A_757_363#_c_1230_n A_923_363# 0.0024545f $X=4.75 $Y=2.295 $X2=-0.19
+ $Y2=1.305
cc_790 N_A_757_363#_c_1231_n A_923_363# 0.00100945f $X=5.56 $Y=2 $X2=-0.19
+ $Y2=1.305
cc_791 N_A_757_363#_c_1235_n A_923_363# 0.00323827f $X=4.835 $Y=2 $X2=-0.19
+ $Y2=1.305
cc_792 N_A_750_97#_c_1294_n A_923_363# 4.09647e-19 $X=7.495 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_793 N_A_750_97#_c_1334_n N_VGND_c_1491_n 0.00996926f $X=7.39 $Y=0.5 $X2=0
+ $Y2=0
cc_794 N_A_750_97#_c_1338_n N_VGND_c_1491_n 0.0110309f $X=7.115 $Y=0.42 $X2=0
+ $Y2=0
cc_795 N_A_750_97#_M1005_s N_VGND_c_1493_n 0.00180769f $X=6.99 $Y=0.235 $X2=0
+ $Y2=0
cc_796 N_A_750_97#_c_1334_n N_VGND_c_1493_n 0.00525789f $X=7.39 $Y=0.5 $X2=0
+ $Y2=0
cc_797 N_A_750_97#_c_1338_n N_VGND_c_1493_n 0.00282232f $X=7.115 $Y=0.42 $X2=0
+ $Y2=0
cc_798 N_A_750_97#_c_1284_n N_A_668_97#_c_1607_n 0.00773981f $X=3.82 $Y=0.92
+ $X2=0 $Y2=0
cc_799 N_A_750_97#_c_1284_n N_A_668_97#_c_1610_n 0.0187718f $X=3.82 $Y=0.92
+ $X2=0 $Y2=0
cc_800 N_A_750_97#_c_1288_n N_A_834_97#_c_1638_n 5.57612e-19 $X=4.165 $Y=1.53
+ $X2=0 $Y2=0
cc_801 N_A_750_97#_c_1284_n N_A_834_97#_c_1640_n 0.0143102f $X=3.82 $Y=0.92
+ $X2=0 $Y2=0
cc_802 N_A_750_97#_c_1285_n N_A_834_97#_c_1640_n 2.20399e-19 $X=3.82 $Y=1.445
+ $X2=0 $Y2=0
cc_803 N_X_c_1428_n N_VGND_c_1492_n 0.018001f $X=9.4 $Y=0.42 $X2=0 $Y2=0
cc_804 N_X_M1020_d N_VGND_c_1493_n 0.00382897f $X=9.265 $Y=0.235 $X2=0 $Y2=0
cc_805 N_X_c_1428_n N_VGND_c_1493_n 0.00993603f $X=9.4 $Y=0.42 $X2=0 $Y2=0
cc_806 N_A_27_47#_c_1438_n N_VGND_M1021_d 0.00159539f $X=1.015 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_807 N_A_27_47#_c_1438_n N_VGND_c_1481_n 0.0159625f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_808 N_A_27_47#_c_1470_p N_VGND_c_1488_n 0.0110686f $X=0.26 $Y=0.425 $X2=0
+ $Y2=0
cc_809 N_A_27_47#_c_1438_n N_VGND_c_1488_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_810 N_A_27_47#_c_1438_n N_VGND_c_1489_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_811 N_A_27_47#_c_1440_n N_VGND_c_1489_n 0.0544788f $X=1.92 $Y=0.34 $X2=0
+ $Y2=0
cc_812 N_A_27_47#_c_1474_p N_VGND_c_1489_n 0.0112984f $X=1.185 $Y=0.34 $X2=0
+ $Y2=0
cc_813 N_A_27_47#_M1021_s N_VGND_c_1493_n 0.00368818f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_814 N_A_27_47#_c_1470_p N_VGND_c_1493_n 0.00641722f $X=0.26 $Y=0.425 $X2=0
+ $Y2=0
cc_815 N_A_27_47#_c_1438_n N_VGND_c_1493_n 0.00988417f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_816 N_A_27_47#_c_1440_n N_VGND_c_1493_n 0.0196628f $X=1.92 $Y=0.34 $X2=0
+ $Y2=0
cc_817 N_A_27_47#_c_1474_p N_VGND_c_1493_n 0.00651108f $X=1.185 $Y=0.34 $X2=0
+ $Y2=0
cc_818 N_A_27_47#_c_1474_p A_193_47# 0.00180745f $X=1.185 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_819 N_VGND_c_1493_n A_193_47# 0.00235053f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_820 N_VGND_c_1493_n N_A_668_97#_M1023_s 0.00172441f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_821 N_VGND_c_1482_n N_A_668_97#_c_1607_n 0.0193861f $X=2.945 $Y=0.64 $X2=0
+ $Y2=0
cc_822 N_VGND_c_1482_n N_A_668_97#_c_1608_n 0.0102674f $X=2.945 $Y=0.64 $X2=0
+ $Y2=0
cc_823 N_VGND_c_1486_n N_A_668_97#_c_1608_n 0.0119809f $X=5.15 $Y=0 $X2=0 $Y2=0
cc_824 N_VGND_c_1493_n N_A_668_97#_c_1608_n 0.00308016f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_825 N_VGND_c_1486_n N_A_668_97#_c_1610_n 0.0894826f $X=5.15 $Y=0 $X2=0 $Y2=0
cc_826 N_VGND_c_1493_n N_A_668_97#_c_1610_n 0.0237524f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_827 N_VGND_c_1493_n N_A_834_97#_M1024_d 0.00206233f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_828 N_VGND_c_1483_n N_A_834_97#_c_1638_n 0.0116663f $X=5.235 $Y=0.38 $X2=0
+ $Y2=0
cc_829 N_VGND_c_1486_n N_A_834_97#_c_1638_n 0.00241057f $X=5.15 $Y=0 $X2=0 $Y2=0
cc_830 N_VGND_c_1490_n N_A_834_97#_c_1638_n 0.00247324f $X=6.01 $Y=0 $X2=0 $Y2=0
cc_831 N_VGND_c_1493_n N_A_834_97#_c_1638_n 0.00528319f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_832 N_VGND_c_1484_n N_A_834_97#_c_1639_n 0.00977026f $X=6.175 $Y=0.38 $X2=0
+ $Y2=0
cc_833 N_VGND_c_1490_n N_A_834_97#_c_1639_n 0.0118607f $X=6.01 $Y=0 $X2=0 $Y2=0
cc_834 N_VGND_c_1493_n N_A_834_97#_c_1639_n 0.00426669f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_835 N_A_668_97#_c_1609_n N_A_834_97#_c_1638_n 0.0146409f $X=4.815 $Y=0.38
+ $X2=0 $Y2=0
cc_836 N_A_668_97#_c_1610_n N_A_834_97#_c_1638_n 0.00907987f $X=4.625 $Y=0.36
+ $X2=0 $Y2=0
cc_837 N_A_668_97#_c_1610_n N_A_834_97#_c_1640_n 0.0114035f $X=4.625 $Y=0.36
+ $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dlclkp_2.pxi.spice
* Created: Tue Sep  1 19:04:37 2020
* 
x_PM_SKY130_FD_SC_HD__DLCLKP_2%CLK N_CLK_c_158_n N_CLK_c_147_n N_CLK_M1018_g
+ N_CLK_c_159_n N_CLK_M1011_g N_CLK_M1001_g N_CLK_M1016_g N_CLK_c_149_n
+ N_CLK_c_161_n CLK N_CLK_c_150_n N_CLK_c_151_n N_CLK_c_152_n N_CLK_c_153_n
+ N_CLK_c_154_n N_CLK_c_155_n N_CLK_c_156_n N_CLK_c_157_n
+ PM_SKY130_FD_SC_HD__DLCLKP_2%CLK
x_PM_SKY130_FD_SC_HD__DLCLKP_2%GATE N_GATE_c_281_n N_GATE_M1015_g N_GATE_c_282_n
+ N_GATE_M1013_g GATE GATE N_GATE_c_287_n PM_SKY130_FD_SC_HD__DLCLKP_2%GATE
x_PM_SKY130_FD_SC_HD__DLCLKP_2%A_193_47# N_A_193_47#_M1012_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1004_g N_A_193_47#_M1005_g N_A_193_47#_c_326_n
+ N_A_193_47#_c_333_n N_A_193_47#_c_327_n N_A_193_47#_c_335_n
+ N_A_193_47#_c_328_n N_A_193_47#_c_329_n N_A_193_47#_c_336_n
+ N_A_193_47#_c_330_n PM_SKY130_FD_SC_HD__DLCLKP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DLCLKP_2%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1011_s
+ N_A_27_47#_c_419_n N_A_27_47#_M1012_g N_A_27_47#_c_420_n N_A_27_47#_M1000_g
+ N_A_27_47#_c_421_n N_A_27_47#_c_422_n N_A_27_47#_c_423_n N_A_27_47#_c_424_n
+ N_A_27_47#_M1003_g N_A_27_47#_c_426_n N_A_27_47#_c_427_n N_A_27_47#_M1020_g
+ N_A_27_47#_c_428_n N_A_27_47#_c_541_p N_A_27_47#_c_429_n N_A_27_47#_c_430_n
+ N_A_27_47#_c_438_n N_A_27_47#_c_439_n N_A_27_47#_c_440_n N_A_27_47#_c_431_n
+ N_A_27_47#_c_432_n N_A_27_47#_c_433_n PM_SKY130_FD_SC_HD__DLCLKP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DLCLKP_2%A_643_307# N_A_643_307#_M1017_d
+ N_A_643_307#_M1019_s N_A_643_307#_M1002_g N_A_643_307#_M1021_g
+ N_A_643_307#_c_554_n N_A_643_307#_M1010_g N_A_643_307#_c_555_n
+ N_A_643_307#_c_556_n N_A_643_307#_M1006_g N_A_643_307#_c_565_n
+ N_A_643_307#_c_639_p N_A_643_307#_c_557_n N_A_643_307#_c_567_n
+ N_A_643_307#_c_558_n N_A_643_307#_c_559_n N_A_643_307#_c_560_n
+ N_A_643_307#_c_568_n PM_SKY130_FD_SC_HD__DLCLKP_2%A_643_307#
x_PM_SKY130_FD_SC_HD__DLCLKP_2%A_477_413# N_A_477_413#_M1003_d
+ N_A_477_413#_M1004_d N_A_477_413#_M1017_g N_A_477_413#_M1019_g
+ N_A_477_413#_c_685_n N_A_477_413#_c_678_n N_A_477_413#_c_672_n
+ N_A_477_413#_c_664_n N_A_477_413#_c_665_n N_A_477_413#_c_666_n
+ N_A_477_413#_c_667_n N_A_477_413#_c_668_n N_A_477_413#_c_669_n
+ N_A_477_413#_c_670_n PM_SKY130_FD_SC_HD__DLCLKP_2%A_477_413#
x_PM_SKY130_FD_SC_HD__DLCLKP_2%A_957_369# N_A_957_369#_M1006_s
+ N_A_957_369#_M1010_d N_A_957_369#_c_754_n N_A_957_369#_M1007_g
+ N_A_957_369#_M1008_g N_A_957_369#_c_755_n N_A_957_369#_M1009_g
+ N_A_957_369#_M1014_g N_A_957_369#_c_756_n N_A_957_369#_c_770_n
+ N_A_957_369#_c_757_n N_A_957_369#_c_758_n N_A_957_369#_c_764_n
+ N_A_957_369#_c_765_n N_A_957_369#_c_759_n N_A_957_369#_c_766_n
+ N_A_957_369#_c_788_n N_A_957_369#_c_760_n N_A_957_369#_c_761_n
+ PM_SKY130_FD_SC_HD__DLCLKP_2%A_957_369#
x_PM_SKY130_FD_SC_HD__DLCLKP_2%VPWR N_VPWR_M1011_d N_VPWR_M1015_s N_VPWR_M1002_d
+ N_VPWR_M1019_d N_VPWR_M1016_d N_VPWR_M1014_d N_VPWR_c_848_n N_VPWR_c_849_n
+ N_VPWR_c_850_n N_VPWR_c_851_n N_VPWR_c_852_n N_VPWR_c_853_n N_VPWR_c_854_n
+ N_VPWR_c_855_n VPWR N_VPWR_c_856_n N_VPWR_c_857_n N_VPWR_c_858_n
+ N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n N_VPWR_c_863_n
+ N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_847_n PM_SKY130_FD_SC_HD__DLCLKP_2%VPWR
x_PM_SKY130_FD_SC_HD__DLCLKP_2%GCLK N_GCLK_M1007_s N_GCLK_M1008_s N_GCLK_c_953_n
+ N_GCLK_c_951_n GCLK GCLK GCLK N_GCLK_c_963_n N_GCLK_c_964_n
+ PM_SKY130_FD_SC_HD__DLCLKP_2%GCLK
x_PM_SKY130_FD_SC_HD__DLCLKP_2%VGND N_VGND_M1018_d N_VGND_M1013_s N_VGND_M1021_d
+ N_VGND_M1001_d N_VGND_M1009_d N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n
+ N_VGND_c_978_n N_VGND_c_979_n N_VGND_c_980_n VGND N_VGND_c_981_n
+ N_VGND_c_982_n N_VGND_c_983_n N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n
+ N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n
+ PM_SKY130_FD_SC_HD__DLCLKP_2%VGND
cc_1 VNB N_CLK_c_147_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_M1001_g 0.0347617f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=0.445
cc_3 VNB N_CLK_c_149_n 0.0236526f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_4 VNB N_CLK_c_150_n 0.0501906f $X=-0.19 $Y=-0.24 $X2=5.15 $Y2=1.19
cc_5 VNB N_CLK_c_151_n 0.00981446f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_6 VNB N_CLK_c_152_n 0.01012f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_7 VNB N_CLK_c_153_n 0.00274722f $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_8 VNB N_CLK_c_154_n 6.94864e-19 $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_9 VNB N_CLK_c_155_n 0.0196229f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_10 VNB N_CLK_c_156_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_11 VNB N_CLK_c_157_n 0.021279f $X=-0.19 $Y=-0.24 $X2=5.32 $Y2=1.27
cc_12 VNB N_GATE_c_281_n 0.0283502f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_13 VNB N_GATE_c_282_n 0.0154525f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_14 VNB GATE 0.0125722f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=1.105
cc_15 VNB N_A_193_47#_M1005_g 0.0212016f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=0.445
cc_16 VNB N_A_193_47#_c_326_n 0.0160308f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=2.165
cc_17 VNB N_A_193_47#_c_327_n 0.00466588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_193_47#_c_328_n 0.00220609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_193_47#_c_329_n 0.00432051f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_20 VNB N_A_193_47#_c_330_n 0.0351767f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_21 VNB N_A_27_47#_c_419_n 0.014637f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_22 VNB N_A_27_47#_c_420_n 0.0125115f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=1.105
cc_23 VNB N_A_27_47#_c_421_n 0.0318145f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=2.165
cc_24 VNB N_A_27_47#_c_422_n 0.0268392f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_25 VNB N_A_27_47#_c_423_n 0.0755917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_424_n 0.00988887f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_27 VNB N_A_27_47#_M1003_g 0.0347402f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_28 VNB N_A_27_47#_c_426_n 0.0177775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_427_n 0.00454503f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_30 VNB N_A_27_47#_c_428_n 0.0052727f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_31 VNB N_A_27_47#_c_429_n 0.00177906f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_32 VNB N_A_27_47#_c_430_n 0.00553431f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_33 VNB N_A_27_47#_c_431_n 7.70731e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_432_n 0.00438392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_433_n 0.0241763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_643_307#_M1021_g 0.0459301f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=0.445
cc_37 VNB N_A_643_307#_c_554_n 0.0417009f $X=-0.19 $Y=-0.24 $X2=5.49 $Y2=1.435
cc_38 VNB N_A_643_307#_c_555_n 0.0278228f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_39 VNB N_A_643_307#_c_556_n 0.0174432f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_40 VNB N_A_643_307#_c_557_n 5.08691e-19 $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_41 VNB N_A_643_307#_c_558_n 0.00430759f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_42 VNB N_A_643_307#_c_559_n 0.00299024f $X=-0.19 $Y=-0.24 $X2=5.32 $Y2=1.27
cc_43 VNB N_A_643_307#_c_560_n 0.00453509f $X=-0.19 $Y=-0.24 $X2=5.375 $Y2=1.435
cc_44 VNB N_A_477_413#_c_664_n 0.00372193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_477_413#_c_665_n 0.00259824f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_46 VNB N_A_477_413#_c_666_n 0.00315607f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_47 VNB N_A_477_413#_c_667_n 0.00682797f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_48 VNB N_A_477_413#_c_668_n 0.0256133f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_49 VNB N_A_477_413#_c_669_n 0.00436469f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_50 VNB N_A_477_413#_c_670_n 0.0201343f $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_51 VNB N_A_957_369#_c_754_n 0.0160981f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_52 VNB N_A_957_369#_c_755_n 0.0215069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_957_369#_c_756_n 7.4909e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_957_369#_c_757_n 0.0126023f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_55 VNB N_A_957_369#_c_758_n 0.0033067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_957_369#_c_759_n 0.00212679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_957_369#_c_760_n 6.0684e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_58 VNB N_A_957_369#_c_761_n 0.0488973f $X=-0.19 $Y=-0.24 $X2=5.32 $Y2=1.27
cc_59 VNB N_VPWR_c_847_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_GCLK_c_951_n 6.42879e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_61 VNB N_VGND_c_975_n 4.16958e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_976_n 0.0099519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_977_n 0.00236436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_978_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_65 VNB N_VGND_c_979_n 0.0104543f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.19
cc_66 VNB N_VGND_c_980_n 0.0345443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_981_n 0.0151256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_982_n 0.0157587f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_69 VNB N_VGND_c_983_n 0.0563377f $X=-0.19 $Y=-0.24 $X2=5.375 $Y2=1.435
cc_70 VNB N_VGND_c_984_n 0.0423061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_985_n 0.0187979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_986_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_987_n 0.00439458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_988_n 0.0035406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_989_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_990_n 0.343507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VPB N_CLK_c_158_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_78 VPB N_CLK_c_159_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_79 VPB N_CLK_M1016_g 0.0378287f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=2.165
cc_80 VPB N_CLK_c_161_n 0.0238508f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_81 VPB N_CLK_c_152_n 0.0153801f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_82 VPB N_CLK_c_153_n 3.42542e-19 $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_83 VPB N_CLK_c_154_n 0.00231958f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_84 VPB N_CLK_c_155_n 0.0107553f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_85 VPB N_CLK_c_157_n 0.0175343f $X=-0.19 $Y=1.305 $X2=5.32 $Y2=1.27
cc_86 VPB N_GATE_c_281_n 0.0321222f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.88
cc_87 VPB N_GATE_M1015_g 0.0227927f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_88 VPB GATE 0.00679153f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=1.105
cc_89 VPB N_GATE_c_287_n 0.00528403f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=2.165
cc_90 VPB N_A_193_47#_M1004_g 0.0219062f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_91 VPB N_A_193_47#_c_326_n 0.0125439f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=2.165
cc_92 VPB N_A_193_47#_c_333_n 0.014084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_93 VPB N_A_193_47#_c_327_n 0.00330024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_193_47#_c_335_n 0.0379744f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_95 VPB N_A_193_47#_c_336_n 0.00726753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_27_47#_M1000_g 0.0415627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_47#_c_426_n 0.0174955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_27_47#_c_427_n 0.00326597f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_99 VPB N_A_27_47#_M1020_g 0.0480975f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.19
cc_100 VPB N_A_27_47#_c_438_n 0.00121249f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_101 VPB N_A_27_47#_c_439_n 0.00647616f $X=-0.19 $Y=1.305 $X2=5.32 $Y2=1.27
cc_102 VPB N_A_27_47#_c_440_n 0.00345702f $X=-0.19 $Y=1.305 $X2=5.375 $Y2=1.435
cc_103 VPB N_A_27_47#_c_431_n 0.00152564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_47#_c_433_n 0.0108291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_643_307#_M1002_g 0.023974f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_106 VPB N_A_643_307#_M1021_g 0.0151639f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=0.445
cc_107 VPB N_A_643_307#_c_554_n 0.00467023f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=1.435
cc_108 VPB N_A_643_307#_M1010_g 0.043187f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=2.165
cc_109 VPB N_A_643_307#_c_565_n 0.00440075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_643_307#_c_557_n 0.00171385f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_111 VPB N_A_643_307#_c_567_n 0.00187855f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_112 VPB N_A_643_307#_c_568_n 0.0476653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_477_413#_M1019_g 0.0232329f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=0.445
cc_114 VPB N_A_477_413#_c_672_n 0.00839419f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_115 VPB N_A_477_413#_c_664_n 0.00291629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_477_413#_c_665_n 2.88203e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_117 VPB N_A_477_413#_c_667_n 0.00225196f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.19
cc_118 VPB N_A_477_413#_c_668_n 0.00617835f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_119 VPB N_A_477_413#_c_669_n 2.00706e-19 $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_120 VPB N_A_957_369#_M1008_g 0.0182514f $X=-0.19 $Y=1.305 $X2=5.49 $Y2=0.445
cc_121 VPB N_A_957_369#_M1014_g 0.0253003f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_122 VPB N_A_957_369#_c_764_n 0.00325238f $X=-0.19 $Y=1.305 $X2=5.15 $Y2=1.19
cc_123 VPB N_A_957_369#_c_765_n 0.00607277f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.19
cc_124 VPB N_A_957_369#_c_766_n 0.00125601f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_125 VPB N_A_957_369#_c_761_n 0.00861025f $X=-0.19 $Y=1.305 $X2=5.32 $Y2=1.27
cc_126 VPB N_VPWR_c_848_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_127 VPB N_VPWR_c_849_n 0.00530537f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_128 VPB N_VPWR_c_850_n 0.00913564f $X=-0.19 $Y=1.305 $X2=5.15 $Y2=1.19
cc_129 VPB N_VPWR_c_851_n 0.0175728f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.19
cc_130 VPB N_VPWR_c_852_n 0.00477384f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_131 VPB N_VPWR_c_853_n 0.00283746f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_132 VPB N_VPWR_c_854_n 0.0104317f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_133 VPB N_VPWR_c_855_n 0.0472986f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_134 VPB N_VPWR_c_856_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.19
cc_135 VPB N_VPWR_c_857_n 0.0155349f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_858_n 0.0400543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_859_n 0.0278771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_860_n 0.0157155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_861_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_862_n 0.00554087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_863_n 0.00574408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_864_n 0.00545601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_865_n 0.00546326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_847_n 0.058381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_GCLK_c_951_n 0.00105438f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_146 N_CLK_c_150_n N_GATE_c_281_n 0.0167008f $X=5.15 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_147 N_CLK_c_150_n GATE 0.0265263f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_148 N_CLK_c_150_n N_GATE_c_287_n 0.015573f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_149 N_CLK_c_150_n N_A_193_47#_c_326_n 0.0314284f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_150 N_CLK_c_150_n N_A_193_47#_c_333_n 0.0138827f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_151 N_CLK_c_150_n N_A_193_47#_c_327_n 0.026832f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_152 N_CLK_c_150_n N_A_193_47#_c_335_n 0.00382482f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_153 N_CLK_c_150_n N_A_193_47#_c_329_n 0.0231277f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_154 N_CLK_c_150_n N_A_193_47#_c_330_n 0.00789047f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_155 N_CLK_c_147_n N_A_27_47#_c_419_n 0.0101063f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_156 N_CLK_c_156_n N_A_27_47#_c_420_n 0.00406396f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_157 N_CLK_c_161_n N_A_27_47#_M1000_g 0.0256048f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_158 N_CLK_c_155_n N_A_27_47#_M1000_g 0.00439288f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_159 N_CLK_c_150_n N_A_27_47#_c_421_n 0.00590074f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_160 N_CLK_c_150_n N_A_27_47#_M1003_g 0.00145143f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_161 N_CLK_c_150_n N_A_27_47#_c_426_n 0.0165582f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_162 N_CLK_c_150_n N_A_27_47#_c_427_n 2.72279e-19 $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_163 N_CLK_c_149_n N_A_27_47#_c_428_n 0.0101063f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_164 N_CLK_c_147_n N_A_27_47#_c_429_n 0.00770412f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_165 N_CLK_c_149_n N_A_27_47#_c_429_n 0.00553647f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_166 N_CLK_c_150_n N_A_27_47#_c_429_n 0.00817564f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_167 N_CLK_c_151_n N_A_27_47#_c_429_n 0.00120578f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_168 N_CLK_c_149_n N_A_27_47#_c_430_n 0.0057713f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_169 N_CLK_c_151_n N_A_27_47#_c_430_n 0.00161409f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_170 N_CLK_c_152_n N_A_27_47#_c_430_n 0.0105869f $X=0.235 $Y=1.19 $X2=0 $Y2=0
cc_171 N_CLK_c_155_n N_A_27_47#_c_430_n 3.38487e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_172 N_CLK_c_159_n N_A_27_47#_c_438_n 0.0107161f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_173 N_CLK_c_161_n N_A_27_47#_c_438_n 0.00220936f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_174 N_CLK_c_150_n N_A_27_47#_c_438_n 0.0067661f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_175 N_CLK_c_151_n N_A_27_47#_c_438_n 0.00108512f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_176 N_CLK_c_158_n N_A_27_47#_c_439_n 8.6641e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_177 N_CLK_c_161_n N_A_27_47#_c_439_n 0.00435948f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_178 N_CLK_c_159_n N_A_27_47#_c_440_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_179 N_CLK_c_161_n N_A_27_47#_c_440_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_180 N_CLK_c_151_n N_A_27_47#_c_440_n 0.00126485f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_181 N_CLK_c_152_n N_A_27_47#_c_440_n 0.0133866f $X=0.235 $Y=1.19 $X2=0 $Y2=0
cc_182 N_CLK_c_155_n N_A_27_47#_c_440_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_183 N_CLK_c_150_n N_A_27_47#_c_431_n 0.0293907f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_184 N_CLK_c_151_n N_A_27_47#_c_431_n 0.00217029f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_185 N_CLK_c_155_n N_A_27_47#_c_431_n 0.00320487f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_186 N_CLK_c_149_n N_A_27_47#_c_432_n 0.00227671f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_187 N_CLK_c_152_n N_A_27_47#_c_432_n 0.0288044f $X=0.235 $Y=1.19 $X2=0 $Y2=0
cc_188 N_CLK_c_156_n N_A_27_47#_c_432_n 0.00146724f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_189 N_CLK_c_150_n N_A_27_47#_c_433_n 0.0137802f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_190 N_CLK_c_151_n N_A_27_47#_c_433_n 4.33045e-19 $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_191 N_CLK_c_152_n N_A_27_47#_c_433_n 9.53587e-19 $X=0.235 $Y=1.19 $X2=0 $Y2=0
cc_192 N_CLK_c_155_n N_A_27_47#_c_433_n 0.0183089f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_193 N_CLK_M1001_g N_A_643_307#_c_554_n 0.00423272f $X=5.49 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_CLK_c_150_n N_A_643_307#_c_554_n 0.00515067f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_195 N_CLK_c_153_n N_A_643_307#_c_554_n 0.00132959f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_196 N_CLK_c_154_n N_A_643_307#_c_554_n 0.00126011f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_197 N_CLK_c_157_n N_A_643_307#_c_554_n 0.0101866f $X=5.32 $Y=1.27 $X2=0 $Y2=0
cc_198 N_CLK_M1016_g N_A_643_307#_M1010_g 0.016147f $X=5.49 $Y=2.165 $X2=0 $Y2=0
cc_199 N_CLK_c_150_n N_A_643_307#_c_555_n 0.0029373f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_200 N_CLK_c_157_n N_A_643_307#_c_555_n 0.00125674f $X=5.32 $Y=1.27 $X2=0
+ $Y2=0
cc_201 N_CLK_M1001_g N_A_643_307#_c_556_n 0.048072f $X=5.49 $Y=0.445 $X2=0 $Y2=0
cc_202 N_CLK_c_150_n N_A_643_307#_c_565_n 0.00312808f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_203 N_CLK_M1016_g N_A_643_307#_c_557_n 4.46469e-19 $X=5.49 $Y=2.165 $X2=0
+ $Y2=0
cc_204 N_CLK_c_150_n N_A_643_307#_c_557_n 0.0257572f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_205 N_CLK_c_153_n N_A_643_307#_c_557_n 0.00111807f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_206 N_CLK_M1016_g N_A_643_307#_c_567_n 9.376e-19 $X=5.49 $Y=2.165 $X2=0 $Y2=0
cc_207 N_CLK_c_150_n N_A_643_307#_c_567_n 0.00836374f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_208 N_CLK_c_150_n N_A_643_307#_c_558_n 0.00121313f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_209 N_CLK_M1001_g N_A_643_307#_c_559_n 4.56376e-19 $X=5.49 $Y=0.445 $X2=0
+ $Y2=0
cc_210 N_CLK_c_150_n N_A_643_307#_c_559_n 0.0239966f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_211 N_CLK_c_153_n N_A_643_307#_c_559_n 0.00150716f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_212 N_CLK_c_154_n N_A_643_307#_c_559_n 0.00767001f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_213 N_CLK_c_157_n N_A_643_307#_c_559_n 0.00117292f $X=5.32 $Y=1.27 $X2=0
+ $Y2=0
cc_214 N_CLK_c_150_n N_A_477_413#_c_678_n 0.00744419f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_215 N_CLK_c_150_n N_A_477_413#_c_664_n 0.0134571f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_216 N_CLK_c_150_n N_A_477_413#_c_665_n 0.0132246f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_217 N_CLK_c_150_n N_A_477_413#_c_667_n 0.0271675f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_218 N_CLK_c_150_n N_A_477_413#_c_668_n 0.00688144f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_219 N_CLK_c_150_n N_A_477_413#_c_669_n 0.0150787f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_220 N_CLK_M1001_g N_A_957_369#_c_754_n 0.0211038f $X=5.49 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_CLK_c_157_n N_A_957_369#_M1008_g 0.0316327f $X=5.32 $Y=1.27 $X2=0 $Y2=0
cc_222 N_CLK_M1016_g N_A_957_369#_c_770_n 0.0111305f $X=5.49 $Y=2.165 $X2=0
+ $Y2=0
cc_223 N_CLK_M1001_g N_A_957_369#_c_757_n 0.014425f $X=5.49 $Y=0.445 $X2=0 $Y2=0
cc_224 N_CLK_c_153_n N_A_957_369#_c_757_n 0.00937027f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_225 N_CLK_c_154_n N_A_957_369#_c_757_n 0.0175451f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_226 N_CLK_c_157_n N_A_957_369#_c_757_n 0.00202596f $X=5.32 $Y=1.27 $X2=0
+ $Y2=0
cc_227 N_CLK_c_150_n N_A_957_369#_c_758_n 0.0113287f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_228 N_CLK_M1016_g N_A_957_369#_c_764_n 0.0159097f $X=5.49 $Y=2.165 $X2=0
+ $Y2=0
cc_229 N_CLK_c_153_n N_A_957_369#_c_764_n 5.38361e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_230 N_CLK_c_154_n N_A_957_369#_c_764_n 0.00638282f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_231 N_CLK_c_157_n N_A_957_369#_c_764_n 4.69573e-19 $X=5.32 $Y=1.27 $X2=0
+ $Y2=0
cc_232 N_CLK_c_150_n N_A_957_369#_c_765_n 0.00553595f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_233 N_CLK_c_153_n N_A_957_369#_c_765_n 0.00337569f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_234 N_CLK_c_154_n N_A_957_369#_c_765_n 0.00631021f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_235 N_CLK_c_157_n N_A_957_369#_c_765_n 0.00197273f $X=5.32 $Y=1.27 $X2=0
+ $Y2=0
cc_236 N_CLK_M1001_g N_A_957_369#_c_759_n 0.00395515f $X=5.49 $Y=0.445 $X2=0
+ $Y2=0
cc_237 N_CLK_c_153_n N_A_957_369#_c_759_n 0.00249539f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_238 N_CLK_c_154_n N_A_957_369#_c_759_n 0.016f $X=5.295 $Y=1.19 $X2=0 $Y2=0
cc_239 N_CLK_M1016_g N_A_957_369#_c_766_n 0.00395515f $X=5.49 $Y=2.165 $X2=0
+ $Y2=0
cc_240 N_CLK_M1001_g N_A_957_369#_c_788_n 0.00212158f $X=5.49 $Y=0.445 $X2=0
+ $Y2=0
cc_241 N_CLK_c_150_n N_A_957_369#_c_788_n 0.0033383f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_242 N_CLK_c_157_n N_A_957_369#_c_760_n 0.00395515f $X=5.32 $Y=1.27 $X2=0
+ $Y2=0
cc_243 N_CLK_M1001_g N_A_957_369#_c_761_n 0.02052f $X=5.49 $Y=0.445 $X2=0 $Y2=0
cc_244 N_CLK_c_154_n N_A_957_369#_c_761_n 2.39322e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_245 N_CLK_c_159_n N_VPWR_c_848_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_246 N_CLK_M1016_g N_VPWR_c_853_n 0.00322532f $X=5.49 $Y=2.165 $X2=0 $Y2=0
cc_247 N_CLK_c_159_n N_VPWR_c_856_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_248 N_CLK_M1016_g N_VPWR_c_859_n 0.00585385f $X=5.49 $Y=2.165 $X2=0 $Y2=0
cc_249 N_CLK_c_159_n N_VPWR_c_847_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_250 N_CLK_M1016_g N_VPWR_c_847_n 0.00695319f $X=5.49 $Y=2.165 $X2=0 $Y2=0
cc_251 N_CLK_c_147_n N_VGND_c_975_n 0.0082568f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_252 N_CLK_c_150_n N_VGND_c_976_n 0.0107817f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_253 N_CLK_c_150_n N_VGND_c_977_n 0.00163791f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_254 N_CLK_M1001_g N_VGND_c_978_n 0.00512205f $X=5.49 $Y=0.445 $X2=0 $Y2=0
cc_255 N_CLK_c_147_n N_VGND_c_981_n 0.00337001f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_256 N_CLK_c_149_n N_VGND_c_981_n 4.4475e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_257 N_CLK_M1001_g N_VGND_c_984_n 0.00585385f $X=5.49 $Y=0.445 $X2=0 $Y2=0
cc_258 N_CLK_c_147_n N_VGND_c_990_n 0.00485988f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_259 N_CLK_M1001_g N_VGND_c_990_n 0.00618632f $X=5.49 $Y=0.445 $X2=0 $Y2=0
cc_260 N_GATE_M1015_g N_A_193_47#_M1004_g 0.0196956f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_261 N_GATE_c_281_n N_A_193_47#_c_326_n 0.00825636f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_262 N_GATE_M1015_g N_A_193_47#_c_326_n 0.00442795f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_263 N_GATE_c_282_n N_A_193_47#_c_326_n 0.00415576f $X=1.91 $Y=1.09 $X2=0
+ $Y2=0
cc_264 N_GATE_c_287_n N_A_193_47#_c_326_n 0.016495f $X=1.985 $Y=1.56 $X2=0 $Y2=0
cc_265 N_GATE_c_281_n N_A_193_47#_c_333_n 0.00256542f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_266 N_GATE_M1015_g N_A_193_47#_c_333_n 0.01366f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_267 GATE N_A_193_47#_c_333_n 0.0186924f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_268 N_GATE_c_287_n N_A_193_47#_c_333_n 0.0284766f $X=1.985 $Y=1.56 $X2=0
+ $Y2=0
cc_269 N_GATE_c_281_n N_A_193_47#_c_327_n 0.00151598f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_270 GATE N_A_193_47#_c_327_n 0.0519273f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_271 N_GATE_c_281_n N_A_193_47#_c_335_n 0.0196956f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_272 GATE N_A_193_47#_c_335_n 8.73251e-19 $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_273 GATE N_A_193_47#_c_328_n 0.0130549f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_274 N_GATE_M1015_g N_A_193_47#_c_336_n 0.00359119f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_275 N_GATE_c_282_n N_A_27_47#_c_422_n 0.0062944f $X=1.91 $Y=1.09 $X2=0 $Y2=0
cc_276 N_GATE_c_282_n N_A_27_47#_c_423_n 0.0104164f $X=1.91 $Y=1.09 $X2=0 $Y2=0
cc_277 GATE N_A_27_47#_c_423_n 0.00557118f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_278 N_GATE_c_281_n N_A_27_47#_M1003_g 0.00293968f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_279 N_GATE_c_282_n N_A_27_47#_M1003_g 0.0177339f $X=1.91 $Y=1.09 $X2=0 $Y2=0
cc_280 GATE N_A_27_47#_M1003_g 0.0167771f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_281 N_GATE_c_281_n N_A_27_47#_c_433_n 0.00324766f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_282 GATE N_A_477_413#_c_678_n 0.00554297f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_283 N_GATE_M1015_g N_VPWR_c_849_n 0.0143344f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_284 N_GATE_M1015_g N_VPWR_c_858_n 0.00245007f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_285 N_GATE_M1015_g N_VPWR_c_847_n 0.00328215f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_286 N_GATE_c_281_n N_VGND_c_976_n 0.00400287f $X=1.83 $Y=1.685 $X2=0 $Y2=0
cc_287 N_GATE_c_282_n N_VGND_c_976_n 0.0012231f $X=1.91 $Y=1.09 $X2=0 $Y2=0
cc_288 GATE N_VGND_c_976_n 0.025038f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_289 N_GATE_c_287_n N_VGND_c_976_n 0.00393464f $X=1.985 $Y=1.56 $X2=0 $Y2=0
cc_290 GATE N_VGND_c_983_n 0.0137319f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_291 N_GATE_c_282_n N_VGND_c_990_n 9.32477e-19 $X=1.91 $Y=1.09 $X2=0 $Y2=0
cc_292 GATE N_VGND_c_990_n 0.00774147f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_293 GATE A_397_119# 0.0141467f $X=1.99 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_294 N_A_193_47#_c_326_n N_A_27_47#_c_419_n 8.4897e-19 $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_295 N_A_193_47#_c_326_n N_A_27_47#_c_420_n 0.0184282f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_296 N_A_193_47#_c_336_n N_A_27_47#_M1000_g 2.19569e-19 $X=1.1 $Y=1.96 $X2=0
+ $Y2=0
cc_297 N_A_193_47#_c_326_n N_A_27_47#_c_421_n 0.0167883f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_298 N_A_193_47#_c_326_n N_A_27_47#_c_422_n 0.00432739f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_299 N_A_193_47#_M1005_g N_A_27_47#_c_423_n 0.0109825f $X=3.185 $Y=0.43 $X2=0
+ $Y2=0
cc_300 N_A_193_47#_c_327_n N_A_27_47#_M1003_g 0.00799435f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_301 N_A_193_47#_c_328_n N_A_27_47#_M1003_g 0.00938487f $X=2.645 $Y=0.9 $X2=0
+ $Y2=0
cc_302 N_A_193_47#_c_330_n N_A_27_47#_M1003_g 0.00902451f $X=3.185 $Y=0.9 $X2=0
+ $Y2=0
cc_303 N_A_193_47#_c_327_n N_A_27_47#_c_426_n 0.00765287f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_304 N_A_193_47#_c_329_n N_A_27_47#_c_426_n 0.00751138f $X=3.06 $Y=0.9 $X2=0
+ $Y2=0
cc_305 N_A_193_47#_c_330_n N_A_27_47#_c_426_n 0.00778651f $X=3.185 $Y=0.9 $X2=0
+ $Y2=0
cc_306 N_A_193_47#_c_327_n N_A_27_47#_c_427_n 0.0039413f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_307 N_A_193_47#_c_335_n N_A_27_47#_c_427_n 0.0169173f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_308 N_A_193_47#_M1004_g N_A_27_47#_M1020_g 0.0177914f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_309 N_A_193_47#_c_333_n N_A_27_47#_M1020_g 0.00173817f $X=2.395 $Y=1.94 $X2=0
+ $Y2=0
cc_310 N_A_193_47#_c_327_n N_A_27_47#_M1020_g 0.00530001f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_311 N_A_193_47#_c_335_n N_A_27_47#_M1020_g 0.0164248f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_312 N_A_193_47#_c_326_n N_A_27_47#_c_429_n 0.00863104f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_313 N_A_193_47#_c_326_n N_A_27_47#_c_438_n 0.0013042f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_314 N_A_193_47#_c_326_n N_A_27_47#_c_439_n 0.0250776f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_315 N_A_193_47#_c_326_n N_A_27_47#_c_431_n 0.0232864f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_316 N_A_193_47#_c_326_n N_A_27_47#_c_432_n 0.0166222f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_317 N_A_193_47#_M1005_g N_A_643_307#_M1021_g 0.0349624f $X=3.185 $Y=0.43
+ $X2=0 $Y2=0
cc_318 N_A_193_47#_c_330_n N_A_643_307#_c_568_n 8.61266e-19 $X=3.185 $Y=0.9
+ $X2=0 $Y2=0
cc_319 N_A_193_47#_M1004_g N_A_477_413#_c_685_n 0.00290984f $X=2.31 $Y=2.275
+ $X2=0 $Y2=0
cc_320 N_A_193_47#_c_333_n N_A_477_413#_c_685_n 0.0100551f $X=2.395 $Y=1.94
+ $X2=0 $Y2=0
cc_321 N_A_193_47#_c_335_n N_A_477_413#_c_685_n 7.93623e-19 $X=2.48 $Y=1.74
+ $X2=0 $Y2=0
cc_322 N_A_193_47#_M1005_g N_A_477_413#_c_678_n 0.00947094f $X=3.185 $Y=0.43
+ $X2=0 $Y2=0
cc_323 N_A_193_47#_c_329_n N_A_477_413#_c_678_n 0.0177012f $X=3.06 $Y=0.9 $X2=0
+ $Y2=0
cc_324 N_A_193_47#_c_330_n N_A_477_413#_c_678_n 0.0044688f $X=3.185 $Y=0.9 $X2=0
+ $Y2=0
cc_325 N_A_193_47#_c_333_n N_A_477_413#_c_672_n 0.00760196f $X=2.395 $Y=1.94
+ $X2=0 $Y2=0
cc_326 N_A_193_47#_c_327_n N_A_477_413#_c_672_n 0.0207723f $X=2.48 $Y=1.74 $X2=0
+ $Y2=0
cc_327 N_A_193_47#_c_330_n N_A_477_413#_c_664_n 4.27554e-19 $X=3.185 $Y=0.9
+ $X2=0 $Y2=0
cc_328 N_A_193_47#_c_327_n N_A_477_413#_c_665_n 0.00577086f $X=2.48 $Y=1.74
+ $X2=0 $Y2=0
cc_329 N_A_193_47#_c_329_n N_A_477_413#_c_665_n 0.010612f $X=3.06 $Y=0.9 $X2=0
+ $Y2=0
cc_330 N_A_193_47#_c_330_n N_A_477_413#_c_665_n 0.00425627f $X=3.185 $Y=0.9
+ $X2=0 $Y2=0
cc_331 N_A_193_47#_M1005_g N_A_477_413#_c_666_n 0.0045695f $X=3.185 $Y=0.43
+ $X2=0 $Y2=0
cc_332 N_A_193_47#_c_329_n N_A_477_413#_c_666_n 0.00815137f $X=3.06 $Y=0.9 $X2=0
+ $Y2=0
cc_333 N_A_193_47#_c_330_n N_A_477_413#_c_669_n 9.68257e-19 $X=3.185 $Y=0.9
+ $X2=0 $Y2=0
cc_334 N_A_193_47#_c_333_n N_VPWR_M1015_s 0.0051328f $X=2.395 $Y=1.94 $X2=0
+ $Y2=0
cc_335 N_A_193_47#_c_336_n N_VPWR_c_848_n 0.0127357f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_336 N_A_193_47#_M1004_g N_VPWR_c_849_n 0.00222571f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_337 N_A_193_47#_c_333_n N_VPWR_c_849_n 0.0235186f $X=2.395 $Y=1.94 $X2=0
+ $Y2=0
cc_338 N_A_193_47#_c_336_n N_VPWR_c_849_n 0.0186826f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_339 N_A_193_47#_c_333_n N_VPWR_c_857_n 0.0028118f $X=2.395 $Y=1.94 $X2=0
+ $Y2=0
cc_340 N_A_193_47#_c_336_n N_VPWR_c_857_n 0.016699f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_341 N_A_193_47#_M1004_g N_VPWR_c_858_n 0.00433717f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_342 N_A_193_47#_c_333_n N_VPWR_c_858_n 0.00977623f $X=2.395 $Y=1.94 $X2=0
+ $Y2=0
cc_343 N_A_193_47#_M1004_g N_VPWR_c_847_n 0.00665706f $X=2.31 $Y=2.275 $X2=0
+ $Y2=0
cc_344 N_A_193_47#_c_333_n N_VPWR_c_847_n 0.0235511f $X=2.395 $Y=1.94 $X2=0
+ $Y2=0
cc_345 N_A_193_47#_c_336_n N_VPWR_c_847_n 0.00973235f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_346 N_A_193_47#_c_333_n A_381_369# 0.00558891f $X=2.395 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_347 N_A_193_47#_c_326_n N_VGND_c_976_n 0.0456749f $X=1.1 $Y=0.425 $X2=0 $Y2=0
cc_348 N_A_193_47#_c_326_n N_VGND_c_982_n 0.0177915f $X=1.1 $Y=0.425 $X2=0 $Y2=0
cc_349 N_A_193_47#_M1005_g N_VGND_c_983_n 0.00384492f $X=3.185 $Y=0.43 $X2=0
+ $Y2=0
cc_350 N_A_193_47#_M1012_d N_VGND_c_990_n 0.00381667f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_351 N_A_193_47#_M1005_g N_VGND_c_990_n 0.00616835f $X=3.185 $Y=0.43 $X2=0
+ $Y2=0
cc_352 N_A_193_47#_c_326_n N_VGND_c_990_n 0.0101048f $X=1.1 $Y=0.425 $X2=0 $Y2=0
cc_353 N_A_193_47#_c_328_n N_VGND_c_990_n 0.00893094f $X=2.645 $Y=0.9 $X2=0
+ $Y2=0
cc_354 N_A_193_47#_c_329_n N_VGND_c_990_n 0.00601035f $X=3.06 $Y=0.9 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_426_n N_A_643_307#_M1021_g 0.00385724f $X=2.855 $Y=1.32
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_M1020_g N_A_643_307#_c_568_n 0.0656786f $X=2.93 $Y=2.275 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_M1020_g N_A_477_413#_c_685_n 0.0146203f $X=2.93 $Y=2.275 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1003_g N_A_477_413#_c_678_n 0.00214477f $X=2.46 $Y=0.54 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_426_n N_A_477_413#_c_672_n 0.00916534f $X=2.855 $Y=1.32
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_M1003_g N_A_477_413#_c_665_n 3.68297e-19 $X=2.46 $Y=0.54 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_426_n N_A_477_413#_c_665_n 0.00145425f $X=2.855 $Y=1.32
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_438_n N_VPWR_M1011_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_363 N_A_27_47#_M1000_g N_VPWR_c_848_n 0.0094125f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_364 N_A_27_47#_c_438_n N_VPWR_c_848_n 0.0155904f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_365 N_A_27_47#_c_440_n N_VPWR_c_848_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_366 N_A_27_47#_M1000_g N_VPWR_c_849_n 0.00181455f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_438_n N_VPWR_c_856_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_440_n N_VPWR_c_856_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_369 N_A_27_47#_M1000_g N_VPWR_c_857_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1020_g N_VPWR_c_858_n 0.00366111f $X=2.93 $Y=2.275 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_M1000_g N_VPWR_c_847_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_M1020_g N_VPWR_c_847_n 0.00560345f $X=2.93 $Y=2.275 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_438_n N_VPWR_c_847_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_440_n N_VPWR_c_847_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_375 N_A_27_47#_c_429_n N_VGND_M1018_d 0.00169549f $X=0.61 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_376 N_A_27_47#_c_419_n N_VGND_c_975_n 0.00728685f $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_377 N_A_27_47#_c_424_n N_VGND_c_975_n 6.21483e-19 $X=1.45 $Y=0.18 $X2=0 $Y2=0
cc_378 N_A_27_47#_c_429_n N_VGND_c_975_n 0.0149823f $X=0.61 $Y=0.7 $X2=0 $Y2=0
cc_379 N_A_27_47#_c_431_n N_VGND_c_975_n 0.00122968f $X=0.755 $Y=1.225 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_433_n N_VGND_c_975_n 5.68744e-19 $X=0.89 $Y=1.225 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_419_n N_VGND_c_976_n 3.94476e-19 $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_382 N_A_27_47#_c_422_n N_VGND_c_976_n 0.00935054f $X=1.375 $Y=0.73 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_423_n N_VGND_c_976_n 0.0231282f $X=2.385 $Y=0.18 $X2=0 $Y2=0
cc_384 N_A_27_47#_M1003_g N_VGND_c_976_n 9.4481e-19 $X=2.46 $Y=0.54 $X2=0 $Y2=0
cc_385 N_A_27_47#_c_541_p N_VGND_c_981_n 0.0110394f $X=0.26 $Y=0.425 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_429_n N_VGND_c_981_n 0.00255672f $X=0.61 $Y=0.7 $X2=0 $Y2=0
cc_387 N_A_27_47#_c_419_n N_VGND_c_982_n 0.0046653f $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_388 N_A_27_47#_c_421_n N_VGND_c_982_n 3.66494e-19 $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_389 N_A_27_47#_c_424_n N_VGND_c_982_n 0.00718072f $X=1.45 $Y=0.18 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_423_n N_VGND_c_983_n 0.0229036f $X=2.385 $Y=0.18 $X2=0 $Y2=0
cc_391 N_A_27_47#_M1018_s N_VGND_c_990_n 0.00367415f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_419_n N_VGND_c_990_n 0.00805453f $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_423_n N_VGND_c_990_n 0.0294157f $X=2.385 $Y=0.18 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_424_n N_VGND_c_990_n 0.0100212f $X=1.45 $Y=0.18 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_541_p N_VGND_c_990_n 0.00641103f $X=0.26 $Y=0.425 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_429_n N_VGND_c_990_n 0.00557795f $X=0.61 $Y=0.7 $X2=0 $Y2=0
cc_397 N_A_643_307#_M1021_g N_A_477_413#_M1019_g 0.011022f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_643_307#_M1010_g N_A_477_413#_M1019_g 0.0322235f $X=4.71 $Y=2.165
+ $X2=0 $Y2=0
cc_399 N_A_643_307#_c_557_n N_A_477_413#_M1019_g 0.00355944f $X=4.542 $Y=1.535
+ $X2=0 $Y2=0
cc_400 N_A_643_307#_c_567_n N_A_477_413#_M1019_g 0.0184685f $X=4.025 $Y=1.7
+ $X2=0 $Y2=0
cc_401 N_A_643_307#_M1002_g N_A_477_413#_c_685_n 0.00338501f $X=3.29 $Y=2.275
+ $X2=0 $Y2=0
cc_402 N_A_643_307#_M1021_g N_A_477_413#_c_678_n 0.00728784f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_643_307#_M1002_g N_A_477_413#_c_672_n 0.0140667f $X=3.29 $Y=2.275
+ $X2=0 $Y2=0
cc_404 N_A_643_307#_M1021_g N_A_477_413#_c_672_n 0.00390654f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_405 N_A_643_307#_c_565_n N_A_477_413#_c_672_n 0.0214954f $X=3.915 $Y=1.7
+ $X2=0 $Y2=0
cc_406 N_A_643_307#_c_568_n N_A_477_413#_c_672_n 0.00742928f $X=3.66 $Y=1.7
+ $X2=0 $Y2=0
cc_407 N_A_643_307#_c_565_n N_A_477_413#_c_664_n 0.00686021f $X=3.915 $Y=1.7
+ $X2=0 $Y2=0
cc_408 N_A_643_307#_c_568_n N_A_477_413#_c_664_n 0.0100115f $X=3.66 $Y=1.7 $X2=0
+ $Y2=0
cc_409 N_A_643_307#_M1021_g N_A_477_413#_c_666_n 0.0133637f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_643_307#_c_560_n N_A_477_413#_c_666_n 0.00989198f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_411 N_A_643_307#_M1021_g N_A_477_413#_c_667_n 0.00399182f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_412 N_A_643_307#_c_554_n N_A_477_413#_c_667_n 3.19628e-19 $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_413 N_A_643_307#_c_565_n N_A_477_413#_c_667_n 0.0120422f $X=3.915 $Y=1.7
+ $X2=0 $Y2=0
cc_414 N_A_643_307#_c_567_n N_A_477_413#_c_667_n 0.0147817f $X=4.025 $Y=1.7
+ $X2=0 $Y2=0
cc_415 N_A_643_307#_c_559_n N_A_477_413#_c_667_n 0.0255776f $X=4.65 $Y=1.16
+ $X2=0 $Y2=0
cc_416 N_A_643_307#_M1021_g N_A_477_413#_c_668_n 0.0195909f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_643_307#_c_554_n N_A_477_413#_c_668_n 0.0212501f $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_418 N_A_643_307#_c_567_n N_A_477_413#_c_668_n 0.00440551f $X=4.025 $Y=1.7
+ $X2=0 $Y2=0
cc_419 N_A_643_307#_c_559_n N_A_477_413#_c_668_n 0.00355944f $X=4.65 $Y=1.16
+ $X2=0 $Y2=0
cc_420 N_A_643_307#_M1021_g N_A_477_413#_c_669_n 0.0120634f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_421 N_A_643_307#_c_565_n N_A_477_413#_c_669_n 0.0104535f $X=3.915 $Y=1.7
+ $X2=0 $Y2=0
cc_422 N_A_643_307#_c_568_n N_A_477_413#_c_669_n 6.84542e-19 $X=3.66 $Y=1.7
+ $X2=0 $Y2=0
cc_423 N_A_643_307#_M1021_g N_A_477_413#_c_670_n 0.019226f $X=3.66 $Y=0.445
+ $X2=0 $Y2=0
cc_424 N_A_643_307#_c_554_n N_A_477_413#_c_670_n 0.00652411f $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_425 N_A_643_307#_c_560_n N_A_477_413#_c_670_n 0.00612822f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_426 N_A_643_307#_c_555_n N_A_957_369#_c_756_n 0.00438336f $X=5.055 $Y=0.805
+ $X2=0 $Y2=0
cc_427 N_A_643_307#_c_556_n N_A_957_369#_c_756_n 0.00371139f $X=5.13 $Y=0.73
+ $X2=0 $Y2=0
cc_428 N_A_643_307#_c_560_n N_A_957_369#_c_756_n 0.00675325f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_429 N_A_643_307#_M1010_g N_A_957_369#_c_770_n 0.00786899f $X=4.71 $Y=2.165
+ $X2=0 $Y2=0
cc_430 N_A_643_307#_c_555_n N_A_957_369#_c_757_n 0.00338698f $X=5.055 $Y=0.805
+ $X2=0 $Y2=0
cc_431 N_A_643_307#_c_554_n N_A_957_369#_c_758_n 7.14018e-19 $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_432 N_A_643_307#_c_555_n N_A_957_369#_c_758_n 0.00750927f $X=5.055 $Y=0.805
+ $X2=0 $Y2=0
cc_433 N_A_643_307#_c_560_n N_A_957_369#_c_758_n 0.00841744f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_434 N_A_643_307#_M1010_g N_A_957_369#_c_765_n 0.00275865f $X=4.71 $Y=2.165
+ $X2=0 $Y2=0
cc_435 N_A_643_307#_c_567_n N_A_957_369#_c_765_n 0.00714245f $X=4.025 $Y=1.7
+ $X2=0 $Y2=0
cc_436 N_A_643_307#_c_555_n N_A_957_369#_c_788_n 0.00372863f $X=5.055 $Y=0.805
+ $X2=0 $Y2=0
cc_437 N_A_643_307#_c_556_n N_A_957_369#_c_788_n 0.00816324f $X=5.13 $Y=0.73
+ $X2=0 $Y2=0
cc_438 N_A_643_307#_c_558_n N_A_957_369#_c_788_n 0.0200453f $X=4.4 $Y=0.45 $X2=0
+ $Y2=0
cc_439 N_A_643_307#_c_567_n N_VPWR_M1019_d 0.00213578f $X=4.025 $Y=1.7 $X2=0
+ $Y2=0
cc_440 N_A_643_307#_M1002_g N_VPWR_c_850_n 0.00467052f $X=3.29 $Y=2.275 $X2=0
+ $Y2=0
cc_441 N_A_643_307#_c_565_n N_VPWR_c_850_n 0.0144253f $X=3.915 $Y=1.7 $X2=0
+ $Y2=0
cc_442 N_A_643_307#_c_639_p N_VPWR_c_850_n 0.0199633f $X=4.02 $Y=2.27 $X2=0
+ $Y2=0
cc_443 N_A_643_307#_c_568_n N_VPWR_c_850_n 0.00709979f $X=3.66 $Y=1.7 $X2=0
+ $Y2=0
cc_444 N_A_643_307#_c_639_p N_VPWR_c_851_n 0.0118127f $X=4.02 $Y=2.27 $X2=0
+ $Y2=0
cc_445 N_A_643_307#_c_554_n N_VPWR_c_852_n 2.18472e-19 $X=4.71 $Y=1.325 $X2=0
+ $Y2=0
cc_446 N_A_643_307#_M1010_g N_VPWR_c_852_n 0.00343634f $X=4.71 $Y=2.165 $X2=0
+ $Y2=0
cc_447 N_A_643_307#_c_567_n N_VPWR_c_852_n 0.0204994f $X=4.025 $Y=1.7 $X2=0
+ $Y2=0
cc_448 N_A_643_307#_M1002_g N_VPWR_c_858_n 0.00563437f $X=3.29 $Y=2.275 $X2=0
+ $Y2=0
cc_449 N_A_643_307#_M1010_g N_VPWR_c_859_n 0.00585385f $X=4.71 $Y=2.165 $X2=0
+ $Y2=0
cc_450 N_A_643_307#_M1019_s N_VPWR_c_847_n 0.00297268f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_A_643_307#_M1002_g N_VPWR_c_847_n 0.0112135f $X=3.29 $Y=2.275 $X2=0
+ $Y2=0
cc_452 N_A_643_307#_M1010_g N_VPWR_c_847_n 0.0115319f $X=4.71 $Y=2.165 $X2=0
+ $Y2=0
cc_453 N_A_643_307#_c_565_n N_VPWR_c_847_n 0.00859146f $X=3.915 $Y=1.7 $X2=0
+ $Y2=0
cc_454 N_A_643_307#_c_639_p N_VPWR_c_847_n 0.00827281f $X=4.02 $Y=2.27 $X2=0
+ $Y2=0
cc_455 N_A_643_307#_c_568_n N_VPWR_c_847_n 0.00167685f $X=3.66 $Y=1.7 $X2=0
+ $Y2=0
cc_456 N_A_643_307#_M1021_g N_VGND_c_977_n 0.00750422f $X=3.66 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_643_307#_M1021_g N_VGND_c_983_n 0.00397712f $X=3.66 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_643_307#_c_554_n N_VGND_c_984_n 0.00399304f $X=4.71 $Y=1.325 $X2=0
+ $Y2=0
cc_459 N_A_643_307#_c_555_n N_VGND_c_984_n 3.02019e-19 $X=5.055 $Y=0.805 $X2=0
+ $Y2=0
cc_460 N_A_643_307#_c_556_n N_VGND_c_984_n 0.00447211f $X=5.13 $Y=0.73 $X2=0
+ $Y2=0
cc_461 N_A_643_307#_c_558_n N_VGND_c_984_n 0.0186302f $X=4.4 $Y=0.45 $X2=0 $Y2=0
cc_462 N_A_643_307#_M1017_d N_VGND_c_990_n 0.00387172f $X=4.265 $Y=0.235 $X2=0
+ $Y2=0
cc_463 N_A_643_307#_M1021_g N_VGND_c_990_n 0.00618418f $X=3.66 $Y=0.445 $X2=0
+ $Y2=0
cc_464 N_A_643_307#_c_554_n N_VGND_c_990_n 0.00516754f $X=4.71 $Y=1.325 $X2=0
+ $Y2=0
cc_465 N_A_643_307#_c_556_n N_VGND_c_990_n 0.00684735f $X=5.13 $Y=0.73 $X2=0
+ $Y2=0
cc_466 N_A_643_307#_c_558_n N_VGND_c_990_n 0.0103005f $X=4.4 $Y=0.45 $X2=0 $Y2=0
cc_467 N_A_477_413#_c_685_n N_VPWR_c_849_n 0.00474258f $X=3.06 $Y=2.34 $X2=0
+ $Y2=0
cc_468 N_A_477_413#_M1019_g N_VPWR_c_850_n 0.00242172f $X=4.23 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_A_477_413#_M1019_g N_VPWR_c_851_n 0.00585385f $X=4.23 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_A_477_413#_M1019_g N_VPWR_c_852_n 0.0021777f $X=4.23 $Y=1.985 $X2=0
+ $Y2=0
cc_471 N_A_477_413#_c_685_n N_VPWR_c_858_n 0.0344605f $X=3.06 $Y=2.34 $X2=0
+ $Y2=0
cc_472 N_A_477_413#_M1004_d N_VPWR_c_847_n 0.00425502f $X=2.385 $Y=2.065 $X2=0
+ $Y2=0
cc_473 N_A_477_413#_M1019_g N_VPWR_c_847_n 0.0121396f $X=4.23 $Y=1.985 $X2=0
+ $Y2=0
cc_474 N_A_477_413#_c_685_n N_VPWR_c_847_n 0.0267056f $X=3.06 $Y=2.34 $X2=0
+ $Y2=0
cc_475 N_A_477_413#_c_685_n A_601_413# 0.00102341f $X=3.06 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_476 N_A_477_413#_c_678_n N_VGND_c_977_n 0.0137306f $X=3.555 $Y=0.475 $X2=0
+ $Y2=0
cc_477 N_A_477_413#_c_666_n N_VGND_c_977_n 0.00358434f $X=3.64 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_477_413#_c_667_n N_VGND_c_977_n 0.00830843f $X=4.095 $Y=1.16 $X2=0
+ $Y2=0
cc_479 N_A_477_413#_c_668_n N_VGND_c_977_n 0.00291445f $X=4.095 $Y=1.16 $X2=0
+ $Y2=0
cc_480 N_A_477_413#_c_670_n N_VGND_c_977_n 0.0102616f $X=4.132 $Y=0.995 $X2=0
+ $Y2=0
cc_481 N_A_477_413#_c_678_n N_VGND_c_983_n 0.0291799f $X=3.555 $Y=0.475 $X2=0
+ $Y2=0
cc_482 N_A_477_413#_c_670_n N_VGND_c_984_n 0.0046653f $X=4.132 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_477_413#_M1003_d N_VGND_c_990_n 0.00392318f $X=2.535 $Y=0.33 $X2=0
+ $Y2=0
cc_484 N_A_477_413#_c_678_n N_VGND_c_990_n 0.0305382f $X=3.555 $Y=0.475 $X2=0
+ $Y2=0
cc_485 N_A_477_413#_c_670_n N_VGND_c_990_n 0.00934473f $X=4.132 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_A_477_413#_c_678_n A_652_47# 0.00632435f $X=3.555 $Y=0.475 $X2=-0.19
+ $Y2=-0.24
cc_487 N_A_957_369#_c_764_n N_VPWR_M1016_d 0.00677965f $X=5.755 $Y=1.81 $X2=0
+ $Y2=0
cc_488 N_A_957_369#_c_766_n N_VPWR_M1016_d 0.00281046f $X=5.84 $Y=1.725 $X2=0
+ $Y2=0
cc_489 N_A_957_369#_M1008_g N_VPWR_c_853_n 0.00836197f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_490 N_A_957_369#_M1014_g N_VPWR_c_853_n 4.9642e-19 $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_A_957_369#_c_764_n N_VPWR_c_853_n 0.0152939f $X=5.755 $Y=1.81 $X2=0
+ $Y2=0
cc_492 N_A_957_369#_M1014_g N_VPWR_c_855_n 0.00626263f $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_957_369#_c_770_n N_VPWR_c_859_n 0.0230652f $X=5.175 $Y=2 $X2=0 $Y2=0
cc_494 N_A_957_369#_M1008_g N_VPWR_c_860_n 0.0046653f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_495 N_A_957_369#_M1014_g N_VPWR_c_860_n 0.005192f $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_957_369#_M1010_d N_VPWR_c_847_n 0.0134269f $X=4.785 $Y=1.845 $X2=0
+ $Y2=0
cc_497 N_A_957_369#_M1008_g N_VPWR_c_847_n 0.00789179f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_A_957_369#_M1014_g N_VPWR_c_847_n 0.00997547f $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_957_369#_c_770_n N_VPWR_c_847_n 0.0126319f $X=5.175 $Y=2 $X2=0 $Y2=0
cc_500 N_A_957_369#_c_764_n N_VPWR_c_847_n 0.00843664f $X=5.755 $Y=1.81 $X2=0
+ $Y2=0
cc_501 N_A_957_369#_M1014_g N_GCLK_c_953_n 0.00158565f $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_502 N_A_957_369#_c_761_n N_GCLK_c_953_n 0.00133324f $X=6.39 $Y=1.16 $X2=0
+ $Y2=0
cc_503 N_A_957_369#_c_754_n N_GCLK_c_951_n 0.00513877f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_957_369#_M1008_g N_GCLK_c_951_n 0.00114665f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_505 N_A_957_369#_c_755_n N_GCLK_c_951_n 0.0111315f $X=6.39 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_957_369#_M1014_g N_GCLK_c_951_n 0.00801433f $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_507 N_A_957_369#_c_757_n N_GCLK_c_951_n 0.0135582f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_508 N_A_957_369#_c_759_n N_GCLK_c_951_n 0.0275571f $X=5.91 $Y=1.16 $X2=0
+ $Y2=0
cc_509 N_A_957_369#_c_766_n N_GCLK_c_951_n 0.0094365f $X=5.84 $Y=1.725 $X2=0
+ $Y2=0
cc_510 N_A_957_369#_c_761_n N_GCLK_c_951_n 0.0258072f $X=6.39 $Y=1.16 $X2=0
+ $Y2=0
cc_511 N_A_957_369#_M1014_g N_GCLK_c_963_n 0.0124369f $X=6.39 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_A_957_369#_c_755_n N_GCLK_c_964_n 0.00458879f $X=6.39 $Y=0.995 $X2=0
+ $Y2=0
cc_513 N_A_957_369#_c_761_n N_GCLK_c_964_n 0.00114811f $X=6.39 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_A_957_369#_c_757_n N_VGND_M1001_d 0.00249767f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_515 N_A_957_369#_c_754_n N_VGND_c_978_n 0.00277568f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_A_957_369#_c_757_n N_VGND_c_978_n 0.0107385f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_517 N_A_957_369#_c_788_n N_VGND_c_978_n 0.00776254f $X=4.92 $Y=0.455 $X2=0
+ $Y2=0
cc_518 N_A_957_369#_c_761_n N_VGND_c_978_n 3.12249e-19 $X=6.39 $Y=1.16 $X2=0
+ $Y2=0
cc_519 N_A_957_369#_c_755_n N_VGND_c_980_n 0.00674434f $X=6.39 $Y=0.995 $X2=0
+ $Y2=0
cc_520 N_A_957_369#_c_788_n N_VGND_c_984_n 0.0158526f $X=4.92 $Y=0.455 $X2=0
+ $Y2=0
cc_521 N_A_957_369#_c_754_n N_VGND_c_985_n 0.00585385f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_522 N_A_957_369#_c_755_n N_VGND_c_985_n 0.00517132f $X=6.39 $Y=0.995 $X2=0
+ $Y2=0
cc_523 N_A_957_369#_M1006_s N_VGND_c_990_n 0.00258814f $X=4.795 $Y=0.235 $X2=0
+ $Y2=0
cc_524 N_A_957_369#_c_754_n N_VGND_c_990_n 0.0076584f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_525 N_A_957_369#_c_755_n N_VGND_c_990_n 0.00992885f $X=6.39 $Y=0.995 $X2=0
+ $Y2=0
cc_526 N_A_957_369#_c_757_n N_VGND_c_990_n 0.0238944f $X=5.755 $Y=0.85 $X2=0
+ $Y2=0
cc_527 N_A_957_369#_c_788_n N_VGND_c_990_n 0.0113132f $X=4.92 $Y=0.455 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_847_n A_381_369# 0.00416624f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_529 N_VPWR_c_847_n A_601_413# 0.00170467f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_530 N_VPWR_c_847_n N_GCLK_M1008_s 0.00389051f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_531 N_VPWR_c_855_n N_GCLK_c_951_n 0.0730626f $X=6.63 $Y=1.66 $X2=0 $Y2=0
cc_532 N_VPWR_c_860_n N_GCLK_c_963_n 0.0152033f $X=6.53 $Y=2.72 $X2=0 $Y2=0
cc_533 N_VPWR_c_847_n N_GCLK_c_963_n 0.00980611f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_534 N_VPWR_c_855_n N_VGND_c_980_n 0.00987441f $X=6.63 $Y=1.66 $X2=0 $Y2=0
cc_535 N_GCLK_c_951_n N_VGND_c_980_n 0.0213856f $X=6.227 $Y=1.495 $X2=0 $Y2=0
cc_536 N_GCLK_c_964_n N_VGND_c_980_n 0.0258553f $X=6.262 $Y=0.425 $X2=0 $Y2=0
cc_537 N_GCLK_c_964_n N_VGND_c_985_n 0.0167319f $X=6.262 $Y=0.425 $X2=0 $Y2=0
cc_538 N_GCLK_M1007_s N_VGND_c_990_n 0.00263828f $X=6.045 $Y=0.235 $X2=0 $Y2=0
cc_539 N_GCLK_c_964_n N_VGND_c_990_n 0.0110716f $X=6.262 $Y=0.425 $X2=0 $Y2=0
cc_540 N_VGND_c_990_n A_652_47# 0.00282597f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_541 N_VGND_c_990_n A_1041_47# 0.00285576f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24

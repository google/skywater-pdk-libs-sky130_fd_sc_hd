# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__inv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.970000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 5.270000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 5.895000 0.905000 ;
        RECT 0.085000 0.905000 0.510000 1.495000 ;
        RECT 0.085000 1.495000 5.895000 1.665000 ;
        RECT 0.680000 0.255000 1.010000 0.715000 ;
        RECT 0.680000 1.665000 1.010000 2.465000 ;
        RECT 1.520000 0.255000 1.850000 0.715000 ;
        RECT 1.520000 1.665000 1.850000 2.465000 ;
        RECT 2.360000 0.255000 2.690000 0.715000 ;
        RECT 2.360000 1.665000 2.690000 2.465000 ;
        RECT 3.200000 0.255000 3.530000 0.715000 ;
        RECT 3.200000 1.665000 3.530000 2.465000 ;
        RECT 4.040000 0.255000 4.370000 0.715000 ;
        RECT 4.040000 1.665000 4.370000 2.465000 ;
        RECT 4.880000 0.255000 5.210000 0.715000 ;
        RECT 4.880000 1.665000 5.210000 2.465000 ;
        RECT 5.545000 0.905000 5.895000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.180000  0.085000 1.350000 0.545000 ;
      RECT 1.180000  1.835000 1.350000 2.635000 ;
      RECT 2.020000  0.085000 2.190000 0.545000 ;
      RECT 2.020000  1.835000 2.190000 2.635000 ;
      RECT 2.860000  0.085000 3.030000 0.545000 ;
      RECT 2.860000  1.835000 3.030000 2.635000 ;
      RECT 3.700000  0.085000 3.870000 0.545000 ;
      RECT 3.700000  1.835000 3.870000 2.635000 ;
      RECT 4.540000  0.085000 4.710000 0.545000 ;
      RECT 4.540000  1.835000 4.710000 2.635000 ;
      RECT 5.555000  0.085000 5.895000 0.545000 ;
      RECT 5.555000  1.835000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_12
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 Y B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.3328e+12p pd=1.271e+07u as=1.08e+12p ps=1.016e+07u
M1001 a_31_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=1.5665e+12p pd=1.652e+07u as=1.40075e+12p ps=1.211e+07u
M1002 VGND A3 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_31_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.51e+11p ps=3.68e+06u
M1004 Y A3 a_449_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.08e+12p ps=1.016e+07u
M1005 a_27_297# A2 a_449_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.3505e+12p pd=1.274e+07u as=0p ps=0u
M1006 Y B1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_449_297# A3 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_31_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_31_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_31_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_31_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_449_297# A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# A2 a_449_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_31_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A1 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A2 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_31_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A3 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_449_297# A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A3 a_449_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A2 a_31_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_449_297# A3 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__einvp_4.spice.SKY130_FD_SC_HD__EINVP_4.pxi
* Created: Thu Aug 27 14:20:50 2020
* 
x_PM_SKY130_FD_SC_HD__EINVP_4%TE N_TE_c_83_n N_TE_M1015_g N_TE_M1011_g
+ N_TE_c_84_n N_TE_c_85_n N_TE_c_86_n N_TE_M1003_g N_TE_c_87_n N_TE_c_88_n
+ N_TE_M1007_g N_TE_c_89_n N_TE_c_90_n N_TE_M1009_g N_TE_c_91_n N_TE_c_92_n
+ N_TE_M1010_g N_TE_c_93_n N_TE_c_94_n N_TE_c_95_n TE TE
+ PM_SKY130_FD_SC_HD__EINVP_4%TE
x_PM_SKY130_FD_SC_HD__EINVP_4%A_27_47# N_A_27_47#_M1015_s N_A_27_47#_M1011_s
+ N_A_27_47#_c_170_n N_A_27_47#_M1000_g N_A_27_47#_c_171_n N_A_27_47#_c_172_n
+ N_A_27_47#_c_173_n N_A_27_47#_M1001_g N_A_27_47#_c_174_n N_A_27_47#_c_175_n
+ N_A_27_47#_M1002_g N_A_27_47#_c_176_n N_A_27_47#_M1006_g N_A_27_47#_c_177_n
+ N_A_27_47#_c_178_n N_A_27_47#_c_165_n N_A_27_47#_c_179_n N_A_27_47#_c_166_n
+ N_A_27_47#_c_167_n N_A_27_47#_c_180_n N_A_27_47#_c_168_n N_A_27_47#_c_169_n
+ N_A_27_47#_c_208_n PM_SKY130_FD_SC_HD__EINVP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVP_4%A N_A_c_270_n N_A_M1013_g N_A_M1004_g N_A_c_271_n
+ N_A_M1014_g N_A_M1005_g N_A_M1016_g N_A_M1008_g N_A_c_274_n N_A_M1017_g
+ N_A_M1012_g A A A PM_SKY130_FD_SC_HD__EINVP_4%A
x_PM_SKY130_FD_SC_HD__EINVP_4%VPWR N_VPWR_M1011_d N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n VPWR N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_345_n N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_356_n PM_SKY130_FD_SC_HD__EINVP_4%VPWR
x_PM_SKY130_FD_SC_HD__EINVP_4%A_215_309# N_A_215_309#_M1000_d
+ N_A_215_309#_M1001_d N_A_215_309#_M1006_d N_A_215_309#_M1005_s
+ N_A_215_309#_M1012_s N_A_215_309#_c_419_n N_A_215_309#_c_424_n
+ N_A_215_309#_c_416_n N_A_215_309#_c_456_n N_A_215_309#_c_430_n
+ N_A_215_309#_c_434_n N_A_215_309#_c_439_n N_A_215_309#_c_463_n
+ N_A_215_309#_c_473_p N_A_215_309#_c_417_n N_A_215_309#_c_418_n
+ N_A_215_309#_c_422_n N_A_215_309#_c_468_n
+ PM_SKY130_FD_SC_HD__EINVP_4%A_215_309#
x_PM_SKY130_FD_SC_HD__EINVP_4%Z N_Z_M1013_d N_Z_M1016_d N_Z_M1004_d N_Z_M1008_d
+ N_Z_c_480_n N_Z_c_481_n N_Z_c_482_n Z Z Z Z N_Z_c_511_n
+ PM_SKY130_FD_SC_HD__EINVP_4%Z
x_PM_SKY130_FD_SC_HD__EINVP_4%VGND N_VGND_M1015_d N_VGND_M1007_d N_VGND_M1010_d
+ N_VGND_c_535_n N_VGND_c_536_n N_VGND_c_537_n VGND N_VGND_c_538_n
+ N_VGND_c_539_n N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n
+ N_VGND_c_544_n N_VGND_c_545_n PM_SKY130_FD_SC_HD__EINVP_4%VGND
x_PM_SKY130_FD_SC_HD__EINVP_4%A_193_47# N_A_193_47#_M1003_s N_A_193_47#_M1009_s
+ N_A_193_47#_M1013_s N_A_193_47#_M1014_s N_A_193_47#_M1017_s
+ N_A_193_47#_c_616_n N_A_193_47#_c_617_n N_A_193_47#_c_620_n
+ N_A_193_47#_c_656_n N_A_193_47#_c_612_n N_A_193_47#_c_613_n
+ N_A_193_47#_c_614_n N_A_193_47#_c_615_n N_A_193_47#_c_624_n
+ PM_SKY130_FD_SC_HD__EINVP_4%A_193_47#
cc_1 VNB N_TE_c_83_n 0.0186243f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_2 VNB N_TE_c_84_n 0.0144728f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=1.035
cc_3 VNB N_TE_c_85_n 0.039391f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.035
cc_4 VNB N_TE_c_86_n 0.0141775f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.96
cc_5 VNB N_TE_c_87_n 0.0152216f $X=-0.19 $Y=-0.24 $X2=1.255 $Y2=1.035
cc_6 VNB N_TE_c_88_n 0.0141947f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.96
cc_7 VNB N_TE_c_89_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=1.035
cc_8 VNB N_TE_c_90_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.96
cc_9 VNB N_TE_c_91_n 0.016072f $X=-0.19 $Y=-0.24 $X2=2.095 $Y2=1.035
cc_10 VNB N_TE_c_92_n 0.018285f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.96
cc_11 VNB N_TE_c_93_n 0.00661167f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.035
cc_12 VNB N_TE_c_94_n 0.0053816f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.035
cc_13 VNB N_TE_c_95_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.035
cc_14 VNB TE 0.0134173f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_27_47#_c_165_n 0.0156742f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_16 VNB N_A_27_47#_c_166_n 0.00753012f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_17 VNB N_A_27_47#_c_167_n 7.10498e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.142
cc_18 VNB N_A_27_47#_c_168_n 0.00764942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_169_n 0.0274244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_c_270_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_21 VNB N_A_c_271_n 0.0155271f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=1.035
cc_22 VNB N_A_M1016_g 0.0173901f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_23 VNB N_A_M1008_g 4.49313e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_24 VNB N_A_c_274_n 0.0864023f $X=-0.19 $Y=-0.24 $X2=2.095 $Y2=1.035
cc_25 VNB N_A_M1017_g 0.0235825f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.96
cc_26 VNB A 0.0189454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_345_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Z_c_480_n 0.0140745f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.96
cc_29 VNB N_VGND_c_535_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_30 VNB N_VGND_c_536_n 3.05427e-19 $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_31 VNB N_VGND_c_537_n 0.00523058f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.96
cc_32 VNB N_VGND_c_538_n 0.014319f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.035
cc_33 VNB N_VGND_c_539_n 0.0123936f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.035
cc_34 VNB N_VGND_c_540_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_541_n 0.0595324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_542_n 0.260684f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_37 VNB N_VGND_c_543_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_544_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_545_n 0.00526505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_612_n 0.00621295f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.56
cc_41 VNB N_A_193_47#_c_613_n 0.0029431f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_42 VNB N_A_193_47#_c_614_n 0.00268471f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_43 VNB N_A_193_47#_c_615_n 0.0136445f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_44 VPB N_TE_M1011_g 0.025505f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB N_TE_c_85_n 0.0104436f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.035
cc_46 VPB TE 0.0127315f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_A_27_47#_c_170_n 0.0174982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_171_n 0.00892157f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.96
cc_49 VPB N_A_27_47#_c_172_n 0.00858091f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_50 VPB N_A_27_47#_c_173_n 0.0140273f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_51 VPB N_A_27_47#_c_174_n 0.00892095f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.96
cc_52 VPB N_A_27_47#_c_175_n 0.0140273f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_53 VPB N_A_27_47#_c_176_n 0.0144646f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.96
cc_54 VPB N_A_27_47#_c_177_n 0.00391059f $X=-0.19 $Y=1.305 $X2=2.095 $Y2=1.035
cc_55 VPB N_A_27_47#_c_178_n 0.0215363f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.56
cc_56 VPB N_A_27_47#_c_179_n 0.0198657f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.142
cc_57 VPB N_A_27_47#_c_180_n 0.0168045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_168_n 0.0139959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_169_n 0.00101273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_M1004_g 0.0187449f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_A_M1005_g 0.0176224f $X=-0.19 $Y=1.305 $X2=1.255 $Y2=1.035
cc_62 VPB N_A_M1008_g 0.0191533f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_63 VPB N_A_c_274_n 0.0122327f $X=-0.19 $Y=1.305 $X2=2.095 $Y2=1.035
cc_64 VPB N_A_M1012_g 0.0263683f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.035
cc_65 VPB N_VPWR_c_346_n 0.0066501f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_66 VPB N_VPWR_c_347_n 3.14017e-19 $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_67 VPB N_VPWR_c_348_n 3.95616e-19 $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.96
cc_68 VPB N_VPWR_c_349_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.035
cc_69 VPB N_VPWR_c_350_n 0.0153895f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.035
cc_70 VPB N_VPWR_c_351_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_352_n 0.0569038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_345_n 0.0537362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_354_n 0.00565587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_355_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_356_n 0.00476819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_215_309#_c_416_n 0.00133077f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_77 VPB N_A_215_309#_c_417_n 0.0101124f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.142
cc_78 VPB N_A_215_309#_c_418_n 0.0439944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_Z_c_481_n 0.0026552f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.035
cc_80 VPB N_Z_c_482_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_81 TE N_A_27_47#_M1011_s 0.00429701f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_82 N_TE_c_89_n N_A_27_47#_c_171_n 0.0147681f $X=1.675 $Y=1.035 $X2=0 $Y2=0
cc_83 N_TE_c_94_n N_A_27_47#_c_172_n 0.0147681f $X=1.33 $Y=1.035 $X2=0 $Y2=0
cc_84 N_TE_c_91_n N_A_27_47#_c_174_n 0.0147681f $X=2.095 $Y=1.035 $X2=0 $Y2=0
cc_85 N_TE_c_95_n N_A_27_47#_c_177_n 0.0147681f $X=1.75 $Y=1.035 $X2=0 $Y2=0
cc_86 N_TE_c_83_n N_A_27_47#_c_166_n 0.0150211f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_87 N_TE_c_84_n N_A_27_47#_c_166_n 3.34655e-19 $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_88 N_TE_c_85_n N_A_27_47#_c_166_n 0.0030701f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_89 N_TE_c_86_n N_A_27_47#_c_166_n 0.00161437f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_90 TE N_A_27_47#_c_166_n 0.0191066f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_91 N_TE_c_83_n N_A_27_47#_c_167_n 0.00680774f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_92 N_TE_c_84_n N_A_27_47#_c_167_n 0.00300693f $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_93 N_TE_c_85_n N_A_27_47#_c_167_n 0.0014487f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_94 N_TE_c_86_n N_A_27_47#_c_167_n 0.00302911f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_95 N_TE_M1011_g N_A_27_47#_c_180_n 0.0379477f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_96 N_TE_c_84_n N_A_27_47#_c_180_n 5.69379e-19 $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_97 N_TE_c_85_n N_A_27_47#_c_180_n 0.00193181f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_98 TE N_A_27_47#_c_180_n 0.0421802f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_99 N_TE_c_87_n N_A_27_47#_c_168_n 0.0139399f $X=1.255 $Y=1.035 $X2=0 $Y2=0
cc_100 N_TE_c_89_n N_A_27_47#_c_168_n 0.0083577f $X=1.675 $Y=1.035 $X2=0 $Y2=0
cc_101 N_TE_c_91_n N_A_27_47#_c_168_n 0.0145953f $X=2.095 $Y=1.035 $X2=0 $Y2=0
cc_102 N_TE_c_93_n N_A_27_47#_c_168_n 0.00686545f $X=0.89 $Y=1.035 $X2=0 $Y2=0
cc_103 N_TE_c_94_n N_A_27_47#_c_168_n 0.0058582f $X=1.33 $Y=1.035 $X2=0 $Y2=0
cc_104 N_TE_c_95_n N_A_27_47#_c_168_n 0.0051004f $X=1.75 $Y=1.035 $X2=0 $Y2=0
cc_105 N_TE_c_91_n N_A_27_47#_c_169_n 0.00670028f $X=2.095 $Y=1.035 $X2=0 $Y2=0
cc_106 N_TE_c_84_n N_A_27_47#_c_208_n 0.0120485f $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_107 N_TE_c_85_n N_A_27_47#_c_208_n 0.0115149f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_108 N_TE_c_93_n N_A_27_47#_c_208_n 0.00442816f $X=0.89 $Y=1.035 $X2=0 $Y2=0
cc_109 TE N_A_27_47#_c_208_n 0.025787f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_110 N_TE_M1011_g N_VPWR_c_346_n 0.0113741f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_111 N_TE_M1011_g N_VPWR_c_349_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_112 N_TE_M1011_g N_VPWR_c_345_n 0.00523707f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_TE_M1011_g N_A_215_309#_c_419_n 0.00545173f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_TE_M1011_g N_A_215_309#_c_416_n 6.87579e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_TE_c_87_n N_A_215_309#_c_416_n 0.00101624f $X=1.255 $Y=1.035 $X2=0
+ $Y2=0
cc_116 N_TE_c_91_n N_A_215_309#_c_422_n 2.11158e-19 $X=2.095 $Y=1.035 $X2=0
+ $Y2=0
cc_117 N_TE_c_83_n N_VGND_c_535_n 0.00856801f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_118 N_TE_c_84_n N_VGND_c_535_n 5.1499e-19 $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_119 N_TE_c_86_n N_VGND_c_535_n 0.00735324f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_120 N_TE_c_88_n N_VGND_c_535_n 5.57248e-19 $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_121 N_TE_c_86_n N_VGND_c_536_n 5.5023e-19 $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_122 N_TE_c_88_n N_VGND_c_536_n 0.00691072f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_123 N_TE_c_90_n N_VGND_c_536_n 0.00685342f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_124 N_TE_c_92_n N_VGND_c_536_n 5.54209e-19 $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_125 N_TE_c_90_n N_VGND_c_537_n 5.54817e-19 $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_126 N_TE_c_92_n N_VGND_c_537_n 0.0079747f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_127 N_TE_c_83_n N_VGND_c_538_n 0.00341689f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_128 N_TE_c_86_n N_VGND_c_539_n 0.0046653f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_129 N_TE_c_88_n N_VGND_c_539_n 0.00341689f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_130 N_TE_c_90_n N_VGND_c_540_n 0.00341689f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_131 N_TE_c_92_n N_VGND_c_540_n 0.00341689f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_132 N_TE_c_83_n N_VGND_c_542_n 0.0050171f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_133 N_TE_c_86_n N_VGND_c_542_n 0.00802193f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_134 N_TE_c_88_n N_VGND_c_542_n 0.00408046f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_135 N_TE_c_90_n N_VGND_c_542_n 0.0040262f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_136 N_TE_c_92_n N_VGND_c_542_n 0.0040262f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_137 N_TE_c_86_n N_A_193_47#_c_616_n 0.0043107f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_138 N_TE_c_88_n N_A_193_47#_c_617_n 0.0103667f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_139 N_TE_c_89_n N_A_193_47#_c_617_n 0.00179137f $X=1.675 $Y=1.035 $X2=0 $Y2=0
cc_140 N_TE_c_90_n N_A_193_47#_c_617_n 0.0104925f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_141 N_TE_c_86_n N_A_193_47#_c_620_n 0.00161811f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_142 N_TE_c_87_n N_A_193_47#_c_620_n 0.00227361f $X=1.255 $Y=1.035 $X2=0 $Y2=0
cc_143 N_TE_c_92_n N_A_193_47#_c_612_n 0.0126397f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_144 N_TE_c_92_n N_A_193_47#_c_613_n 0.00356665f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_145 N_TE_c_91_n N_A_193_47#_c_624_n 0.00186022f $X=2.095 $Y=1.035 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_178_n N_A_M1004_g 0.0169217f $X=2.67 $Y=1.395 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_168_n N_A_c_274_n 0.00353496f $X=2.61 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_169_n N_A_c_274_n 0.0169217f $X=2.61 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_180_n N_VPWR_M1011_d 0.00535662f $X=0.687 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_27_47#_c_170_n N_VPWR_c_346_n 0.00230982f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_180_n N_VPWR_c_346_n 0.0238531f $X=0.687 $Y=1.785 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_170_n N_VPWR_c_347_n 0.0109235f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_173_n N_VPWR_c_347_n 0.0104025f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_175_n N_VPWR_c_347_n 6.14905e-19 $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_173_n N_VPWR_c_348_n 6.16465e-19 $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_175_n N_VPWR_c_348_n 0.0104025f $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_176_n N_VPWR_c_348_n 0.0141295f $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_179_n N_VPWR_c_349_n 0.0176305f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_170_n N_VPWR_c_350_n 0.0046653f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_173_n N_VPWR_c_351_n 0.0046653f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_175_n N_VPWR_c_351_n 0.0046653f $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_176_n N_VPWR_c_352_n 0.00349454f $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1011_s N_VPWR_c_345_n 0.00238524f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_170_n N_VPWR_c_345_n 0.00934473f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_173_n N_VPWR_c_345_n 0.00789179f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_175_n N_VPWR_c_345_n 0.00789179f $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_176_n N_VPWR_c_345_n 0.00622848f $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_179_n N_VPWR_c_345_n 0.00986266f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_180_n N_VPWR_c_345_n 0.00671954f $X=0.687 $Y=1.785 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_180_n N_A_215_309#_c_419_n 0.0168242f $X=0.687 $Y=1.785
+ $X2=0 $Y2=0
cc_171 N_A_27_47#_c_170_n N_A_215_309#_c_424_n 0.0155912f $X=1.41 $Y=1.47 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_171_n N_A_215_309#_c_424_n 0.00197697f $X=1.755 $Y=1.395
+ $X2=0 $Y2=0
cc_173 N_A_27_47#_c_173_n N_A_215_309#_c_424_n 0.0142192f $X=1.83 $Y=1.47 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_168_n N_A_215_309#_c_424_n 0.0323847f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_180_n N_A_215_309#_c_416_n 0.0132199f $X=0.687 $Y=1.785
+ $X2=0 $Y2=0
cc_176 N_A_27_47#_c_168_n N_A_215_309#_c_416_n 0.0143803f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_175_n N_A_215_309#_c_430_n 0.0143019f $X=2.25 $Y=1.47 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_176_n N_A_215_309#_c_430_n 0.0133206f $X=2.67 $Y=1.47 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_178_n N_A_215_309#_c_430_n 0.0021442f $X=2.67 $Y=1.395 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_168_n N_A_215_309#_c_430_n 0.0459386f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_176_n N_A_215_309#_c_434_n 0.00446602f $X=2.67 $Y=1.47 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_174_n N_A_215_309#_c_422_n 0.00209962f $X=2.175 $Y=1.395
+ $X2=0 $Y2=0
cc_183 N_A_27_47#_c_168_n N_A_215_309#_c_422_n 0.0106208f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_178_n Z 6.97699e-19 $X=2.67 $Y=1.395 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_168_n Z 0.027927f $X=2.61 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_169_n Z 2.33571e-19 $X=2.61 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_178_n Z 5.5131e-19 $X=2.67 $Y=1.395 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_166_n N_VGND_M1015_d 0.00310523f $X=0.597 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_27_47#_c_167_n N_VGND_M1015_d 9.5711e-19 $X=0.597 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_27_47#_c_166_n N_VGND_c_535_n 0.00918217f $X=0.597 $Y=0.825 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_208_n N_VGND_c_535_n 0.004225f $X=0.687 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_165_n N_VGND_c_538_n 0.0173297f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_166_n N_VGND_c_538_n 0.00235711f $X=0.597 $Y=0.825 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1015_s N_VGND_c_542_n 0.00230206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_165_n N_VGND_c_542_n 0.00980382f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_166_n N_VGND_c_542_n 0.00499131f $X=0.597 $Y=0.825 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_168_n N_A_193_47#_c_617_n 0.0408222f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_166_n N_A_193_47#_c_620_n 0.00897896f $X=0.597 $Y=0.825
+ $X2=0 $Y2=0
cc_199 N_A_27_47#_c_168_n N_A_193_47#_c_620_n 0.0135368f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_178_n N_A_193_47#_c_612_n 7.32088e-19 $X=2.67 $Y=1.395 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_168_n N_A_193_47#_c_612_n 0.0720037f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_169_n N_A_193_47#_c_612_n 0.00705672f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_168_n N_A_193_47#_c_624_n 0.0132296f $X=2.61 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_A_M1004_g N_VPWR_c_348_n 0.00108764f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_M1004_g N_VPWR_c_352_n 0.00357877f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_M1005_g N_VPWR_c_352_n 0.00357877f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_M1008_g N_VPWR_c_352_n 0.00357877f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_M1012_g N_VPWR_c_352_n 0.00357877f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_M1004_g N_VPWR_c_345_n 0.00538183f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_M1005_g N_VPWR_c_345_n 0.00522516f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_M1008_g N_VPWR_c_345_n 0.00522516f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_M1012_g N_VPWR_c_345_n 0.00631565f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_M1004_g N_A_215_309#_c_430_n 0.00151659f $X=3.145 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_M1004_g N_A_215_309#_c_434_n 0.00464905f $X=3.145 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_M1004_g N_A_215_309#_c_439_n 0.0112448f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_M1005_g N_A_215_309#_c_439_n 0.0112143f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_M1008_g N_A_215_309#_c_417_n 0.0112878f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_M1012_g N_A_215_309#_c_417_n 0.0112878f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_c_274_n N_A_215_309#_c_418_n 0.00515666f $X=4.405 $Y=1.015 $X2=0
+ $Y2=0
cc_220 N_A_M1012_g N_A_215_309#_c_418_n 0.00629935f $X=4.405 $Y=1.985 $X2=0
+ $Y2=0
cc_221 A N_A_215_309#_c_418_n 0.0376052f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A_c_271_n N_Z_c_480_n 0.00662588f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_M1016_g N_Z_c_480_n 0.00955084f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_c_274_n N_Z_c_480_n 0.00729715f $X=4.405 $Y=1.015 $X2=0 $Y2=0
cc_225 N_A_M1017_g N_Z_c_480_n 0.0118735f $X=4.405 $Y=0.56 $X2=0 $Y2=0
cc_226 A N_Z_c_480_n 0.0845534f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_227 N_A_M1005_g N_Z_c_481_n 0.00792131f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_M1008_g N_Z_c_481_n 0.0107189f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_c_274_n N_Z_c_481_n 0.00202711f $X=4.405 $Y=1.015 $X2=0 $Y2=0
cc_230 A N_Z_c_481_n 0.020892f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_231 N_A_M1005_g N_Z_c_482_n 5.55259e-19 $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A_M1008_g N_Z_c_482_n 0.00821596f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A_c_274_n N_Z_c_482_n 0.00206069f $X=4.405 $Y=1.015 $X2=0 $Y2=0
cc_234 N_A_M1012_g N_Z_c_482_n 0.00874816f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_235 A N_Z_c_482_n 0.0270809f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_236 N_A_c_270_n Z 0.0113088f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_M1004_g Z 0.00368663f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A_c_271_n Z 0.00721077f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_M1005_g Z 0.00403311f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_M1016_g Z 9.23891e-19 $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_241 N_A_M1008_g Z 8.07324e-19 $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A_c_274_n Z 0.0233987f $X=4.405 $Y=1.015 $X2=0 $Y2=0
cc_243 A Z 0.0204219f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_244 N_A_M1004_g Z 0.00349612f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_M1005_g Z 0.00435499f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_M1004_g N_Z_c_511_n 0.00613722f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_M1005_g N_Z_c_511_n 0.00700222f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_M1008_g N_Z_c_511_n 5.53432e-19 $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_c_274_n N_Z_c_511_n 3.13877e-19 $X=4.405 $Y=1.015 $X2=0 $Y2=0
cc_250 N_A_c_270_n N_VGND_c_537_n 0.00297242f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_270_n N_VGND_c_541_n 0.00357877f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_271_n N_VGND_c_541_n 0.00357877f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_M1016_g N_VGND_c_541_n 0.00357877f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_M1017_g N_VGND_c_541_n 0.00357877f $X=4.405 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A_c_270_n N_VGND_c_542_n 0.00664112f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_c_271_n N_VGND_c_542_n 0.00522516f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A_M1016_g N_VGND_c_542_n 0.00522516f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A_M1017_g N_VGND_c_542_n 0.00631565f $X=4.405 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_c_270_n N_A_193_47#_c_615_n 0.0141663f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_c_271_n N_A_193_47#_c_615_n 0.00866372f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_M1016_g N_A_193_47#_c_615_n 0.00866705f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_c_274_n N_A_193_47#_c_615_n 3.01257e-19 $X=4.405 $Y=1.015 $X2=0 $Y2=0
cc_263 N_A_M1017_g N_A_193_47#_c_615_n 0.00866705f $X=4.405 $Y=0.56 $X2=0 $Y2=0
cc_264 N_VPWR_c_345_n N_A_215_309#_M1000_d 0.00386369f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_265 N_VPWR_c_345_n N_A_215_309#_M1001_d 0.00562358f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_345_n N_A_215_309#_M1006_d 0.00535913f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_345_n N_A_215_309#_M1005_s 0.0021521f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_345_n N_A_215_309#_M1012_s 0.00209324f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_346_n N_A_215_309#_c_419_n 0.0240954f $X=0.68 $Y=2.34 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_350_n N_A_215_309#_c_419_n 0.0144177f $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_345_n N_A_215_309#_c_419_n 0.00801045f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_272 N_VPWR_M1000_s N_A_215_309#_c_424_n 0.00318028f $X=1.485 $Y=1.545 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_347_n N_A_215_309#_c_424_n 0.0170258f $X=1.62 $Y=2.02 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_351_n N_A_215_309#_c_456_n 0.0113958f $X=2.295 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_345_n N_A_215_309#_c_456_n 0.00646998f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_M1002_s N_A_215_309#_c_430_n 0.00328966f $X=2.325 $Y=1.545 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_348_n N_A_215_309#_c_430_n 0.0193111f $X=2.46 $Y=2.02 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_348_n N_A_215_309#_c_434_n 0.0296995f $X=2.46 $Y=2.02 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_352_n N_A_215_309#_c_439_n 0.037199f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_345_n N_A_215_309#_c_439_n 0.0243735f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_348_n N_A_215_309#_c_463_n 0.0141244f $X=2.46 $Y=2.02 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_352_n N_A_215_309#_c_463_n 0.0119545f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_345_n N_A_215_309#_c_463_n 0.006547f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_c_352_n N_A_215_309#_c_417_n 0.0672109f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_345_n N_A_215_309#_c_417_n 0.0405749f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_352_n N_A_215_309#_c_468_n 0.0114668f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_345_n N_A_215_309#_c_468_n 0.006547f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_345_n N_Z_M1004_d 0.00216833f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_345_n N_Z_M1008_d 0.00216833f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_290 N_A_215_309#_c_439_n N_Z_M1004_d 0.00312752f $X=3.69 $Y=2.38 $X2=0 $Y2=0
cc_291 N_A_215_309#_c_417_n N_Z_M1008_d 0.00312348f $X=4.53 $Y=2.38 $X2=0 $Y2=0
cc_292 N_A_215_309#_M1005_s N_Z_c_481_n 0.00165831f $X=3.64 $Y=1.485 $X2=0 $Y2=0
cc_293 N_A_215_309#_c_473_p N_Z_c_481_n 0.0126919f $X=3.775 $Y=1.96 $X2=0 $Y2=0
cc_294 N_A_215_309#_c_417_n N_Z_c_482_n 0.015949f $X=4.53 $Y=2.38 $X2=0 $Y2=0
cc_295 N_A_215_309#_c_418_n N_Z_c_482_n 0.00886584f $X=4.752 $Y=2.295 $X2=0
+ $Y2=0
cc_296 N_A_215_309#_c_430_n Z 0.00471238f $X=2.825 $Y=1.64 $X2=0 $Y2=0
cc_297 N_A_215_309#_c_430_n N_Z_c_511_n 0.00813072f $X=2.825 $Y=1.64 $X2=0 $Y2=0
cc_298 N_A_215_309#_c_434_n N_Z_c_511_n 0.0265852f $X=2.91 $Y=1.96 $X2=0 $Y2=0
cc_299 N_A_215_309#_c_439_n N_Z_c_511_n 0.0156199f $X=3.69 $Y=2.38 $X2=0 $Y2=0
cc_300 N_Z_M1013_d N_VGND_c_542_n 0.00216833f $X=3.22 $Y=0.235 $X2=0 $Y2=0
cc_301 N_Z_M1016_d N_VGND_c_542_n 0.00216833f $X=4.06 $Y=0.235 $X2=0 $Y2=0
cc_302 N_Z_c_480_n N_A_193_47#_M1014_s 0.00338736f $X=4.195 $Y=0.76 $X2=0 $Y2=0
cc_303 N_Z_c_480_n N_A_193_47#_M1017_s 0.00533714f $X=4.195 $Y=0.76 $X2=0 $Y2=0
cc_304 N_Z_M1013_d N_A_193_47#_c_615_n 0.00304479f $X=3.22 $Y=0.235 $X2=0 $Y2=0
cc_305 N_Z_M1016_d N_A_193_47#_c_615_n 0.00305599f $X=4.06 $Y=0.235 $X2=0 $Y2=0
cc_306 N_Z_c_480_n N_A_193_47#_c_615_n 0.0784481f $X=4.195 $Y=0.76 $X2=0 $Y2=0
cc_307 Z N_A_193_47#_c_615_n 0.0201274f $X=3.39 $Y=0.765 $X2=0 $Y2=0
cc_308 N_VGND_c_542_n N_A_193_47#_M1003_s 0.00498236f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_309 N_VGND_c_542_n N_A_193_47#_M1009_s 0.00254582f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_542_n N_A_193_47#_M1013_s 0.00210127f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_542_n N_A_193_47#_M1014_s 0.00215227f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_542_n N_A_193_47#_M1017_s 0.00225742f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_535_n N_A_193_47#_c_616_n 0.0155846f $X=0.68 $Y=0.36 $X2=0 $Y2=0
cc_314 N_VGND_c_539_n N_A_193_47#_c_616_n 0.011459f $X=1.375 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_542_n N_A_193_47#_c_616_n 0.00644035f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_M1007_d N_A_193_47#_c_617_n 0.00297022f $X=1.405 $Y=0.235 $X2=0
+ $Y2=0
cc_317 N_VGND_c_536_n N_A_193_47#_c_617_n 0.0160613f $X=1.54 $Y=0.36 $X2=0 $Y2=0
cc_318 N_VGND_c_539_n N_A_193_47#_c_617_n 0.00232396f $X=1.375 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_540_n N_A_193_47#_c_617_n 0.00232396f $X=2.215 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_542_n N_A_193_47#_c_617_n 0.00970544f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_540_n N_A_193_47#_c_656_n 0.0112554f $X=2.215 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_542_n N_A_193_47#_c_656_n 0.00644035f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_M1010_d N_A_193_47#_c_612_n 0.00522868f $X=2.245 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_VGND_c_537_n N_A_193_47#_c_612_n 0.0214727f $X=2.38 $Y=0.36 $X2=0 $Y2=0
cc_325 N_VGND_c_540_n N_A_193_47#_c_612_n 0.00232396f $X=2.215 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_541_n N_A_193_47#_c_612_n 0.0031369f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_542_n N_A_193_47#_c_612_n 0.0106541f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_537_n N_A_193_47#_c_613_n 0.00154657f $X=2.38 $Y=0.36 $X2=0
+ $Y2=0
cc_329 N_VGND_c_537_n N_A_193_47#_c_614_n 0.0178768f $X=2.38 $Y=0.36 $X2=0 $Y2=0
cc_330 N_VGND_c_541_n N_A_193_47#_c_614_n 0.0196468f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_331 N_VGND_c_542_n N_A_193_47#_c_614_n 0.0109256f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_332 N_VGND_c_541_n N_A_193_47#_c_615_n 0.11167f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_542_n N_A_193_47#_c_615_n 0.0701989f $X=4.83 $Y=0 $X2=0 $Y2=0

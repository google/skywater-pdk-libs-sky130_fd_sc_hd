* File: sky130_fd_sc_hd__and3b_1.spice
* Created: Thu Aug 27 14:07:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and3b_1.spice.pex"
.subckt sky130_fd_sc_hd__and3b_1  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_A_109_93#_M1008_d N_A_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.10785 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_296_53# N_A_109_93#_M1005_g N_A_209_311#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.107825 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 A_368_53# N_B_M1006_g A_296_53# VNB NSHORT L=0.15 W=0.42 AD=0.05355
+ AS=0.0441 PD=0.675 PS=0.63 NRD=20.712 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g A_368_53# VNB NSHORT L=0.15 W=0.42
+ AD=0.0959916 AS=0.05355 PD=0.84785 PS=0.675 NRD=44.28 NRS=20.712 M=1 R=2.8
+ SA=75000.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_209_311#_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.148558 PD=1.82 PS=1.31215 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_109_93#_M1004_d N_A_N_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1087 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_109_93#_M1003_g N_A_209_311#_M1003_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1085 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_209_311#_M1000_d N_B_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.074375 AS=0.0567 PD=0.815 PS=0.69 NRD=21.0987 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_A_209_311#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0841331 AS=0.074375 PD=0.789718 PS=0.815 NRD=68.1423 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1007_d N_A_209_311#_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.200317 PD=2.52 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__and3b_1.spice.SKY130_FD_SC_HD__AND3B_1.pxi"
*
.ends
*
*

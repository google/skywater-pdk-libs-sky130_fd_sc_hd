* File: sky130_fd_sc_hd__o211ai_4.pxi.spice
* Created: Tue Sep  1 19:20:59 2020
* 
x_PM_SKY130_FD_SC_HD__O211AI_4%A1 N_A1_c_106_n N_A1_M1006_g N_A1_M1008_g
+ N_A1_c_107_n N_A1_M1009_g N_A1_M1013_g N_A1_c_108_n N_A1_M1019_g N_A1_M1017_g
+ N_A1_M1029_g N_A1_M1031_g N_A1_c_109_n N_A1_c_124_p N_A1_c_110_n N_A1_c_111_n
+ A1 N_A1_c_132_p N_A1_c_112_n N_A1_c_113_n PM_SKY130_FD_SC_HD__O211AI_4%A1
x_PM_SKY130_FD_SC_HD__O211AI_4%A2 N_A2_c_224_n N_A2_M1005_g N_A2_c_230_n
+ N_A2_M1007_g N_A2_c_225_n N_A2_M1014_g N_A2_c_231_n N_A2_M1010_g N_A2_c_226_n
+ N_A2_M1018_g N_A2_c_232_n N_A2_M1021_g N_A2_c_227_n N_A2_M1028_g N_A2_c_233_n
+ N_A2_M1027_g A2 N_A2_c_228_n N_A2_c_229_n PM_SKY130_FD_SC_HD__O211AI_4%A2
x_PM_SKY130_FD_SC_HD__O211AI_4%B1 N_B1_c_301_n N_B1_M1002_g N_B1_M1001_g
+ N_B1_c_302_n N_B1_M1026_g N_B1_M1003_g N_B1_c_303_n N_B1_M1012_g N_B1_M1011_g
+ N_B1_M1023_g N_B1_M1025_g N_B1_c_331_p N_B1_c_304_n N_B1_c_305_n B1
+ N_B1_c_306_n N_B1_c_307_n N_B1_c_308_n N_B1_c_309_n
+ PM_SKY130_FD_SC_HD__O211AI_4%B1
x_PM_SKY130_FD_SC_HD__O211AI_4%C1 N_C1_c_417_n N_C1_M1016_g N_C1_M1000_g
+ N_C1_c_418_n N_C1_M1020_g N_C1_M1004_g N_C1_c_419_n N_C1_M1022_g N_C1_M1024_g
+ N_C1_c_420_n N_C1_M1015_g N_C1_M1030_g C1 N_C1_c_421_n
+ PM_SKY130_FD_SC_HD__O211AI_4%C1
x_PM_SKY130_FD_SC_HD__O211AI_4%VPWR N_VPWR_M1008_d N_VPWR_M1013_d N_VPWR_M1029_d
+ N_VPWR_M1003_d N_VPWR_M1000_d N_VPWR_M1024_d N_VPWR_M1023_d N_VPWR_c_497_n
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n
+ N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n VPWR N_VPWR_c_511_n
+ N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_516_n
+ N_VPWR_c_496_n PM_SKY130_FD_SC_HD__O211AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O211AI_4%A_110_297# N_A_110_297#_M1008_s
+ N_A_110_297#_M1017_s N_A_110_297#_M1010_s N_A_110_297#_M1027_s
+ N_A_110_297#_c_623_n N_A_110_297#_c_646_n N_A_110_297#_c_629_n
+ N_A_110_297#_c_631_n PM_SKY130_FD_SC_HD__O211AI_4%A_110_297#
x_PM_SKY130_FD_SC_HD__O211AI_4%Y N_Y_M1016_d N_Y_M1022_d N_Y_M1007_d N_Y_M1021_d
+ N_Y_M1001_s N_Y_M1011_s N_Y_M1004_s N_Y_M1030_s N_Y_c_663_n N_Y_c_677_n
+ N_Y_c_678_n N_Y_c_679_n N_Y_c_704_n N_Y_c_665_n N_Y_c_658_n N_Y_c_657_n Y
+ N_Y_c_667_n PM_SKY130_FD_SC_HD__O211AI_4%Y
x_PM_SKY130_FD_SC_HD__O211AI_4%A_27_47# N_A_27_47#_M1006_d N_A_27_47#_M1009_d
+ N_A_27_47#_M1005_d N_A_27_47#_M1018_d N_A_27_47#_M1031_d N_A_27_47#_M1026_s
+ N_A_27_47#_M1025_s N_A_27_47#_c_765_n N_A_27_47#_c_796_n N_A_27_47#_c_778_n
+ N_A_27_47#_c_781_n N_A_27_47#_c_812_n N_A_27_47#_c_766_n N_A_27_47#_c_767_n
+ N_A_27_47#_c_768_n N_A_27_47#_c_785_n N_A_27_47#_c_786_n N_A_27_47#_c_769_n
+ N_A_27_47#_c_789_n N_A_27_47#_c_770_n N_A_27_47#_c_771_n N_A_27_47#_c_772_n
+ PM_SKY130_FD_SC_HD__O211AI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O211AI_4%VGND N_VGND_M1006_s N_VGND_M1019_s N_VGND_M1014_s
+ N_VGND_M1028_s N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n N_VGND_c_908_n
+ N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n
+ N_VGND_c_914_n VGND N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n
+ N_VGND_c_918_n PM_SKY130_FD_SC_HD__O211AI_4%VGND
x_PM_SKY130_FD_SC_HD__O211AI_4%A_806_47# N_A_806_47#_M1002_d N_A_806_47#_M1020_s
+ N_A_806_47#_c_1029_n PM_SKY130_FD_SC_HD__O211AI_4%A_806_47#
cc_1 VNB N_A1_c_106_n 0.0213945f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A1_c_107_n 0.015805f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_A1_c_108_n 0.0162114f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_4 VNB N_A1_c_109_n 0.0091186f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_A1_c_110_n 0.00113785f $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=1.16
cc_6 VNB N_A1_c_111_n 0.0260601f $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=1.16
cc_7 VNB N_A1_c_112_n 0.0550772f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.16
cc_8 VNB N_A1_c_113_n 0.0168629f $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=0.995
cc_9 VNB N_A2_c_224_n 0.0163088f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_10 VNB N_A2_c_225_n 0.0160041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_226_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_12 VNB N_A2_c_227_n 0.0162948f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.985
cc_13 VNB N_A2_c_228_n 0.00191239f $X=-0.19 $Y=-0.24 $X2=3.49 $Y2=1.515
cc_14 VNB N_A2_c_229_n 0.0644386f $X=-0.19 $Y=-0.24 $X2=3.49 $Y2=1.16
cc_15 VNB N_B1_c_301_n 0.0167177f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_16 VNB N_B1_c_302_n 0.0162054f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_17 VNB N_B1_c_303_n 0.0163495f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_18 VNB N_B1_c_304_n 5.01549e-19 $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=1.16
cc_19 VNB N_B1_c_305_n 0.0243404f $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=1.16
cc_20 VNB N_B1_c_306_n 0.0452091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B1_c_307_n 0.0199297f $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=1.325
cc_22 VNB N_B1_c_308_n 0.00276098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B1_c_309_n 0.00356456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C1_c_417_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_25 VNB N_C1_c_418_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_26 VNB N_C1_c_419_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_27 VNB N_C1_c_420_n 0.0167026f $X=-0.19 $Y=-0.24 $X2=3.485 $Y2=1.325
cc_28 VNB N_C1_c_421_n 0.0648698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_496_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_657_n 0.0198554f $X=-0.19 $Y=-0.24 $X2=1.245 $Y2=1.16
cc_31 VNB N_A_27_47#_c_765_n 0.00431558f $X=-0.19 $Y=-0.24 $X2=3.485 $Y2=1.325
cc_32 VNB N_A_27_47#_c_766_n 0.00224113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_767_n 0.00837836f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.16
cc_34 VNB N_A_27_47#_c_768_n 0.00472633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_769_n 4.96561e-19 $X=-0.19 $Y=-0.24 $X2=3.505 $Y2=1.325
cc_36 VNB N_A_27_47#_c_770_n 0.00171161f $X=-0.19 $Y=-0.24 $X2=1.187 $Y2=1.53
cc_37 VNB N_A_27_47#_c_771_n 0.0208627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_772_n 0.0124137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_905_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_40 VNB N_VGND_c_906_n 0.00354152f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.985
cc_41 VNB N_VGND_c_907_n 3.22457e-19 $X=-0.19 $Y=-0.24 $X2=3.485 $Y2=1.985
cc_42 VNB N_VGND_c_908_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=0.56
cc_43 VNB N_VGND_c_909_n 0.0151902f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.202
cc_44 VNB N_VGND_c_910_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_45 VNB N_VGND_c_911_n 0.0156274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_912_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=3.35 $Y2=1.6
cc_47 VNB N_VGND_c_913_n 0.0123154f $X=-0.19 $Y=-0.24 $X2=3.49 $Y2=1.515
cc_48 VNB N_VGND_c_914_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=3.49 $Y2=1.16
cc_49 VNB N_VGND_c_915_n 0.0159537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_916_n 0.105297f $X=-0.19 $Y=-0.24 $X2=1.187 $Y2=1.6
cc_51 VNB N_VGND_c_917_n 0.373734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_918_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_A1_M1008_g 0.0259007f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_54 VPB N_A1_M1013_g 0.017817f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_55 VPB N_A1_M1017_g 0.0181566f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_56 VPB N_A1_M1029_g 0.0179366f $X=-0.19 $Y=1.305 $X2=3.485 $Y2=1.985
cc_57 VPB N_A1_c_109_n 0.00517698f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_58 VPB N_A1_c_110_n 0.00290629f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.16
cc_59 VPB N_A1_c_111_n 0.00654746f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.16
cc_60 VPB N_A1_c_112_n 0.00883016f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.16
cc_61 VPB N_A2_c_230_n 0.0164258f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_62 VPB N_A2_c_231_n 0.0162054f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.56
cc_63 VPB N_A2_c_232_n 0.016204f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=0.56
cc_64 VPB N_A2_c_233_n 0.01642f $X=-0.19 $Y=1.305 $X2=3.485 $Y2=1.325
cc_65 VPB N_A2_c_228_n 7.05409e-19 $X=-0.19 $Y=1.305 $X2=3.49 $Y2=1.515
cc_66 VPB N_A2_c_229_n 0.0203981f $X=-0.19 $Y=1.305 $X2=3.49 $Y2=1.16
cc_67 VPB N_B1_M1001_g 0.0183904f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_68 VPB N_B1_M1003_g 0.0171638f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_69 VPB N_B1_M1011_g 0.0171234f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_70 VPB N_B1_M1023_g 0.0223957f $X=-0.19 $Y=1.305 $X2=3.485 $Y2=1.985
cc_71 VPB N_B1_c_304_n 0.00306156f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.16
cc_72 VPB N_B1_c_305_n 0.00480298f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.16
cc_73 VPB N_B1_c_306_n 0.00832232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B1_c_308_n 0.00496449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B1_c_309_n 0.00271392f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_C1_M1000_g 0.0185674f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_77 VPB N_C1_M1004_g 0.0181261f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_78 VPB N_C1_M1024_g 0.0181272f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.985
cc_79 VPB N_C1_M1030_g 0.0184798f $X=-0.19 $Y=1.305 $X2=3.495 $Y2=0.56
cc_80 VPB C1 0.00709655f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_81 VPB N_C1_c_421_n 0.0114398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_497_n 0.0107202f $X=-0.19 $Y=1.305 $X2=3.485 $Y2=1.325
cc_83 VPB N_VPWR_c_498_n 0.0379377f $X=-0.19 $Y=1.305 $X2=3.485 $Y2=1.985
cc_84 VPB N_VPWR_c_499_n 4.06069e-19 $X=-0.19 $Y=1.305 $X2=3.495 $Y2=0.56
cc_85 VPB N_VPWR_c_500_n 0.00252303f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_86 VPB N_VPWR_c_501_n 3.09901e-19 $X=-0.19 $Y=1.305 $X2=3.49 $Y2=1.515
cc_87 VPB N_VPWR_c_502_n 0.0118594f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.16
cc_88 VPB N_VPWR_c_503_n 3.02679e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_504_n 3.95476e-19 $X=-0.19 $Y=1.305 $X2=1.245 $Y2=1.16
cc_90 VPB N_VPWR_c_505_n 0.0128205f $X=-0.19 $Y=1.305 $X2=1.245 $Y2=1.16
cc_91 VPB N_VPWR_c_506_n 0.0136265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_507_n 0.0523073f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.325
cc_93 VPB N_VPWR_c_508_n 0.0040697f $X=-0.19 $Y=1.305 $X2=1.187 $Y2=1.16
cc_94 VPB N_VPWR_c_509_n 0.0129196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_510_n 0.00436029f $X=-0.19 $Y=1.305 $X2=1.187 $Y2=1.202
cc_96 VPB N_VPWR_c_511_n 0.0149927f $X=-0.19 $Y=1.305 $X2=1.187 $Y2=1.6
cc_97 VPB N_VPWR_c_512_n 0.0117235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_513_n 0.0233778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_514_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_515_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_516_n 0.00442675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_496_n 0.0452394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_Y_c_658_n 0.0266072f $X=-0.19 $Y=1.305 $X2=1.245 $Y2=1.16
cc_104 VPB N_Y_c_657_n 0.00159252f $X=-0.19 $Y=1.305 $X2=1.245 $Y2=1.16
cc_105 VPB Y 0.0207561f $X=-0.19 $Y=1.305 $X2=1.245 $Y2=1.16
cc_106 N_A1_c_108_n N_A2_c_224_n 0.0284954f $X=1.335 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A1_M1017_g N_A2_c_230_n 0.0284954f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A1_c_124_p N_A2_c_230_n 0.0121907f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_109 N_A1_c_124_p N_A2_c_231_n 0.010446f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_110 N_A1_c_124_p N_A2_c_232_n 0.0104926f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_111 N_A1_c_113_n N_A2_c_227_n 0.0252793f $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_c_124_p N_A2_c_233_n 0.010446f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_113 N_A1_c_124_p N_A2_c_228_n 0.0917809f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_114 N_A1_c_110_n N_A2_c_228_n 0.0224261f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A1_c_111_n N_A2_c_228_n 0.00155774f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_c_132_p N_A2_c_228_n 0.0140188f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A1_c_112_n N_A2_c_228_n 0.00115693f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A1_M1029_g N_A2_c_229_n 0.0451359f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A1_c_124_p N_A2_c_229_n 0.00717248f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_120 N_A1_c_110_n N_A2_c_229_n 0.00462885f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A1_c_111_n N_A2_c_229_n 0.021402f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A1_c_132_p N_A2_c_229_n 0.00233113f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A1_c_112_n N_A2_c_229_n 0.0284954f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A1_c_113_n N_B1_c_301_n 0.0210245f $X=3.505 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_125 N_A1_M1029_g N_B1_M1001_g 0.0375208f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A1_c_124_p N_B1_M1001_g 0.00195545f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_127 N_A1_c_110_n N_B1_M1001_g 0.00128836f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A1_c_110_n N_B1_c_306_n 3.2456e-19 $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A1_c_111_n N_B1_c_306_n 0.0206161f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_M1029_g N_B1_c_308_n 2.93401e-19 $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_c_110_n N_B1_c_308_n 0.0347784f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A1_c_111_n N_B1_c_308_n 0.00218633f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A1_c_110_n N_B1_c_309_n 0.00301223f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A1_c_132_p N_VPWR_M1013_d 0.00218345f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A1_c_124_p N_VPWR_M1029_d 0.00278501f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_136 N_A1_c_110_n N_VPWR_M1029_d 4.41398e-19 $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_M1008_g N_VPWR_c_498_n 0.00574377f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_M1008_g N_VPWR_c_499_n 0.00106903f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_M1013_g N_VPWR_c_499_n 0.00784974f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_M1017_g N_VPWR_c_499_n 0.0073891f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_M1029_g N_VPWR_c_500_n 0.00286483f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A1_M1017_g N_VPWR_c_507_n 0.00351072f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A1_M1029_g N_VPWR_c_507_n 0.00418369f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A1_M1008_g N_VPWR_c_511_n 0.00585385f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1013_g N_VPWR_c_511_n 0.00351072f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1008_g N_VPWR_c_496_n 0.0115115f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_M1013_g N_VPWR_c_496_n 0.00411677f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A1_M1017_g N_VPWR_c_496_n 0.00414308f $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A1_M1029_g N_VPWR_c_496_n 0.00585583f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A1_c_124_p N_A_110_297#_M1017_s 0.00543081f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_151 N_A1_c_124_p N_A_110_297#_M1010_s 0.00330122f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_152 N_A1_c_124_p N_A_110_297#_M1027_s 0.00766992f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_153 N_A1_c_110_n N_A_110_297#_M1027_s 3.70432e-19 $X=3.505 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A1_M1013_g N_A_110_297#_c_623_n 0.0112986f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A1_M1017_g N_A_110_297#_c_623_n 0.0101703f $X=1.335 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A1_c_109_n N_A_110_297#_c_623_n 0.00420181f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_157 N_A1_c_124_p N_A_110_297#_c_623_n 0.00994603f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_158 N_A1_c_132_p N_A_110_297#_c_623_n 0.0190872f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_c_112_n N_A_110_297#_c_623_n 3.31404e-19 $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A1_M1029_g N_A_110_297#_c_629_n 0.00250134f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A1_c_124_p N_A_110_297#_c_629_n 0.00280123f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_162 N_A1_c_109_n N_A_110_297#_c_631_n 0.00684462f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_163 N_A1_c_112_n N_A_110_297#_c_631_n 5.81512e-19 $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A1_c_124_p N_Y_M1007_d 0.00330122f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_165 N_A1_c_124_p N_Y_M1021_d 0.00330122f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_166 N_A1_M1017_g N_Y_c_663_n 4.52533e-19 $X=1.335 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_c_124_p N_Y_c_663_n 0.0830965f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_168 N_A1_M1029_g N_Y_c_665_n 0.00745179f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A1_c_124_p N_Y_c_665_n 0.0125836f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_170 N_A1_M1029_g N_Y_c_667_n 0.0069938f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A1_c_111_n N_Y_c_667_n 0.00120879f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A1_c_106_n N_A_27_47#_c_765_n 0.0127311f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_107_n N_A_27_47#_c_765_n 0.01245f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_109_n N_A_27_47#_c_765_n 0.0421759f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A1_c_132_p N_A_27_47#_c_765_n 0.00474248f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A1_c_112_n N_A_27_47#_c_765_n 0.00249616f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A1_c_110_n N_A_27_47#_c_778_n 0.0138653f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A1_c_111_n N_A_27_47#_c_778_n 0.00254845f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A1_c_113_n N_A_27_47#_c_778_n 0.0106643f $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_113_n N_A_27_47#_c_781_n 3.27348e-19 $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_108_n N_A_27_47#_c_768_n 0.010776f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_124_p N_A_27_47#_c_768_n 0.0071519f $X=3.35 $Y=1.6 $X2=0 $Y2=0
cc_183 N_A1_c_132_p N_A_27_47#_c_768_n 0.0124947f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A1_c_108_n N_A_27_47#_c_785_n 2.19873e-19 $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A1_c_113_n N_A_27_47#_c_786_n 4.25317e-19 $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A1_c_108_n N_A_27_47#_c_769_n 0.00200012f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_113_n N_A_27_47#_c_769_n 0.0024487f $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_107_n N_A_27_47#_c_789_n 0.00422671f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_108_n N_A_27_47#_c_789_n 0.00209019f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A1_c_132_p N_A_27_47#_c_789_n 9.06457e-19 $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A1_c_107_n N_A_27_47#_c_770_n 0.00160224f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_108_n N_A_27_47#_c_770_n 0.00150782f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_132_p N_A_27_47#_c_770_n 0.0176035f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A1_c_112_n N_A_27_47#_c_770_n 0.00253413f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A1_c_106_n N_VGND_c_905_n 0.01411f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_107_n N_VGND_c_905_n 0.0078413f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_108_n N_VGND_c_905_n 0.00101736f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_108_n N_VGND_c_906_n 0.00152327f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_113_n N_VGND_c_908_n 0.0067518f $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_107_n N_VGND_c_909_n 0.0035231f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_108_n N_VGND_c_909_n 0.00433717f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A1_c_106_n N_VGND_c_915_n 0.0035231f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_113_n N_VGND_c_916_n 0.0038055f $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_106_n N_VGND_c_917_n 0.00510533f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A1_c_107_n N_VGND_c_917_n 0.00413686f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A1_c_108_n N_VGND_c_917_n 0.00495538f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_c_113_n N_VGND_c_917_n 0.00374445f $X=3.505 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A2_c_230_n N_VPWR_c_499_n 0.00121908f $X=1.765 $Y=1.375 $X2=0 $Y2=0
cc_209 N_A2_c_230_n N_VPWR_c_507_n 0.00357877f $X=1.765 $Y=1.375 $X2=0 $Y2=0
cc_210 N_A2_c_231_n N_VPWR_c_507_n 0.00357877f $X=2.195 $Y=1.375 $X2=0 $Y2=0
cc_211 N_A2_c_232_n N_VPWR_c_507_n 0.00357877f $X=2.625 $Y=1.375 $X2=0 $Y2=0
cc_212 N_A2_c_233_n N_VPWR_c_507_n 0.00357877f $X=3.055 $Y=1.375 $X2=0 $Y2=0
cc_213 N_A2_c_230_n N_VPWR_c_496_n 0.00534514f $X=1.765 $Y=1.375 $X2=0 $Y2=0
cc_214 N_A2_c_231_n N_VPWR_c_496_n 0.00527894f $X=2.195 $Y=1.375 $X2=0 $Y2=0
cc_215 N_A2_c_232_n N_VPWR_c_496_n 0.00527894f $X=2.625 $Y=1.375 $X2=0 $Y2=0
cc_216 N_A2_c_233_n N_VPWR_c_496_n 0.00530427f $X=3.055 $Y=1.375 $X2=0 $Y2=0
cc_217 N_A2_c_230_n N_A_110_297#_c_629_n 0.0107771f $X=1.765 $Y=1.375 $X2=0
+ $Y2=0
cc_218 N_A2_c_231_n N_A_110_297#_c_629_n 0.00816381f $X=2.195 $Y=1.375 $X2=0
+ $Y2=0
cc_219 N_A2_c_232_n N_A_110_297#_c_629_n 0.00821592f $X=2.625 $Y=1.375 $X2=0
+ $Y2=0
cc_220 N_A2_c_233_n N_A_110_297#_c_629_n 0.00821592f $X=3.055 $Y=1.375 $X2=0
+ $Y2=0
cc_221 N_A2_c_230_n N_Y_c_663_n 0.00437939f $X=1.765 $Y=1.375 $X2=0 $Y2=0
cc_222 N_A2_c_231_n N_Y_c_663_n 0.0105629f $X=2.195 $Y=1.375 $X2=0 $Y2=0
cc_223 N_A2_c_232_n N_Y_c_663_n 0.0105629f $X=2.625 $Y=1.375 $X2=0 $Y2=0
cc_224 N_A2_c_233_n N_Y_c_663_n 0.0104941f $X=3.055 $Y=1.375 $X2=0 $Y2=0
cc_225 N_A2_c_224_n N_A_27_47#_c_796_n 0.00252062f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A2_c_225_n N_A_27_47#_c_796_n 0.0113837f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A2_c_226_n N_A_27_47#_c_796_n 0.0113837f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_227_n N_A_27_47#_c_796_n 0.00164133f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A2_c_228_n N_A_27_47#_c_796_n 0.0672087f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A2_c_229_n N_A_27_47#_c_796_n 0.00748111f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_231 N_A2_c_224_n N_A_27_47#_c_768_n 0.00731508f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A2_c_228_n N_A_27_47#_c_768_n 0.00618622f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A2_c_224_n N_A_27_47#_c_785_n 0.00280332f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_227_n N_A_27_47#_c_786_n 0.00921008f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_224_n N_A_27_47#_c_769_n 0.00356497f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A2_c_225_n N_A_27_47#_c_769_n 0.00305544f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A2_c_226_n N_A_27_47#_c_769_n 0.00305544f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A2_c_227_n N_A_27_47#_c_769_n 0.00306494f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A2_c_224_n N_A_27_47#_c_789_n 2.0792e-19 $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_224_n N_VGND_c_906_n 0.00207974f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A2_c_224_n N_VGND_c_907_n 0.00109579f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A2_c_225_n N_VGND_c_907_n 0.0078976f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A2_c_226_n N_VGND_c_907_n 0.00748051f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A2_c_227_n N_VGND_c_907_n 0.00104544f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A2_c_226_n N_VGND_c_908_n 0.00104544f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A2_c_227_n N_VGND_c_908_n 0.00748967f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A2_c_224_n N_VGND_c_911_n 0.00429337f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A2_c_225_n N_VGND_c_911_n 0.0035231f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A2_c_226_n N_VGND_c_913_n 0.0035231f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A2_c_227_n N_VGND_c_913_n 0.0035231f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A2_c_224_n N_VGND_c_917_n 0.00495923f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A2_c_225_n N_VGND_c_917_n 0.00341787f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A2_c_226_n N_VGND_c_917_n 0.00341787f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A2_c_227_n N_VGND_c_917_n 0.00341787f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_255 N_B1_c_303_n N_C1_c_417_n 0.0340492f $X=4.815 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_256 N_B1_M1011_g N_C1_M1000_g 0.0340492f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B1_c_331_p N_C1_M1000_g 0.0149047f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_258 N_B1_c_331_p N_C1_M1004_g 0.0103677f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_259 N_B1_c_331_p N_C1_M1024_g 0.0103677f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_260 N_B1_c_307_n N_C1_c_420_n 0.0345564f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B1_M1023_g N_C1_M1030_g 0.0432628f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B1_c_331_p N_C1_M1030_g 0.0142939f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_263 N_B1_c_304_n N_C1_M1030_g 0.00279207f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_c_331_p C1 0.0696674f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_265 N_B1_c_304_n C1 0.0104854f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B1_c_305_n C1 7.07237e-19 $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B1_c_306_n C1 2.09507e-19 $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B1_c_309_n C1 0.0127619f $X=4.975 $Y=1.34 $X2=0 $Y2=0
cc_269 N_B1_c_331_p N_C1_c_421_n 0.00179982f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_270 N_B1_c_304_n N_C1_c_421_n 0.00156121f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B1_c_305_n N_C1_c_421_n 0.0221532f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_306_n N_C1_c_421_n 0.0340492f $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B1_c_309_n N_C1_c_421_n 0.00972946f $X=4.975 $Y=1.34 $X2=0 $Y2=0
cc_274 N_B1_c_309_n N_VPWR_M1003_d 0.00184669f $X=4.975 $Y=1.34 $X2=0 $Y2=0
cc_275 N_B1_c_331_p N_VPWR_M1000_d 0.00309215f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_276 N_B1_c_331_p N_VPWR_M1024_d 0.00312412f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_277 N_B1_M1001_g N_VPWR_c_500_n 0.00767323f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1003_g N_VPWR_c_500_n 0.00138479f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_M1001_g N_VPWR_c_501_n 0.00105652f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B1_M1003_g N_VPWR_c_501_n 0.00775841f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B1_M1011_g N_VPWR_c_501_n 0.00755691f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B1_M1011_g N_VPWR_c_502_n 0.00351072f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_283 N_B1_M1011_g N_VPWR_c_503_n 0.00104745f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B1_M1023_g N_VPWR_c_504_n 0.00209959f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B1_M1023_g N_VPWR_c_506_n 0.00888872f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_286 N_B1_M1001_g N_VPWR_c_509_n 0.00418493f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_287 N_B1_M1003_g N_VPWR_c_509_n 0.00351072f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_288 N_B1_M1023_g N_VPWR_c_513_n 0.00422112f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_289 N_B1_M1001_g N_VPWR_c_496_n 0.00487066f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_290 N_B1_M1003_g N_VPWR_c_496_n 0.00411677f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_291 N_B1_M1011_g N_VPWR_c_496_n 0.00411763f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_292 N_B1_M1023_g N_VPWR_c_496_n 0.0072343f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_293 N_B1_c_331_p N_Y_M1011_s 0.00619908f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_294 N_B1_c_309_n N_Y_M1011_s 7.29311e-19 $X=4.975 $Y=1.34 $X2=0 $Y2=0
cc_295 N_B1_c_331_p N_Y_M1004_s 0.00312412f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_296 N_B1_c_331_p N_Y_M1030_s 0.00750015f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_297 N_B1_c_307_n N_Y_c_677_n 0.00229246f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B1_c_307_n N_Y_c_678_n 0.00348426f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_304_n N_Y_c_679_n 0.0102076f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_300 N_B1_c_305_n N_Y_c_679_n 0.00220272f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B1_c_307_n N_Y_c_679_n 0.0138791f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B1_M1001_g N_Y_c_665_n 2.55386e-19 $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_303 N_B1_M1023_g N_Y_c_657_n 0.00271557f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_304 N_B1_c_304_n N_Y_c_657_n 0.0379564f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_305 N_B1_c_305_n N_Y_c_657_n 0.00754311f $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_306 N_B1_c_307_n N_Y_c_657_n 0.00608305f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_M1003_g Y 0.0116082f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_308 N_B1_M1011_g Y 0.0115863f $X=4.815 $Y=1.985 $X2=0 $Y2=0
cc_309 N_B1_M1023_g Y 0.0213536f $X=6.915 $Y=1.985 $X2=0 $Y2=0
cc_310 N_B1_c_331_p Y 0.0117161f $X=6.83 $Y=1.6 $X2=0 $Y2=0
cc_311 N_B1_c_305_n Y 8.75512e-19 $X=6.915 $Y=1.16 $X2=0 $Y2=0
cc_312 N_B1_c_306_n Y 8.54516e-19 $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_313 N_B1_c_309_n Y 0.137438f $X=4.975 $Y=1.34 $X2=0 $Y2=0
cc_314 N_B1_M1001_g N_Y_c_667_n 0.0115403f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_315 N_B1_c_308_n N_Y_c_667_n 0.0153926f $X=4.26 $Y=1.34 $X2=0 $Y2=0
cc_316 N_B1_c_308_n N_A_27_47#_c_778_n 0.00205362f $X=4.26 $Y=1.34 $X2=0 $Y2=0
cc_317 N_B1_c_301_n N_A_27_47#_c_812_n 0.00938584f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_302_n N_A_27_47#_c_812_n 0.00756577f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B1_c_303_n N_A_27_47#_c_812_n 0.0059805f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_320 N_B1_c_308_n N_A_27_47#_c_812_n 0.00251253f $X=4.26 $Y=1.34 $X2=0 $Y2=0
cc_321 N_B1_c_307_n N_A_27_47#_c_766_n 0.00335865f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B1_c_301_n N_A_27_47#_c_769_n 0.00228237f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B1_c_302_n N_A_27_47#_c_769_n 0.00199894f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B1_c_303_n N_A_27_47#_c_769_n 0.00228446f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_325 N_B1_c_307_n N_A_27_47#_c_769_n 0.00284618f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B1_c_308_n N_A_27_47#_c_769_n 0.00570535f $X=4.26 $Y=1.34 $X2=0 $Y2=0
cc_327 N_B1_c_307_n N_A_27_47#_c_771_n 8.38249e-19 $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B1_c_307_n N_A_27_47#_c_772_n 9.94574e-19 $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B1_c_301_n N_VGND_c_908_n 0.00112406f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B1_c_301_n N_VGND_c_916_n 0.00357877f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B1_c_302_n N_VGND_c_916_n 0.00357877f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B1_c_303_n N_VGND_c_916_n 0.00357877f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B1_c_307_n N_VGND_c_916_n 0.00404461f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B1_c_301_n N_VGND_c_917_n 0.00492027f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B1_c_302_n N_VGND_c_917_n 0.00478374f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B1_c_303_n N_VGND_c_917_n 0.0047846f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B1_c_307_n N_VGND_c_917_n 0.0063646f $X=6.915 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B1_c_301_n N_A_806_47#_c_1029_n 0.00265506f $X=3.955 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_B1_c_302_n N_A_806_47#_c_1029_n 0.00872107f $X=4.385 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_B1_c_303_n N_A_806_47#_c_1029_n 0.0107784f $X=4.815 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_B1_c_306_n N_A_806_47#_c_1029_n 0.00446133f $X=4.815 $Y=1.16 $X2=0
+ $Y2=0
cc_342 N_B1_c_308_n N_A_806_47#_c_1029_n 0.0575102f $X=4.26 $Y=1.34 $X2=0 $Y2=0
cc_343 N_C1_M1000_g N_VPWR_c_501_n 0.00103591f $X=5.235 $Y=1.985 $X2=0 $Y2=0
cc_344 N_C1_M1000_g N_VPWR_c_502_n 0.00337001f $X=5.235 $Y=1.985 $X2=0 $Y2=0
cc_345 N_C1_M1000_g N_VPWR_c_503_n 0.00778794f $X=5.235 $Y=1.985 $X2=0 $Y2=0
cc_346 N_C1_M1004_g N_VPWR_c_503_n 0.00775994f $X=5.655 $Y=1.985 $X2=0 $Y2=0
cc_347 N_C1_M1024_g N_VPWR_c_503_n 0.0010441f $X=6.075 $Y=1.985 $X2=0 $Y2=0
cc_348 N_C1_M1004_g N_VPWR_c_504_n 0.00104438f $X=5.655 $Y=1.985 $X2=0 $Y2=0
cc_349 N_C1_M1024_g N_VPWR_c_504_n 0.00775994f $X=6.075 $Y=1.985 $X2=0 $Y2=0
cc_350 N_C1_M1030_g N_VPWR_c_504_n 0.00947076f $X=6.495 $Y=1.985 $X2=0 $Y2=0
cc_351 N_C1_M1004_g N_VPWR_c_512_n 0.00337001f $X=5.655 $Y=1.985 $X2=0 $Y2=0
cc_352 N_C1_M1024_g N_VPWR_c_512_n 0.00337001f $X=6.075 $Y=1.985 $X2=0 $Y2=0
cc_353 N_C1_M1030_g N_VPWR_c_513_n 0.00322931f $X=6.495 $Y=1.985 $X2=0 $Y2=0
cc_354 N_C1_M1000_g N_VPWR_c_496_n 0.00397658f $X=5.235 $Y=1.985 $X2=0 $Y2=0
cc_355 N_C1_M1004_g N_VPWR_c_496_n 0.00394833f $X=5.655 $Y=1.985 $X2=0 $Y2=0
cc_356 N_C1_M1024_g N_VPWR_c_496_n 0.00394833f $X=6.075 $Y=1.985 $X2=0 $Y2=0
cc_357 N_C1_M1030_g N_VPWR_c_496_n 0.00383553f $X=6.495 $Y=1.985 $X2=0 $Y2=0
cc_358 N_C1_c_417_n N_Y_c_677_n 0.00307758f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_359 N_C1_c_418_n N_Y_c_677_n 0.00717095f $X=5.655 $Y=0.995 $X2=0 $Y2=0
cc_360 N_C1_c_419_n N_Y_c_677_n 0.00717095f $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_361 N_C1_c_420_n N_Y_c_677_n 0.00877277f $X=6.495 $Y=0.995 $X2=0 $Y2=0
cc_362 C1 N_Y_c_677_n 0.00324806f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_363 N_C1_c_421_n N_Y_c_677_n 0.00142423f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_364 N_C1_c_419_n N_Y_c_678_n 0.00105938f $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_365 N_C1_c_420_n N_Y_c_678_n 0.00544982f $X=6.495 $Y=0.995 $X2=0 $Y2=0
cc_366 N_C1_c_419_n N_Y_c_704_n 2.11895e-19 $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_367 N_C1_c_420_n N_Y_c_704_n 0.00484835f $X=6.495 $Y=0.995 $X2=0 $Y2=0
cc_368 N_C1_M1000_g Y 0.0114731f $X=5.235 $Y=1.985 $X2=0 $Y2=0
cc_369 N_C1_M1004_g Y 0.0114731f $X=5.655 $Y=1.985 $X2=0 $Y2=0
cc_370 N_C1_M1024_g Y 0.0114731f $X=6.075 $Y=1.985 $X2=0 $Y2=0
cc_371 N_C1_M1030_g Y 0.0114301f $X=6.495 $Y=1.985 $X2=0 $Y2=0
cc_372 N_C1_c_417_n N_A_27_47#_c_812_n 6.02163e-19 $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_373 N_C1_c_417_n N_A_27_47#_c_769_n 0.0033487f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_374 N_C1_c_418_n N_A_27_47#_c_769_n 0.00201201f $X=5.655 $Y=0.995 $X2=0 $Y2=0
cc_375 N_C1_c_419_n N_A_27_47#_c_769_n 0.00201201f $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_376 N_C1_c_420_n N_A_27_47#_c_769_n 0.0056229f $X=6.495 $Y=0.995 $X2=0 $Y2=0
cc_377 C1 N_A_27_47#_c_769_n 0.00732371f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_378 N_C1_c_421_n N_A_27_47#_c_769_n 0.00188106f $X=6.495 $Y=1.16 $X2=0 $Y2=0
cc_379 N_C1_c_417_n N_VGND_c_916_n 0.00412276f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_380 N_C1_c_418_n N_VGND_c_916_n 0.00361001f $X=5.655 $Y=0.995 $X2=0 $Y2=0
cc_381 N_C1_c_419_n N_VGND_c_916_n 0.00361001f $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_382 N_C1_c_420_n N_VGND_c_916_n 0.00360994f $X=6.495 $Y=0.995 $X2=0 $Y2=0
cc_383 N_C1_c_417_n N_VGND_c_917_n 0.00495007f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_384 N_C1_c_418_n N_VGND_c_917_n 0.00473164f $X=5.655 $Y=0.995 $X2=0 $Y2=0
cc_385 N_C1_c_419_n N_VGND_c_917_n 0.00473164f $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_386 N_C1_c_420_n N_VGND_c_917_n 0.00488265f $X=6.495 $Y=0.995 $X2=0 $Y2=0
cc_387 N_C1_c_417_n N_A_806_47#_c_1029_n 0.0161813f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_388 N_C1_c_418_n N_A_806_47#_c_1029_n 0.00914325f $X=5.655 $Y=0.995 $X2=0
+ $Y2=0
cc_389 N_C1_c_419_n N_A_806_47#_c_1029_n 0.007672f $X=6.075 $Y=0.995 $X2=0 $Y2=0
cc_390 C1 N_A_806_47#_c_1029_n 0.032575f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_391 N_C1_c_421_n N_A_806_47#_c_1029_n 0.00417921f $X=6.495 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_496_n N_A_110_297#_M1008_s 0.00311082f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_393 N_VPWR_c_496_n N_A_110_297#_M1017_s 0.00239971f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_496_n N_A_110_297#_M1010_s 0.00223258f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_496_n N_A_110_297#_M1027_s 0.00223258f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_M1013_d N_A_110_297#_c_623_n 0.00367112f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_499_n N_A_110_297#_c_623_n 0.0158375f $X=1.12 $Y=2.36 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_507_n N_A_110_297#_c_623_n 0.0025909f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_511_n N_A_110_297#_c_623_n 0.00269405f $X=0.955 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_496_n N_A_110_297#_c_623_n 0.0103519f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_507_n N_A_110_297#_c_646_n 0.0119601f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_496_n N_A_110_297#_c_646_n 0.00687765f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_507_n N_A_110_297#_c_629_n 0.0989961f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_496_n N_A_110_297#_c_629_n 0.0640639f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_511_n N_A_110_297#_c_631_n 0.00457776f $X=0.955 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_496_n N_A_110_297#_c_631_n 0.00686321f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_496_n N_Y_M1007_d 0.00224864f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_496_n N_Y_M1021_d 0.00224864f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_496_n N_Y_M1001_s 0.00320715f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_496_n N_Y_M1011_s 0.00307577f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_496_n N_Y_M1004_s 0.00307577f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_496_n N_Y_M1030_s 0.00307577f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_c_496_n N_Y_c_663_n 0.00416708f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_507_n N_Y_c_665_n 6.14891e-19 $X=3.615 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_M1023_d N_Y_c_658_n 0.00394416f $X=6.99 $Y=1.485 $X2=0 $Y2=0
cc_416 N_VPWR_M1003_d Y 0.0033902f $X=4.46 $Y=1.485 $X2=0 $Y2=0
cc_417 N_VPWR_M1000_d Y 0.00315804f $X=5.31 $Y=1.485 $X2=0 $Y2=0
cc_418 N_VPWR_M1024_d Y 0.00319039f $X=6.15 $Y=1.485 $X2=0 $Y2=0
cc_419 N_VPWR_M1023_d Y 0.0331671f $X=6.99 $Y=1.485 $X2=0 $Y2=0
cc_420 N_VPWR_c_501_n Y 0.0163189f $X=4.6 $Y=2.36 $X2=0 $Y2=0
cc_421 N_VPWR_c_502_n Y 0.0083745f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_c_503_n Y 0.0162695f $X=5.445 $Y=2.36 $X2=0 $Y2=0
cc_423 N_VPWR_c_504_n Y 0.0166335f $X=6.285 $Y=2.36 $X2=0 $Y2=0
cc_424 N_VPWR_c_506_n Y 0.0252336f $X=7.52 $Y=2.36 $X2=0 $Y2=0
cc_425 N_VPWR_c_509_n Y 0.00631693f $X=4.435 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_c_512_n Y 0.00828666f $X=6.12 $Y=2.72 $X2=0 $Y2=0
cc_427 N_VPWR_c_513_n Y 0.0150977f $X=7.355 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_496_n Y 0.0695918f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_429 N_VPWR_M1029_d N_Y_c_667_n 0.00822541f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_430 N_VPWR_c_500_n N_Y_c_667_n 0.0162461f $X=3.72 $Y=2.36 $X2=0 $Y2=0
cc_431 N_VPWR_c_507_n N_Y_c_667_n 0.0017323f $X=3.615 $Y=2.72 $X2=0 $Y2=0
cc_432 N_VPWR_c_509_n N_Y_c_667_n 0.00218329f $X=4.435 $Y=2.72 $X2=0 $Y2=0
cc_433 N_VPWR_c_496_n N_Y_c_667_n 0.00811531f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_434 N_A_110_297#_c_629_n N_Y_M1007_d 0.00333945f $X=3.27 $Y=2.36 $X2=0.475
+ $Y2=0.56
cc_435 N_A_110_297#_c_629_n N_Y_M1021_d 0.00333945f $X=3.27 $Y=2.36 $X2=0.475
+ $Y2=1.325
cc_436 N_A_110_297#_M1010_s N_Y_c_663_n 0.00337918f $X=2.27 $Y=1.485 $X2=0 $Y2=0
cc_437 N_A_110_297#_M1027_s N_Y_c_663_n 0.00327214f $X=3.13 $Y=1.485 $X2=0 $Y2=0
cc_438 N_A_110_297#_c_629_n N_Y_c_663_n 0.0807669f $X=3.27 $Y=2.36 $X2=0 $Y2=0
cc_439 N_Y_c_679_n N_A_27_47#_M1025_s 0.0141187f $X=7.17 $Y=0.74 $X2=0 $Y2=0
cc_440 N_Y_c_657_n N_A_27_47#_M1025_s 0.0033607f $X=7.425 $Y=1.34 $X2=0 $Y2=0
cc_441 N_Y_c_677_n N_A_27_47#_c_812_n 0.004097f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_442 N_Y_c_677_n N_A_27_47#_c_766_n 0.00880632f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_443 N_Y_c_678_n N_A_27_47#_c_766_n 0.00129806f $X=6.65 $Y=0.655 $X2=0 $Y2=0
cc_444 N_Y_c_679_n N_A_27_47#_c_766_n 0.0210046f $X=7.17 $Y=0.74 $X2=0 $Y2=0
cc_445 N_Y_M1016_d N_A_27_47#_c_769_n 0.00195079f $X=5.31 $Y=0.235 $X2=0 $Y2=0
cc_446 N_Y_M1022_d N_A_27_47#_c_769_n 0.00306981f $X=6.15 $Y=0.235 $X2=0 $Y2=0
cc_447 N_Y_c_677_n N_A_27_47#_c_769_n 0.0293204f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_448 N_Y_c_678_n N_A_27_47#_c_769_n 0.0170874f $X=6.65 $Y=0.655 $X2=0 $Y2=0
cc_449 N_Y_c_679_n N_A_27_47#_c_769_n 0.0183128f $X=7.17 $Y=0.74 $X2=0 $Y2=0
cc_450 N_Y_c_677_n N_VGND_c_916_n 0.0738943f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_451 N_Y_c_679_n N_VGND_c_916_n 0.00321471f $X=7.17 $Y=0.74 $X2=0 $Y2=0
cc_452 N_Y_M1016_d N_VGND_c_917_n 0.00121737f $X=5.31 $Y=0.235 $X2=0 $Y2=0
cc_453 N_Y_M1022_d N_VGND_c_917_n 0.00121737f $X=6.15 $Y=0.235 $X2=0 $Y2=0
cc_454 N_Y_c_677_n N_VGND_c_917_n 0.0135794f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_455 N_Y_c_677_n N_A_806_47#_M1020_s 0.00232151f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_456 N_Y_M1016_d N_A_806_47#_c_1029_n 0.00323238f $X=5.31 $Y=0.235 $X2=0 $Y2=0
cc_457 N_Y_c_677_n N_A_806_47#_c_1029_n 0.0395983f $X=6.565 $Y=0.36 $X2=0 $Y2=0
cc_458 N_Y_c_677_n A_978_47# 0.0030005f $X=6.565 $Y=0.36 $X2=-0.19 $Y2=-0.24
cc_459 N_Y_c_678_n A_978_47# 0.00275744f $X=6.65 $Y=0.655 $X2=-0.19 $Y2=-0.24
cc_460 N_Y_c_679_n A_978_47# 0.00378718f $X=7.17 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_461 N_Y_c_704_n A_978_47# 0.00475485f $X=6.735 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_462 N_A_27_47#_c_765_n N_VGND_M1006_s 0.0017606f $X=1.025 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_463 N_A_27_47#_c_768_n N_VGND_M1019_s 0.00158929f $X=1.775 $Y=0.765 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_769_n N_VGND_M1019_s 0.00270346f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_465 N_A_27_47#_c_796_n N_VGND_M1014_s 0.0032959f $X=3.01 $Y=0.745 $X2=0 $Y2=0
cc_466 N_A_27_47#_c_769_n N_VGND_M1014_s 0.00201521f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_467 N_A_27_47#_c_778_n N_VGND_M1028_s 0.00776529f $X=3.605 $Y=0.71 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_769_n N_VGND_M1028_s 0.00208718f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_469 N_A_27_47#_c_765_n N_VGND_c_905_n 0.0156621f $X=1.025 $Y=0.765 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_789_n N_VGND_c_905_n 0.00165084f $X=1.3 $Y=0.51 $X2=0 $Y2=0
cc_471 N_A_27_47#_c_770_n N_VGND_c_905_n 9.59647e-19 $X=1.155 $Y=0.51 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_768_n N_VGND_c_906_n 0.0109253f $X=1.775 $Y=0.765 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_769_n N_VGND_c_906_n 0.00872737f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_474 N_A_27_47#_c_789_n N_VGND_c_906_n 0.00131174f $X=1.3 $Y=0.51 $X2=0 $Y2=0
cc_475 N_A_27_47#_c_770_n N_VGND_c_906_n 0.00248803f $X=1.155 $Y=0.51 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_796_n N_VGND_c_907_n 0.0149288f $X=3.01 $Y=0.745 $X2=0 $Y2=0
cc_477 N_A_27_47#_c_769_n N_VGND_c_907_n 0.00769506f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_478 N_A_27_47#_c_781_n N_VGND_c_908_n 0.00723147f $X=3.835 $Y=0.355 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_786_n N_VGND_c_908_n 0.0147053f $X=3.13 $Y=0.745 $X2=0 $Y2=0
cc_480 N_A_27_47#_c_769_n N_VGND_c_908_n 0.00763013f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_481 N_A_27_47#_c_765_n N_VGND_c_909_n 0.00259536f $X=1.025 $Y=0.765 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_768_n N_VGND_c_909_n 0.00251741f $X=1.775 $Y=0.765 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_769_n N_VGND_c_909_n 4.86291e-19 $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_484 N_A_27_47#_c_789_n N_VGND_c_909_n 8.48275e-19 $X=1.3 $Y=0.51 $X2=0 $Y2=0
cc_485 N_A_27_47#_c_770_n N_VGND_c_909_n 0.00700829f $X=1.155 $Y=0.51 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_768_n N_VGND_c_911_n 0.00152824f $X=1.775 $Y=0.765 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_785_n N_VGND_c_911_n 0.00671444f $X=1.795 $Y=0.765 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_769_n N_VGND_c_911_n 0.0018386f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_489 N_A_27_47#_c_796_n N_VGND_c_913_n 0.00761956f $X=3.01 $Y=0.745 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_769_n N_VGND_c_913_n 0.00158683f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_491 N_A_27_47#_c_765_n N_VGND_c_915_n 0.00259536f $X=1.025 $Y=0.765 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_767_n N_VGND_c_915_n 0.00453599f $X=0.355 $Y=0.72 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_c_778_n N_VGND_c_916_n 0.00236478f $X=3.605 $Y=0.71 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_781_n N_VGND_c_916_n 0.0147597f $X=3.835 $Y=0.355 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_812_n N_VGND_c_916_n 0.0598905f $X=4.6 $Y=0.365 $X2=0 $Y2=0
cc_496 N_A_27_47#_c_766_n N_VGND_c_916_n 0.0237013f $X=7.51 $Y=0.395 $X2=0 $Y2=0
cc_497 N_A_27_47#_c_769_n N_VGND_c_916_n 0.00463578f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_498 N_A_27_47#_c_771_n N_VGND_c_916_n 5.08791e-19 $X=7.595 $Y=0.51 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_772_n N_VGND_c_916_n 0.00838914f $X=7.595 $Y=0.395 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_M1006_d N_VGND_c_917_n 0.00344766f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_M1009_d N_VGND_c_917_n 0.00151771f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_M1005_d N_VGND_c_917_n 0.00165029f $X=1.84 $Y=0.235 $X2=0
+ $Y2=0
cc_503 N_A_27_47#_M1018_d N_VGND_c_917_n 0.00165029f $X=2.7 $Y=0.235 $X2=0 $Y2=0
cc_504 N_A_27_47#_M1031_d N_VGND_c_917_n 0.00145272f $X=3.57 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_M1026_s N_VGND_c_917_n 0.00126013f $X=4.46 $Y=0.235 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_M1025_s N_VGND_c_917_n 0.00184732f $X=7.04 $Y=0.235 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_765_n N_VGND_c_917_n 0.00985019f $X=1.025 $Y=0.765 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_781_n N_VGND_c_917_n 0.00244609f $X=3.835 $Y=0.355 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_c_812_n N_VGND_c_917_n 0.00998032f $X=4.6 $Y=0.365 $X2=0 $Y2=0
cc_510 N_A_27_47#_c_766_n N_VGND_c_917_n 0.00493677f $X=7.51 $Y=0.395 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_767_n N_VGND_c_917_n 0.00630153f $X=0.355 $Y=0.72 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_c_769_n N_VGND_c_917_n 0.521812f $X=7.45 $Y=0.51 $X2=0 $Y2=0
cc_513 N_A_27_47#_c_789_n N_VGND_c_917_n 0.0297622f $X=1.3 $Y=0.51 $X2=0 $Y2=0
cc_514 N_A_27_47#_c_770_n N_VGND_c_917_n 8.86502e-19 $X=1.155 $Y=0.51 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_c_771_n N_VGND_c_917_n 0.0288358f $X=7.595 $Y=0.51 $X2=0 $Y2=0
cc_516 N_A_27_47#_c_772_n N_VGND_c_917_n 0.00152175f $X=7.595 $Y=0.395 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_812_n N_A_806_47#_M1002_d 0.00240054f $X=4.6 $Y=0.365
+ $X2=-0.19 $Y2=-0.24
cc_518 N_A_27_47#_c_769_n N_A_806_47#_M1002_d 0.00200859f $X=7.45 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_519 N_A_27_47#_c_769_n N_A_806_47#_M1020_s 0.00193634f $X=7.45 $Y=0.51 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_M1026_s N_A_806_47#_c_1029_n 0.00318278f $X=4.46 $Y=0.235
+ $X2=0 $Y2=0
cc_521 N_A_27_47#_c_812_n N_A_806_47#_c_1029_n 0.0419342f $X=4.6 $Y=0.365 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_769_n N_A_806_47#_c_1029_n 0.0614601f $X=7.45 $Y=0.51 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_c_769_n A_1314_47# 0.00331135f $X=7.45 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_524 N_A_27_47#_c_769_n A_978_47# 0.00201338f $X=7.45 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_525 N_VGND_c_917_n N_A_806_47#_M1002_d 0.0012692f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_526 N_VGND_c_917_n N_A_806_47#_M1020_s 0.00122645f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_916_n N_A_806_47#_c_1029_n 0.00500307f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_917_n A_1314_47# 0.00156226f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_529 N_VGND_c_917_n A_978_47# 0.00168555f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_530 N_A_806_47#_c_1029_n A_1314_47# 0.00762341f $X=5.865 $Y=0.725 $X2=0.475
+ $Y2=0.995

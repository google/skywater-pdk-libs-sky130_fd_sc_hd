# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__ebufn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.355000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 1.075000 1.240000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.601000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.495000 3.595000 2.465000 ;
        RECT 3.125000 0.255000 3.595000 0.825000 ;
        RECT 3.255000 0.825000 3.595000 1.495000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.445000 ;
        RECT 2.195000  0.085000 2.955000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.515000 2.175000 0.845000 2.635000 ;
        RECT 1.440000 2.175000 1.805000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.280000 0.345000 0.615000 ;
      RECT 0.085000 0.615000 1.185000 0.825000 ;
      RECT 0.085000 1.785000 0.740000 2.005000 ;
      RECT 0.085000 2.005000 0.345000 2.465000 ;
      RECT 0.525000 0.825000 0.740000 1.785000 ;
      RECT 1.015000 0.255000 2.025000 0.465000 ;
      RECT 1.015000 0.465000 1.185000 0.615000 ;
      RECT 1.015000 1.800000 1.805000 2.005000 ;
      RECT 1.015000 2.005000 1.270000 2.460000 ;
      RECT 1.355000 0.635000 1.685000 0.885000 ;
      RECT 1.410000 0.885000 1.685000 1.075000 ;
      RECT 1.410000 1.075000 2.535000 1.325000 ;
      RECT 1.410000 1.325000 1.805000 1.800000 ;
      RECT 1.855000 0.465000 2.025000 0.735000 ;
      RECT 1.855000 0.735000 2.955000 0.905000 ;
      RECT 2.705000 0.905000 2.955000 0.995000 ;
      RECT 2.705000 0.995000 3.085000 1.325000 ;
  END
END sky130_fd_sc_hd__ebufn_1

* File: sky130_fd_sc_hd__dlrtp_1.pex.spice
* Created: Thu Aug 27 14:17:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRTP_1%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.36043e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r47 19 20 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.205 $Y=1.19
+ $X2=0.205 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r49 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%A_27_47# 1 2 9 13 15 17 19 23 29 31 32 33 38
+ 41 43 46 47 50 53 54 58
c147 54 0 2.31569e-20 $X=2.53 $Y=1.53
c148 53 0 6.27501e-20 $X=2.53 $Y=1.53
c149 15 0 1.28491e-19 $X=2.725 $Y=1.69
c150 13 0 2.68021e-20 $X=0.89 $Y=2.135
c151 9 0 2.68021e-20 $X=0.89 $Y=0.445
r152 60 62 25.1791 $w=2.68e-07 $l=1.4e-07 $layer=POLY_cond $X=2.67 $Y=1.38
+ $X2=2.67 $Y2=1.52
r153 54 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r154 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.53
+ $X2=2.53 $Y2=1.53
r155 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.53
+ $X2=0.69 $Y2=1.53
r156 47 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.53
+ $X2=0.69 $Y2=1.53
r157 46 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.53
+ $X2=2.53 $Y2=1.53
r158 46 47 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.385 $Y=1.53
+ $X2=0.835 $Y2=1.53
r159 45 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=1.795
+ $X2=0.69 $Y2=1.53
r160 44 50 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.69 $Y=1.4
+ $X2=0.69 $Y2=1.53
r161 42 58 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=0.75 $Y=1.235
+ $X2=0.89 $Y2=1.235
r162 41 44 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.235
+ $X2=0.72 $Y2=1.4
r163 41 43 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.235
+ $X2=0.72 $Y2=1.07
r164 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.235 $X2=0.75 $Y2=1.235
r165 35 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=0.805
+ $X2=0.69 $Y2=1.07
r166 34 38 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r167 33 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.69 $Y2=1.795
r168 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.345 $Y2=1.88
r169 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.69 $Y2=0.805
r170 31 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.345 $Y2=0.72
r171 27 32 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.345 $Y2=0.72
r172 27 29 7.92208 $w=1.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.257 $Y2=0.51
r173 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.195 $Y=1.305
+ $X2=3.195 $Y2=0.445
r174 20 60 16.3317 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.805 $Y=1.38
+ $X2=2.67 $Y2=1.38
r175 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.12 $Y=1.38
+ $X2=3.195 $Y2=1.305
r176 19 20 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.12 $Y=1.38
+ $X2=2.805 $Y2=1.38
r177 15 62 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=2.725 $Y=1.69
+ $X2=2.67 $Y2=1.52
r178 15 17 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.725 $Y=1.69
+ $X2=2.725 $Y2=2.305
r179 11 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r180 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r181 7 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r182 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r183 2 38 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r184 1 29 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%D 2 5 9 13 15 19 22
c49 19 0 1.04465e-19 $X=1.6 $Y=1.04
c50 13 0 1.43123e-19 $X=1.83 $Y=1.64
r51 21 22 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.66 $Y=1.04
+ $X2=1.83 $Y2=1.04
r52 18 21 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.6 $Y=1.04 $X2=1.66
+ $Y2=1.04
r53 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.04 $X2=1.6 $Y2=1.04
r54 15 19 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.6 $Y=1.19 $X2=1.6
+ $Y2=1.04
r55 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.66 $Y=1.64
+ $X2=1.83 $Y2=1.64
r56 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.715
+ $X2=1.83 $Y2=1.64
r57 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.83 $Y=1.715 $X2=1.83
+ $Y2=2.165
r58 3 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r59 3 5 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
r60 2 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.66 $Y=1.565
+ $X2=1.66 $Y2=1.64
r61 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.205
+ $X2=1.66 $Y2=1.04
r62 1 2 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.66 $Y=1.205 $X2=1.66
+ $Y2=1.565
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%A_299_47# 1 2 7 9 12 16 18 20 21 24 27 34
c85 34 0 1.04465e-19 $X=2.25 $Y=0.93
r86 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=0.93 $X2=2.25 $Y2=0.93
r87 27 29 10.8065 $w=1.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.607 $Y=0.51
+ $X2=1.607 $Y2=0.7
r88 21 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.495
+ $X2=2.03 $Y2=1.58
r89 20 33 8.95599 $w=3.21e-07 $l=2.13014e-07 $layer=LI1_cond $X=2.03 $Y=1.095
+ $X2=2.14 $Y2=0.93
r90 20 21 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.03 $Y=1.095 $X2=2.03
+ $Y2=1.495
r91 19 29 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.607 $Y2=0.7
r92 18 33 8.74143 $w=3.21e-07 $l=3.1265e-07 $layer=LI1_cond $X=1.945 $Y=0.7
+ $X2=2.14 $Y2=0.93
r93 18 19 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.945 $Y=0.7
+ $X2=1.705 $Y2=0.7
r94 14 24 27.5968 $w=1.68e-07 $l=4.23e-07 $layer=LI1_cond $X=1.607 $Y=1.58
+ $X2=2.03 $Y2=1.58
r95 14 16 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=1.607 $Y=1.665
+ $X2=1.607 $Y2=1.99
r96 10 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.095
+ $X2=2.25 $Y2=0.93
r97 10 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=1.095
+ $X2=2.25 $Y2=2.165
r98 7 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.765
+ $X2=2.25 $Y2=0.93
r99 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.765 $X2=2.25
+ $Y2=0.445
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r101 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%A_193_47# 1 2 9 12 16 19 20 24 26 28 29 32
+ 35 39 45 51
c120 51 0 6.27501e-20 $X=3.125 $Y=1.815
c121 45 0 2.31569e-20 $X=3.245 $Y=1.8
c122 28 0 1.28491e-19 $X=2.865 $Y=1.87
c123 26 0 2.26849e-19 $X=3.125 $Y=0.93
c124 20 0 8.72205e-20 $X=1.125 $Y=1.795
c125 16 0 5.59029e-20 $X=1.1 $Y=0.51
r126 43 51 2.12342 $w=3.16e-07 $l=5.5e-08 $layer=LI1_cond $X=3.18 $Y=1.815
+ $X2=3.125 $Y2=1.815
r127 42 45 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=3.18 $Y=1.8
+ $X2=3.245 $Y2=1.8
r128 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.8 $X2=3.18 $Y2=1.8
r129 36 51 4.43987 $w=3.16e-07 $l=1.15e-07 $layer=LI1_cond $X=3.01 $Y=1.815
+ $X2=3.125 $Y2=1.815
r130 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.01 $Y=1.87
+ $X2=3.01 $Y2=1.87
r131 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r132 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r133 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.865 $Y=1.87
+ $X2=3.01 $Y2=1.87
r134 28 29 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.865 $Y=1.87
+ $X2=1.295 $Y2=1.87
r135 24 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=0.93
+ $X2=2.775 $Y2=0.765
r136 23 26 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.775 $Y=0.93
+ $X2=3.125 $Y2=0.93
r137 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.775
+ $Y=0.93 $X2=2.775 $Y2=0.93
r138 20 32 3.92878 $w=2.18e-07 $l=7.5e-08 $layer=LI1_cond $X=1.125 $Y=1.795
+ $X2=1.125 $Y2=1.87
r139 20 21 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=1.125 $Y=1.795
+ $X2=1.125 $Y2=1.685
r140 19 51 2.35055 $w=2.4e-07 $l=1.8e-07 $layer=LI1_cond $X=3.125 $Y=1.635
+ $X2=3.125 $Y2=1.815
r141 18 26 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=1.095
+ $X2=3.125 $Y2=0.93
r142 18 19 25.93 $w=2.38e-07 $l=5.4e-07 $layer=LI1_cond $X=3.125 $Y=1.095
+ $X2=3.125 $Y2=1.635
r143 16 21 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r144 10 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.245 $Y=1.935
+ $X2=3.245 $Y2=1.8
r145 10 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.245 $Y=1.935
+ $X2=3.245 $Y2=2.305
r146 9 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.765 $Y=0.445
+ $X2=2.765 $Y2=0.765
r147 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r148 1 16 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%A_711_21# 1 2 9 11 14 18 21 23 24 28 31 34
+ 37 39 43 44 47 49 50 59
c109 49 0 1.19e-19 $X=5.47 $Y=1.16
c110 24 0 1.34791e-19 $X=3.65 $Y=0.905
c111 11 0 9.20582e-20 $X=3.67 $Y=1.535
r112 53 55 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.67 $Y=1.7
+ $X2=3.81 $Y2=1.7
r113 50 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.16
+ $X2=5.47 $Y2=1.325
r114 50 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.16
+ $X2=5.47 $Y2=0.995
r115 49 52 7.12114 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=5.4 $Y=1.16
+ $X2=5.4 $Y2=1.325
r116 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.16 $X2=5.47 $Y2=1.16
r117 46 47 6.2995 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=4.815 $Y=1.685
+ $X2=4.965 $Y2=1.685
r118 44 46 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=4.795 $Y=1.685
+ $X2=4.815 $Y2=1.685
r119 42 44 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=4.46 $Y=1.685
+ $X2=4.795 $Y2=1.685
r120 42 43 3.78243 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.46 $Y=1.685
+ $X2=4.345 $Y2=1.685
r121 39 41 14.6716 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=4.385 $Y=0.38
+ $X2=4.385 $Y2=0.805
r122 37 52 9.42908 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=5.355 $Y=1.505
+ $X2=5.355 $Y2=1.325
r123 34 37 6.82087 $w=2.3e-07 $l=1.60857e-07 $layer=LI1_cond $X=5.245 $Y=1.62
+ $X2=5.355 $Y2=1.505
r124 34 47 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.245 $Y=1.62
+ $X2=4.965 $Y2=1.62
r125 31 42 3.35874 $w=2.3e-07 $l=1.8e-07 $layer=LI1_cond $X=4.46 $Y=1.505
+ $X2=4.46 $Y2=1.685
r126 31 41 35.0744 $w=2.28e-07 $l=7e-07 $layer=LI1_cond $X=4.46 $Y=1.505
+ $X2=4.46 $Y2=0.805
r127 28 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.9 $Y=1.7 $X2=3.81
+ $Y2=1.7
r128 27 43 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.9 $Y=1.7
+ $X2=4.345 $Y2=1.7
r129 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9
+ $Y=1.7 $X2=3.9 $Y2=1.7
r130 23 24 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=3.65 $Y=0.755
+ $X2=3.65 $Y2=0.905
r131 21 60 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.51 $Y=1.985
+ $X2=5.51 $Y2=1.325
r132 18 59 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.51 $Y=0.56
+ $X2=5.51 $Y2=0.995
r133 12 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.865
+ $X2=3.81 $Y2=1.7
r134 12 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.81 $Y=1.865
+ $X2=3.81 $Y2=2.275
r135 11 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.535
+ $X2=3.67 $Y2=1.7
r136 11 24 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.67 $Y=1.535
+ $X2=3.67 $Y2=0.905
r137 9 23 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=3.63 $Y=0.445
+ $X2=3.63 $Y2=0.755
r138 2 46 300 $w=1.7e-07 $l=3.44674e-07 $layer=licon1_PDIFF $count=2 $X=4.645
+ $Y=1.485 $X2=4.815 $Y2=1.755
r139 1 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.235
+ $Y=0.235 $X2=4.36 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%A_560_425# 1 2 7 9 12 14 15 16 20 25 27 30
+ 33
c86 33 0 1.25684e-19 $X=3.415 $Y=0.995
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.16 $X2=4.09 $Y2=1.16
r88 28 33 0.89609 $w=3.3e-07 $l=2.80624e-07 $layer=LI1_cond $X=3.625 $Y=1.16
+ $X2=3.415 $Y2=0.995
r89 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.625 $Y=1.16
+ $X2=4.09 $Y2=1.16
r90 26 33 8.61065 $w=1.7e-07 $l=3.87492e-07 $layer=LI1_cond $X=3.54 $Y=1.325
+ $X2=3.415 $Y2=0.995
r91 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.54 $Y=1.325
+ $X2=3.54 $Y2=2.255
r92 25 33 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=0.995
+ $X2=3.415 $Y2=0.995
r93 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.5 $Y=0.535 $X2=3.5
+ $Y2=0.995
r94 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=0.45
+ $X2=3.5 $Y2=0.535
r95 20 22 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.415 $Y=0.45
+ $X2=2.98 $Y2=0.45
r96 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.455 $Y=2.34
+ $X2=3.54 $Y2=2.255
r97 16 18 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.455 $Y=2.34
+ $X2=2.975 $Y2=2.34
r98 14 31 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=4.495 $Y=1.16
+ $X2=4.09 $Y2=1.16
r99 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.495 $Y=1.16
+ $X2=4.57 $Y2=1.16
r100 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.325
+ $X2=4.57 $Y2=1.16
r101 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.57 $Y=1.325
+ $X2=4.57 $Y2=1.985
r102 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=0.995
+ $X2=4.57 $Y2=1.16
r103 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.57 $Y=0.995
+ $X2=4.57 $Y2=0.56
r104 2 18 600 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=2.125 $X2=2.975 $Y2=2.34
r105 1 22 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.235 $X2=2.98 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%RESET_B 3 6 8 9 10 15 16 17
r36 16 26 6.83261 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.91 $Y=1.16
+ $X2=4.91 $Y2=0.995
r37 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.99 $Y=1.16
+ $X2=4.99 $Y2=1.325
r38 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.99 $Y=1.16
+ $X2=4.99 $Y2=0.995
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.16 $X2=4.99 $Y2=1.16
r40 10 16 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=4.91 $Y=1.19 $X2=4.91
+ $Y2=1.16
r41 9 26 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.86 $Y=0.85 $X2=4.86
+ $Y2=0.995
r42 8 9 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.86 $Y=0.51 $X2=4.86
+ $Y2=0.85
r43 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.985
+ $X2=5.05 $Y2=1.325
r44 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.56 $X2=5.05
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%VPWR 1 2 3 4 15 19 23 26 29 32 34 39 51 57
+ 58 61 64 67
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r91 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r92 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r93 58 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r94 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r95 55 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.3 $Y2=2.72
r96 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.75 $Y2=2.72
r97 54 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r99 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.3 $Y2=2.72
r100 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=4.83 $Y2=2.72
r101 50 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r103 47 50 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 47 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r105 46 49 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 44 64 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.245 $Y=2.72
+ $X2=2.1 $Y2=2.72
r108 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=2.72
+ $X2=2.53 $Y2=2.72
r109 43 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 43 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r113 40 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 39 64 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.1 $Y2=2.72
r115 39 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r117 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r118 32 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r120 30 53 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.445 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 29 49 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.93 $Y=2.72 $X2=3.91
+ $Y2=2.72
r122 29 30 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=4.187 $Y=2.72
+ $X2=4.445 $Y2=2.72
r123 26 29 9.75443 $w=5.13e-07 $l=4.2e-07 $layer=LI1_cond $X=4.187 $Y=2.3
+ $X2=4.187 $Y2=2.72
r124 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635 $X2=5.3
+ $Y2=2.72
r125 21 23 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2
r126 17 64 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.635
+ $X2=2.1 $Y2=2.72
r127 17 19 25.2345 $w=2.88e-07 $l=6.35e-07 $layer=LI1_cond $X=2.1 $Y=2.635
+ $X2=2.1 $Y2=2
r128 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r129 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r130 4 23 300 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.485 $X2=5.3 $Y2=2
r131 3 26 300 $w=1.7e-07 $l=5.80732e-07 $layer=licon1_PDIFF $count=2 $X=3.885
+ $Y=2.065 $X2=4.36 $Y2=2.3
r132 2 19 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r133 1 15 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%Q 1 2 9 10 11 19 30
r17 28 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.81 $Y=0.745
+ $X2=5.81 $Y2=1.67
r18 16 19 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.765 $Y=1.8
+ $X2=5.765 $Y2=1.835
r19 10 16 0.354598 $w=2.58e-07 $l=8e-09 $layer=LI1_cond $X=5.765 $Y=1.792
+ $X2=5.765 $Y2=1.8
r20 10 30 6.78766 $w=2.58e-07 $l=1.22e-07 $layer=LI1_cond $X=5.765 $Y=1.792
+ $X2=5.765 $Y2=1.67
r21 10 11 14.7601 $w=2.58e-07 $l=3.33e-07 $layer=LI1_cond $X=5.765 $Y=1.877
+ $X2=5.765 $Y2=2.21
r22 10 19 1.86164 $w=2.58e-07 $l=4.2e-08 $layer=LI1_cond $X=5.765 $Y=1.877
+ $X2=5.765 $Y2=1.835
r23 9 28 11.3641 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=5.752 $Y=0.51
+ $X2=5.752 $Y2=0.745
r24 2 19 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=1.835
r25 1 9 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_1%VGND 1 2 3 4 15 19 23 27 29 31 36 41 49 56
+ 57 60 63 66 69
c94 57 0 2.71124e-20 $X=5.75 $Y=0
r95 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r96 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r97 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r98 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r99 57 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r100 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r101 54 69 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.297
+ $Y2=0
r102 54 56 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.75
+ $Y2=0
r103 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r104 53 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r105 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r106 50 66 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=3.89
+ $Y2=0
r107 50 52 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=4.83 $Y2=0
r108 49 69 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.297 $Y2=0
r109 49 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=4.83 $Y2=0
r110 48 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r111 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r112 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r113 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r114 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r115 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r116 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r117 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r118 41 66 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.89
+ $Y2=0
r119 41 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=0
+ $X2=3.45 $Y2=0
r120 40 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r121 40 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r122 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r123 37 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r124 37 39 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r125 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r126 36 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r127 31 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r128 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r129 29 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r130 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r131 25 69 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.297 $Y=0.085
+ $X2=5.297 $Y2=0
r132 25 27 18.803 $w=2.83e-07 $l=4.65e-07 $layer=LI1_cond $X=5.297 $Y=0.085
+ $X2=5.297 $Y2=0.55
r133 21 66 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=0.085
+ $X2=3.89 $Y2=0
r134 21 23 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.89 $Y=0.085
+ $X2=3.89 $Y2=0.445
r135 17 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r136 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r137 13 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r138 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r139 4 27 182 $w=1.7e-07 $l=3.92874e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.3 $Y2=0.55
r140 3 23 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.235 $X2=3.84 $Y2=0.445
r141 2 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r142 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__and2_2.pex.spice
* Created: Tue Sep  1 18:56:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND2_2%A 3 7 9 10 11 19 21
r35 17 24 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=0.465 $Y=1.2 $X2=0.4
+ $Y2=1.2
r36 16 19 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.465 $Y=1.16
+ $X2=0.66 $Y2=1.16
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.465
+ $Y=1.16 $X2=0.465 $Y2=1.16
r38 11 17 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.69 $Y=1.2
+ $X2=0.465 $Y2=1.2
r39 10 21 7.50003 $w=3.13e-07 $l=2.05e-07 $layer=LI1_cond $X=0.242 $Y=1.53
+ $X2=0.242 $Y2=1.325
r40 9 21 3.06294 $w=3.15e-07 $l=1.25e-07 $layer=LI1_cond $X=0.242 $Y=1.2
+ $X2=0.242 $Y2=1.325
r41 9 24 3.87155 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=0.242 $Y=1.2 $X2=0.4
+ $Y2=1.2
r42 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.66 $Y=1.325
+ $X2=0.66 $Y2=1.16
r43 5 7 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.66 $Y=1.325 $X2=0.66
+ $Y2=2.065
r44 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.66 $Y=0.995
+ $X2=0.66 $Y2=1.16
r45 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.66 $Y=0.995 $X2=0.66
+ $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_2%B 3 7 9 12
r35 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.17 $Y2=1.325
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.17 $Y2=0.995
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r38 7 15 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.08 $Y=2.065
+ $X2=1.08 $Y2=1.325
r39 3 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.08 $Y=0.585
+ $X2=1.08 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_2%A_61_75# 1 2 7 9 12 14 16 19 22 23 24 27 29
+ 30 33 35 36 37 38
r95 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.16 $X2=1.71 $Y2=1.16
r96 39 41 18.2479 $w=2.34e-07 $l=3.5e-07 $layer=LI1_cond $X=1.65 $Y=0.81
+ $X2=1.65 $Y2=1.16
r97 37 41 9.53671 $w=2.34e-07 $l=1.92678e-07 $layer=LI1_cond $X=1.59 $Y=1.325
+ $X2=1.65 $Y2=1.16
r98 37 38 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.59 $Y=1.325
+ $X2=1.59 $Y2=1.575
r99 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.66
+ $X2=1.59 $Y2=1.575
r100 35 36 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.505 $Y=1.66
+ $X2=1.035 $Y2=1.66
r101 31 36 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.885 $Y=1.745
+ $X2=1.035 $Y2=1.66
r102 31 33 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.885 $Y=1.745
+ $X2=0.885 $Y2=2.13
r103 29 39 1.95941 $w=1.9e-07 $l=1.45e-07 $layer=LI1_cond $X=1.505 $Y=0.81
+ $X2=1.65 $Y2=0.81
r104 29 30 51.9522 $w=1.88e-07 $l=8.9e-07 $layer=LI1_cond $X=1.505 $Y=0.81
+ $X2=0.615 $Y2=0.81
r105 25 30 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.45 $Y=0.715
+ $X2=0.615 $Y2=0.81
r106 25 27 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.45 $Y=0.715
+ $X2=0.45 $Y2=0.52
r107 23 42 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.085 $Y=1.16
+ $X2=1.71 $Y2=1.16
r108 23 24 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.085 $Y=1.16
+ $X2=2.16 $Y2=1.16
r109 21 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.695 $Y=1.16
+ $X2=1.71 $Y2=1.16
r110 21 22 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.695 $Y=1.16
+ $X2=1.62 $Y2=1.16
r111 17 24 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.325
+ $X2=2.16 $Y2=1.16
r112 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.16 $Y=1.325
+ $X2=2.16 $Y2=1.985
r113 14 24 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=0.995
+ $X2=2.16 $Y2=1.16
r114 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.16 $Y=0.995
+ $X2=2.16 $Y2=0.56
r115 10 22 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.325
+ $X2=1.62 $Y2=1.16
r116 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.62 $Y=1.325
+ $X2=1.62 $Y2=1.985
r117 7 22 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=0.995
+ $X2=1.62 $Y2=1.16
r118 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.62 $Y=0.995
+ $X2=1.62 $Y2=0.56
r119 2 33 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=1.855 $X2=0.87 $Y2=2.13
r120 1 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.305
+ $Y=0.375 $X2=0.45 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_2%VPWR 1 2 3 12 16 18 20 25 26 28 29 30 38 44
r39 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r40 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 38 43 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.572 $Y2=2.72
r43 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 37 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 30 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 30 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r48 28 36 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.41 $Y2=2.72
r50 27 40 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.575 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=2.72
+ $X2=1.41 $Y2=2.72
r52 25 33 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.285 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 25 26 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.285 $Y=2.72
+ $X2=0.425 $Y2=2.72
r54 24 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 24 26 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.425 $Y2=2.72
r56 20 23 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=1.66
+ $X2=2.53 $Y2=2.34
r57 18 43 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.53 $Y=2.635
+ $X2=2.572 $Y2=2.72
r58 18 23 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.53 $Y=2.635
+ $X2=2.53 $Y2=2.34
r59 14 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=2.635
+ $X2=1.41 $Y2=2.72
r60 14 16 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.41 $Y=2.635
+ $X2=1.41 $Y2=2
r61 10 26 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.425 $Y=2.635
+ $X2=0.425 $Y2=2.72
r62 10 12 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=0.425 $Y=2.635
+ $X2=0.425 $Y2=2.13
r63 3 23 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.485 $X2=2.47 $Y2=2.34
r64 3 20 400 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.485 $X2=2.47 $Y2=1.66
r65 2 16 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=1.155
+ $Y=1.855 $X2=1.41 $Y2=2
r66 1 12 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.855 $X2=0.45 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_2%X 1 2 7 11 12 13 14 15 16 25 36
r31 36 40 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=2.09 $Y=1.87 $X2=2.09
+ $Y2=1.915
r32 16 42 5.5817 $w=4.48e-07 $l=2.1e-07 $layer=LI1_cond $X=1.99 $Y=2.21 $X2=1.99
+ $Y2=2
r33 15 42 1.72767 $w=4.48e-07 $l=6.5e-08 $layer=LI1_cond $X=1.99 $Y=1.935
+ $X2=1.99 $Y2=2
r34 15 40 2.87587 $w=4.48e-07 $l=2e-08 $layer=LI1_cond $X=1.99 $Y=1.935 $X2=1.99
+ $Y2=1.915
r35 15 36 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=2.09 $Y=1.85 $X2=2.09
+ $Y2=1.87
r36 14 15 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.09 $Y=1.53
+ $X2=2.09 $Y2=1.85
r37 13 14 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.09 $Y=1.19
+ $X2=2.09 $Y2=1.53
r38 12 13 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.09 $Y=0.85
+ $X2=2.09 $Y2=1.19
r39 11 25 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=2.09 $Y=0.4 $X2=2.09
+ $Y2=0.545
r40 11 12 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.09 $Y=0.57
+ $X2=2.09 $Y2=0.85
r41 11 25 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.09 $Y=0.57
+ $X2=2.09 $Y2=0.545
r42 7 11 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=1.965 $Y=0.4 $X2=2.09
+ $Y2=0.4
r43 7 9 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.965 $Y=0.4 $X2=1.83
+ $Y2=0.4
r44 2 42 300 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.485 $X2=1.93 $Y2=2
r45 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.235 $X2=1.83 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_2%VGND 1 2 9 11 13 16 17 18 27 33
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r36 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r37 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r38 27 32 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.572
+ $Y2=0
r39 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.07
+ $Y2=0
r40 26 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r41 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r42 21 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r43 18 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r44 18 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r45 16 25 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.15
+ $Y2=0
r46 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.37
+ $Y2=0
r47 15 29 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=2.07
+ $Y2=0
r48 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.37
+ $Y2=0
r49 11 32 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.572 $Y2=0
r50 11 13 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0.38
r51 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=0.085
+ $X2=1.37 $Y2=0
r52 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.37 $Y=0.085
+ $X2=1.37 $Y2=0.38
r53 2 13 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=2.235
+ $Y=0.235 $X2=2.47 $Y2=0.38
r54 1 9 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.375 $X2=1.41 $Y2=0.38
.ends


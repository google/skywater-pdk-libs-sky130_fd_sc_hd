* File: sky130_fd_sc_hd__inv_12.pex.spice
* Created: Thu Aug 27 14:22:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_12%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 57 59 62 64 66 69 71 73 76 78 80 83 85 86 87 88 89 90
+ 91 92 93 94 123
r236 121 123 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.045 $Y=1.16
+ $X2=5.255 $Y2=1.16
r237 119 121 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.835 $Y=1.16
+ $X2=5.045 $Y2=1.16
r238 118 119 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.415 $Y=1.16
+ $X2=4.835 $Y2=1.16
r239 117 118 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.995 $Y=1.16
+ $X2=4.415 $Y2=1.16
r240 116 117 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.575 $Y=1.16
+ $X2=3.995 $Y2=1.16
r241 115 116 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.155 $Y=1.16
+ $X2=3.575 $Y2=1.16
r242 114 115 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=3.155 $Y2=1.16
r243 113 114 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.315 $Y=1.16
+ $X2=2.735 $Y2=1.16
r244 112 113 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.895 $Y=1.16
+ $X2=2.315 $Y2=1.16
r245 111 112 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.475 $Y=1.16
+ $X2=1.895 $Y2=1.16
r246 110 111 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=1.475 $Y2=1.16
r247 108 110 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.845 $Y=1.16
+ $X2=1.055 $Y2=1.16
r248 108 109 26.4145 $w=1.7e-07 $l=9.35e-07 $layer=licon1_POLY $count=5 $X=0.845
+ $Y=1.16 $X2=0.845 $Y2=1.16
r249 105 108 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.635 $Y=1.16
+ $X2=0.845 $Y2=1.16
r250 94 121 26.4145 $w=1.7e-07 $l=9.35e-07 $layer=licon1_POLY $count=5 $X=5.045
+ $Y=1.16 $X2=5.045 $Y2=1.16
r251 93 94 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=4.67 $Y=1.2
+ $X2=5.045 $Y2=1.2
r252 92 93 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.29 $Y=1.2
+ $X2=4.67 $Y2=1.2
r253 91 92 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=3.83 $Y=1.2 $X2=4.29
+ $Y2=1.2
r254 90 91 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=3.45 $Y=1.2
+ $X2=3.83 $Y2=1.2
r255 89 90 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=1.2 $X2=3.45
+ $Y2=1.2
r256 88 89 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=1.2 $X2=2.99
+ $Y2=1.2
r257 87 88 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=1.2 $X2=2.53
+ $Y2=1.2
r258 86 87 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=2.07
+ $Y2=1.2
r259 85 86 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.61
+ $Y2=1.2
r260 85 109 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=1.15 $Y=1.2
+ $X2=0.845 $Y2=1.2
r261 81 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.255 $Y=1.325
+ $X2=5.255 $Y2=1.16
r262 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.255 $Y=1.325
+ $X2=5.255 $Y2=1.985
r263 78 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.255 $Y=0.995
+ $X2=5.255 $Y2=1.16
r264 78 80 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.255 $Y=0.995
+ $X2=5.255 $Y2=0.56
r265 74 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.325
+ $X2=4.835 $Y2=1.16
r266 74 76 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.835 $Y=1.325
+ $X2=4.835 $Y2=1.985
r267 71 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=0.995
+ $X2=4.835 $Y2=1.16
r268 71 73 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.835 $Y=0.995
+ $X2=4.835 $Y2=0.56
r269 67 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.325
+ $X2=4.415 $Y2=1.16
r270 67 69 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.415 $Y=1.325
+ $X2=4.415 $Y2=1.985
r271 64 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=0.995
+ $X2=4.415 $Y2=1.16
r272 64 66 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.415 $Y=0.995
+ $X2=4.415 $Y2=0.56
r273 60 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.325
+ $X2=3.995 $Y2=1.16
r274 60 62 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.995 $Y=1.325
+ $X2=3.995 $Y2=1.985
r275 57 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=0.995
+ $X2=3.995 $Y2=1.16
r276 57 59 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.995 $Y=0.995
+ $X2=3.995 $Y2=0.56
r277 53 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.325
+ $X2=3.575 $Y2=1.16
r278 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.575 $Y=1.325
+ $X2=3.575 $Y2=1.985
r279 50 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=1.16
r280 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=0.56
r281 46 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=1.325
+ $X2=3.155 $Y2=1.16
r282 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.155 $Y=1.325
+ $X2=3.155 $Y2=1.985
r283 43 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=0.995
+ $X2=3.155 $Y2=1.16
r284 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.155 $Y=0.995
+ $X2=3.155 $Y2=0.56
r285 39 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.325
+ $X2=2.735 $Y2=1.16
r286 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.735 $Y=1.325
+ $X2=2.735 $Y2=1.985
r287 36 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=1.16
r288 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=0.56
r289 32 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.16
r290 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.985
r291 29 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=1.16
r292 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=0.56
r293 25 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.325
+ $X2=1.895 $Y2=1.16
r294 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.895 $Y=1.325
+ $X2=1.895 $Y2=1.985
r295 22 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=1.16
r296 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=0.56
r297 18 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.325
+ $X2=1.475 $Y2=1.16
r298 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.475 $Y=1.325
+ $X2=1.475 $Y2=1.985
r299 15 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=1.16
r300 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.56
r301 11 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.325
+ $X2=1.055 $Y2=1.16
r302 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.055 $Y=1.325
+ $X2=1.055 $Y2=1.985
r303 8 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=1.16
r304 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r305 4 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.325
+ $X2=0.635 $Y2=1.16
r306 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.635 $Y=1.325
+ $X2=0.635 $Y2=1.985
r307 1 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=1.16
r308 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_12%VPWR 1 2 3 4 5 6 7 22 24 28 30 34 38 42 46 48
+ 50 52 53 55 56 58 59 61 62 63 79 87 91
r93 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r94 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r95 82 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r96 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r97 79 90 4.90987 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=5.555 $Y=2.72
+ $X2=5.767 $Y2=2.72
r98 79 81 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.555 $Y=2.72
+ $X2=5.29 $Y2=2.72
r99 78 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r100 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r101 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r102 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r103 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r104 72 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r105 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 69 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.72
+ $X2=2.105 $Y2=2.72
r107 69 71 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=2.72
+ $X2=2.53 $Y2=2.72
r108 68 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r110 65 84 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=0.255 $Y2=2.72
r111 65 67 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 63 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r113 63 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r114 61 77 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.54 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.72
+ $X2=4.625 $Y2=2.72
r116 60 81 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.71 $Y=2.72
+ $X2=5.29 $Y2=2.72
r117 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=2.72
+ $X2=4.625 $Y2=2.72
r118 58 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=2.72
+ $X2=3.785 $Y2=2.72
r120 57 77 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.87 $Y=2.72 $X2=4.37
+ $Y2=2.72
r121 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=2.72
+ $X2=3.785 $Y2=2.72
r122 55 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.86 $Y=2.72
+ $X2=2.53 $Y2=2.72
r123 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=2.72
+ $X2=2.945 $Y2=2.72
r124 54 74 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.03 $Y=2.72
+ $X2=3.45 $Y2=2.72
r125 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.72
+ $X2=2.945 $Y2=2.72
r126 52 67 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=2.72 $X2=1.15
+ $Y2=2.72
r127 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.72
+ $X2=1.265 $Y2=2.72
r128 48 90 2.94129 $w=3.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.725 $Y=2.635
+ $X2=5.767 $Y2=2.72
r129 48 50 21.5236 $w=3.38e-07 $l=6.35e-07 $layer=LI1_cond $X=5.725 $Y=2.635
+ $X2=5.725 $Y2=2
r130 44 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=2.635
+ $X2=4.625 $Y2=2.72
r131 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.625 $Y=2.635
+ $X2=4.625 $Y2=2
r132 40 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=2.635
+ $X2=3.785 $Y2=2.72
r133 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.785 $Y=2.635
+ $X2=3.785 $Y2=2
r134 36 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2.72
r135 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2
r136 32 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2.72
r137 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2
r138 31 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=2.72
+ $X2=1.265 $Y2=2.72
r139 30 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=2.72
+ $X2=2.105 $Y2=2.72
r140 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.02 $Y=2.72
+ $X2=1.35 $Y2=2.72
r141 26 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2.72
r142 26 28 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2
r143 22 84 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.255 $Y2=2.72
r144 22 24 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.382 $Y2=2
r145 7 50 300 $w=1.7e-07 $l=6.82697e-07 $layer=licon1_PDIFF $count=2 $X=5.33
+ $Y=1.485 $X2=5.72 $Y2=2
r146 6 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.485 $X2=4.625 $Y2=2
r147 5 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.65
+ $Y=1.485 $X2=3.785 $Y2=2
r148 4 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.485 $X2=2.945 $Y2=2
r149 3 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=1.485 $X2=2.105 $Y2=2
r150 2 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.485 $X2=1.265 $Y2=2
r151 1 24 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=1.485 $X2=0.425 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__INV_12%Y 1 2 3 4 5 6 7 8 9 10 11 12 39 43 45 46 47
+ 48 51 55 57 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 105 107 118 120 121
+ 123 124 126 127 129 130 132 135 136
r243 134 136 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.72 $Y=1.495
+ $X2=5.72 $Y2=1.19
r244 133 136 9.38418 $w=3.48e-07 $l=2.85e-07 $layer=LI1_cond $X=5.72 $Y=0.905
+ $X2=5.72 $Y2=1.19
r245 114 135 8.27047 $w=4.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.297 $Y=1.495
+ $X2=0.297 $Y2=1.19
r246 114 117 35.7519 $w=1.68e-07 $l=5.48e-07 $layer=LI1_cond $X=0.297 $Y=1.58
+ $X2=0.845 $Y2=1.58
r247 110 135 7.72815 $w=4.23e-07 $l=2.85e-07 $layer=LI1_cond $X=0.297 $Y=0.905
+ $X2=0.297 $Y2=1.19
r248 108 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=1.58
+ $X2=5.045 $Y2=1.58
r249 107 134 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.545 $Y=1.58
+ $X2=5.72 $Y2=1.495
r250 107 108 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.545 $Y=1.58
+ $X2=5.21 $Y2=1.58
r251 106 130 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0.81
+ $X2=5.045 $Y2=0.81
r252 105 133 7.62524 $w=1.9e-07 $l=2.17371e-07 $layer=LI1_cond $X=5.545 $Y=0.81
+ $X2=5.72 $Y2=0.905
r253 105 106 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=5.545 $Y=0.81
+ $X2=5.21 $Y2=0.81
r254 101 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=1.665
+ $X2=5.045 $Y2=1.58
r255 101 103 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.045 $Y=1.665
+ $X2=5.045 $Y2=2.34
r256 97 130 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.045 $Y=0.715
+ $X2=5.045 $Y2=0.81
r257 97 99 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.045 $Y=0.715
+ $X2=5.045 $Y2=0.38
r258 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=1.58
+ $X2=4.205 $Y2=1.58
r259 95 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=1.58
+ $X2=5.045 $Y2=1.58
r260 95 96 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.88 $Y=1.58
+ $X2=4.37 $Y2=1.58
r261 94 127 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=0.81
+ $X2=4.205 $Y2=0.81
r262 93 130 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=0.81
+ $X2=5.045 $Y2=0.81
r263 93 94 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=4.88 $Y=0.81
+ $X2=4.37 $Y2=0.81
r264 89 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=1.665
+ $X2=4.205 $Y2=1.58
r265 89 91 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.205 $Y=1.665
+ $X2=4.205 $Y2=2.34
r266 85 127 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.205 $Y=0.715
+ $X2=4.205 $Y2=0.81
r267 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.205 $Y=0.715
+ $X2=4.205 $Y2=0.38
r268 84 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=1.58
+ $X2=3.365 $Y2=1.58
r269 83 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=1.58
+ $X2=4.205 $Y2=1.58
r270 83 84 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.04 $Y=1.58
+ $X2=3.53 $Y2=1.58
r271 82 124 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=0.81
+ $X2=3.365 $Y2=0.81
r272 81 127 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=0.81
+ $X2=4.205 $Y2=0.81
r273 81 82 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=4.04 $Y=0.81
+ $X2=3.53 $Y2=0.81
r274 77 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=1.665
+ $X2=3.365 $Y2=1.58
r275 77 79 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.365 $Y=1.665
+ $X2=3.365 $Y2=2.34
r276 73 124 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.365 $Y=0.715
+ $X2=3.365 $Y2=0.81
r277 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.365 $Y=0.715
+ $X2=3.365 $Y2=0.38
r278 72 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.58
+ $X2=2.525 $Y2=1.58
r279 71 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=1.58
+ $X2=3.365 $Y2=1.58
r280 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.2 $Y=1.58
+ $X2=2.69 $Y2=1.58
r281 70 121 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.81
+ $X2=2.525 $Y2=0.81
r282 69 124 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=0.81
+ $X2=3.365 $Y2=0.81
r283 69 70 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=3.2 $Y=0.81
+ $X2=2.69 $Y2=0.81
r284 65 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.665
+ $X2=2.525 $Y2=1.58
r285 65 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.525 $Y=1.665
+ $X2=2.525 $Y2=2.34
r286 61 121 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.525 $Y=0.715
+ $X2=2.525 $Y2=0.81
r287 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.525 $Y=0.715
+ $X2=2.525 $Y2=0.38
r288 60 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=1.58
+ $X2=1.685 $Y2=1.58
r289 59 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=1.58
+ $X2=2.525 $Y2=1.58
r290 59 60 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.36 $Y=1.58
+ $X2=1.85 $Y2=1.58
r291 58 118 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0.81
+ $X2=1.685 $Y2=0.81
r292 57 121 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0.81
+ $X2=2.525 $Y2=0.81
r293 57 58 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=2.36 $Y=0.81
+ $X2=1.85 $Y2=0.81
r294 53 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.58
r295 53 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.34
r296 49 118 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=1.685 $Y=0.715
+ $X2=1.685 $Y2=0.81
r297 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.685 $Y=0.715
+ $X2=1.685 $Y2=0.38
r298 48 117 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.58
+ $X2=0.845 $Y2=1.58
r299 47 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=1.685 $Y2=1.58
r300 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=1.01 $Y2=1.58
r301 45 118 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0.81
+ $X2=1.685 $Y2=0.81
r302 45 46 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=1.52 $Y=0.81
+ $X2=1.01 $Y2=0.81
r303 43 117 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.845 $Y=2.34
+ $X2=0.845 $Y2=1.665
r304 37 46 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0.81
+ $X2=1.01 $Y2=0.81
r305 37 110 31.9885 $w=1.88e-07 $l=5.48e-07 $layer=LI1_cond $X=0.845 $Y=0.81
+ $X2=0.297 $Y2=0.81
r306 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.845 $Y=0.715
+ $X2=0.845 $Y2=0.38
r307 12 132 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.485 $X2=5.045 $Y2=1.66
r308 12 103 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.485 $X2=5.045 $Y2=2.34
r309 11 129 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.07
+ $Y=1.485 $X2=4.205 $Y2=1.66
r310 11 91 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.07
+ $Y=1.485 $X2=4.205 $Y2=2.34
r311 10 126 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.485 $X2=3.365 $Y2=1.66
r312 10 79 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.485 $X2=3.365 $Y2=2.34
r313 9 123 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.525 $Y2=1.66
r314 9 67 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.525 $Y2=2.34
r315 8 120 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.685 $Y2=1.66
r316 8 55 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.685 $Y2=2.34
r317 7 117 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.485 $X2=0.845 $Y2=1.66
r318 7 43 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.485 $X2=0.845 $Y2=2.34
r319 6 99 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.235 $X2=5.045 $Y2=0.38
r320 5 87 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.07
+ $Y=0.235 $X2=4.205 $Y2=0.38
r321 4 75 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.23
+ $Y=0.235 $X2=3.365 $Y2=0.38
r322 3 63 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.39
+ $Y=0.235 $X2=2.525 $Y2=0.38
r323 2 51 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.235 $X2=1.685 $Y2=0.38
r324 1 39 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.71
+ $Y=0.235 $X2=0.845 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__INV_12%VGND 1 2 3 4 5 6 7 22 24 28 30 34 38 42 46 48
+ 50 52 53 55 56 58 59 61 62 63 79 87 91
r109 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r110 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r111 82 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r112 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r113 79 90 4.90987 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=5.555 $Y=0
+ $X2=5.767 $Y2=0
r114 79 81 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.555 $Y=0
+ $X2=5.29 $Y2=0
r115 78 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r116 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r117 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r118 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r119 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r120 72 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r121 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r122 69 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.105
+ $Y2=0
r123 69 71 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.53
+ $Y2=0
r124 68 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r125 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r126 65 84 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r127 65 67 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=1.15
+ $Y2=0
r128 63 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r129 63 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r130 61 77 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.37
+ $Y2=0
r131 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.625
+ $Y2=0
r132 60 81 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.71 $Y=0 $X2=5.29
+ $Y2=0
r133 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=0 $X2=4.625
+ $Y2=0
r134 58 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.45
+ $Y2=0
r135 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.785
+ $Y2=0
r136 57 77 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=4.37
+ $Y2=0
r137 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.785
+ $Y2=0
r138 55 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.53
+ $Y2=0
r139 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.945
+ $Y2=0
r140 54 74 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.45
+ $Y2=0
r141 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.945
+ $Y2=0
r142 52 67 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.15
+ $Y2=0
r143 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.265
+ $Y2=0
r144 48 90 2.94129 $w=3.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.725 $Y=0.085
+ $X2=5.767 $Y2=0
r145 48 50 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=5.725 $Y=0.085
+ $X2=5.725 $Y2=0.38
r146 44 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0
r147 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0.38
r148 40 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0
r149 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0.38
r150 36 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0
r151 36 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.38
r152 32 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r153 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.38
r154 31 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.265
+ $Y2=0
r155 30 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0 $X2=2.105
+ $Y2=0
r156 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=1.35
+ $Y2=0
r157 26 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=0.085
+ $X2=1.265 $Y2=0
r158 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.265 $Y=0.085
+ $X2=1.265 $Y2=0.38
r159 22 84 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.255 $Y2=0
r160 22 24 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.382 $Y2=0.38
r161 7 50 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=5.33
+ $Y=0.235 $X2=5.72 $Y2=0.38
r162 6 46 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.235 $X2=4.625 $Y2=0.38
r163 5 42 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.785 $Y2=0.38
r164 4 38 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.945 $Y2=0.38
r165 3 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.105 $Y2=0.38
r166 2 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.265 $Y2=0.38
r167 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.38
.ends


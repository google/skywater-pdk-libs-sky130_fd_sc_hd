* File: sky130_fd_sc_hd__clkinv_8.spice
* Created: Tue Sep  1 19:01:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkinv_8.pex.spice"
.subckt sky130_fd_sc_hd__clkinv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.2 A=0.063
+ P=1.14 MULT=1
MM1002 N_Y_M1001_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.8 A=0.063
+ P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.3 A=0.063
+ P=1.14 MULT=1
MM1008 N_Y_M1005_d N_A_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75001.9 A=0.063
+ P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9 SB=75001.5 A=0.063
+ P=1.14 MULT=1
MM1011 N_Y_M1009_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75001.1 A=0.063
+ P=1.14 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1017 N_Y_M1016_d N_A_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75004.8 A=0.15
+ P=2.3 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.1375 PD=1.27 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75004.4
+ A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.1375 PD=1.27 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75004 A=0.15
+ P=2.3 MULT=1
MM1006 N_Y_M1004_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75003.5
+ A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75003.1
+ A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1007_d N_A_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75002.7
+ A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1013 N_Y_M1012_d N_A_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1014 N_Y_M1014_d N_A_M1014_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1014_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1019 N_Y_M1018_d N_A_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__clkinv_8.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__ha_2.spice.SKY130_FD_SC_HD__HA_2.pxi
* Created: Thu Aug 27 14:22:05 2020
* 
x_PM_SKY130_FD_SC_HD__HA_2%A_79_21# N_A_79_21#_M1012_s N_A_79_21#_M1005_d
+ N_A_79_21#_c_92_n N_A_79_21#_M1015_g N_A_79_21#_M1004_g N_A_79_21#_c_93_n
+ N_A_79_21#_M1016_g N_A_79_21#_M1010_g N_A_79_21#_c_94_n N_A_79_21#_c_95_n
+ N_A_79_21#_c_96_n N_A_79_21#_c_97_n N_A_79_21#_c_122_p N_A_79_21#_c_105_p
+ N_A_79_21#_c_98_n N_A_79_21#_c_99_n PM_SKY130_FD_SC_HD__HA_2%A_79_21#
x_PM_SKY130_FD_SC_HD__HA_2%A_342_199# N_A_342_199#_M1013_s N_A_342_199#_M1009_d
+ N_A_342_199#_M1005_g N_A_342_199#_M1012_g N_A_342_199#_c_168_n
+ N_A_342_199#_M1002_g N_A_342_199#_M1000_g N_A_342_199#_c_169_n
+ N_A_342_199#_M1006_g N_A_342_199#_M1008_g N_A_342_199#_c_170_n
+ N_A_342_199#_c_171_n N_A_342_199#_c_197_n N_A_342_199#_c_199_n
+ N_A_342_199#_c_172_n N_A_342_199#_c_173_n N_A_342_199#_c_174_n
+ N_A_342_199#_c_250_p N_A_342_199#_c_227_p N_A_342_199#_c_175_n
+ N_A_342_199#_c_183_n N_A_342_199#_c_234_p N_A_342_199#_c_176_n
+ PM_SKY130_FD_SC_HD__HA_2%A_342_199#
x_PM_SKY130_FD_SC_HD__HA_2%B N_B_M1003_g N_B_M1011_g N_B_c_303_n N_B_c_310_n
+ N_B_M1009_g N_B_c_304_n N_B_M1013_g N_B_c_305_n B B N_B_c_307_n N_B_c_313_n
+ N_B_c_314_n N_B_c_315_n PM_SKY130_FD_SC_HD__HA_2%B
x_PM_SKY130_FD_SC_HD__HA_2%A N_A_c_379_n N_A_M1017_g N_A_c_380_n N_A_M1007_g
+ N_A_M1014_g N_A_M1001_g A A N_A_c_383_n N_A_c_384_n PM_SKY130_FD_SC_HD__HA_2%A
x_PM_SKY130_FD_SC_HD__HA_2%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1007_d
+ N_VPWR_M1001_d N_VPWR_M1008_s N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n
+ N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_459_n VPWR N_VPWR_c_460_n
+ N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n
+ N_VPWR_c_466_n N_VPWR_c_453_n PM_SKY130_FD_SC_HD__HA_2%VPWR
x_PM_SKY130_FD_SC_HD__HA_2%SUM N_SUM_M1015_s N_SUM_M1004_s SUM SUM SUM SUM SUM
+ SUM N_SUM_c_538_n SUM SUM PM_SKY130_FD_SC_HD__HA_2%SUM
x_PM_SKY130_FD_SC_HD__HA_2%COUT N_COUT_M1002_d N_COUT_M1000_d N_COUT_c_557_n
+ N_COUT_c_559_n N_COUT_c_555_n COUT COUT COUT N_COUT_c_567_n N_COUT_c_570_n
+ PM_SKY130_FD_SC_HD__HA_2%COUT
x_PM_SKY130_FD_SC_HD__HA_2%VGND N_VGND_M1015_d N_VGND_M1016_d N_VGND_M1011_d
+ N_VGND_M1014_d N_VGND_M1006_s N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n
+ N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n VGND
+ N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n N_VGND_c_586_n
+ N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n PM_SKY130_FD_SC_HD__HA_2%VGND
x_PM_SKY130_FD_SC_HD__HA_2%A_389_47# N_A_389_47#_M1012_d N_A_389_47#_M1017_d
+ N_A_389_47#_c_677_n N_A_389_47#_c_658_n N_A_389_47#_c_659_n
+ N_A_389_47#_c_665_n PM_SKY130_FD_SC_HD__HA_2%A_389_47#
cc_1 VNB N_A_79_21#_c_92_n 0.0223279f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_93_n 0.0200913f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.995
cc_3 VNB N_A_79_21#_c_94_n 0.0116115f $X=-0.19 $Y=-0.24 $X2=1.42 $Y2=1.16
cc_4 VNB N_A_79_21#_c_95_n 0.0629369f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_5 VNB N_A_79_21#_c_96_n 0.00964267f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.075
cc_6 VNB N_A_79_21#_c_97_n 0.00125104f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=2.205
cc_7 VNB N_A_79_21#_c_98_n 0.0103009f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=0.51
cc_8 VNB N_A_79_21#_c_99_n 0.00195951f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.16
cc_9 VNB N_A_342_199#_M1012_g 0.0326946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_342_199#_c_168_n 0.0170517f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.56
cc_11 VNB N_A_342_199#_c_169_n 0.0223279f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_12 VNB N_A_342_199#_c_170_n 0.00138473f $X=-0.19 $Y=-0.24 $X2=2.055 $Y2=2.29
cc_13 VNB N_A_342_199#_c_171_n 0.0263526f $X=-0.19 $Y=-0.24 $X2=2.055 $Y2=2.29
cc_14 VNB N_A_342_199#_c_172_n 0.00118612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_342_199#_c_173_n 0.00829257f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_16 VNB N_A_342_199#_c_174_n 8.28664e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_342_199#_c_175_n 0.00594101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_342_199#_c_176_n 0.0509254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_M1011_g 0.0322068f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_B_c_303_n 0.020525f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_21 VNB N_B_c_304_n 0.0172037f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.995
cc_22 VNB N_B_c_305_n 0.0266851f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.985
cc_23 VNB B 0.00480754f $X=-0.19 $Y=-0.24 $X2=1.42 $Y2=1.16
cc_24 VNB N_B_c_307_n 0.0186354f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.075
cc_25 VNB N_A_c_379_n 0.0175235f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=0.235
cc_26 VNB N_A_c_380_n 0.0546964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_M1014_g 0.0349984f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_28 VNB A 0.0175793f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.56
cc_29 VNB N_A_c_383_n 0.0219773f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=2.205
cc_30 VNB N_A_c_384_n 0.00202406f $X=-0.19 $Y=-0.24 $X2=2.055 $Y2=2.29
cc_31 VNB N_VPWR_c_453_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB SUM 0.00205656f $X=-0.19 $Y=-0.24 $X2=1.59 $Y2=2.29
cc_33 VNB N_COUT_c_555_n 0.00179388f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_34 VNB N_VGND_c_575_n 0.0111236f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.56
cc_35 VNB N_VGND_c_576_n 0.00845804f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.985
cc_36 VNB N_VGND_c_577_n 0.0060017f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_37 VNB N_VGND_c_578_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.675
cc_38 VNB N_VGND_c_579_n 0.00513775f $X=-0.19 $Y=-0.24 $X2=1.59 $Y2=2.29
cc_39 VNB N_VGND_c_580_n 0.0111236f $X=-0.19 $Y=-0.24 $X2=2.055 $Y2=2.29
cc_40 VNB N_VGND_c_581_n 0.00845804f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.51
cc_41 VNB N_VGND_c_582_n 0.0188312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_583_n 0.0287637f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_43 VNB N_VGND_c_584_n 0.0425615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_585_n 0.0188312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_586_n 0.00375078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_587_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_588_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_589_n 0.301379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_389_47#_c_658_n 0.00555527f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_50 VNB N_A_389_47#_c_659_n 0.00791132f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_51 VPB N_A_79_21#_M1004_g 0.0263924f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_52 VPB N_A_79_21#_M1010_g 0.0231298f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.985
cc_53 VPB N_A_79_21#_c_95_n 0.0144714f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_54 VPB N_A_79_21#_c_97_n 0.011113f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=2.205
cc_55 VPB N_A_342_199#_M1005_g 0.0430964f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_56 VPB N_A_342_199#_M1000_g 0.0195145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_342_199#_M1008_g 0.0263924f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.075
cc_58 VPB N_A_342_199#_c_170_n 0.00942154f $X=-0.19 $Y=1.305 $X2=2.055 $Y2=2.29
cc_59 VPB N_A_342_199#_c_171_n 0.00612068f $X=-0.19 $Y=1.305 $X2=2.055 $Y2=2.29
cc_60 VPB N_A_342_199#_c_175_n 0.00199884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_342_199#_c_183_n 0.00219138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_342_199#_c_176_n 0.00966569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B_M1003_g 0.0341019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_B_c_303_n 0.00290926f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_65 VPB N_B_c_310_n 0.018537f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_66 VPB B 8.93051e-19 $X=-0.19 $Y=1.305 $X2=1.42 $Y2=1.16
cc_67 VPB N_B_c_307_n 0.0132099f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.075
cc_68 VPB N_B_c_313_n 0.0118224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_B_c_314_n 0.0429383f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=0.51
cc_70 VPB N_B_c_315_n 0.0027266f $X=-0.19 $Y=1.305 $X2=1.66 $Y2=0.51
cc_71 VPB N_A_c_380_n 0.00469083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_M1007_g 0.0433878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_M1001_g 0.0381634f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.995
cc_74 VPB A 0.00477671f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.56
cc_75 VPB N_A_c_383_n 0.0124602f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=2.205
cc_76 VPB N_VPWR_c_454_n 0.0110977f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.56
cc_77 VPB N_VPWR_c_455_n 0.00512364f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.985
cc_78 VPB N_VPWR_c_456_n 0.00483809f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_79 VPB N_VPWR_c_457_n 0.00208414f $X=-0.19 $Y=1.305 $X2=1.59 $Y2=2.29
cc_80 VPB N_VPWR_c_458_n 0.0110977f $X=-0.19 $Y=1.305 $X2=2.055 $Y2=2.29
cc_81 VPB N_VPWR_c_459_n 0.00451915f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=0.51
cc_82 VPB N_VPWR_c_460_n 0.018777f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_83 VPB N_VPWR_c_461_n 0.0142926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_462_n 0.0158669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_463_n 0.00372488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_464_n 0.0410079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_465_n 0.0149234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_466_n 0.00507461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_453_n 0.0469552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB SUM 0.00299561f $X=-0.19 $Y=1.305 $X2=1.59 $Y2=2.29
cc_91 VPB N_COUT_c_555_n 0.00261475f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_92 N_A_79_21#_c_97_n N_A_342_199#_M1005_g 0.0109503f $X=1.505 $Y=2.205 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_105_p N_A_342_199#_M1005_g 0.00982513f $X=2.055 $Y=2.29 $X2=0
+ $Y2=0
cc_94 N_A_79_21#_c_96_n N_A_342_199#_M1012_g 0.00893994f $X=1.505 $Y=1.075 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_98_n N_A_342_199#_M1012_g 4.49111e-19 $X=1.66 $Y=0.51 $X2=0
+ $Y2=0
cc_96 N_A_79_21#_c_96_n N_A_342_199#_c_170_n 0.00568393f $X=1.505 $Y=1.075 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_c_97_n N_A_342_199#_c_170_n 0.045158f $X=1.505 $Y=2.205 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_99_n N_A_342_199#_c_170_n 0.0136441f $X=1.505 $Y=1.16 $X2=0
+ $Y2=0
cc_99 N_A_79_21#_c_95_n N_A_342_199#_c_171_n 0.00668568f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_96_n N_A_342_199#_c_171_n 7.0804e-19 $X=1.505 $Y=1.075 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_c_97_n N_A_342_199#_c_171_n 7.0804e-19 $X=1.505 $Y=2.205 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_98_n N_A_342_199#_c_171_n 0.00120572f $X=1.66 $Y=0.51 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_c_99_n N_A_342_199#_c_171_n 0.00165735f $X=1.505 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_79_21#_M1005_d N_A_342_199#_c_197_n 0.00749068f $X=1.92 $Y=1.845
+ $X2=0 $Y2=0
cc_105 N_A_79_21#_c_105_p N_A_342_199#_c_197_n 0.0121596f $X=2.055 $Y=2.29 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_c_105_p N_A_342_199#_c_199_n 0.0103096f $X=2.055 $Y=2.29 $X2=0
+ $Y2=0
cc_107 N_A_79_21#_c_105_p N_B_M1003_g 0.00413799f $X=2.055 $Y=2.29 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_105_p N_A_M1007_g 5.24173e-19 $X=2.055 $Y=2.29 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_97_n N_VPWR_M1010_d 0.0102227f $X=1.505 $Y=2.205 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_122_p N_VPWR_M1010_d 0.00520436f $X=1.59 $Y=2.29 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_105_p N_VPWR_M1010_d 0.00603148f $X=2.055 $Y=2.29 $X2=0
+ $Y2=0
cc_112 N_A_79_21#_M1004_g N_VPWR_c_455_n 0.00472699f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_79_21#_M1010_g N_VPWR_c_456_n 0.00442456f $X=0.93 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_79_21#_c_94_n N_VPWR_c_456_n 0.0104923f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_95_n N_VPWR_c_456_n 0.00466049f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_97_n N_VPWR_c_456_n 0.0510412f $X=1.505 $Y=2.205 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_122_p N_VPWR_c_456_n 0.0139598f $X=1.59 $Y=2.29 $X2=0 $Y2=0
cc_118 N_A_79_21#_M1004_g N_VPWR_c_460_n 0.00585385f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_79_21#_M1010_g N_VPWR_c_460_n 0.00543342f $X=0.93 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_79_21#_c_122_p N_VPWR_c_464_n 0.00750156f $X=1.59 $Y=2.29 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_105_p N_VPWR_c_464_n 0.022136f $X=2.055 $Y=2.29 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_105_p N_VPWR_c_465_n 0.00475651f $X=2.055 $Y=2.29 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_M1005_d N_VPWR_c_453_n 0.00224151f $X=1.92 $Y=1.845 $X2=0
+ $Y2=0
cc_124 N_A_79_21#_M1004_g N_VPWR_c_453_n 0.0115186f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_79_21#_M1010_g N_VPWR_c_453_n 0.010934f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_122_p N_VPWR_c_453_n 0.00622661f $X=1.59 $Y=2.29 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_105_p N_VPWR_c_453_n 0.0211574f $X=2.055 $Y=2.29 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_93_n SUM 0.0032123f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_79_21#_M1010_g SUM 0.0032678f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_79_21#_M1010_g SUM 0.007823f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_93_n N_SUM_c_538_n 0.00409685f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_92_n SUM 0.00295274f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_79_21#_M1004_g SUM 0.00430721f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_93_n SUM 0.00148828f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_79_21#_M1010_g SUM 0.00236575f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_94_n SUM 0.0129844f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_95_n SUM 0.0326808f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_96_n SUM 0.00542253f $X=1.505 $Y=1.075 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_97_n SUM 0.00779359f $X=1.505 $Y=2.205 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_92_n N_VGND_c_576_n 0.00472699f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_93_n N_VGND_c_577_n 0.00442456f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_94_n N_VGND_c_577_n 0.0137319f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_95_n N_VGND_c_577_n 0.00488398f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_96_n N_VGND_c_577_n 0.0156913f $X=1.505 $Y=1.075 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_98_n N_VGND_c_577_n 0.0259068f $X=1.66 $Y=0.51 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_92_n N_VGND_c_582_n 0.00585385f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_93_n N_VGND_c_582_n 0.00543728f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_98_n N_VGND_c_583_n 0.013655f $X=1.66 $Y=0.51 $X2=0 $Y2=0
cc_149 N_A_79_21#_M1012_s N_VGND_c_589_n 0.00390713f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_150 N_A_79_21#_c_92_n N_VGND_c_589_n 0.0115186f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_93_n N_VGND_c_589_n 0.0109354f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_98_n N_VGND_c_589_n 0.0116462f $X=1.66 $Y=0.51 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_96_n N_A_389_47#_c_659_n 0.00598365f $X=1.505 $Y=1.075 $X2=0
+ $Y2=0
cc_154 N_A_79_21#_c_98_n N_A_389_47#_c_659_n 0.00121593f $X=1.66 $Y=0.51 $X2=0
+ $Y2=0
cc_155 N_A_342_199#_c_197_n N_B_M1003_g 0.0159398f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_156 N_A_342_199#_M1012_g N_B_M1011_g 0.0262586f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_342_199#_c_170_n N_B_M1011_g 3.38346e-19 $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_342_199#_c_171_n N_B_M1011_g 0.00512073f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_342_199#_c_197_n N_B_c_310_n 0.0140856f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_160 N_A_342_199#_c_172_n N_B_c_304_n 0.00230203f $X=3.545 $Y=0.51 $X2=0 $Y2=0
cc_161 N_A_342_199#_c_173_n N_B_c_304_n 0.00451667f $X=4.295 $Y=0.8 $X2=0 $Y2=0
cc_162 N_A_342_199#_c_173_n N_B_c_305_n 0.00576518f $X=4.295 $Y=0.8 $X2=0 $Y2=0
cc_163 N_A_342_199#_c_174_n N_B_c_305_n 0.00989613f $X=3.63 $Y=0.8 $X2=0 $Y2=0
cc_164 N_A_342_199#_c_170_n B 0.0147191f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_342_199#_c_171_n B 9.47274e-19 $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_342_199#_M1005_g N_B_c_307_n 0.0414551f $X=1.845 $Y=2.165 $X2=0 $Y2=0
cc_167 N_A_342_199#_c_170_n N_B_c_307_n 0.00629321f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_342_199#_c_171_n N_B_c_307_n 0.0142701f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_342_199#_c_197_n N_B_c_307_n 6.78521e-19 $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_170 N_A_342_199#_c_197_n N_B_c_313_n 0.0643296f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_171 N_A_342_199#_c_197_n N_B_c_314_n 0.0075391f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_172 N_A_342_199#_M1005_g N_B_c_315_n 2.96137e-19 $X=1.845 $Y=2.165 $X2=0
+ $Y2=0
cc_173 N_A_342_199#_c_170_n N_B_c_315_n 0.012184f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_342_199#_c_197_n N_B_c_315_n 0.0220465f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_175 N_A_342_199#_c_172_n N_A_c_379_n 2.76564e-19 $X=3.545 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_342_199#_c_174_n N_A_c_380_n 5.00359e-19 $X=3.63 $Y=0.8 $X2=0 $Y2=0
cc_177 N_A_342_199#_c_197_n N_A_M1007_g 0.0138095f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_178 N_A_342_199#_c_168_n N_A_M1014_g 0.0196549f $X=4.59 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_342_199#_c_173_n N_A_M1014_g 0.0159716f $X=4.295 $Y=0.8 $X2=0 $Y2=0
cc_180 N_A_342_199#_c_175_n N_A_M1014_g 0.00608428f $X=4.38 $Y=1.325 $X2=0 $Y2=0
cc_181 N_A_342_199#_c_176_n N_A_M1014_g 0.0204223f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_342_199#_c_227_p N_A_M1001_g 0.0159329f $X=4.295 $Y=1.94 $X2=0 $Y2=0
cc_183 N_A_342_199#_c_197_n A 0.00482028f $X=3.81 $Y=1.94 $X2=0 $Y2=0
cc_184 N_A_342_199#_c_173_n A 0.0135181f $X=4.295 $Y=0.8 $X2=0 $Y2=0
cc_185 N_A_342_199#_c_174_n A 0.012949f $X=3.63 $Y=0.8 $X2=0 $Y2=0
cc_186 N_A_342_199#_c_227_p A 0.00293961f $X=4.295 $Y=1.94 $X2=0 $Y2=0
cc_187 N_A_342_199#_c_175_n A 0.00576444f $X=4.38 $Y=1.325 $X2=0 $Y2=0
cc_188 N_A_342_199#_c_183_n A 0.0188346f $X=4.38 $Y=1.855 $X2=0 $Y2=0
cc_189 N_A_342_199#_c_234_p A 0.013878f $X=3.895 $Y=1.94 $X2=0 $Y2=0
cc_190 N_A_342_199#_M1000_g N_A_c_383_n 0.0282491f $X=4.59 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_342_199#_c_173_n N_A_c_383_n 0.00139454f $X=4.295 $Y=0.8 $X2=0 $Y2=0
cc_192 N_A_342_199#_c_183_n N_A_c_383_n 0.00690616f $X=4.38 $Y=1.855 $X2=0 $Y2=0
cc_193 N_A_342_199#_c_234_p N_A_c_383_n 8.4874e-19 $X=3.895 $Y=1.94 $X2=0 $Y2=0
cc_194 N_A_342_199#_c_173_n N_A_c_384_n 0.0187786f $X=4.295 $Y=0.8 $X2=0 $Y2=0
cc_195 N_A_342_199#_c_175_n N_A_c_384_n 0.0106648f $X=4.38 $Y=1.325 $X2=0 $Y2=0
cc_196 N_A_342_199#_c_197_n N_VPWR_M1007_d 0.0153144f $X=3.81 $Y=1.94 $X2=0
+ $Y2=0
cc_197 N_A_342_199#_c_227_p N_VPWR_M1001_d 0.0049013f $X=4.295 $Y=1.94 $X2=0
+ $Y2=0
cc_198 N_A_342_199#_c_183_n N_VPWR_M1001_d 0.00621938f $X=4.38 $Y=1.855 $X2=0
+ $Y2=0
cc_199 N_A_342_199#_M1005_g N_VPWR_c_456_n 0.00534062f $X=1.845 $Y=2.165 $X2=0
+ $Y2=0
cc_200 N_A_342_199#_M1000_g N_VPWR_c_457_n 0.00883088f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_342_199#_M1008_g N_VPWR_c_457_n 6.44697e-19 $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_A_342_199#_c_227_p N_VPWR_c_457_n 0.0167679f $X=4.295 $Y=1.94 $X2=0
+ $Y2=0
cc_203 N_A_342_199#_M1008_g N_VPWR_c_459_n 0.00332104f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_342_199#_c_197_n N_VPWR_c_461_n 0.00205996f $X=3.81 $Y=1.94 $X2=0
+ $Y2=0
cc_205 N_A_342_199#_c_250_p N_VPWR_c_461_n 0.00673756f $X=3.895 $Y=2.19 $X2=0
+ $Y2=0
cc_206 N_A_342_199#_c_227_p N_VPWR_c_461_n 0.00284087f $X=4.295 $Y=1.94 $X2=0
+ $Y2=0
cc_207 N_A_342_199#_M1000_g N_VPWR_c_462_n 0.0046653f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_342_199#_M1008_g N_VPWR_c_462_n 0.00585385f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_342_199#_M1005_g N_VPWR_c_464_n 0.00375986f $X=1.845 $Y=2.165 $X2=0
+ $Y2=0
cc_210 N_A_342_199#_c_197_n N_VPWR_c_464_n 0.0086359f $X=3.81 $Y=1.94 $X2=0
+ $Y2=0
cc_211 N_A_342_199#_c_197_n N_VPWR_c_465_n 0.0492167f $X=3.81 $Y=1.94 $X2=0
+ $Y2=0
cc_212 N_A_342_199#_c_250_p N_VPWR_c_465_n 0.0117111f $X=3.895 $Y=2.19 $X2=0
+ $Y2=0
cc_213 N_A_342_199#_M1009_d N_VPWR_c_453_n 0.00293334f $X=3.75 $Y=1.845 $X2=0
+ $Y2=0
cc_214 N_A_342_199#_M1005_g N_VPWR_c_453_n 0.00668517f $X=1.845 $Y=2.165 $X2=0
+ $Y2=0
cc_215 N_A_342_199#_M1000_g N_VPWR_c_453_n 0.00807415f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_342_199#_M1008_g N_VPWR_c_453_n 0.0115984f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_342_199#_c_197_n N_VPWR_c_453_n 0.0236524f $X=3.81 $Y=1.94 $X2=0
+ $Y2=0
cc_218 N_A_342_199#_c_250_p N_VPWR_c_453_n 0.00602802f $X=3.895 $Y=2.19 $X2=0
+ $Y2=0
cc_219 N_A_342_199#_c_227_p N_VPWR_c_453_n 0.00664813f $X=4.295 $Y=1.94 $X2=0
+ $Y2=0
cc_220 N_A_342_199#_c_197_n A_468_369# 0.00862175f $X=3.81 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_342_199#_c_168_n N_COUT_c_557_n 0.00361485f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_342_199#_c_176_n N_COUT_c_557_n 0.00149139f $X=5.05 $Y=1.16 $X2=0
+ $Y2=0
cc_223 N_A_342_199#_c_176_n N_COUT_c_559_n 0.00147396f $X=5.05 $Y=1.16 $X2=0
+ $Y2=0
cc_224 N_A_342_199#_c_168_n N_COUT_c_555_n 0.00116399f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_342_199#_M1000_g N_COUT_c_555_n 0.00170159f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_342_199#_c_169_n N_COUT_c_555_n 0.00281758f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_342_199#_M1008_g N_COUT_c_555_n 0.00501951f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_342_199#_c_175_n N_COUT_c_555_n 0.0303257f $X=4.38 $Y=1.325 $X2=0
+ $Y2=0
cc_229 N_A_342_199#_c_183_n N_COUT_c_555_n 0.00897386f $X=4.38 $Y=1.855 $X2=0
+ $Y2=0
cc_230 N_A_342_199#_c_176_n N_COUT_c_555_n 0.0270372f $X=5.05 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_342_199#_c_168_n N_COUT_c_567_n 0.00493456f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_342_199#_c_173_n N_VGND_M1014_d 0.00140691f $X=4.295 $Y=0.8 $X2=0
+ $Y2=0
cc_233 N_A_342_199#_c_175_n N_VGND_M1014_d 0.00223361f $X=4.38 $Y=1.325 $X2=0
+ $Y2=0
cc_234 N_A_342_199#_M1012_g N_VGND_c_577_n 0.00468029f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_A_342_199#_M1012_g N_VGND_c_578_n 0.00155517f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_236 N_A_342_199#_c_168_n N_VGND_c_579_n 0.00287759f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_342_199#_c_173_n N_VGND_c_579_n 0.00481848f $X=4.295 $Y=0.8 $X2=0
+ $Y2=0
cc_238 N_A_342_199#_c_175_n N_VGND_c_579_n 0.0140595f $X=4.38 $Y=1.325 $X2=0
+ $Y2=0
cc_239 N_A_342_199#_c_176_n N_VGND_c_579_n 2.60901e-19 $X=5.05 $Y=1.16 $X2=0
+ $Y2=0
cc_240 N_A_342_199#_c_169_n N_VGND_c_581_n 0.00472699f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_342_199#_M1012_g N_VGND_c_583_n 0.00585385f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_242 N_A_342_199#_c_172_n N_VGND_c_584_n 0.00721428f $X=3.545 $Y=0.51 $X2=0
+ $Y2=0
cc_243 N_A_342_199#_c_173_n N_VGND_c_584_n 0.00851686f $X=4.295 $Y=0.8 $X2=0
+ $Y2=0
cc_244 N_A_342_199#_c_168_n N_VGND_c_585_n 0.00543728f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_342_199#_c_169_n N_VGND_c_585_n 0.00585385f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_342_199#_M1013_s N_VGND_c_589_n 0.00286228f $X=3.42 $Y=0.235 $X2=0
+ $Y2=0
cc_247 N_A_342_199#_M1012_g N_VGND_c_589_n 0.0122169f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_248 N_A_342_199#_c_168_n N_VGND_c_589_n 0.00976597f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_342_199#_c_169_n N_VGND_c_589_n 0.0115186f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_342_199#_c_172_n N_VGND_c_589_n 0.00611891f $X=3.545 $Y=0.51 $X2=0
+ $Y2=0
cc_251 N_A_342_199#_c_173_n N_VGND_c_589_n 0.0143392f $X=4.295 $Y=0.8 $X2=0
+ $Y2=0
cc_252 N_A_342_199#_c_175_n N_VGND_c_589_n 7.42202e-19 $X=4.38 $Y=1.325 $X2=0
+ $Y2=0
cc_253 N_A_342_199#_c_172_n N_A_389_47#_c_658_n 0.0033249f $X=3.545 $Y=0.51
+ $X2=0 $Y2=0
cc_254 N_A_342_199#_c_174_n N_A_389_47#_c_658_n 0.00391993f $X=3.63 $Y=0.8 $X2=0
+ $Y2=0
cc_255 N_A_342_199#_M1012_g N_A_389_47#_c_659_n 0.00183499f $X=1.87 $Y=0.445
+ $X2=0 $Y2=0
cc_256 N_A_342_199#_c_172_n N_A_389_47#_c_665_n 0.0101661f $X=3.545 $Y=0.51
+ $X2=0 $Y2=0
cc_257 N_B_M1011_g N_A_c_379_n 0.0211639f $X=2.29 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_258 N_B_M1011_g N_A_c_380_n 0.00733841f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_259 N_B_c_303_n N_A_c_380_n 0.0139446f $X=3.49 $Y=1.355 $X2=0 $Y2=0
cc_260 N_B_c_305_n N_A_c_380_n 0.00671923f $X=3.755 $Y=0.81 $X2=0 $Y2=0
cc_261 B N_A_c_380_n 0.00655679f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_262 N_B_c_307_n N_A_c_380_n 0.0203161f $X=2.395 $Y=1.26 $X2=0 $Y2=0
cc_263 N_B_c_313_n N_A_c_380_n 0.00726461f $X=3.43 $Y=1.52 $X2=0 $Y2=0
cc_264 N_B_M1003_g N_A_M1007_g 0.0371957f $X=2.265 $Y=2.165 $X2=0 $Y2=0
cc_265 N_B_c_303_n N_A_M1007_g 0.00140216f $X=3.49 $Y=1.355 $X2=0 $Y2=0
cc_266 N_B_c_310_n N_A_M1007_g 0.00665793f $X=3.675 $Y=1.745 $X2=0 $Y2=0
cc_267 N_B_c_313_n N_A_M1007_g 0.01723f $X=3.43 $Y=1.52 $X2=0 $Y2=0
cc_268 N_B_c_314_n N_A_M1007_g 0.0112337f $X=3.49 $Y=1.55 $X2=0 $Y2=0
cc_269 N_B_c_303_n N_A_M1014_g 0.00334809f $X=3.49 $Y=1.355 $X2=0 $Y2=0
cc_270 N_B_c_304_n N_A_M1014_g 0.0489227f $X=3.755 $Y=0.735 $X2=0 $Y2=0
cc_271 N_B_c_313_n N_A_M1001_g 8.33208e-19 $X=3.43 $Y=1.52 $X2=0 $Y2=0
cc_272 N_B_c_314_n N_A_M1001_g 0.0307905f $X=3.49 $Y=1.55 $X2=0 $Y2=0
cc_273 N_B_c_303_n A 0.0125404f $X=3.49 $Y=1.355 $X2=0 $Y2=0
cc_274 N_B_c_305_n A 0.00254958f $X=3.755 $Y=0.81 $X2=0 $Y2=0
cc_275 B A 0.0137085f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_276 N_B_c_313_n A 0.0790947f $X=3.43 $Y=1.52 $X2=0 $Y2=0
cc_277 N_B_c_314_n A 0.00658547f $X=3.49 $Y=1.55 $X2=0 $Y2=0
cc_278 N_B_c_303_n N_A_c_383_n 0.0176486f $X=3.49 $Y=1.355 $X2=0 $Y2=0
cc_279 N_B_c_305_n N_A_c_383_n 0.00363872f $X=3.755 $Y=0.81 $X2=0 $Y2=0
cc_280 N_B_c_310_n N_VPWR_c_461_n 0.00317293f $X=3.675 $Y=1.745 $X2=0 $Y2=0
cc_281 N_B_M1003_g N_VPWR_c_464_n 0.00422171f $X=2.265 $Y=2.165 $X2=0 $Y2=0
cc_282 N_B_M1003_g N_VPWR_c_465_n 0.00199618f $X=2.265 $Y=2.165 $X2=0 $Y2=0
cc_283 N_B_c_310_n N_VPWR_c_465_n 0.0100755f $X=3.675 $Y=1.745 $X2=0 $Y2=0
cc_284 N_B_M1003_g N_VPWR_c_453_n 0.00619671f $X=2.265 $Y=2.165 $X2=0 $Y2=0
cc_285 N_B_c_310_n N_VPWR_c_453_n 0.00387254f $X=3.675 $Y=1.745 $X2=0 $Y2=0
cc_286 N_B_M1011_g N_VGND_c_578_n 0.00853463f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_287 N_B_M1011_g N_VGND_c_583_n 0.00339367f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_288 N_B_c_304_n N_VGND_c_584_n 0.00436487f $X=3.755 $Y=0.735 $X2=0 $Y2=0
cc_289 N_B_c_305_n N_VGND_c_584_n 0.00155105f $X=3.755 $Y=0.81 $X2=0 $Y2=0
cc_290 N_B_M1011_g N_VGND_c_589_n 0.00401529f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_291 N_B_c_304_n N_VGND_c_589_n 0.007316f $X=3.755 $Y=0.735 $X2=0 $Y2=0
cc_292 N_B_c_305_n N_VGND_c_589_n 0.0012507f $X=3.755 $Y=0.81 $X2=0 $Y2=0
cc_293 N_B_M1011_g N_A_389_47#_c_658_n 0.0137182f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_294 N_B_c_304_n N_A_389_47#_c_658_n 3.48618e-19 $X=3.755 $Y=0.735 $X2=0 $Y2=0
cc_295 N_B_c_305_n N_A_389_47#_c_658_n 6.47077e-19 $X=3.755 $Y=0.81 $X2=0 $Y2=0
cc_296 B N_A_389_47#_c_658_n 0.0223308f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_297 N_B_c_307_n N_A_389_47#_c_658_n 0.00181786f $X=2.395 $Y=1.26 $X2=0 $Y2=0
cc_298 N_B_c_313_n N_A_389_47#_c_658_n 0.0049701f $X=3.43 $Y=1.52 $X2=0 $Y2=0
cc_299 N_A_M1001_g N_VPWR_c_457_n 0.00161704f $X=4.115 $Y=2.165 $X2=0 $Y2=0
cc_300 N_A_M1001_g N_VPWR_c_461_n 0.00433717f $X=4.115 $Y=2.165 $X2=0 $Y2=0
cc_301 N_A_M1007_g N_VPWR_c_464_n 0.00317293f $X=2.815 $Y=2.165 $X2=0 $Y2=0
cc_302 N_A_M1007_g N_VPWR_c_465_n 0.0129568f $X=2.815 $Y=2.165 $X2=0 $Y2=0
cc_303 N_A_M1001_g N_VPWR_c_465_n 8.50365e-19 $X=4.115 $Y=2.165 $X2=0 $Y2=0
cc_304 N_A_M1007_g N_VPWR_c_453_n 0.00411949f $X=2.815 $Y=2.165 $X2=0 $Y2=0
cc_305 N_A_M1001_g N_VPWR_c_453_n 0.00602978f $X=4.115 $Y=2.165 $X2=0 $Y2=0
cc_306 N_A_M1014_g N_COUT_c_567_n 8.09418e-19 $X=4.115 $Y=0.445 $X2=0 $Y2=0
cc_307 N_A_c_379_n N_VGND_c_578_n 0.0112612f $X=2.71 $Y=0.735 $X2=0 $Y2=0
cc_308 N_A_M1014_g N_VGND_c_579_n 0.00302106f $X=4.115 $Y=0.445 $X2=0 $Y2=0
cc_309 N_A_c_379_n N_VGND_c_584_n 0.00339367f $X=2.71 $Y=0.735 $X2=0 $Y2=0
cc_310 N_A_c_380_n N_VGND_c_584_n 3.81503e-19 $X=2.815 $Y=1.305 $X2=0 $Y2=0
cc_311 N_A_M1014_g N_VGND_c_584_n 0.00436487f $X=4.115 $Y=0.445 $X2=0 $Y2=0
cc_312 N_A_c_379_n N_VGND_c_589_n 0.00536411f $X=2.71 $Y=0.735 $X2=0 $Y2=0
cc_313 N_A_M1014_g N_VGND_c_589_n 0.00586581f $X=4.115 $Y=0.445 $X2=0 $Y2=0
cc_314 N_A_c_379_n N_A_389_47#_c_658_n 0.00706861f $X=2.71 $Y=0.735 $X2=0 $Y2=0
cc_315 N_A_c_380_n N_A_389_47#_c_658_n 0.0132747f $X=2.815 $Y=1.305 $X2=0 $Y2=0
cc_316 A N_A_389_47#_c_658_n 0.0118158f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_317 N_VPWR_c_453_n N_SUM_M1004_s 0.00285715f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_460_n SUM 0.0147117f $X=1.055 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_c_453_n SUM 0.0121088f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_c_453_n A_468_369# 0.00502228f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_321 N_VPWR_c_453_n N_COUT_M1000_d 0.00467225f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_c_462_n N_COUT_c_570_n 0.0118479f $X=5.145 $Y=2.72 $X2=0 $Y2=0
cc_323 N_VPWR_c_453_n N_COUT_c_570_n 0.00931197f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_c_455_n N_VGND_c_576_n 0.00695811f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_325 N_VPWR_c_459_n N_VGND_c_581_n 0.00695811f $X=5.26 $Y=1.66 $X2=0 $Y2=0
cc_326 N_SUM_c_538_n N_VGND_c_582_n 0.0139874f $X=0.72 $Y=0.4 $X2=0 $Y2=0
cc_327 N_SUM_M1015_s N_VGND_c_589_n 0.00286985f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_328 N_SUM_c_538_n N_VGND_c_589_n 0.0120073f $X=0.72 $Y=0.4 $X2=0 $Y2=0
cc_329 N_COUT_c_567_n N_VGND_c_585_n 0.0139366f $X=4.8 $Y=0.4 $X2=0 $Y2=0
cc_330 N_COUT_M1002_d N_VGND_c_589_n 0.00286985f $X=4.665 $Y=0.235 $X2=0 $Y2=0
cc_331 N_COUT_c_567_n N_VGND_c_589_n 0.0119907f $X=4.8 $Y=0.4 $X2=0 $Y2=0
cc_332 N_VGND_c_589_n N_A_389_47#_M1012_d 0.00416801f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_333 N_VGND_c_589_n N_A_389_47#_M1017_d 0.003754f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_c_583_n N_A_389_47#_c_677_n 0.00701792f $X=2.335 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_589_n N_A_389_47#_c_677_n 0.00608739f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_M1011_d N_A_389_47#_c_658_n 0.00159539f $X=2.365 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_VGND_c_578_n N_A_389_47#_c_658_n 0.0159625f $X=2.5 $Y=0.38 $X2=0 $Y2=0
cc_338 N_VGND_c_583_n N_A_389_47#_c_658_n 0.00243651f $X=2.335 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_584_n N_A_389_47#_c_658_n 0.00243651f $X=4.215 $Y=0 $X2=0 $Y2=0
cc_340 N_VGND_c_589_n N_A_389_47#_c_658_n 0.00990569f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_584_n N_A_389_47#_c_665_n 0.00713694f $X=4.215 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_589_n N_A_389_47#_c_665_n 0.00608739f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_589_n A_766_47# 0.00269901f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a311o_2.spice
* Created: Thu Aug 27 14:04:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a311o_2.spice.pex"
.subckt sky130_fd_sc_hd__a311o_2  VNB VPB A3 A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_79_21#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_79_21#_M1012_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.156 AS=0.08775 PD=1.13 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1002 A_319_47# N_A3_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65 AD=0.1105
+ AS=0.156 PD=0.99 PS=1.13 NRD=21.228 NRS=23.076 M=1 R=4.33333 SA=75001.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1009 A_417_47# N_A2_M1009_g A_319_47# VNB NSHORT L=0.15 W=0.65 AD=0.12025
+ AS=0.1105 PD=1.02 PS=0.99 NRD=23.988 NRS=21.228 M=1 R=4.33333 SA=75001.7
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1001 N_A_79_21#_M1001_d N_A1_M1001_g A_417_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.13325 AS=0.12025 PD=1.06 PS=1.02 NRD=23.988 NRS=23.988 M=1 R=4.33333
+ SA=75002.2 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g N_A_79_21#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.13975 AS=0.13325 PD=1.08 PS=1.06 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1006 N_A_79_21#_M1006_d N_C1_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.13975 PD=1.82 PS=1.08 NRD=0 NRS=12.912 M=1 R=4.33333 SA=75003.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_79_21#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_79_21#_M1010_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.24 AS=0.135 PD=1.48 PS=1.27 NRD=27.5603 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003 A=0.15 P=2.3 MULT=1
MM1011 N_A_319_297#_M1011_d N_A3_M1011_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.17 AS=0.24 PD=1.34 PS=1.48 NRD=3.9203 NRS=11.8003 M=1 R=6.66667
+ SA=75001.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_319_297#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.185 AS=0.17 PD=1.37 PS=1.34 NRD=12.7853 NRS=7.8603 M=1 R=6.66667
+ SA=75001.7 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1013 N_A_319_297#_M1013_d N_A1_M1013_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.185 PD=1.42 PS=1.37 NRD=22.6353 NRS=4.9053 M=1 R=6.66667
+ SA=75002.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1003 A_635_297# N_B1_M1003_g N_A_319_297#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.21 PD=1.42 PS=1.42 NRD=30.5153 NRS=4.9053 M=1 R=6.66667
+ SA=75002.8 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_A_79_21#_M1000_d N_C1_M1000_g A_635_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.21 PD=2.52 PS=1.42 NRD=0 NRS=30.5153 M=1 R=6.66667 SA=75003.4 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__a311o_2.spice.SKY130_FD_SC_HD__A311O_2.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a21oi_1.spice.pex
* Created: Thu Aug 27 14:01:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21OI_1%B1 1 3 6 8 9 16
r29 13 16 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.49 $Y2=1.16
r30 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r31 8 9 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.215 $Y=0.85
+ $X2=0.215 $Y2=1.16
r32 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r34 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_1%A1 3 6 8 9 10 15 17
r39 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.16
+ $X2=0.945 $Y2=1.325
r40 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.16
+ $X2=0.945 $Y2=0.995
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=1.16 $X2=0.945 $Y2=1.16
r42 10 16 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=0.945 $Y2=1.16
r43 10 19 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.15 $Y2=0.995
r44 9 19 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.15 $Y=0.85 $X2=1.15
+ $Y2=0.995
r45 8 9 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.15 $Y=0.51 $X2=1.15
+ $Y2=0.85
r46 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.92 $Y=1.985
+ $X2=0.92 $Y2=1.325
r47 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.92 $Y=0.56 $X2=0.92
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_1%A2 1 3 6 8 13
r27 10 13 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.365 $Y=1.16
+ $X2=1.575 $Y2=1.16
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.16 $X2=1.575 $Y2=1.16
r29 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.985
r31 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_1%Y 1 2 8 15 17 18 19 20
r29 19 20 16.7628 $w=2.73e-07 $l=4e-07 $layer=LI1_cond $X=0.232 $Y=1.81
+ $X2=0.232 $Y2=2.21
r30 17 18 9.81941 $w=2.23e-07 $l=1.8e-07 $layer=LI1_cond $X=0.67 $Y=0.645
+ $X2=0.67 $Y2=0.825
r31 13 19 5.23838 $w=2.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.232 $Y=1.685
+ $X2=0.232 $Y2=1.81
r32 13 15 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.232 $Y=1.59
+ $X2=0.592 $Y2=1.59
r33 11 17 5.15111 $w=2.25e-07 $l=9.5e-08 $layer=LI1_cond $X=0.722 $Y=0.55
+ $X2=0.722 $Y2=0.645
r34 8 15 1.24516 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=0.592 $Y=1.495
+ $X2=0.592 $Y2=1.59
r35 8 18 42.4623 $w=1.73e-07 $l=6.7e-07 $layer=LI1_cond $X=0.592 $Y=1.495
+ $X2=0.592 $Y2=0.825
r36 2 19 300 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=1.485 $X2=0.275 $Y2=1.81
r37 1 11 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_1%A_113_297# 1 2 7 8 9 11
r29 9 17 4.33442 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=1.58 $Y=2.025 $X2=1.58
+ $Y2=1.775
r30 9 11 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.58 $Y=2.025
+ $X2=1.58 $Y2=2.33
r31 8 15 9.70455 $w=2.2e-07 $l=2.43926e-07 $layer=LI1_cond $X=0.87 $Y=1.775
+ $X2=0.705 $Y2=1.95
r32 7 17 2.86072 $w=5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=1.775 $X2=1.58
+ $Y2=1.775
r33 7 8 13.0373 $w=4.98e-07 $l=5.45e-07 $layer=LI1_cond $X=1.415 $Y=1.775
+ $X2=0.87 $Y2=1.775
r34 2 17 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.485 $X2=1.58 $Y2=1.65
r35 2 11 400 $w=1.7e-07 $l=9.12318e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.485 $X2=1.58 $Y2=2.33
r36 1 15 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.705 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_1%VPWR 1 6 8 10 17 18 21
r28 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 15 21 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.137 $Y2=2.72
r32 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.61 $Y2=2.72
r33 13 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r35 10 21 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.04 $Y=2.72
+ $X2=1.137 $Y2=2.72
r36 10 12 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.04 $Y=2.72
+ $X2=0.69 $Y2=2.72
r37 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 4 21 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.137 $Y=2.635
+ $X2=1.137 $Y2=2.72
r39 4 6 15.641 $w=1.93e-07 $l=2.75e-07 $layer=LI1_cond $X=1.137 $Y=2.635
+ $X2=1.137 $Y2=2.36
r40 1 6 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.135 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_1%VGND 1 2 7 9 11 13 15 17 27
r30 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r31 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r32 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r33 18 23 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r34 18 20 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=1.15
+ $Y2=0
r35 17 26 4.50146 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.642
+ $Y2=0
r36 17 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.15
+ $Y2=0
r37 15 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r38 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r39 11 26 3.01621 $w=3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.595 $Y=0.085
+ $X2=1.642 $Y2=0
r40 11 13 17.0946 $w=2.98e-07 $l=4.45e-07 $layer=LI1_cond $X=1.595 $Y=0.085
+ $X2=1.595 $Y2=0.53
r41 7 23 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r42 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r43 2 13 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.58 $Y2=0.53
r44 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends


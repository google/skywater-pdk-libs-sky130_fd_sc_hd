# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__clkdlybuf4s18_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.560000 1.290000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 0.270000 3.150000 0.640000 ;
        RECT 2.715000 1.420000 3.180000 1.525000 ;
        RECT 2.715000 1.525000 3.150000 2.465000 ;
        RECT 2.965000 0.640000 3.150000 0.780000 ;
        RECT 2.965000 0.780000 3.180000 0.945000 ;
        RECT 3.010000 0.945000 3.180000 1.420000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.585000  0.085000 0.915000 0.565000 ;
        RECT 2.165000  0.085000 2.535000 0.565000 ;
        RECT 3.320000  0.085000 3.595000 0.645000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.600000 1.800000 0.930000 2.635000 ;
        RECT 2.130000 1.800000 2.545000 2.635000 ;
        RECT 3.320000 1.625000 3.595000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.270000 0.415000 0.735000 ;
      RECT 0.085000 0.735000 1.055000 0.905000 ;
      RECT 0.085000 1.460000 1.055000 1.630000 ;
      RECT 0.085000 1.630000 0.430000 2.465000 ;
      RECT 0.730000 0.905000 1.055000 1.460000 ;
      RECT 1.110000 1.800000 1.440000 2.465000 ;
      RECT 1.160000 0.270000 1.440000 0.600000 ;
      RECT 1.270000 0.600000 1.440000 1.075000 ;
      RECT 1.270000 1.075000 2.205000 1.255000 ;
      RECT 1.270000 1.255000 1.440000 1.800000 ;
      RECT 1.630000 0.270000 1.960000 0.735000 ;
      RECT 1.630000 0.735000 2.545000 0.905000 ;
      RECT 1.630000 1.460000 2.545000 1.630000 ;
      RECT 1.630000 1.630000 1.960000 2.465000 ;
      RECT 2.375000 0.905000 2.545000 1.075000 ;
      RECT 2.375000 1.075000 2.840000 1.245000 ;
      RECT 2.375000 1.245000 2.545000 1.460000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_2
END LIBRARY

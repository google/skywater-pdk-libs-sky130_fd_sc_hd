* File: sky130_fd_sc_hd__lpflow_isobufsrc_8.spice
* Created: Thu Aug 27 14:25:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_isobufsrc_8.spice.pex"
.subckt sky130_fd_sc_hd__lpflow_isobufsrc_8  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1023 N_A_123_297#_M1023_d N_A_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75007.7 A=0.0975 P=1.6 MULT=1
MM1025 N_A_123_297#_M1023_d N_A_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.19825 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75007.2 A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1002_d N_A_123_297#_M1002_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.19825 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75006.5 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1002_d N_A_123_297#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.8
+ SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_123_297#_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1007_d N_A_123_297#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75005.2 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1013_d N_A_123_297#_M1013_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1028 N_X_M1013_d N_A_123_297#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1032 N_X_M1032_d N_A_123_297#_M1032_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.9
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1035 N_X_M1032_d N_A_123_297#_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.3
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1035_s N_SLEEP_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_SLEEP_M1006_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.1
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1006_d N_SLEEP_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.6
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_SLEEP_M1015_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1015_d N_SLEEP_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.4
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_SLEEP_M1018_g N_X_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.8
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1018_d N_SLEEP_M1019_g N_X_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_SLEEP_M1021_g N_X_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_123_297#_M1010_d N_A_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1029 N_A_123_297#_M1010_d N_A_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_321_297#_M1000_d N_A_123_297#_M1000_g N_VPWR_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75006.5 A=0.15 P=2.3 MULT=1
MM1001 N_A_321_297#_M1001_d N_A_123_297#_M1001_g N_VPWR_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75006.1 A=0.15 P=2.3 MULT=1
MM1014 N_A_321_297#_M1001_d N_A_123_297#_M1014_g N_VPWR_M1014_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75005.7 A=0.15 P=2.3 MULT=1
MM1022 N_A_321_297#_M1022_d N_A_123_297#_M1022_g N_VPWR_M1014_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.5 SB=75005.2 A=0.15 P=2.3 MULT=1
MM1024 N_A_321_297#_M1022_d N_A_123_297#_M1024_g N_VPWR_M1024_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75004.8 A=0.15 P=2.3 MULT=1
MM1026 N_A_321_297#_M1026_d N_A_123_297#_M1026_g N_VPWR_M1024_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75004.4 A=0.15 P=2.3 MULT=1
MM1027 N_A_321_297#_M1026_d N_A_123_297#_M1027_g N_VPWR_M1027_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75004 A=0.15 P=2.3 MULT=1
MM1033 N_A_321_297#_M1033_d N_A_123_297#_M1033_g N_VPWR_M1027_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.1 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1004_d N_SLEEP_M1004_g N_A_321_297#_M1033_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1004_d N_SLEEP_M1011_g N_A_321_297#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1012 N_X_M1012_d N_SLEEP_M1012_g N_A_321_297#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1017 N_X_M1012_d N_SLEEP_M1017_g N_A_321_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1020 N_X_M1020_d N_SLEEP_M1020_g N_A_321_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1030 N_X_M1020_d N_SLEEP_M1030_g N_A_321_297#_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.7
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1031 N_X_M1031_d N_SLEEP_M1031_g N_A_321_297#_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1034 N_X_M1031_d N_SLEEP_M1034_g N_A_321_297#_M1034_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX36_noxref VNB VPB NWDIODE A=14.6376 P=21.45
*
.include "sky130_fd_sc_hd__lpflow_isobufsrc_8.spice.SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8.pxi"
*
.ends
*
*

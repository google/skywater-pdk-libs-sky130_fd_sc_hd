# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.400000 1.075000 1.410000 1.330000 ;
        RECT 0.965000 1.330000 1.410000 1.515000 ;
        RECT 0.965000 1.515000 3.630000 1.685000 ;
        RECT 3.350000 0.995000 3.630000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705000 1.075000 3.180000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.800000 0.995000 4.975000 1.410000 ;
        RECT 4.260000 1.410000 4.975000 1.515000 ;
        RECT 4.260000 1.515000 7.000000 1.685000 ;
        RECT 6.830000 0.995000 7.000000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.370000 1.075000 6.440000 1.345000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.001000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 1.855000 7.680000 2.025000 ;
        RECT 1.805000 2.025000 3.470000 2.105000 ;
        RECT 4.045000 2.025000 7.680000 2.105000 ;
        RECT 5.280000 0.270000 6.735000 0.450000 ;
        RECT 6.565000 0.450000 6.735000 0.655000 ;
        RECT 6.565000 0.655000 7.350000 0.825000 ;
        RECT 7.170000 0.825000 7.350000 1.340000 ;
        RECT 7.170000 1.340000 7.680000 1.855000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  1.665000 0.385000 2.635000 ;
      RECT 0.155000  0.535000 0.355000 0.625000 ;
      RECT 0.155000  0.625000 1.240000 0.695000 ;
      RECT 0.155000  0.695000 3.835000 0.795000 ;
      RECT 0.155000  0.795000 3.130000 0.865000 ;
      RECT 0.155000  0.865000 1.795000 0.905000 ;
      RECT 0.525000  0.085000 0.855000 0.445000 ;
      RECT 0.555000  1.860000 0.775000 1.935000 ;
      RECT 0.555000  1.935000 1.635000 2.105000 ;
      RECT 0.555000  2.105000 0.775000 2.190000 ;
      RECT 0.955000  2.275000 1.285000 2.635000 ;
      RECT 1.025000  0.425000 1.240000 0.625000 ;
      RECT 1.455000  2.105000 1.635000 2.275000 ;
      RECT 1.455000  2.275000 3.435000 2.465000 ;
      RECT 1.465000  0.085000 1.635000 0.525000 ;
      RECT 1.775000  0.625000 3.835000 0.695000 ;
      RECT 2.245000  0.085000 2.575000 0.445000 ;
      RECT 3.105000  0.085000 3.435000 0.445000 ;
      RECT 3.605000  0.255000 4.920000 0.455000 ;
      RECT 3.605000  0.455000 3.835000 0.625000 ;
      RECT 3.615000  2.195000 3.885000 2.635000 ;
      RECT 4.005000  0.635000 6.170000 0.815000 ;
      RECT 4.435000  2.275000 4.765000 2.635000 ;
      RECT 5.280000  2.275000 5.610000 2.635000 ;
      RECT 6.120000  2.275000 6.455000 2.635000 ;
      RECT 6.980000  0.310000 7.680000 0.480000 ;
      RECT 7.355000  2.275000 7.685000 2.635000 ;
      RECT 7.510000  0.480000 7.680000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.425000 1.240000 0.595000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.510000  0.425000 7.680000 0.595000 ;
    LAYER met1 ;
      RECT 1.010000 0.395000 1.300000 0.440000 ;
      RECT 1.010000 0.440000 7.740000 0.580000 ;
      RECT 1.010000 0.580000 1.300000 0.625000 ;
      RECT 7.450000 0.395000 7.740000 0.440000 ;
      RECT 7.450000 0.580000 7.740000 0.625000 ;
  END
END sky130_fd_sc_hd__o211ai_4
END LIBRARY

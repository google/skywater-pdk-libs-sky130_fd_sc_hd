* NGSPICE file created from sky130_fd_sc_hd__nor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
M1000 VPWR A a_193_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u
M1001 a_193_297# B a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1002 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=3.445e+11p ps=3.66e+06u
M1003 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_109_297# C Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1005 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


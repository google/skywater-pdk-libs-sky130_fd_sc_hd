* File: sky130_fd_sc_hd__a31oi_1.spice.pex
* Created: Thu Aug 27 14:04:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A31OI_1%A3 1 3 6 8 14
r23 11 14 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r24 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r25 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r26 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r27 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r28 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%A2 3 6 8 9 10 15 17
c39 15 0 1.83054e-19 $X=0.89 $Y=1.16
c40 6 0 1.1986e-20 $X=0.89 $Y=1.985
r41 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r43 10 16 0.776928 $w=4.43e-07 $l=3e-08 $layer=LI1_cond $X=0.832 $Y=1.19
+ $X2=0.832 $Y2=1.16
r44 9 16 8.02825 $w=4.43e-07 $l=3.1e-07 $layer=LI1_cond $X=0.832 $Y=0.85
+ $X2=0.832 $Y2=1.16
r45 8 9 8.80518 $w=4.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.832 $Y=0.51
+ $X2=0.832 $Y2=0.85
r46 4 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r47 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r48 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.83 $Y=0.56 $X2=0.83
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%A1 3 6 10 11 13 16 21
c42 21 0 1.15177e-19 $X=1.362 $Y=1.555
r43 13 21 10.8434 $w=2.18e-07 $l=2.07e-07 $layer=LI1_cond $X=1.155 $Y=1.555
+ $X2=1.362 $Y2=1.555
r44 11 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.37 $Y2=1.325
r45 11 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.37 $Y2=0.995
r46 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r47 8 21 1.7811 $w=1.85e-07 $l=1.1e-07 $layer=LI1_cond $X=1.362 $Y=1.445
+ $X2=1.362 $Y2=1.555
r48 8 10 17.086 $w=1.83e-07 $l=2.85e-07 $layer=LI1_cond $X=1.362 $Y=1.445
+ $X2=1.362 $Y2=1.16
r49 6 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.345 $Y=1.985
+ $X2=1.345 $Y2=1.325
r50 3 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.345 $Y=0.56
+ $X2=1.345 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%B1 1 3 6 8 13
c28 6 0 1.15177e-19 $X=1.82 $Y=1.985
r29 10 13 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=2.06 $Y2=1.16
r30 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r31 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.325
+ $X2=1.82 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.82 $Y=1.325 $X2=1.82
+ $Y2=1.985
r33 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.82 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%VPWR 1 2 7 9 15 17 19 26 27 33
r40 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r41 27 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r44 24 26 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 20 30 4.79676 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=2.72 $X2=0.21
+ $Y2=2.72
r48 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.42 $Y=2.72 $X2=0.69
+ $Y2=2.72
r49 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r50 19 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 17 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r54 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2.34
r55 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=2.34
r56 7 30 2.96942 $w=3.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.21 $Y2=2.72
r57 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=2.34
r58 2 15 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r59 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r60 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%A_109_297# 1 2 9 11 12 15
c21 12 0 1.83054e-19 $X=0.765 $Y=1.92
r22 13 15 12.5488 $w=2.23e-07 $l=2.45e-07 $layer=LI1_cond $X=1.582 $Y=2.005
+ $X2=1.582 $Y2=2.25
r23 11 13 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.47 $Y=1.92
+ $X2=1.582 $Y2=2.005
r24 11 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.47 $Y=1.92
+ $X2=0.765 $Y2=1.92
r25 7 12 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.677 $Y=2.005
+ $X2=0.765 $Y2=1.92
r26 7 9 15.5273 $w=1.73e-07 $l=2.45e-07 $layer=LI1_cond $X=0.677 $Y=2.005
+ $X2=0.677 $Y2=2.25
r27 2 15 600 $w=1.7e-07 $l=8.29759e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.485 $X2=1.555 $Y2=2.25
r28 1 9 600 $w=1.7e-07 $l=8.29759e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%Y 1 2 9 12 14 18 21 22
c39 14 0 1.35623e-19 $X=1.587 $Y=0.825
c40 12 0 1.1986e-20 $X=1.71 $Y=1.495
r41 22 30 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=2.042 $Y=2.21
+ $X2=2.042 $Y2=2.34
r42 21 22 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.042 $Y=1.87
+ $X2=2.042 $Y2=2.21
r43 18 21 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=2.042 $Y=1.665
+ $X2=2.042 $Y2=1.87
r44 15 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.71 $Y=1.58
+ $X2=2.04 $Y2=1.58
r45 13 14 7.10376 $w=4.03e-07 $l=1.1e-07 $layer=LI1_cond $X=1.587 $Y=0.715
+ $X2=1.587 $Y2=0.825
r46 12 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.495
+ $X2=1.71 $Y2=1.58
r47 12 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.71 $Y=1.495
+ $X2=1.71 $Y2=0.825
r48 9 13 9.53255 $w=4.03e-07 $l=3.35e-07 $layer=LI1_cond $X=1.582 $Y=0.38
+ $X2=1.582 $Y2=0.715
r49 2 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.04 $Y2=2.34
r50 2 18 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.04 $Y2=1.66
r51 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.235 $X2=1.555 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A31OI_1%VGND 1 2 7 9 11 13 15 17 30
c32 17 0 1.35623e-19 $X=1.955 $Y=0
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r34 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r35 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r36 21 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r37 20 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r38 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r39 18 26 4.89275 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r40 18 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.69
+ $Y2=0
r41 17 29 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=2.127
+ $Y2=0
r42 17 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.61
+ $Y2=0
r43 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r44 15 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r45 11 29 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.127 $Y2=0
r46 11 13 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0.4
r47 7 26 2.95841 $w=3.4e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.215 $Y2=0
r48 7 9 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r49 2 13 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.04 $Y2=0.4
r50 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends


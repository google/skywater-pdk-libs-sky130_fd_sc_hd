* File: sky130_fd_sc_hd__nand3_4.pex.spice
* Created: Thu Aug 27 14:29:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND3_4%C 3 7 11 15 19 23 25 27 31 33 34 35 36
c90 36 0 1.88146e-19 $X=1.615 $Y=1.19
r91 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r92 42 44 34.1782 $w=2.75e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r93 36 49 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.52 $Y2=1.175
r94 35 49 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.52 $Y2=1.175
r95 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.155 $Y2=1.175
r96 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r97 33 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r98 25 48 36.8073 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.52 $Y2=1.16
r99 25 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r100 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r101 17 48 36.8073 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r102 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r103 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r104 9 17 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r105 9 44 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.47 $Y2=1.16
r106 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r107 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r108 5 44 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r109 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.985
r110 1 44 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r111 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%B 3 7 11 15 19 23 27 31 33 34 35 36 51
c86 51 0 1.88146e-19 $X=3.41 $Y=1.16
r87 49 51 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.2 $Y=1.16 $X2=3.41
+ $Y2=1.16
r88 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.16 $X2=3.2 $Y2=1.16
r89 47 49 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.99 $Y=1.16 $X2=3.2
+ $Y2=1.16
r90 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16 $X2=2.99
+ $Y2=1.16
r91 44 46 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.36 $Y=1.16
+ $X2=2.57 $Y2=1.16
r92 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r93 41 44 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.36 $Y2=1.16
r94 36 50 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.455 $Y=1.175
+ $X2=3.2 $Y2=1.175
r95 35 50 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=3.2 $Y2=1.175
r96 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.995 $Y2=1.175
r97 34 45 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.36 $Y2=1.175
r98 33 45 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=2.36 $Y2=1.175
r99 29 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r100 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r101 25 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r102 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r103 21 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r104 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r105 17 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r106 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r107 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r108 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r109 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r110 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r111 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r112 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r113 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r114 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%A 3 7 11 15 19 23 27 31 33 34 35 36 41 52
r74 50 52 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.4 $Y=1.16 $X2=5.61
+ $Y2=1.16
r75 48 50 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.19 $Y=1.16 $X2=5.4
+ $Y2=1.16
r76 47 48 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16 $X2=5.19
+ $Y2=1.16
r77 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.35 $Y=1.16 $X2=4.77
+ $Y2=1.16
r78 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.11
+ $Y=1.16 $X2=4.11 $Y2=1.16
r79 41 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.275 $Y=1.16
+ $X2=4.35 $Y2=1.16
r80 41 43 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.275 $Y=1.16
+ $X2=4.11 $Y2=1.16
r81 36 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.4 $Y=1.16
+ $X2=5.4 $Y2=1.16
r82 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.855 $Y=1.175
+ $X2=5.315 $Y2=1.175
r83 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.855 $Y2=1.175
r84 34 44 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.11 $Y2=1.175
r85 33 44 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=4.11 $Y2=1.175
r86 29 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.16
r87 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.985
r88 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=1.16
r89 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=0.56
r90 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.16
r91 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.985
r92 17 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=1.16
r93 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=0.56
r94 13 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.16
r95 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.985
r96 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=1.16
r97 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=0.56
r98 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.16
r99 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.295 $X2=4.35
+ $Y2=1.985
r100 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r101 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%VPWR 1 2 3 4 5 6 7 8 25 27 33 37 41 45 50 52
+ 56 59 60 62 63 65 66 67 68 69 81 91 92 98 101
r94 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r95 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 92 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r97 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r98 89 101 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=6 $Y=2.72 $X2=5.867
+ $Y2=2.72
r99 89 91 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6 $Y=2.72 $X2=6.21
+ $Y2=2.72
r100 88 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 88 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r102 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r103 85 98 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=3.88 $Y2=2.72
r104 85 87 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.83 $Y2=2.72
r105 84 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 81 98 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.88 $Y2=2.72
r108 81 83 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r109 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r110 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r111 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 71 95 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r116 71 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 69 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 69 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r119 67 87 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.83 $Y2=2.72
r120 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.98 $Y2=2.72
r121 65 79 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.78 $Y2=2.72
r123 64 83 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.45 $Y2=2.72
r124 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.78 $Y2=2.72
r125 62 76 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r126 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r127 61 79 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r128 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r129 59 73 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r131 58 76 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r132 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r133 54 101 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.867 $Y=2.635
+ $X2=5.867 $Y2=2.72
r134 54 56 27.6151 $w=2.63e-07 $l=6.35e-07 $layer=LI1_cond $X=5.867 $Y=2.635
+ $X2=5.867 $Y2=2
r135 53 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.98 $Y2=2.72
r136 52 101 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.867 $Y2=2.72
r137 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.065 $Y2=2.72
r138 48 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r139 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2
r140 43 98 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.72
r141 43 45 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2
r142 39 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r143 39 41 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r144 35 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r145 35 37 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r146 31 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r147 31 33 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r148 27 30 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r149 25 95 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r150 25 30 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r151 8 56 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2
r152 7 50 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2
r153 6 45 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=4.015
+ $Y=1.485 $X2=4.14 $Y2=2
r154 5 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2
r155 4 41 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r156 3 37 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r157 2 33 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r158 1 30 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r159 1 27 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%Y 1 2 3 4 5 6 7 8 25 27 29 33 35 39 41 45 47
+ 51 53 57 62 64 66 68 71 72 73 74 82
r133 90 93 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.78
+ $X2=5.4 $Y2=0.78
r134 73 74 9.41096 $w=3.98e-07 $l=2.55e-07 $layer=LI1_cond $X=6.24 $Y=1.19
+ $X2=6.24 $Y2=1.445
r135 72 82 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=6.24 $Y=0.78
+ $X2=6.24 $Y2=0.905
r136 72 93 22.9041 $w=3.88e-07 $l=7.25e-07 $layer=LI1_cond $X=6.125 $Y=0.78
+ $X2=5.4 $Y2=0.78
r137 72 73 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.24 $Y=0.92
+ $X2=6.24 $Y2=1.19
r138 72 82 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.24 $Y=0.92
+ $X2=6.24 $Y2=0.905
r139 69 74 17.8211 $w=3.88e-07 $l=5.6e-07 $layer=LI1_cond $X=5.565 $Y=1.555
+ $X2=6.125 $Y2=1.555
r140 69 71 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=1.555
+ $X2=5.4 $Y2=1.555
r141 55 71 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.4 $Y=1.665
+ $X2=5.4 $Y2=1.555
r142 55 57 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.4 $Y=1.665
+ $X2=5.4 $Y2=2.34
r143 54 68 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=1.555
+ $X2=4.56 $Y2=1.555
r144 53 71 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=1.555
+ $X2=5.4 $Y2=1.555
r145 53 54 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=5.235 $Y=1.555
+ $X2=4.725 $Y2=1.555
r146 49 68 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.555
r147 49 51 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=2.34
r148 48 66 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=1.555
+ $X2=3.2 $Y2=1.555
r149 47 68 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.555
+ $X2=4.56 $Y2=1.555
r150 47 48 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=4.395 $Y=1.555
+ $X2=3.365 $Y2=1.555
r151 43 66 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.2 $Y=1.665
+ $X2=3.2 $Y2=1.555
r152 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.2 $Y=1.665
+ $X2=3.2 $Y2=2.34
r153 42 64 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=1.555
+ $X2=2.36 $Y2=1.555
r154 41 66 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.555
+ $X2=3.2 $Y2=1.555
r155 41 42 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=3.035 $Y=1.555
+ $X2=2.525 $Y2=1.555
r156 37 64 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=1.555
r157 37 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=2.34
r158 36 62 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.555
+ $X2=1.52 $Y2=1.555
r159 35 64 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=2.36 $Y2=1.555
r160 35 36 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=1.685 $Y2=1.555
r161 31 62 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.555
r162 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r163 30 60 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.555
+ $X2=0.68 $Y2=1.555
r164 29 62 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=1.52 $Y2=1.555
r165 29 30 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=0.845 $Y2=1.555
r166 25 60 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.555
r167 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r168 8 71 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.66
r169 8 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=2.34
r170 7 68 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.66
r171 7 51 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.34
r172 6 66 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.66
r173 6 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.34
r174 5 64 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.66
r175 5 39 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.34
r176 4 62 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r177 4 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r178 3 60 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r179 3 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r180 2 93 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.74
r181 1 90 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%A_27_47# 1 2 3 4 5 18 20 21 24 32 35 36 39
+ 40 42 43
r85 42 43 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0.78
+ $X2=3.455 $Y2=0.78
r86 40 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.945 $Y=0.82
+ $X2=3.455 $Y2=0.82
r87 38 40 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0.78
+ $X2=2.945 $Y2=0.78
r88 38 39 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0.78
+ $X2=2.615 $Y2=0.78
r89 36 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.105 $Y=0.82
+ $X2=2.615 $Y2=0.82
r90 34 36 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0.78
+ $X2=2.105 $Y2=0.78
r91 34 35 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0.78
+ $X2=1.775 $Y2=0.78
r92 27 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0.82
+ $X2=1.1 $Y2=0.82
r93 27 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.265 $Y=0.82
+ $X2=1.775 $Y2=0.82
r94 22 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.735 $X2=1.1
+ $Y2=0.82
r95 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.735 $X2=1.1
+ $Y2=0.4
r96 20 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=1.1 $Y2=0.82
r97 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=0.425 $Y2=0.82
r98 16 21 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r99 16 18 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.4
r100 5 42 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.74
r101 4 38 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.74
r102 3 34 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.74
r103 2 24 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r104 1 18 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%VGND 1 2 9 13 16 17 19 20 21 34 35
r72 34 35 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r73 32 35 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=6.21
+ $Y2=0
r74 31 34 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=6.21
+ $Y2=0
r75 31 32 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r76 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r77 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r78 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r79 21 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r80 19 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.15
+ $Y2=0
r81 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.52
+ $Y2=0
r82 18 31 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.61
+ $Y2=0
r83 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.52
+ $Y2=0
r84 16 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r85 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r86 15 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.15
+ $Y2=0
r87 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r88 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r89 11 13 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r90 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r91 7 9 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r92 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r93 1 9 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_4%A_445_47# 1 2 3 4 5 26
r32 24 26 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=4.98 $Y=0.37
+ $X2=5.82 $Y2=0.37
r33 22 24 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.37
+ $X2=4.98 $Y2=0.37
r34 20 22 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.2 $Y=0.37 $X2=4.14
+ $Y2=0.37
r35 17 20 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.37 $X2=3.2
+ $Y2=0.37
r36 5 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.4
r37 4 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.4
r38 3 22 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.4
r39 2 20 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.4
r40 1 17 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__a32oi_1.spice
* Created: Thu Aug 27 14:05:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a32oi_1.spice.pex"
.subckt sky130_fd_sc_hd__a32oi_1  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 A_109_47# N_B2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.169 PD=0.88 PS=1.82 NRD=11.076 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75002
+ A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.15275
+ AS=0.07475 PD=1.12 PS=0.88 NRD=2.76 NRS=11.076 M=1 R=4.33333 SA=75000.6
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1003 A_309_47# N_A1_M1003_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.65 AD=0.0715
+ AS=0.15275 PD=0.87 PS=1.12 NRD=10.152 NRS=32.304 M=1 R=4.33333 SA=75001.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1004 A_383_47# N_A2_M1004_g A_309_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.0715 PD=0.98 PS=0.87 NRD=20.304 NRS=10.152 M=1 R=4.33333 SA=75001.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A3_M1009_g A_383_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333 SA=75002 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_B2_M1006_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1001 N_A_27_297#_M1001_d N_B1_M1001_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.215 AS=0.135 PD=1.43 PS=1.27 NRD=30.535 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_27_297#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.215 PD=1.27 PS=1.43 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1005 N_A_27_297#_M1005_d N_A2_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A3_M1002_g N_A_27_297#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0.9653 M=1 R=6.66667 SA=75002
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a32oi_1.spice.SKY130_FD_SC_HD__A32OI_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__clkbuf_2.pxi.spice
* Created: Tue Sep  1 19:00:10 2020
* 
x_PM_SKY130_FD_SC_HD__CLKBUF_2%A N_A_M1001_g N_A_c_39_n N_A_M1002_g A A
+ PM_SKY130_FD_SC_HD__CLKBUF_2%A
x_PM_SKY130_FD_SC_HD__CLKBUF_2%A_27_47# N_A_27_47#_M1001_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_66_n N_A_27_47#_M1003_g N_A_27_47#_c_71_n N_A_27_47#_M1000_g
+ N_A_27_47#_c_67_n N_A_27_47#_M1004_g N_A_27_47#_c_72_n N_A_27_47#_M1005_g
+ N_A_27_47#_c_68_n N_A_27_47#_c_74_n N_A_27_47#_c_83_n N_A_27_47#_c_75_n
+ N_A_27_47#_c_69_n N_A_27_47#_c_70_n N_A_27_47#_c_77_n
+ PM_SKY130_FD_SC_HD__CLKBUF_2%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKBUF_2%VPWR N_VPWR_M1002_d N_VPWR_M1005_s N_VPWR_c_126_n
+ N_VPWR_c_127_n N_VPWR_c_128_n VPWR N_VPWR_c_129_n N_VPWR_c_130_n
+ N_VPWR_c_131_n N_VPWR_c_125_n PM_SKY130_FD_SC_HD__CLKBUF_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKBUF_2%X N_X_M1003_d N_X_M1000_d N_X_c_156_n N_X_c_178_n
+ X X X X X PM_SKY130_FD_SC_HD__CLKBUF_2%X
x_PM_SKY130_FD_SC_HD__CLKBUF_2%VGND N_VGND_M1001_d N_VGND_M1004_s N_VGND_c_191_n
+ N_VGND_c_192_n N_VGND_c_193_n VGND N_VGND_c_194_n N_VGND_c_195_n
+ N_VGND_c_196_n N_VGND_c_197_n PM_SKY130_FD_SC_HD__CLKBUF_2%VGND
cc_1 VNB N_A_M1001_g 0.0270129f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_c_39_n 0.0330091f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.395
cc_3 VNB A 0.00608165f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_4 VNB N_A_27_47#_c_66_n 0.0156271f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_5 VNB N_A_27_47#_c_67_n 0.0174297f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_6 VNB N_A_27_47#_c_68_n 0.0329771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_69_n 0.0624951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_70_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_VPWR_c_125_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_X_c_156_n 3.57995e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_11 VNB X 0.0126029f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.85
cc_12 VNB X 0.0204789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_191_n 0.00468168f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_14 VNB N_VGND_c_192_n 0.0102408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_193_n 0.013519f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_16 VNB N_VGND_c_194_n 0.0168654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_195_n 0.014857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_196_n 0.0052624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_197_n 0.122794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VPB N_A_c_39_n 0.0291972f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.395
cc_21 VPB A 0.00123468f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_22 VPB N_A_27_47#_c_71_n 0.0152786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB N_A_27_47#_c_72_n 0.0177838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_A_27_47#_c_68_n 0.00902172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A_27_47#_c_74_n 0.0297332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_47#_c_75_n 5.27187e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_27_47#_c_69_n 0.0121081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_c_77_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_126_n 0.00217145f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_30 VPB N_VPWR_c_127_n 0.0102423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_128_n 0.0144976f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_32 VPB N_VPWR_c_129_n 0.0154253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_130_n 0.0143966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_131_n 0.00510842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_125_n 0.0428703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB X 0.00737155f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_37 VPB X 0.0215462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 N_A_M1001_g N_A_27_47#_c_66_n 0.0164192f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_39 N_A_c_39_n N_A_27_47#_c_71_n 0.0185097f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_40 N_A_M1001_g N_A_27_47#_c_68_n 0.00979399f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_41 N_A_c_39_n N_A_27_47#_c_68_n 0.0149128f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_42 A N_A_27_47#_c_68_n 0.0438413f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_43 N_A_c_39_n N_A_27_47#_c_83_n 0.01729f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_44 A N_A_27_47#_c_83_n 0.0259259f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_45 N_A_c_39_n N_A_27_47#_c_75_n 0.00119671f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_46 A N_A_27_47#_c_75_n 0.0246972f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_47 N_A_c_39_n N_A_27_47#_c_69_n 0.0322061f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_48 A N_A_27_47#_c_69_n 0.00565351f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_49 N_A_c_39_n N_VPWR_c_126_n 0.0134352f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_50 N_A_c_39_n N_VPWR_c_129_n 0.00486043f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_51 N_A_c_39_n N_VPWR_c_125_n 0.00927066f $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_52 A X 0.00492153f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_53 A X 0.00519615f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_54 N_A_M1001_g N_VGND_c_191_n 0.00317144f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_55 N_A_c_39_n N_VGND_c_191_n 4.71188e-19 $X=0.475 $Y=1.395 $X2=0 $Y2=0
cc_56 A N_VGND_c_191_n 0.0168184f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_M1001_g N_VGND_c_194_n 0.00465542f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_58 A N_VGND_c_194_n 0.00180873f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VGND_c_197_n 0.00771383f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_60 A N_VGND_c_197_n 0.00384383f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A_27_47#_c_83_n N_VPWR_M1002_d 0.00538844f $X=0.965 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_62 N_A_27_47#_c_71_n N_VPWR_c_126_n 0.00166775f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_63 N_A_27_47#_c_83_n N_VPWR_c_126_n 0.0174317f $X=0.965 $Y=1.58 $X2=0 $Y2=0
cc_64 N_A_27_47#_c_71_n N_VPWR_c_128_n 5.99443e-19 $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_65 N_A_27_47#_c_72_n N_VPWR_c_128_n 0.00858985f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_66 N_A_27_47#_c_74_n N_VPWR_c_129_n 0.015543f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_67 N_A_27_47#_c_71_n N_VPWR_c_130_n 0.00585385f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_68 N_A_27_47#_c_72_n N_VPWR_c_130_n 0.00345652f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_69 N_A_27_47#_M1002_s N_VPWR_c_125_n 0.00375137f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_70 N_A_27_47#_c_71_n N_VPWR_c_125_n 0.010776f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_71 N_A_27_47#_c_72_n N_VPWR_c_125_n 0.00409556f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_72 N_A_27_47#_c_74_n N_VPWR_c_125_n 0.0101702f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_73 N_A_27_47#_c_83_n N_X_M1000_d 0.00298074f $X=0.965 $Y=1.58 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_69_n N_X_c_156_n 6.13678e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_66_n X 0.00291318f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_67_n X 0.00702038f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_75_n X 0.013238f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_69_n X 0.0170488f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_72_n X 0.0149933f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_83_n X 0.00992463f $X=0.965 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_69_n X 3.44464e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_71_n X 0.0012162f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_72_n X 0.0165999f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_83_n X 0.0140678f $X=0.965 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_75_n X 0.03713f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_69_n X 0.0244793f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_66_n N_VGND_c_191_n 0.00152531f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_66_n N_VGND_c_193_n 5.45981e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_67_n N_VGND_c_193_n 0.00813915f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_70_n N_VGND_c_194_n 0.017242f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_66_n N_VGND_c_195_n 0.00585385f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_67_n N_VGND_c_195_n 0.00341689f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1001_s N_VGND_c_197_n 0.00400903f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_66_n N_VGND_c_197_n 0.0106812f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_67_n N_VGND_c_197_n 0.0039829f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_70_n N_VGND_c_197_n 0.00981906f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_97 N_VPWR_c_125_n N_X_M1000_d 0.00361236f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_98 N_VPWR_c_130_n N_X_c_178_n 0.009677f $X=1.415 $Y=2.72 $X2=0 $Y2=0
cc_99 N_VPWR_c_125_n N_X_c_178_n 0.00684471f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_100 N_VPWR_M1005_s X 0.00351259f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_101 N_VPWR_c_128_n X 0.0184681f $X=1.58 $Y=2.295 $X2=0 $Y2=0
cc_102 N_VPWR_c_130_n X 0.0021695f $X=1.415 $Y=2.72 $X2=0 $Y2=0
cc_103 N_VPWR_c_125_n X 0.00537675f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_104 N_VPWR_M1005_s X 0.00223862f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_105 X N_VGND_c_193_n 0.0214173f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_106 N_X_c_156_n N_VGND_c_195_n 0.0122263f $X=1.16 $Y=0.42 $X2=0 $Y2=0
cc_107 X N_VGND_c_195_n 0.00275256f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_108 N_X_M1003_d N_VGND_c_197_n 0.0028269f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_109 N_X_c_156_n N_VGND_c_197_n 0.00771386f $X=1.16 $Y=0.42 $X2=0 $Y2=0
cc_110 X N_VGND_c_197_n 0.00550683f $X=1.525 $Y=0.765 $X2=0 $Y2=0

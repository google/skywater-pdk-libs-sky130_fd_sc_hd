* File: sky130_fd_sc_hd__nor3b_2.spice.pex
* Created: Thu Aug 27 14:32:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR3B_2%A 1 3 6 8 10 13 15 16 24
r40 22 24 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.645 $Y=1.16
+ $X2=0.91 $Y2=1.16
r41 19 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.645 $Y2=1.16
r42 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r43 15 16 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.645 $Y2=1.18
r44 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r45 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r46 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r47 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r48 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r50 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%B 1 3 6 8 10 13 15 16 17 26
r45 24 26 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.525 $Y=1.16
+ $X2=1.75 $Y2=1.16
r46 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.16 $X2=1.525 $Y2=1.16
r47 21 24 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.525 $Y2=1.16
r48 16 17 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=2.075 $Y=1.18
+ $X2=2.555 $Y2=1.18
r49 15 16 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=2.075 $Y2=1.18
r50 15 25 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=1.525 $Y2=1.18
r51 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r52 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r53 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r54 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r55 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r56 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325 $X2=1.33
+ $Y2=1.985
r57 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995 $X2=1.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%A_531_21# 1 2 7 9 12 14 16 19 21 24 27 31 34
+ 36 37
r62 39 41 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=3.15 $Y2=1.16
r63 36 37 11.2584 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=3.867 $Y=1.705
+ $X2=3.867 $Y2=1.455
r64 31 33 11.0961 $w=3.53e-07 $l=2.45e-07 $layer=LI1_cond $X=3.867 $Y=0.66
+ $X2=3.867 $Y2=0.905
r65 28 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.775 $Y=1.285
+ $X2=3.775 $Y2=1.18
r66 28 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.775 $Y=1.285
+ $X2=3.775 $Y2=1.455
r67 27 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.775 $Y=1.075
+ $X2=3.775 $Y2=1.18
r68 27 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.775 $Y=1.075
+ $X2=3.775 $Y2=0.905
r69 24 41 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.4 $Y=1.16 $X2=3.15
+ $Y2=1.16
r70 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.16 $X2=3.4 $Y2=1.16
r71 21 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=1.18
+ $X2=3.775 $Y2=1.18
r72 21 23 15.316 $w=2.08e-07 $l=2.9e-07 $layer=LI1_cond $X=3.69 $Y=1.18 $X2=3.4
+ $Y2=1.18
r73 17 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.16
r74 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.985
r75 14 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=1.16
r76 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=0.56
r77 10 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.16
r78 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.985
r79 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=0.995
+ $X2=2.73 $Y2=1.16
r80 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.995 $X2=2.73
+ $Y2=0.56
r81 2 36 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.485 $X2=3.92 $Y2=1.705
r82 1 31 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.465 $X2=3.92 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%C_N 3 6 8 11 13
r27 11 14 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.192 $Y=1.16
+ $X2=4.192 $Y2=1.325
r28 11 13 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.192 $Y=1.16
+ $X2=4.192 $Y2=0.995
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=1.16 $X2=4.195 $Y2=1.16
r30 8 12 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=4.37 $Y=1.18
+ $X2=4.195 $Y2=1.18
r31 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.13 $Y=1.695
+ $X2=4.13 $Y2=1.325
r32 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.13 $Y=0.675
+ $X2=4.13 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%A_27_297# 1 2 3 10 12 14 18 20 27 29
r35 21 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.54
+ $X2=1.12 $Y2=1.54
r36 20 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.96 $Y2=1.54
r37 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.245 $Y2=1.54
r38 16 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=1.54
r39 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=2.3
r40 15 25 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.247 $Y2=1.54
r41 14 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=1.12 $Y2=1.54
r42 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=0.405 $Y2=1.54
r43 10 25 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=1.54
r44 10 12 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.247 $Y=1.625
+ $X2=0.247 $Y2=2.3
r45 3 29 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r46 2 27 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r47 2 18 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r48 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r49 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%VPWR 1 2 9 11 13 15 17 22 31 35
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r52 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r54 28 29 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r55 26 29 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 25 28 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 25 26 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 23 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r60 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 22 34 3.98688 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.215 $Y=2.72
+ $X2=4.407 $Y2=2.72
r62 22 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.215 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 17 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r64 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 11 34 3.15628 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=4.34 $Y=2.635
+ $X2=4.407 $Y2=2.72
r68 11 13 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=4.34 $Y=2.635
+ $X2=4.34 $Y2=1.705
r69 7 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r70 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r71 2 13 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=1.705
r72 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%A_281_297# 1 2 3 12 14 15 18 20 22 24 27
c37 18 0 1.49843e-19 $X=2.52 $Y=1.62
r38 22 29 2.91961 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.357 $Y=2.295
+ $X2=3.357 $Y2=2.38
r39 22 24 31.751 $w=2.43e-07 $l=6.75e-07 $layer=LI1_cond $X=3.357 $Y=2.295
+ $X2=3.357 $Y2=1.62
r40 21 27 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.645 $Y=2.38
+ $X2=2.51 $Y2=2.38
r41 20 29 4.1905 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=3.235 $Y=2.38
+ $X2=3.357 $Y2=2.38
r42 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.235 $Y=2.38
+ $X2=2.645 $Y2=2.38
r43 16 27 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.295
+ $X2=2.51 $Y2=2.38
r44 16 18 28.8111 $w=2.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.51 $Y=2.295
+ $X2=2.51 $Y2=1.62
r45 14 27 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=2.51 $Y2=2.38
r46 14 15 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=1.665 $Y2=2.38
r47 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.665 $Y2=2.38
r48 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.54 $Y2=1.96
r49 3 29 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=2.3
r50 3 24 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=1.62
r51 2 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.485 $X2=2.52 $Y2=2.3
r52 2 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.485 $X2=2.52 $Y2=1.62
r53 1 12 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%Y 1 2 3 4 15 17 18 21 23 27 29 31 32 35
c71 23 0 1.49843e-19 $X=2.775 $Y=0.815
r72 32 35 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.94 $Y=0.51 $X2=2.94
+ $Y2=0.39
r73 30 32 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.94 $Y=0.725
+ $X2=2.94 $Y2=0.51
r74 30 31 3.41797 $w=2.9e-07 $l=9e-08 $layer=LI1_cond $X=2.94 $Y=0.725 $X2=2.94
+ $Y2=0.815
r75 25 31 3.41797 $w=2.9e-07 $l=9e-08 $layer=LI1_cond $X=2.94 $Y=0.905 $X2=2.94
+ $Y2=0.815
r76 25 27 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=2.94 $Y=0.905
+ $X2=2.94 $Y2=1.62
r77 24 29 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r78 23 31 3.10432 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=2.94 $Y2=0.815
r79 23 24 65.9293 $w=1.78e-07 $l=1.07e-06 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=1.705 $Y2=0.815
r80 19 29 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725 $X2=1.54
+ $Y2=0.815
r81 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r82 17 29 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r83 17 18 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r84 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r85 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725 $X2=0.7
+ $Y2=0.39
r86 4 27 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=1.62
r87 3 35 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.235 $X2=2.94 $Y2=0.39
r88 2 21 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r89 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_2%VGND 1 2 3 4 5 6 19 21 25 29 31 33 36 37 39
+ 40 41 55 64 70 73
r68 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r69 69 70 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0.235
+ $X2=2.605 $Y2=0.235
r70 66 69 8.40993 $w=6.38e-07 $l=4.5e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.52 $Y2=0.235
r71 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r72 63 66 2.05576 $w=6.38e-07 $l=1.1e-07 $layer=LI1_cond $X=1.96 $Y=0.235
+ $X2=2.07 $Y2=0.235
r73 63 64 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.235
+ $X2=1.875 $Y2=0.235
r74 58 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r75 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r76 55 72 4.40761 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.407
+ $Y2=0
r77 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=3.91
+ $Y2=0
r78 54 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r79 54 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r80 53 70 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.605
+ $Y2=0
r81 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r82 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r83 49 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.875
+ $Y2=0
r84 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r85 46 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r86 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r87 43 60 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r88 43 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r89 41 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r90 41 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r91 39 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=2.99
+ $Y2=0
r92 39 40 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.377
+ $Y2=0
r93 38 57 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=3.91
+ $Y2=0
r94 38 40 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=3.377
+ $Y2=0
r95 36 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r96 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r97 35 49 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.61
+ $Y2=0
r98 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r99 31 72 3.03023 $w=2.9e-07 $l=1.05924e-07 $layer=LI1_cond $X=4.36 $Y=0.085
+ $X2=4.407 $Y2=0
r100 31 33 22.8502 $w=2.88e-07 $l=5.75e-07 $layer=LI1_cond $X=4.36 $Y=0.085
+ $X2=4.36 $Y2=0.66
r101 27 40 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.377 $Y=0.085
+ $X2=3.377 $Y2=0
r102 27 29 16.5011 $w=2.03e-07 $l=3.05e-07 $layer=LI1_cond $X=3.377 $Y=0.085
+ $X2=3.377 $Y2=0.39
r103 23 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r104 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r105 19 60 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r106 19 21 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r107 6 33 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.465 $X2=4.34 $Y2=0.66
r108 5 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.225
+ $Y=0.235 $X2=3.36 $Y2=0.39
r109 4 69 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.52 $Y2=0.39
r110 3 63 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r111 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r112 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__nand4b_1.spice.pex
* Created: Thu Aug 27 14:30:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4B_1%A_N 3 6 8 11 13
r31 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r34 8 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.51
+ $Y2=1.16
r35 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.6 $Y=1.695 $X2=0.6
+ $Y2=1.325
r36 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.545 $Y=0.675
+ $X2=0.545 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%D 3 6 8 11 13
c35 13 0 1.60027e-19 $X=1.05 $Y=0.995
r36 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=1.05 $Y2=1.325
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=1.05 $Y2=0.995
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r39 8 12 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.05
+ $Y2=1.16
r40 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.085 $Y=1.985
+ $X2=1.085 $Y2=1.325
r41 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.085 $Y=0.56
+ $X2=1.085 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%C 3 6 8 9 13 15
r38 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.16
+ $X2=1.59 $Y2=1.325
r39 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.16
+ $X2=1.59 $Y2=0.995
r40 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.59
+ $Y=1.16 $X2=1.59 $Y2=1.16
r41 8 9 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=1.63 $Y=0.85 $X2=1.63
+ $Y2=1.16
r42 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.505 $Y=1.985
+ $X2=1.505 $Y2=1.325
r43 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.505 $Y=0.56
+ $X2=1.505 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%B 3 6 8 9 13 15
r39 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=1.16 $X2=2.1
+ $Y2=1.325
r40 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=1.16 $X2=2.1
+ $Y2=0.995
r41 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.1 $Y=1.16
+ $X2=2.1 $Y2=1.16
r42 8 9 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.055 $Y=0.85
+ $X2=2.055 $Y2=1.16
r43 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.04 $Y=1.985
+ $X2=2.04 $Y2=1.325
r44 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.04 $Y=0.56 $X2=2.04
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%A_41_93# 1 2 9 12 15 16 18 21 26 30 32 39
+ 40 43
c84 18 0 1.60027e-19 $X=2.355 $Y=0.51
r85 40 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.67 $Y2=1.325
r86 40 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.67 $Y2=0.995
r87 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.16 $X2=2.67 $Y2=1.16
r88 36 39 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.44 $Y=1.16
+ $X2=2.67 $Y2=1.16
r89 32 34 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=1.245 $Y=0.51
+ $X2=1.245 $Y2=0.74
r90 27 30 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.17 $Y=1.76
+ $X2=0.39 $Y2=1.76
r91 25 26 7.96465 $w=3.78e-07 $l=1.45e-07 $layer=LI1_cond $X=0.33 $Y=0.635
+ $X2=0.475 $Y2=0.635
r92 22 25 4.85239 $w=3.78e-07 $l=1.6e-07 $layer=LI1_cond $X=0.17 $Y=0.635
+ $X2=0.33 $Y2=0.635
r93 21 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=0.995
+ $X2=2.44 $Y2=1.16
r94 20 21 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.44 $Y=0.595 $X2=2.44
+ $Y2=0.995
r95 19 32 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.335 $Y=0.51 $X2=1.245
+ $Y2=0.51
r96 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.355 $Y=0.51
+ $X2=2.44 $Y2=0.595
r97 18 19 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.355 $Y=0.51
+ $X2=1.335 $Y2=0.51
r98 16 34 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=0.74 $X2=1.245
+ $Y2=0.74
r99 16 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=0.74
+ $X2=0.475 $Y2=0.74
r100 15 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.595
+ $X2=0.17 $Y2=1.76
r101 14 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.635
r102 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.595
r103 12 44 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.58 $Y=1.985
+ $X2=2.58 $Y2=1.325
r104 9 43 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.58 $Y=0.56
+ $X2=2.58 $Y2=0.995
r105 2 30 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.485 $X2=0.39 $Y2=1.76
r106 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.465 $X2=0.33 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%VPWR 1 2 3 12 18 22 25 26 28 29 31 32 33 46
+ 47
c42 3 0 1.15679e-19 $X=2.655 $Y=1.485
r43 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 44 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 37 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 33 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 31 43 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.53 $Y2=2.72
r52 31 32 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.812 $Y2=2.72
r53 30 46 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.92 $Y=2.72 $X2=2.99
+ $Y2=2.72
r54 30 32 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.92 $Y=2.72
+ $X2=2.812 $Y2=2.72
r55 28 40 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.63 $Y=2.72 $X2=1.61
+ $Y2=2.72
r56 28 29 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.63 $Y=2.72
+ $X2=1.772 $Y2=2.72
r57 27 43 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 27 29 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.772 $Y2=2.72
r59 25 36 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.71 $Y=2.72 $X2=0.69
+ $Y2=2.72
r60 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.71 $Y=2.72
+ $X2=0.835 $Y2=2.72
r61 24 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=0.835 $Y2=2.72
r63 20 32 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.812 $Y=2.635
+ $X2=2.812 $Y2=2.72
r64 20 22 34.0373 $w=2.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.812 $Y=2.635
+ $X2=2.812 $Y2=2
r65 16 29 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.772 $Y=2.635
+ $X2=1.772 $Y2=2.72
r66 16 18 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=1.772 $Y=2.635
+ $X2=1.772 $Y2=2
r67 12 15 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.835 $Y=1.66
+ $X2=0.835 $Y2=2
r68 10 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=2.635
+ $X2=0.835 $Y2=2.72
r69 10 15 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.835 $Y=2.635
+ $X2=0.835 $Y2=2
r70 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.655
+ $Y=1.485 $X2=2.79 $Y2=2
r71 2 18 300 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.485 $X2=1.775 $Y2=2
r72 1 15 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=0.675
+ $Y=1.485 $X2=0.875 $Y2=2
r73 1 12 600 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.485 $X2=0.875 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%Y 1 2 3 10 12 14 18 20 23 27 28 31
c46 23 0 1.15679e-19 $X=3.03 $Y=1.495
r47 28 35 11.4137 $w=4.38e-07 $l=3.15e-07 $layer=LI1_cond $X=2.915 $Y=0.51
+ $X2=2.915 $Y2=0.825
r48 28 31 3.40495 $w=4.38e-07 $l=1.3e-07 $layer=LI1_cond $X=2.915 $Y=0.51
+ $X2=2.915 $Y2=0.38
r49 23 35 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=3.03 $Y=1.495
+ $X2=3.03 $Y2=0.825
r50 21 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=1.58
+ $X2=2.25 $Y2=1.58
r51 20 23 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=3.03 $Y2=1.495
r52 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=2.415 $Y2=1.58
r53 16 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=1.665
+ $X2=2.25 $Y2=1.58
r54 16 18 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.25 $Y=1.665
+ $X2=2.25 $Y2=2.335
r55 15 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=1.58
+ $X2=1.295 $Y2=1.58
r56 14 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=1.58
+ $X2=2.25 $Y2=1.58
r57 14 15 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.085 $Y=1.58
+ $X2=1.46 $Y2=1.58
r58 10 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=1.665
+ $X2=1.295 $Y2=1.58
r59 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.295 $Y=1.665
+ $X2=1.295 $Y2=2.34
r60 3 27 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.485 $X2=2.25 $Y2=1.655
r61 3 18 400 $w=1.7e-07 $l=9.15014e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.485 $X2=2.25 $Y2=2.335
r62 2 25 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.485 $X2=1.295 $Y2=1.66
r63 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.485 $X2=1.295 $Y2=2.34
r64 1 31 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=2.655
+ $Y=0.235 $X2=2.86 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_1%VGND 1 8 10 17 18 21
r34 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r35 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r36 15 18 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r37 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r38 14 17 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r39 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r40 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.82
+ $Y2=0
r41 12 14 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r42 10 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=0.085 $X2=0.82
+ $Y2=0
r44 6 8 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0.38
r45 1 8 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.465 $X2=0.82 $Y2=0.38
.ends


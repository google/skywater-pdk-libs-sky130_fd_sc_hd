* File: sky130_fd_sc_hd__and4_4.spice
* Created: Thu Aug 27 14:08:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4_4.spice.pex"
.subckt sky130_fd_sc_hd__and4_4  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1014 A_109_47# N_A_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.079625 AS=0.169 PD=0.895 PS=1.82 NRD=12.456 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1007 A_188_47# N_B_M1007_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.108875
+ AS=0.079625 PD=0.985 PS=0.895 NRD=20.76 NRS=12.456 M=1 R=4.33333 SA=75000.6
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1002 A_285_47# N_C_M1002_g A_188_47# VNB NSHORT L=0.15 W=0.65 AD=0.141375
+ AS=0.108875 PD=1.085 PS=0.985 NRD=30 NRS=20.76 M=1 R=4.33333 SA=75001.1
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_D_M1009_g A_285_47# VNB NSHORT L=0.15 W=0.65 AD=0.105625
+ AS=0.141375 PD=0.975 PS=1.085 NRD=7.38 NRS=30 M=1 R=4.33333 SA=75001.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.105625 PD=0.92 PS=0.975 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75002.1 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1001_d N_A_27_47#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1010_d N_A_27_47#_M1010_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1010_d N_A_27_47#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_27_47#_M1012_d N_A_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_27_47#_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.135 PD=1.31 PS=1.27 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_47#_M1008_d N_C_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.215 AS=0.155 PD=1.43 PS=1.31 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75001.1
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_D_M1013_g N_A_27_47#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.215 PD=1.33 PS=1.43 NRD=8.8453 NRS=30.535 M=1 R=6.66667
+ SA=75001.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1013_d N_A_27_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75002.1
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_47#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1003_d N_A_27_47#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_27_47#_M1011_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__and4_4.spice.SKY130_FD_SC_HD__AND4_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a311o_4.spice
* Created: Thu Aug 27 14:04:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a311o_4.spice.pex"
.subckt sky130_fd_sc_hd__a311o_4  VNB VPB C1 B1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_C1_M1013_g N_A_109_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1027_d N_C1_M1027_g N_A_109_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1027_d N_B1_M1018_g N_A_109_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_B1_M1019_g N_A_109_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1019_d N_A_109_47#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.09425 PD=0.92 PS=0.94 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75001.9
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_109_47#_M1011_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.09425 PD=0.92 PS=0.94 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1011_d N_A_109_47#_M1015_g N_X_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_A_109_47#_M1025_g N_X_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.21125 AS=0.08775 PD=1.3 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 N_A_861_47#_M1002_d N_A3_M1002_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.21125 PD=0.92 PS=1.3 NRD=0 NRS=6.456 M=1 R=4.33333 SA=75003.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_861_47#_M1002_d N_A3_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_1059_47#_M1000_d N_A2_M1000_g N_A_861_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1003 N_A_1059_47#_M1003_d N_A2_M1003_g N_A_861_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1004 N_A_1059_47#_M1003_d N_A1_M1004_g N_A_109_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_A_1059_47#_M1006_d N_A1_M1006_g N_A_109_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_297#_M1005_d N_C1_M1005_g N_A_109_47#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1020 N_A_27_297#_M1020_d N_C1_M1020_g N_A_109_47#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1001 N_A_277_297#_M1001_d N_B1_M1001_g N_A_27_297#_M1020_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1026 N_A_277_297#_M1001_d N_B1_M1026_g N_A_27_297#_M1026_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_109_47#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_A_109_47#_M1016_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1016_d N_A_109_47#_M1017_g N_X_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_A_109_47#_M1024_g N_X_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1024_d N_A3_M1008_g N_A_277_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A3_M1012_g N_A_277_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1012_d N_A2_M1021_g N_A_277_297#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_A2_M1023_g N_A_277_297#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.325 AS=0.135 PD=1.65 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1023_d N_A1_M1014_g N_A_277_297#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.325 AS=0.135 PD=1.65 PS=1.27 NRD=73.8553 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_A1_M1022_g N_A_277_297#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=12.4227 P=18.69
*
.include "sky130_fd_sc_hd__a311o_4.spice.SKY130_FD_SC_HD__A311O_4.pxi"
*
.ends
*
*

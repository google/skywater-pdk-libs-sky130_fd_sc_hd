* File: sky130_fd_sc_hd__a31o_1.pxi.spice
* Created: Tue Sep  1 18:55:01 2020
* 
x_PM_SKY130_FD_SC_HD__A31O_1%A_80_21# N_A_80_21#_M1006_d N_A_80_21#_M1009_d
+ N_A_80_21#_M1002_g N_A_80_21#_M1005_g N_A_80_21#_c_60_n N_A_80_21#_c_73_p
+ N_A_80_21#_c_120_p N_A_80_21#_c_85_p N_A_80_21#_c_61_n N_A_80_21#_c_62_n
+ N_A_80_21#_c_63_n N_A_80_21#_c_86_p N_A_80_21#_c_69_n N_A_80_21#_c_64_n
+ N_A_80_21#_c_65_n PM_SKY130_FD_SC_HD__A31O_1%A_80_21#
x_PM_SKY130_FD_SC_HD__A31O_1%A3 N_A3_M1004_g N_A3_M1008_g A3 A3 N_A3_c_141_n
+ N_A3_c_142_n N_A3_c_143_n PM_SKY130_FD_SC_HD__A31O_1%A3
x_PM_SKY130_FD_SC_HD__A31O_1%A2 N_A2_M1001_g N_A2_M1003_g A2 A2 N_A2_c_178_n
+ N_A2_c_179_n N_A2_c_180_n PM_SKY130_FD_SC_HD__A31O_1%A2
x_PM_SKY130_FD_SC_HD__A31O_1%A1 N_A1_M1006_g N_A1_M1000_g A1 A1 N_A1_c_213_n
+ N_A1_c_214_n N_A1_c_215_n PM_SKY130_FD_SC_HD__A31O_1%A1
x_PM_SKY130_FD_SC_HD__A31O_1%B1 N_B1_M1007_g N_B1_M1009_g B1 B1 N_B1_c_250_n
+ N_B1_c_251_n PM_SKY130_FD_SC_HD__A31O_1%B1
x_PM_SKY130_FD_SC_HD__A31O_1%X N_X_M1002_s N_X_M1005_s N_X_c_277_n N_X_c_280_n
+ N_X_c_278_n X X X N_X_c_279_n PM_SKY130_FD_SC_HD__A31O_1%X
x_PM_SKY130_FD_SC_HD__A31O_1%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_298_n
+ N_VPWR_c_299_n VPWR N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n
+ N_VPWR_c_297_n N_VPWR_c_304_n N_VPWR_c_305_n PM_SKY130_FD_SC_HD__A31O_1%VPWR
x_PM_SKY130_FD_SC_HD__A31O_1%A_209_297# N_A_209_297#_M1008_d
+ N_A_209_297#_M1000_d N_A_209_297#_c_344_n N_A_209_297#_c_347_n
+ N_A_209_297#_c_348_n N_A_209_297#_c_355_n N_A_209_297#_c_366_n
+ PM_SKY130_FD_SC_HD__A31O_1%A_209_297#
x_PM_SKY130_FD_SC_HD__A31O_1%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_c_369_n
+ N_VGND_c_370_n VGND N_VGND_c_371_n N_VGND_c_372_n N_VGND_c_373_n
+ N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n PM_SKY130_FD_SC_HD__A31O_1%VGND
cc_1 VNB N_A_80_21#_c_60_n 0.00205417f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_2 VNB N_A_80_21#_c_61_n 0.0101465f $X=-0.19 $Y=-0.24 $X2=2.79 $Y2=0.74
cc_3 VNB N_A_80_21#_c_62_n 0.0239534f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_4 VNB N_A_80_21#_c_63_n 0.00208902f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_5 VNB N_A_80_21#_c_64_n 0.0224965f $X=-0.19 $Y=-0.24 $X2=2.732 $Y2=1.825
cc_6 VNB N_A_80_21#_c_65_n 0.0200709f $X=-0.19 $Y=-0.24 $X2=0.537 $Y2=0.995
cc_7 VNB N_A3_c_141_n 0.0205104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A3_c_142_n 0.00368411f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.825
cc_9 VNB N_A3_c_143_n 0.0173008f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_10 VNB N_A2_c_178_n 0.0205555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_179_n 0.00366597f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.825
cc_12 VNB N_A2_c_180_n 0.0174901f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_13 VNB N_A1_c_213_n 0.0205753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_214_n 0.00355186f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.825
cc_15 VNB N_A1_c_215_n 0.0175802f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_16 VNB B1 0.00420804f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_17 VNB N_B1_c_250_n 0.0262606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_c_251_n 0.0202857f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_19 VNB N_X_c_277_n 0.00638732f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_20 VNB N_X_c_278_n 0.0227807f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.825
cc_21 VNB N_X_c_279_n 0.013624f $X=-0.19 $Y=-0.24 $X2=2.79 $Y2=0.74
cc_22 VNB N_VPWR_c_297_n 0.136896f $X=-0.19 $Y=-0.24 $X2=2.14 $Y2=0.74
cc_23 VNB N_VGND_c_369_n 0.00277135f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_24 VNB N_VGND_c_370_n 0.0149911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_371_n 0.0182515f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=0.74
cc_26 VNB N_VGND_c_372_n 0.0402435f $X=-0.19 $Y=-0.24 $X2=2.79 $Y2=0.74
cc_27 VNB N_VGND_c_373_n 0.0146906f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_28 VNB N_VGND_c_374_n 0.189151f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_29 VNB N_VGND_c_375_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_376_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=2.732 $Y2=1.91
cc_31 VPB N_A_80_21#_M1005_g 0.0230726f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_32 VPB N_A_80_21#_c_62_n 0.00549446f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_33 VPB N_A_80_21#_c_63_n 9.47497e-19 $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_34 VPB N_A_80_21#_c_69_n 0.0263626f $X=-0.19 $Y=1.305 $X2=2.67 $Y2=1.91
cc_35 VPB N_A_80_21#_c_64_n 0.0221634f $X=-0.19 $Y=1.305 $X2=2.732 $Y2=1.825
cc_36 VPB N_A3_M1008_g 0.0195924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A3 9.49913e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_38 VPB N_A3_c_141_n 0.00474451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A2_M1003_g 0.0193569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A2_c_178_n 0.00452009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A2_c_179_n 0.00112587f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.825
cc_42 VPB N_A1_M1000_g 0.0194612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A1_c_213_n 0.00453676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A1_c_214_n 0.00117037f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.825
cc_45 VPB N_B1_M1009_g 0.0239379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB B1 0.00166406f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_47 VPB N_B1_c_250_n 0.0049054f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_X_c_280_n 0.00638732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_X_c_278_n 0.0124167f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.825
cc_50 VPB X 0.0267831f $X=-0.19 $Y=1.305 $X2=1.975 $Y2=0.74
cc_51 VPB N_VPWR_c_298_n 0.00460743f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_52 VPB N_VPWR_c_299_n 0.00508424f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.995
cc_53 VPB N_VPWR_c_300_n 0.0182237f $X=-0.19 $Y=1.305 $X2=2.14 $Y2=0.4
cc_54 VPB N_VPWR_c_301_n 0.0182782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_302_n 0.039579f $X=-0.19 $Y=1.305 $X2=2.14 $Y2=0.74
cc_56 VPB N_VPWR_c_297_n 0.052692f $X=-0.19 $Y=1.305 $X2=2.14 $Y2=0.74
cc_57 VPB N_VPWR_c_304_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.732 $Y2=1.825
cc_58 VPB N_VPWR_c_305_n 0.00631953f $X=-0.19 $Y=1.305 $X2=0.537 $Y2=0.995
cc_59 N_A_80_21#_M1005_g N_A3_M1008_g 0.010387f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_60 N_A_80_21#_M1005_g A3 8.1503e-19 $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_73_p N_A3_c_141_n 6.51071e-19 $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_62_n N_A3_c_141_n 0.0201932f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_63_n N_A3_c_141_n 0.00198104f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_73_p N_A3_c_142_n 0.02142f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_62_n N_A3_c_142_n 3.16507e-19 $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_63_n N_A3_c_142_n 0.0258073f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_60_n N_A3_c_143_n 0.00379389f $X=0.68 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_73_p N_A3_c_143_n 0.0130549f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_65_n N_A3_c_143_n 0.0220662f $X=0.537 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_73_p N_A2_c_178_n 7.21566e-19 $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_73_p N_A2_c_179_n 0.0201593f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_73_p N_A2_c_180_n 0.0139217f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_85_p N_A2_c_180_n 0.00160503f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_86_p N_A1_c_213_n 7.62589e-19 $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_73_p N_A1_c_214_n 0.00596871f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_86_p N_A1_c_214_n 0.0133444f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_73_p N_A1_c_215_n 0.0106251f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_85_p N_A1_c_215_n 0.00651874f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_86_p N_A1_c_215_n 5.61078e-19 $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_64_n N_B1_M1009_g 0.0050266f $X=2.732 $Y=1.825 $X2=0 $Y2=0
cc_81 N_A_80_21#_M1009_d B1 0.00279395f $X=2.475 $Y=1.485 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_61_n B1 0.0168425f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_69_n B1 0.00775461f $X=2.67 $Y=1.91 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_64_n B1 0.0506399f $X=2.732 $Y=1.825 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_61_n N_B1_c_250_n 7.21566e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_69_n N_B1_c_250_n 3.02704e-19 $X=2.67 $Y=1.91 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_64_n N_B1_c_250_n 0.00217704f $X=2.732 $Y=1.825 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_61_n N_B1_c_251_n 0.0131761f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_64_n N_B1_c_251_n 0.00495664f $X=2.732 $Y=1.825 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_65_n N_X_c_277_n 0.00291861f $X=0.537 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_80_21#_M1005_g N_X_c_280_n 0.00287883f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_60_n N_X_c_278_n 0.00606252f $X=0.68 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_63_n N_X_c_278_n 0.0248653f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_65_n N_X_c_278_n 0.0163624f $X=0.537 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_80_21#_M1005_g X 0.00722251f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_65_n N_X_c_279_n 0.00518935f $X=0.537 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_80_21#_M1005_g N_VPWR_c_298_n 0.00293462f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_98 N_A_80_21#_c_73_p N_VPWR_c_298_n 0.00209429f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_62_n N_VPWR_c_298_n 0.00180684f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_63_n N_VPWR_c_298_n 0.0138324f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_80_21#_M1005_g N_VPWR_c_300_n 0.00550269f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_102 N_A_80_21#_c_69_n N_VPWR_c_302_n 0.0196627f $X=2.67 $Y=1.91 $X2=0 $Y2=0
cc_103 N_A_80_21#_M1009_d N_VPWR_c_297_n 0.00365159f $X=2.475 $Y=1.485 $X2=0
+ $Y2=0
cc_104 N_A_80_21#_M1005_g N_VPWR_c_297_n 0.0108358f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_105 N_A_80_21#_c_69_n N_VPWR_c_297_n 0.0158336f $X=2.67 $Y=1.91 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_60_n N_VGND_M1002_d 6.67963e-19 $X=0.68 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_80_21#_c_73_p N_VGND_M1002_d 0.00225732f $X=1.975 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_80_21#_c_120_p N_VGND_M1002_d 0.00260473f $X=0.765 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_80_21#_c_61_n N_VGND_M1007_d 0.0111922f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_64_n N_VGND_M1007_d 7.68922e-19 $X=2.732 $Y=1.825 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_c_73_p N_VGND_c_369_n 0.00761378f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_120_p N_VGND_c_369_n 0.0127713f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_62_n N_VGND_c_369_n 2.81605e-19 $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_65_n N_VGND_c_369_n 0.00430087f $X=0.537 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_c_61_n N_VGND_c_370_n 0.0209899f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_65_n N_VGND_c_371_n 0.0055043f $X=0.537 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_73_p N_VGND_c_372_n 0.0154232f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_85_p N_VGND_c_372_n 0.0140581f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_61_n N_VGND_c_372_n 0.00251419f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_61_n N_VGND_c_373_n 0.00301183f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_80_21#_M1006_d N_VGND_c_374_n 0.00275175f $X=1.995 $Y=0.235 $X2=0
+ $Y2=0
cc_122 N_A_80_21#_c_73_p N_VGND_c_374_n 0.02799f $X=1.975 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_120_p N_VGND_c_374_n 7.70209e-19 $X=0.765 $Y=0.74 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_85_p N_VGND_c_374_n 0.0119805f $X=2.14 $Y=0.4 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_61_n N_VGND_c_374_n 0.00999022f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_65_n N_VGND_c_374_n 0.0109196f $X=0.537 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_73_p A_209_47# 0.00764369f $X=1.975 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_128 N_A_80_21#_c_73_p A_303_47# 0.00845612f $X=1.975 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A3_M1008_g N_A2_M1003_g 0.0205759f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_130 A3 N_A2_M1003_g 0.00210073f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_131 N_A3_c_141_n N_A2_c_178_n 0.0201884f $X=1.02 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A3_c_142_n N_A2_c_178_n 0.00210073f $X=1.02 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A3_M1008_g N_A2_c_179_n 2.91261e-19 $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A3_c_141_n N_A2_c_179_n 3.23502e-19 $X=1.02 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A3_c_142_n N_A2_c_179_n 0.0492492f $X=1.02 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A3_c_143_n N_A2_c_180_n 0.0366407f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A3_c_143_n N_X_c_279_n 5.4882e-19 $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A3_M1008_g N_VPWR_c_298_n 0.00162346f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A3_M1008_g N_VPWR_c_301_n 0.00572337f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A3_M1008_g N_VPWR_c_297_n 0.010633f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_141 A3 N_A_209_297#_M1008_d 0.00302948f $X=1.07 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_142 N_A3_M1008_g N_A_209_297#_c_344_n 0.00176304f $X=0.97 $Y=1.985 $X2=0
+ $Y2=0
cc_143 A3 N_A_209_297#_c_344_n 0.0129912f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_144 N_A3_c_141_n N_A_209_297#_c_344_n 3.34527e-19 $X=1.02 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A3_M1008_g N_A_209_297#_c_347_n 0.00412949f $X=0.97 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A3_c_143_n N_VGND_c_369_n 0.0101254f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A3_c_143_n N_VGND_c_372_n 0.00341689f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A3_c_143_n N_VGND_c_374_n 0.00417721f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_M1003_g N_A1_M1000_g 0.0329813f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A2_c_178_n N_A1_c_213_n 0.0202395f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_c_179_n N_A1_c_213_n 0.00429923f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A2_M1003_g N_A1_c_214_n 2.99415e-19 $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A2_c_178_n N_A1_c_214_n 3.39451e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_c_179_n N_A1_c_214_n 0.045554f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_180_n N_A1_c_215_n 0.035658f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_c_179_n N_VPWR_M1003_d 0.00295022f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_M1003_g N_VPWR_c_299_n 0.00208463f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A2_M1003_g N_VPWR_c_301_n 0.00437059f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A2_M1003_g N_VPWR_c_297_n 0.00617519f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A2_M1003_g N_A_209_297#_c_348_n 0.0119341f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A2_c_178_n N_A_209_297#_c_348_n 3.48199e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A2_c_179_n N_A_209_297#_c_348_n 0.0178298f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A2_c_180_n N_VGND_c_369_n 0.00218126f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_180_n N_VGND_c_372_n 0.00428022f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_180_n N_VGND_c_374_n 0.00625078f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_M1000_g N_B1_M1009_g 0.0203059f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_M1000_g B1 3.10428e-19 $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A1_c_213_n B1 3.55259e-19 $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A1_c_214_n B1 0.0418543f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A1_c_213_n N_B1_c_250_n 0.0202959f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A1_c_214_n N_B1_c_250_n 0.00427215f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A1_c_215_n N_B1_c_251_n 0.0102221f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_M1000_g N_VPWR_c_299_n 0.00348446f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_VPWR_c_302_n 0.00437059f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A1_M1000_g N_VPWR_c_297_n 0.00619843f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A1_c_214_n N_A_209_297#_M1000_d 0.00276155f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A1_M1000_g N_A_209_297#_c_348_n 0.0119647f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A1_c_213_n N_A_209_297#_c_348_n 2.08409e-19 $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A1_c_214_n N_A_209_297#_c_348_n 0.00931861f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A1_c_214_n N_A_209_297#_c_355_n 0.00747889f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A1_c_215_n N_VGND_c_372_n 0.00421711f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_215_n N_VGND_c_374_n 0.00613475f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B1_M1009_g N_VPWR_c_302_n 0.00585385f $X=2.4 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1009_g N_VPWR_c_297_n 0.0122361f $X=2.4 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_c_251_n N_VGND_c_370_n 0.00495855f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_251_n N_VGND_c_372_n 0.00427293f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_251_n N_VGND_c_374_n 0.00706845f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_188 X N_VPWR_c_300_n 0.0167669f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_189 N_X_M1005_s N_VPWR_c_297_n 0.00215706f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_190 X N_VPWR_c_297_n 0.0121989f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_191 N_X_c_279_n N_VGND_c_371_n 0.0162614f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_192 N_X_M1002_s N_VGND_c_374_n 0.00216172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_193 N_X_c_279_n N_VGND_c_374_n 0.012122f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_194 N_VPWR_c_297_n N_A_209_297#_M1008_d 0.00298875f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_195 N_VPWR_c_297_n N_A_209_297#_M1000_d 0.00306213f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_299_n N_A_209_297#_c_347_n 0.0161081f $X=1.68 $Y=2.25 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_301_n N_A_209_297#_c_347_n 0.0115771f $X=1.515 $Y=2.72 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_297_n N_A_209_297#_c_347_n 0.00921846f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_199 N_VPWR_M1003_d N_A_209_297#_c_348_n 0.00691181f $X=1.515 $Y=1.485 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_299_n N_A_209_297#_c_348_n 0.0169069f $X=1.68 $Y=2.25 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_301_n N_A_209_297#_c_348_n 0.00276328f $X=1.515 $Y=2.72 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_302_n N_A_209_297#_c_348_n 0.00276328f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_297_n N_A_209_297#_c_348_n 0.0119122f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_299_n N_A_209_297#_c_366_n 0.0161081f $X=1.68 $Y=2.25 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_302_n N_A_209_297#_c_366_n 0.0116427f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_297_n N_A_209_297#_c_366_n 0.00927173f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_207 N_VGND_c_374_n A_209_47# 0.00382975f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_208 N_VGND_c_374_n A_303_47# 0.00394943f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

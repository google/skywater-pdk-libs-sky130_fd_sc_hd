* File: sky130_fd_sc_hd__dfxbp_2.pxi.spice
* Created: Thu Aug 27 14:15:44 2020
* 
x_PM_SKY130_FD_SC_HD__DFXBP_2%CLK N_CLK_c_205_n N_CLK_c_209_n N_CLK_c_206_n
+ N_CLK_M1028_g N_CLK_c_210_n N_CLK_M1017_g N_CLK_c_211_n CLK
+ PM_SKY130_FD_SC_HD__DFXBP_2%CLK
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_27_47# N_A_27_47#_M1028_s N_A_27_47#_M1017_s
+ N_A_27_47#_M1020_g N_A_27_47#_M1000_g N_A_27_47#_M1009_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1024_g N_A_27_47#_c_247_n N_A_27_47#_M1004_g N_A_27_47#_c_470_p
+ N_A_27_47#_c_249_n N_A_27_47#_c_250_n N_A_27_47#_c_262_n N_A_27_47#_c_369_p
+ N_A_27_47#_c_251_n N_A_27_47#_c_252_n N_A_27_47#_c_253_n N_A_27_47#_c_254_n
+ N_A_27_47#_c_265_n N_A_27_47#_c_266_n N_A_27_47#_c_267_n N_A_27_47#_c_268_n
+ N_A_27_47#_c_337_p N_A_27_47#_c_269_n N_A_27_47#_c_270_n N_A_27_47#_c_255_n
+ N_A_27_47#_c_272_n N_A_27_47#_c_256_n N_A_27_47#_c_257_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DFXBP_2%D N_D_M1006_g N_D_M1023_g D N_D_c_489_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%D
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_193_47# N_A_193_47#_M1020_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1012_g N_A_193_47#_c_529_n N_A_193_47#_M1016_g
+ N_A_193_47#_c_531_n N_A_193_47#_M1031_g N_A_193_47#_M1018_g
+ N_A_193_47#_c_532_n N_A_193_47#_c_533_n N_A_193_47#_c_541_n
+ N_A_193_47#_c_542_n N_A_193_47#_c_543_n N_A_193_47#_c_544_n
+ N_A_193_47#_c_589_n N_A_193_47#_c_534_n N_A_193_47#_c_535_n
+ N_A_193_47#_c_536_n N_A_193_47#_c_548_n N_A_193_47#_c_537_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_634_159# N_A_634_159#_M1013_d
+ N_A_634_159#_M1008_d N_A_634_159#_M1029_g N_A_634_159#_M1026_g
+ N_A_634_159#_c_710_n N_A_634_159#_c_733_n N_A_634_159#_c_711_n
+ N_A_634_159#_c_750_p N_A_634_159#_c_712_n N_A_634_159#_c_723_n
+ N_A_634_159#_c_713_n N_A_634_159#_c_714_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_634_159#
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_466_413# N_A_466_413#_M1009_d
+ N_A_466_413#_M1012_d N_A_466_413#_c_798_n N_A_466_413#_M1008_g
+ N_A_466_413#_M1013_g N_A_466_413#_c_799_n N_A_466_413#_c_800_n
+ N_A_466_413#_c_801_n N_A_466_413#_c_802_n N_A_466_413#_c_818_n
+ N_A_466_413#_c_824_n N_A_466_413#_c_803_n N_A_466_413#_c_808_n
+ N_A_466_413#_c_809_n N_A_466_413#_c_810_n N_A_466_413#_c_804_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_466_413#
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_1059_315# N_A_1059_315#_M1015_s
+ N_A_1059_315#_M1025_s N_A_1059_315#_M1007_g N_A_1059_315#_M1011_g
+ N_A_1059_315#_M1014_g N_A_1059_315#_c_919_n N_A_1059_315#_M1021_g
+ N_A_1059_315#_M1019_g N_A_1059_315#_c_920_n N_A_1059_315#_M1022_g
+ N_A_1059_315#_c_921_n N_A_1059_315#_c_922_n N_A_1059_315#_c_923_n
+ N_A_1059_315#_M1002_g N_A_1059_315#_M1010_g N_A_1059_315#_c_924_n
+ N_A_1059_315#_c_925_n N_A_1059_315#_c_926_n N_A_1059_315#_c_939_n
+ N_A_1059_315#_c_940_n N_A_1059_315#_c_941_n N_A_1059_315#_c_942_n
+ N_A_1059_315#_c_943_n N_A_1059_315#_c_927_n N_A_1059_315#_c_928_n
+ N_A_1059_315#_c_944_n N_A_1059_315#_c_929_n N_A_1059_315#_c_946_n
+ N_A_1059_315#_c_930_n N_A_1059_315#_c_964_p
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_1059_315#
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_891_413# N_A_891_413#_M1031_d
+ N_A_891_413#_M1024_d N_A_891_413#_M1025_g N_A_891_413#_c_1065_n
+ N_A_891_413#_M1015_g N_A_891_413#_c_1066_n N_A_891_413#_c_1067_n
+ N_A_891_413#_c_1076_n N_A_891_413#_c_1079_n N_A_891_413#_c_1068_n
+ N_A_891_413#_c_1074_n N_A_891_413#_c_1069_n N_A_891_413#_c_1070_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_891_413#
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_1589_47# N_A_1589_47#_M1002_s
+ N_A_1589_47#_M1010_s N_A_1589_47#_c_1147_n N_A_1589_47#_M1003_g
+ N_A_1589_47#_M1027_g N_A_1589_47#_c_1148_n N_A_1589_47#_M1005_g
+ N_A_1589_47#_M1030_g N_A_1589_47#_c_1155_n N_A_1589_47#_c_1156_n
+ N_A_1589_47#_c_1149_n N_A_1589_47#_c_1150_n N_A_1589_47#_c_1151_n
+ N_A_1589_47#_c_1158_n N_A_1589_47#_c_1179_n N_A_1589_47#_c_1152_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_1589_47#
x_PM_SKY130_FD_SC_HD__DFXBP_2%VPWR N_VPWR_M1017_d N_VPWR_M1023_s N_VPWR_M1029_d
+ N_VPWR_M1007_d N_VPWR_M1025_d N_VPWR_M1019_d N_VPWR_M1010_d N_VPWR_M1030_d
+ N_VPWR_c_1225_n N_VPWR_c_1226_n N_VPWR_c_1227_n N_VPWR_c_1228_n
+ N_VPWR_c_1229_n N_VPWR_c_1230_n N_VPWR_c_1231_n N_VPWR_c_1232_n
+ N_VPWR_c_1233_n N_VPWR_c_1234_n N_VPWR_c_1235_n N_VPWR_c_1236_n
+ N_VPWR_c_1237_n N_VPWR_c_1238_n N_VPWR_c_1239_n N_VPWR_c_1240_n
+ N_VPWR_c_1241_n VPWR N_VPWR_c_1242_n N_VPWR_c_1243_n N_VPWR_c_1244_n
+ N_VPWR_c_1245_n N_VPWR_c_1246_n N_VPWR_c_1247_n N_VPWR_c_1248_n
+ N_VPWR_c_1224_n PM_SKY130_FD_SC_HD__DFXBP_2%VPWR
x_PM_SKY130_FD_SC_HD__DFXBP_2%A_381_47# N_A_381_47#_M1006_d N_A_381_47#_M1023_d
+ N_A_381_47#_c_1373_n N_A_381_47#_c_1376_n N_A_381_47#_c_1371_n
+ N_A_381_47#_c_1372_n N_A_381_47#_c_1375_n N_A_381_47#_c_1387_n
+ PM_SKY130_FD_SC_HD__DFXBP_2%A_381_47#
x_PM_SKY130_FD_SC_HD__DFXBP_2%Q N_Q_M1021_s N_Q_M1014_s N_Q_c_1427_n
+ N_Q_c_1425_n N_Q_c_1438_n Q N_Q_c_1444_n PM_SKY130_FD_SC_HD__DFXBP_2%Q
x_PM_SKY130_FD_SC_HD__DFXBP_2%Q_N N_Q_N_M1003_s N_Q_N_M1027_s N_Q_N_c_1466_n
+ N_Q_N_c_1463_n Q_N N_Q_N_c_1464_n Q_N PM_SKY130_FD_SC_HD__DFXBP_2%Q_N
x_PM_SKY130_FD_SC_HD__DFXBP_2%VGND N_VGND_M1028_d N_VGND_M1006_s N_VGND_M1026_d
+ N_VGND_M1011_d N_VGND_M1015_d N_VGND_M1022_d N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_c_1483_n N_VGND_c_1484_n N_VGND_c_1485_n N_VGND_c_1486_n
+ N_VGND_c_1487_n N_VGND_c_1488_n N_VGND_c_1489_n N_VGND_c_1490_n
+ N_VGND_c_1491_n N_VGND_c_1492_n N_VGND_c_1493_n N_VGND_c_1494_n
+ N_VGND_c_1495_n N_VGND_c_1496_n N_VGND_c_1497_n VGND N_VGND_c_1498_n
+ N_VGND_c_1499_n N_VGND_c_1500_n N_VGND_c_1501_n N_VGND_c_1502_n
+ N_VGND_c_1503_n N_VGND_c_1504_n N_VGND_c_1505_n N_VGND_c_1506_n
+ N_VGND_c_1507_n PM_SKY130_FD_SC_HD__DFXBP_2%VGND
cc_1 VNB N_CLK_c_205_n 0.0577303f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.325
cc_2 VNB N_CLK_c_206_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0187424f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1020_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_5 VNB N_A_27_47#_M1009_g 0.0201185f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_A_27_47#_c_247_n 0.0139254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1004_g 0.0468453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_249_n 0.00174761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_250_n 0.00642437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_251_n 0.00246672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_252_n 0.00476174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_253_n 0.028129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_254_n 0.00413669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_255_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_256_n 0.00991732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_257_n 0.00554756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1006_g 0.0510188f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_18 VNB D 0.0148295f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_19 VNB N_A_193_47#_c_529_n 0.0150433f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_20 VNB N_A_193_47#_M1016_g 0.0410877f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_21 VNB N_A_193_47#_c_531_n 0.0181685f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_22 VNB N_A_193_47#_c_532_n 0.00392862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_193_47#_c_533_n 0.0306268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_193_47#_c_534_n 0.00250297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_c_535_n 0.0103947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_536_n 0.00328545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_537_n 0.0131782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_634_159#_M1029_g 0.0135419f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_29 VNB N_A_634_159#_M1026_g 0.0196396f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_30 VNB N_A_634_159#_c_710_n 0.00301483f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_31 VNB N_A_634_159#_c_711_n 0.00253803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_634_159#_c_712_n 0.00185702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_634_159#_c_713_n 0.00302393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_634_159#_c_714_n 0.0330642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_466_413#_c_798_n 0.0118387f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_36 VNB N_A_466_413#_c_799_n 0.0153956f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_37 VNB N_A_466_413#_c_800_n 0.0132021f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_38 VNB N_A_466_413#_c_801_n 0.00937197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_466_413#_c_802_n 8.51874e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_466_413#_c_803_n 0.00500789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_466_413#_c_804_n 0.00203506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_1059_315#_M1011_g 0.0491605f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_43 VNB N_A_1059_315#_c_919_n 0.016217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_1059_315#_c_920_n 0.0196899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_1059_315#_c_921_n 0.0520616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1059_315#_c_922_n 0.0289124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1059_315#_c_923_n 0.00961911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1059_315#_c_924_n 0.0179129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1059_315#_c_925_n 0.0111966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1059_315#_c_926_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1059_315#_c_927_n 0.00409052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1059_315#_c_928_n 0.00159557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1059_315#_c_929_n 0.00373683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1059_315#_c_930_n 0.00294971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_891_413#_c_1065_n 0.0201807f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_56 VNB N_A_891_413#_c_1066_n 0.0425915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_891_413#_c_1067_n 0.00868625f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_58 VNB N_A_891_413#_c_1068_n 0.00702319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_891_413#_c_1069_n 0.00755581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_891_413#_c_1070_n 0.002763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1589_47#_c_1147_n 0.0166962f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_62 VNB N_A_1589_47#_c_1148_n 0.0209917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1589_47#_c_1149_n 0.00504231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1589_47#_c_1150_n 0.00299916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1589_47#_c_1151_n 0.00378506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1589_47#_c_1152_n 0.0512674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VPWR_c_1224_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_381_47#_c_1371_n 0.00302607f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_69 VNB N_A_381_47#_c_1372_n 0.00471007f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_70 VNB N_Q_c_1425_n 0.00107771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_Q_N_c_1463_n 4.71558e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_72 VNB N_Q_N_c_1464_n 0.00103074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1483_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1484_n 0.00815485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1485_n 0.002903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1486_n 0.00495442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1487_n 0.00412995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1488_n 0.00417678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1489_n 0.0043628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1490_n 0.01004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1491_n 0.0337939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1492_n 0.0486029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1493_n 0.00401403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1494_n 0.0214543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1495_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1496_n 0.0181932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1497_n 0.00324414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1498_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1499_n 0.0165423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1500_n 0.0442602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1501_n 0.0239951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1502_n 0.0154896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1503_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1504_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1505_n 0.00569971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1506_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1507_n 0.478709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VPB N_CLK_c_205_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.325
cc_99 VPB N_CLK_c_209_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_100 VPB N_CLK_c_210_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_101 VPB N_CLK_c_211_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_102 VPB CLK 0.0177397f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_103 VPB N_A_27_47#_M1000_g 0.0363957f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_104 VPB N_A_27_47#_M1001_g 0.0194139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_M1024_g 0.0337518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_47#_c_247_n 0.0198013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_47#_c_262_n 0.00164133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_c_251_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_c_254_n 0.00294199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_c_265_n 0.00356676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_266_n 0.0146795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_c_267_n 0.00167498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_27_47#_c_268_n 8.93482e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_27_47#_c_269_n 0.00927855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_270_n 0.00408403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_255_n 0.0116518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_272_n 0.027052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_c_256_n 0.0214134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_257_n 0.00376433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_D_M1006_g 0.00138392f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_121 VPB N_D_M1023_g 0.0372175f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_122 VPB D 0.00524197f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_123 VPB N_D_c_489_n 0.0483462f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_124 VPB N_A_193_47#_M1012_g 0.0401277f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_125 VPB N_A_193_47#_c_529_n 0.0146132f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_126 VPB N_A_193_47#_M1018_g 0.0210305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_193_47#_c_541_n 0.0103414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_193_47#_c_542_n 0.00544274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_193_47#_c_543_n 0.0161262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_193_47#_c_544_n 0.00124024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_193_47#_c_534_n 0.00678993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_193_47#_c_535_n 0.0183158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_193_47#_c_536_n 0.00299446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_193_47#_c_548_n 0.0265183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_193_47#_c_537_n 0.0106408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_634_159#_M1029_g 0.0524393f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_137 VPB N_A_634_159#_c_713_n 0.00217667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_466_413#_M1008_g 0.0224299f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_139 VPB N_A_466_413#_c_801_n 0.018904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_466_413#_c_802_n 0.00681499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_466_413#_c_808_n 0.00401864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_466_413#_c_809_n 0.00132049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_466_413#_c_810_n 0.00156001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_466_413#_c_804_n 0.00457166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_1059_315#_M1007_g 0.0241837f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_146 VPB N_A_1059_315#_M1011_g 0.0176141f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_147 VPB N_A_1059_315#_M1014_g 0.0187898f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_148 VPB N_A_1059_315#_M1019_g 0.0226685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_1059_315#_c_921_n 0.0276548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_1059_315#_c_922_n 0.0062547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_1059_315#_M1010_g 0.0252571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_1059_315#_c_926_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_1059_315#_c_939_n 0.0126366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_1059_315#_c_940_n 0.0130917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_1059_315#_c_941_n 0.0116311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_1059_315#_c_942_n 0.0408399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_1059_315#_c_943_n 0.00735054f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_1059_315#_c_944_n 0.00231284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_1059_315#_c_929_n 0.00346808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_1059_315#_c_946_n 0.00102121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_891_413#_M1025_g 0.0233469f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_162 VPB N_A_891_413#_c_1066_n 0.0155556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_891_413#_c_1067_n 0.00108521f $X=-0.19 $Y=1.305 $X2=0.327
+ $Y2=1.16
cc_164 VPB N_A_891_413#_c_1074_n 0.00703062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_891_413#_c_1069_n 0.00302752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1589_47#_M1027_g 0.019727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1589_47#_M1030_g 0.0253014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1589_47#_c_1155_n 0.00282264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_1589_47#_c_1156_n 0.00651067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1589_47#_c_1150_n 0.00399301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_1589_47#_c_1158_n 0.00544737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1589_47#_c_1152_n 0.0108905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1225_n 0.00105771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1226_n 0.00820812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1227_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1228_n 0.0107474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1229_n 0.00411841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1230_n 0.0042033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1231_n 0.00658407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1232_n 0.0100108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1233_n 0.0422235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1234_n 0.0494152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1235_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1236_n 0.044979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1237_n 0.00603258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1238_n 0.0203381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1239_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1240_n 0.0184312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1241_n 0.00334019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1242_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1243_n 0.0162996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1244_n 0.0243358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1245_n 0.0180594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1246_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1247_n 0.00506592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1248_n 0.00410625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1224_n 0.0708186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_381_47#_c_1373_n 2.53606e-19 $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_199 VPB N_A_381_47#_c_1372_n 0.00370682f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_200 VPB N_A_381_47#_c_1375_n 0.00296152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_Q_c_1425_n 0.00199028f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_Q_N_c_1464_n 0.00151302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 N_CLK_c_205_n N_A_27_47#_M1020_g 0.00510767f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_204 N_CLK_c_206_n N_A_27_47#_M1020_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_205 CLK N_A_27_47#_M1020_g 3.09846e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_206 N_CLK_c_209_n N_A_27_47#_M1000_g 0.00531917f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_207 N_CLK_c_211_n N_A_27_47#_M1000_g 0.0276478f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_208 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_209 N_CLK_c_205_n N_A_27_47#_c_249_n 0.00787672f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_210 N_CLK_c_206_n N_A_27_47#_c_249_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_211 CLK N_A_27_47#_c_249_n 0.00736322f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_212 N_CLK_c_205_n N_A_27_47#_c_250_n 0.00639426f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_213 CLK N_A_27_47#_c_250_n 0.0144136f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_214 N_CLK_c_210_n N_A_27_47#_c_262_n 0.0128144f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_215 N_CLK_c_211_n N_A_27_47#_c_262_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_216 CLK N_A_27_47#_c_262_n 0.00728212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_217 N_CLK_c_205_n N_A_27_47#_c_251_n 0.00466159f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_218 N_CLK_c_209_n N_A_27_47#_c_251_n 7.09762e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_219 N_CLK_c_211_n N_A_27_47#_c_251_n 0.00440146f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_220 CLK N_A_27_47#_c_251_n 0.0511527f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_221 N_CLK_c_205_n N_A_27_47#_c_265_n 2.26313e-19 $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_222 N_CLK_c_210_n N_A_27_47#_c_265_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_223 N_CLK_c_211_n N_A_27_47#_c_265_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_224 CLK N_A_27_47#_c_265_n 0.0153364f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_225 N_CLK_c_210_n N_A_27_47#_c_267_n 0.00101667f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_226 N_CLK_c_205_n N_A_27_47#_c_255_n 0.0169285f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_227 CLK N_A_27_47#_c_255_n 0.00161876f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_228 N_CLK_c_210_n N_VPWR_c_1225_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_229 N_CLK_c_210_n N_VPWR_c_1242_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_230 N_CLK_c_210_n N_VPWR_c_1224_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_231 N_CLK_c_206_n N_VGND_c_1483_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_232 N_CLK_c_205_n N_VGND_c_1498_n 4.74473e-19 $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_233 N_CLK_c_206_n N_VGND_c_1498_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_234 N_CLK_c_206_n N_VGND_c_1507_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_235 N_A_27_47#_M1009_g N_D_M1006_g 0.011413f $X=2.39 $Y=0.415 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_252_n N_D_M1006_g 2.41107e-19 $X=2.57 $Y=0.845 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_253_n N_D_M1006_g 0.0106161f $X=2.38 $Y=0.87 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_254_n N_D_M1006_g 6.39744e-19 $X=2.655 $Y=1.655 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_266_n N_D_M1023_g 0.00400813f $X=2.67 $Y=1.87 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_266_n D 0.00506217f $X=2.67 $Y=1.87 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_266_n N_D_c_489_n 0.00164848f $X=2.67 $Y=1.87 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_255_n N_D_c_489_n 0.00766286f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_266_n N_A_193_47#_M1000_d 0.00105035f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_254_n N_A_193_47#_M1012_g 6.96305e-19 $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_245 N_A_27_47#_c_266_n N_A_193_47#_M1012_g 0.00581536f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_269_n N_A_193_47#_M1012_g 0.00279586f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_272_n N_A_193_47#_M1012_g 0.024974f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_252_n N_A_193_47#_c_529_n 7.84575e-19 $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_254_n N_A_193_47#_c_529_n 0.0124732f $X=2.655 $Y=1.655 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_269_n N_A_193_47#_c_529_n 0.00141049f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_272_n N_A_193_47#_c_529_n 0.020457f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1009_g N_A_193_47#_M1016_g 0.0176128f $X=2.39 $Y=0.415 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_252_n N_A_193_47#_M1016_g 0.00162274f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_253_n N_A_193_47#_M1016_g 0.0115319f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_254_n N_A_193_47#_M1016_g 0.00482947f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_256 N_A_27_47#_M1004_g N_A_193_47#_c_531_n 0.0149277f $X=5.01 $Y=0.415 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1024_g N_A_193_47#_M1018_g 0.0177205f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1004_g N_A_193_47#_c_532_n 0.00705204f $X=5.01 $Y=0.415 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_256_n N_A_193_47#_c_532_n 9.61914e-19 $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1004_g N_A_193_47#_c_533_n 0.0213226f $X=5.01 $Y=0.415 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_256_n N_A_193_47#_c_533_n 0.0204589f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_257_n N_A_193_47#_c_533_n 5.64291e-19 $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_266_n N_A_193_47#_c_541_n 0.0717579f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1000_g N_A_193_47#_c_542_n 0.00496481f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_251_n N_A_193_47#_c_542_n 0.00662493f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_266 N_A_27_47#_c_266_n N_A_193_47#_c_542_n 0.0260848f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_247_n N_A_193_47#_c_543_n 0.00316727f $X=4.935 $Y=1.32 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_252_n N_A_193_47#_c_543_n 0.00384011f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_254_n N_A_193_47#_c_543_n 0.0122753f $X=2.655 $Y=1.655 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_266_n N_A_193_47#_c_543_n 0.017766f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_268_n N_A_193_47#_c_543_n 0.102076f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_337_p N_A_193_47#_c_543_n 0.0257765f $X=2.96 $Y=1.87 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_269_n N_A_193_47#_c_543_n 0.00669423f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_270_n N_A_193_47#_c_543_n 0.026031f $X=4.385 $Y=1.87 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_272_n N_A_193_47#_c_543_n 0.00145041f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_256_n N_A_193_47#_c_543_n 0.00523342f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_257_n N_A_193_47#_c_543_n 0.0150724f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_252_n N_A_193_47#_c_544_n 0.00207033f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_253_n N_A_193_47#_c_544_n 2.23087e-19 $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_254_n N_A_193_47#_c_544_n 0.00253246f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_266_n N_A_193_47#_c_544_n 0.026464f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_257_n N_A_193_47#_c_589_n 6.19759e-19 $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1024_g N_A_193_47#_c_534_n 0.0016378f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_247_n N_A_193_47#_c_534_n 0.0169257f $X=4.935 $Y=1.32 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1004_g N_A_193_47#_c_534_n 0.00640774f $X=5.01 $Y=0.415 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_270_n N_A_193_47#_c_534_n 0.00786261f $X=4.385 $Y=1.87 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_256_n N_A_193_47#_c_534_n 0.00345899f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_257_n N_A_193_47#_c_534_n 0.051468f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_252_n N_A_193_47#_c_535_n 0.00105611f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_253_n N_A_193_47#_c_535_n 0.0212537f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_254_n N_A_193_47#_c_535_n 0.00246225f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_266_n N_A_193_47#_c_535_n 4.12072e-19 $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_252_n N_A_193_47#_c_536_n 0.0144031f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_253_n N_A_193_47#_c_536_n 0.00126202f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_254_n N_A_193_47#_c_536_n 0.0374587f $X=2.655 $Y=1.655 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_266_n N_A_193_47#_c_536_n 0.00639021f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_269_n N_A_193_47#_c_536_n 0.00542444f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_272_n N_A_193_47#_c_536_n 3.63869e-19 $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1024_g N_A_193_47#_c_548_n 0.0130792f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_247_n N_A_193_47#_c_548_n 0.0224153f $X=4.935 $Y=1.32 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_257_n N_A_193_47#_c_548_n 6.57469e-19 $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1020_g N_A_193_47#_c_537_n 0.0226423f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_249_n N_A_193_47#_c_537_n 0.0125576f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_369_p N_A_193_47#_c_537_n 0.0082461f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_251_n N_A_193_47#_c_537_n 0.0683411f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_266_n N_A_193_47#_c_537_n 0.0153552f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_267_n N_A_193_47#_c_537_n 0.00241547f $X=0.86 $Y=1.87 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_268_n N_A_634_159#_M1008_d 0.00201378f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1001_g N_A_634_159#_M1029_g 0.0245145f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_254_n N_A_634_159#_M1029_g 0.00171004f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_268_n N_A_634_159#_M1029_g 0.00244796f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_269_n N_A_634_159#_M1029_g 0.00243934f $X=2.815 $Y=1.87
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_272_n N_A_634_159#_M1029_g 0.0205969f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_268_n N_A_634_159#_c_723_n 0.00261642f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_M1024_g N_A_634_159#_c_713_n 0.00420906f $X=4.38 $Y=2.275
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_268_n N_A_634_159#_c_713_n 0.0130552f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_270_n N_A_634_159#_c_713_n 0.00283183f $X=4.385 $Y=1.87
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_c_256_n N_A_634_159#_c_713_n 0.00209722f $X=4.375 $Y=1.32
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_257_n N_A_634_159#_c_713_n 0.0508796f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_256_n N_A_466_413#_c_798_n 0.0165206f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_257_n N_A_466_413#_c_798_n 3.51062e-19 $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_M1024_g N_A_466_413#_M1008_g 0.0247799f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_268_n N_A_466_413#_M1008_g 0.00324412f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_257_n N_A_466_413#_M1008_g 8.16982e-19 $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_268_n N_A_466_413#_c_801_n 2.40114e-19 $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_M1001_g N_A_466_413#_c_818_n 0.00870465f $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_266_n N_A_466_413#_c_818_n 0.00598509f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_268_n N_A_466_413#_c_818_n 0.004788f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_337_p N_A_466_413#_c_818_n 0.00111365f $X=2.96 $Y=1.87 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_269_n N_A_466_413#_c_818_n 0.0322466f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_272_n N_A_466_413#_c_818_n 7.1695e-19 $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_M1009_g N_A_466_413#_c_824_n 0.00387559f $X=2.39 $Y=0.415
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_252_n N_A_466_413#_c_824_n 0.0197404f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_253_n N_A_466_413#_c_824_n 0.00155178f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_M1009_g N_A_466_413#_c_803_n 8.47674e-19 $X=2.39 $Y=0.415
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_252_n N_A_466_413#_c_803_n 0.0173602f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_254_n N_A_466_413#_c_803_n 0.0252666f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_268_n N_A_466_413#_c_808_n 0.00158456f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_269_n N_A_466_413#_c_808_n 0.00132833f $X=2.815 $Y=1.87
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_254_n N_A_466_413#_c_809_n 0.0134794f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_269_n N_A_466_413#_c_809_n 0.0117702f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_272_n N_A_466_413#_c_809_n 2.6825e-19 $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_M1001_g N_A_466_413#_c_810_n 9.36024e-19 $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_c_254_n N_A_466_413#_c_810_n 0.0018075f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_268_n N_A_466_413#_c_810_n 0.0127304f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_337_p N_A_466_413#_c_810_n 4.44641e-19 $X=2.96 $Y=1.87 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_269_n N_A_466_413#_c_810_n 0.0269253f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_272_n N_A_466_413#_c_810_n 5.28921e-19 $X=2.825 $Y=1.74
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_254_n N_A_466_413#_c_804_n 0.00156136f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_268_n N_A_466_413#_c_804_n 0.00178543f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_M1004_g N_A_1059_315#_M1011_g 0.0425652f $X=5.01 $Y=0.415
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_M1024_g N_A_891_413#_c_1076_n 0.00281529f $X=4.38 $Y=2.275
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_270_n N_A_891_413#_c_1076_n 0.00210372f $X=4.385 $Y=1.87
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_257_n N_A_891_413#_c_1076_n 0.0022468f $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_M1004_g N_A_891_413#_c_1079_n 0.0141499f $X=5.01 $Y=0.415
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_M1004_g N_A_891_413#_c_1068_n 0.00515031f $X=5.01 $Y=0.415
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_247_n N_A_891_413#_c_1074_n 6.71564e-19 $X=4.935 $Y=1.32
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_M1004_g N_A_891_413#_c_1070_n 0.00301916f $X=5.01 $Y=0.415
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_369_p N_VPWR_M1017_d 6.91013e-19 $X=0.725 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_360 N_A_27_47#_c_267_n N_VPWR_M1017_d 0.00182035f $X=0.86 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_361 N_A_27_47#_c_268_n N_VPWR_M1029_d 0.00522581f $X=4.24 $Y=1.87 $X2=0 $Y2=0
cc_362 N_A_27_47#_M1000_g N_VPWR_c_1225_n 0.0082523f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_262_n N_VPWR_c_1225_n 0.00319791f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_369_p N_VPWR_c_1225_n 0.0133497f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_265_n N_VPWR_c_1225_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_366 N_A_27_47#_c_267_n N_VPWR_c_1225_n 0.00337045f $X=0.86 $Y=1.87 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_M1000_g N_VPWR_c_1226_n 0.00189262f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_266_n N_VPWR_c_1226_n 0.00518847f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_268_n N_VPWR_c_1227_n 0.00950843f $X=4.24 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1001_g N_VPWR_c_1234_n 0.0037886f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_M1024_g N_VPWR_c_1236_n 0.00430107f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_257_n N_VPWR_c_1236_n 0.00157744f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_262_n N_VPWR_c_1242_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_265_n N_VPWR_c_1242_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_375 N_A_27_47#_M1000_g N_VPWR_c_1243_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_M1000_g N_VPWR_c_1224_n 0.00534972f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_M1001_g N_VPWR_c_1224_n 0.00563311f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_M1024_g N_VPWR_c_1224_n 0.0057371f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_262_n N_VPWR_c_1224_n 0.00402226f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_265_n N_VPWR_c_1224_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_266_n N_VPWR_c_1224_n 0.0879363f $X=2.67 $Y=1.87 $X2=0 $Y2=0
cc_382 N_A_27_47#_c_267_n N_VPWR_c_1224_n 0.0145392f $X=0.86 $Y=1.87 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_268_n N_VPWR_c_1224_n 0.060469f $X=4.24 $Y=1.87 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_337_p N_VPWR_c_1224_n 0.0144739f $X=2.96 $Y=1.87 $X2=0 $Y2=0
cc_385 N_A_27_47#_c_270_n N_VPWR_c_1224_n 0.0159329f $X=4.385 $Y=1.87 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_257_n N_VPWR_c_1224_n 0.00100625f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_M1009_g N_A_381_47#_c_1376_n 0.00393136f $X=2.39 $Y=0.415
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_252_n N_A_381_47#_c_1371_n 0.00551543f $X=2.57 $Y=0.845
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_253_n N_A_381_47#_c_1371_n 2.3327e-19 $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_252_n N_A_381_47#_c_1372_n 0.00940942f $X=2.57 $Y=0.845
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_253_n N_A_381_47#_c_1372_n 0.00100695f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_254_n N_A_381_47#_c_1372_n 0.00542297f $X=2.655 $Y=1.655
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_266_n N_A_381_47#_c_1372_n 0.00974994f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_269_n N_A_381_47#_c_1372_n 0.00481141f $X=2.815 $Y=1.87
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_266_n N_A_381_47#_c_1375_n 0.0136242f $X=2.67 $Y=1.87 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_337_p N_A_381_47#_c_1375_n 2.75481e-19 $X=2.96 $Y=1.87 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_269_n N_A_381_47#_c_1375_n 0.00395909f $X=2.815 $Y=1.87
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_M1009_g N_A_381_47#_c_1387_n 0.00144307f $X=2.39 $Y=0.415
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_249_n N_VGND_M1028_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_400 N_A_27_47#_M1020_g N_VGND_c_1483_n 0.0078844f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_249_n N_VGND_c_1483_n 0.0170164f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_402 N_A_27_47#_c_255_n N_VGND_c_1483_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_M1020_g N_VGND_c_1484_n 0.00310005f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_M1004_g N_VGND_c_1492_n 0.0037981f $X=5.01 $Y=0.415 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_470_p N_VGND_c_1498_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_249_n N_VGND_c_1498_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_M1020_g N_VGND_c_1499_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_M1009_g N_VGND_c_1500_n 0.00415447f $X=2.39 $Y=0.415 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_252_n N_VGND_c_1500_n 0.00253275f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_c_253_n N_VGND_c_1500_n 0.00134958f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_M1028_s N_VGND_c_1507_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_M1020_g N_VGND_c_1507_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_M1009_g N_VGND_c_1507_n 0.00636524f $X=2.39 $Y=0.415 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_M1004_g N_VGND_c_1507_n 0.00579f $X=5.01 $Y=0.415 $X2=0 $Y2=0
cc_415 N_A_27_47#_c_470_p N_VGND_c_1507_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_249_n N_VGND_c_1507_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_252_n N_VGND_c_1507_n 0.00474506f $X=2.57 $Y=0.845 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_253_n N_VGND_c_1507_n 0.00232804f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_419 N_D_c_489_n N_A_193_47#_M1012_g 0.0344137f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_420 D N_A_193_47#_c_541_n 0.0242394f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_421 N_D_c_489_n N_A_193_47#_c_541_n 0.00764469f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_422 D N_A_193_47#_c_542_n 0.00276875f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_423 N_D_M1006_g N_A_193_47#_c_535_n 0.0174319f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_424 N_D_M1006_g N_A_193_47#_c_536_n 8.29261e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_425 N_D_c_489_n N_A_193_47#_c_536_n 5.41323e-19 $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_426 N_D_M1006_g N_A_193_47#_c_537_n 0.00322876f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_427 N_D_M1023_g N_A_193_47#_c_537_n 0.00687078f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_428 D N_A_193_47#_c_537_n 0.0727432f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_429 N_D_c_489_n N_A_193_47#_c_537_n 9.27942e-19 $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_430 N_D_M1023_g N_VPWR_c_1226_n 0.00451231f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_431 D N_VPWR_c_1226_n 0.00339786f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_432 N_D_c_489_n N_VPWR_c_1226_n 0.00294108f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_433 N_D_M1023_g N_VPWR_c_1234_n 0.00485948f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_434 N_D_M1023_g N_VPWR_c_1224_n 0.0070625f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_435 N_D_M1023_g N_A_381_47#_c_1373_n 0.0070545f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_436 N_D_M1006_g N_A_381_47#_c_1376_n 0.00350922f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_437 N_D_M1006_g N_A_381_47#_c_1371_n 0.00477479f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_438 D N_A_381_47#_c_1371_n 0.0683394f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_439 N_D_M1006_g N_A_381_47#_c_1372_n 0.0128307f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_440 N_D_M1023_g N_A_381_47#_c_1372_n 0.0068119f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_441 N_D_c_489_n N_A_381_47#_c_1372_n 0.00783483f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_442 N_D_M1023_g N_A_381_47#_c_1375_n 0.00557195f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_443 N_D_M1006_g N_A_381_47#_c_1387_n 0.00233054f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_444 N_D_M1006_g N_VGND_c_1484_n 0.0044954f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_445 D N_VGND_c_1484_n 0.0170306f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_446 D N_VGND_c_1499_n 0.00144897f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_447 N_D_M1006_g N_VGND_c_1500_n 0.00488602f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_448 N_D_M1006_g N_VGND_c_1507_n 0.00943922f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_449 D N_VGND_c_1507_n 0.00327398f $X=1.445 $Y=1.105 $X2=0 $Y2=0
cc_450 N_A_193_47#_c_529_n N_A_634_159#_M1029_g 0.0173021f $X=2.81 $Y=1.29 $X2=0
+ $Y2=0
cc_451 N_A_193_47#_c_543_n N_A_634_159#_M1029_g 0.00240096f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_452 N_A_193_47#_M1016_g N_A_634_159#_M1026_g 0.0232924f $X=2.885 $Y=0.415
+ $X2=0 $Y2=0
cc_453 N_A_193_47#_c_543_n N_A_634_159#_c_710_n 0.00701802f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_454 N_A_193_47#_c_531_n N_A_634_159#_c_733_n 0.00362005f $X=4.48 $Y=0.705
+ $X2=0 $Y2=0
cc_455 N_A_193_47#_c_532_n N_A_634_159#_c_733_n 0.00240286f $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_456 N_A_193_47#_M1016_g N_A_634_159#_c_711_n 3.52512e-19 $X=2.885 $Y=0.415
+ $X2=0 $Y2=0
cc_457 N_A_193_47#_c_543_n N_A_634_159#_c_711_n 0.00115477f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_458 N_A_193_47#_c_532_n N_A_634_159#_c_712_n 0.0124661f $X=4.59 $Y=0.87 $X2=0
+ $Y2=0
cc_459 N_A_193_47#_c_533_n N_A_634_159#_c_712_n 0.00244688f $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_460 N_A_193_47#_c_534_n N_A_634_159#_c_712_n 0.0011821f $X=4.82 $Y=1.53 $X2=0
+ $Y2=0
cc_461 N_A_193_47#_c_543_n N_A_634_159#_c_713_n 0.015392f $X=4.675 $Y=1.53 $X2=0
+ $Y2=0
cc_462 N_A_193_47#_c_534_n N_A_634_159#_c_713_n 0.00707472f $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_463 N_A_193_47#_M1016_g N_A_634_159#_c_714_n 0.0173021f $X=2.885 $Y=0.415
+ $X2=0 $Y2=0
cc_464 N_A_193_47#_c_534_n N_A_466_413#_c_798_n 6.79435e-19 $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_465 N_A_193_47#_c_543_n N_A_466_413#_M1008_g 0.00174404f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_466 N_A_193_47#_c_531_n N_A_466_413#_c_799_n 0.011709f $X=4.48 $Y=0.705 $X2=0
+ $Y2=0
cc_467 N_A_193_47#_c_532_n N_A_466_413#_c_799_n 3.35082e-19 $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_468 N_A_193_47#_c_533_n N_A_466_413#_c_800_n 0.011709f $X=4.59 $Y=0.87 $X2=0
+ $Y2=0
cc_469 N_A_193_47#_c_534_n N_A_466_413#_c_800_n 3.45909e-19 $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_470 N_A_193_47#_c_543_n N_A_466_413#_c_801_n 9.40522e-19 $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_471 N_A_193_47#_c_543_n N_A_466_413#_c_802_n 0.00133421f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_472 N_A_193_47#_c_536_n N_A_466_413#_c_818_n 7.18938e-19 $X=2.28 $Y=1.35
+ $X2=0 $Y2=0
cc_473 N_A_193_47#_c_529_n N_A_466_413#_c_824_n 0.00133503f $X=2.81 $Y=1.29
+ $X2=0 $Y2=0
cc_474 N_A_193_47#_M1016_g N_A_466_413#_c_824_n 0.0124233f $X=2.885 $Y=0.415
+ $X2=0 $Y2=0
cc_475 N_A_193_47#_c_529_n N_A_466_413#_c_803_n 0.00229374f $X=2.81 $Y=1.29
+ $X2=0 $Y2=0
cc_476 N_A_193_47#_M1016_g N_A_466_413#_c_803_n 0.0138754f $X=2.885 $Y=0.415
+ $X2=0 $Y2=0
cc_477 N_A_193_47#_c_543_n N_A_466_413#_c_808_n 0.0122057f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_478 N_A_193_47#_c_529_n N_A_466_413#_c_809_n 0.00166382f $X=2.81 $Y=1.29
+ $X2=0 $Y2=0
cc_479 N_A_193_47#_c_543_n N_A_466_413#_c_809_n 0.00935699f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_480 N_A_193_47#_c_543_n N_A_466_413#_c_810_n 0.0041284f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_481 N_A_193_47#_c_543_n N_A_466_413#_c_804_n 0.0215551f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_482 N_A_193_47#_c_532_n N_A_1059_315#_M1011_g 3.15846e-19 $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_483 N_A_193_47#_M1018_g N_A_1059_315#_c_942_n 0.0200851f $X=4.8 $Y=2.275
+ $X2=0 $Y2=0
cc_484 N_A_193_47#_c_534_n N_A_1059_315#_c_942_n 7.03497e-19 $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_485 N_A_193_47#_c_548_n N_A_1059_315#_c_942_n 0.0137111f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_486 N_A_193_47#_M1018_g N_A_891_413#_c_1076_n 0.00914972f $X=4.8 $Y=2.275
+ $X2=0 $Y2=0
cc_487 N_A_193_47#_c_543_n N_A_891_413#_c_1076_n 0.00392926f $X=4.675 $Y=1.53
+ $X2=0 $Y2=0
cc_488 N_A_193_47#_c_589_n N_A_891_413#_c_1076_n 0.00102192f $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_489 N_A_193_47#_c_534_n N_A_891_413#_c_1076_n 0.0197136f $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_490 N_A_193_47#_c_548_n N_A_891_413#_c_1076_n 0.0030041f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_491 N_A_193_47#_c_531_n N_A_891_413#_c_1079_n 0.00256259f $X=4.48 $Y=0.705
+ $X2=0 $Y2=0
cc_492 N_A_193_47#_c_532_n N_A_891_413#_c_1079_n 0.0294378f $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_493 N_A_193_47#_c_533_n N_A_891_413#_c_1079_n 0.00107404f $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_494 N_A_193_47#_c_532_n N_A_891_413#_c_1068_n 0.0223409f $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_495 N_A_193_47#_M1018_g N_A_891_413#_c_1074_n 0.00365921f $X=4.8 $Y=2.275
+ $X2=0 $Y2=0
cc_496 N_A_193_47#_c_589_n N_A_891_413#_c_1074_n 0.00168323f $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_497 N_A_193_47#_c_534_n N_A_891_413#_c_1074_n 0.0495221f $X=4.82 $Y=1.53
+ $X2=0 $Y2=0
cc_498 N_A_193_47#_c_548_n N_A_891_413#_c_1074_n 0.00182086f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_499 N_A_193_47#_c_532_n N_A_891_413#_c_1070_n 0.0277807f $X=4.59 $Y=0.87
+ $X2=0 $Y2=0
cc_500 N_A_193_47#_c_537_n N_VPWR_c_1225_n 0.0127254f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_501 N_A_193_47#_c_537_n N_VPWR_c_1226_n 0.0174675f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_502 N_A_193_47#_c_543_n N_VPWR_c_1227_n 5.88241e-19 $X=4.675 $Y=1.53 $X2=0
+ $Y2=0
cc_503 N_A_193_47#_M1012_g N_VPWR_c_1234_n 0.00585385f $X=2.255 $Y=2.275 $X2=0
+ $Y2=0
cc_504 N_A_193_47#_M1018_g N_VPWR_c_1236_n 0.00383564f $X=4.8 $Y=2.275 $X2=0
+ $Y2=0
cc_505 N_A_193_47#_c_537_n N_VPWR_c_1243_n 0.0131202f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_506 N_A_193_47#_M1012_g N_VPWR_c_1224_n 0.00659322f $X=2.255 $Y=2.275 $X2=0
+ $Y2=0
cc_507 N_A_193_47#_M1018_g N_VPWR_c_1224_n 0.00576282f $X=4.8 $Y=2.275 $X2=0
+ $Y2=0
cc_508 N_A_193_47#_c_537_n N_VPWR_c_1224_n 0.00335714f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_509 N_A_193_47#_c_537_n N_A_381_47#_c_1373_n 0.00327515f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_510 N_A_193_47#_c_537_n N_A_381_47#_c_1376_n 0.00309965f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_511 N_A_193_47#_c_537_n N_A_381_47#_c_1371_n 0.00907577f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_512 N_A_193_47#_M1012_g N_A_381_47#_c_1372_n 0.00218414f $X=2.255 $Y=2.275
+ $X2=0 $Y2=0
cc_513 N_A_193_47#_c_541_n N_A_381_47#_c_1372_n 0.0169549f $X=2.155 $Y=1.53
+ $X2=0 $Y2=0
cc_514 N_A_193_47#_c_544_n N_A_381_47#_c_1372_n 0.00241524f $X=2.445 $Y=1.53
+ $X2=0 $Y2=0
cc_515 N_A_193_47#_c_535_n N_A_381_47#_c_1372_n 0.00162494f $X=2.28 $Y=1.29
+ $X2=0 $Y2=0
cc_516 N_A_193_47#_c_536_n N_A_381_47#_c_1372_n 0.0430896f $X=2.28 $Y=1.35 $X2=0
+ $Y2=0
cc_517 N_A_193_47#_M1012_g N_A_381_47#_c_1375_n 0.00251259f $X=2.255 $Y=2.275
+ $X2=0 $Y2=0
cc_518 N_A_193_47#_c_541_n N_A_381_47#_c_1375_n 7.34738e-19 $X=2.155 $Y=1.53
+ $X2=0 $Y2=0
cc_519 N_A_193_47#_c_535_n N_A_381_47#_c_1387_n 0.00121425f $X=2.28 $Y=1.29
+ $X2=0 $Y2=0
cc_520 N_A_193_47#_c_536_n N_A_381_47#_c_1387_n 0.00164458f $X=2.28 $Y=1.35
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_c_537_n N_VGND_c_1484_n 0.0114765f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_522 N_A_193_47#_M1016_g N_VGND_c_1485_n 0.0018559f $X=2.885 $Y=0.415 $X2=0
+ $Y2=0
cc_523 N_A_193_47#_c_531_n N_VGND_c_1492_n 0.00525217f $X=4.48 $Y=0.705 $X2=0
+ $Y2=0
cc_524 N_A_193_47#_c_532_n N_VGND_c_1492_n 2.78187e-19 $X=4.59 $Y=0.87 $X2=0
+ $Y2=0
cc_525 N_A_193_47#_c_537_n N_VGND_c_1499_n 0.00799435f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_526 N_A_193_47#_M1016_g N_VGND_c_1500_n 0.00379747f $X=2.885 $Y=0.415 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_M1020_d N_VGND_c_1507_n 0.0048343f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_528 N_A_193_47#_M1016_g N_VGND_c_1507_n 0.00575924f $X=2.885 $Y=0.415 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_c_531_n N_VGND_c_1507_n 0.00962915f $X=4.48 $Y=0.705 $X2=0
+ $Y2=0
cc_530 N_A_193_47#_c_532_n N_VGND_c_1507_n 0.00130853f $X=4.59 $Y=0.87 $X2=0
+ $Y2=0
cc_531 N_A_193_47#_c_537_n N_VGND_c_1507_n 0.00671652f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_532 N_A_634_159#_c_713_n N_A_466_413#_c_798_n 0.00595764f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_533 N_A_634_159#_M1029_g N_A_466_413#_M1008_g 0.0141558f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_534 N_A_634_159#_c_723_n N_A_466_413#_M1008_g 0.00378805f $X=4.115 $Y=2.3
+ $X2=0 $Y2=0
cc_535 N_A_634_159#_c_713_n N_A_466_413#_M1008_g 0.0120712f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_536 N_A_634_159#_M1026_g N_A_466_413#_c_799_n 0.0119448f $X=3.38 $Y=0.445
+ $X2=0 $Y2=0
cc_537 N_A_634_159#_c_710_n N_A_466_413#_c_799_n 0.00465161f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_538 N_A_634_159#_c_733_n N_A_466_413#_c_799_n 0.00666448f $X=4.035 $Y=0.765
+ $X2=0 $Y2=0
cc_539 N_A_634_159#_c_750_p N_A_466_413#_c_799_n 0.00425242f $X=4.19 $Y=0.45
+ $X2=0 $Y2=0
cc_540 N_A_634_159#_c_712_n N_A_466_413#_c_799_n 0.00299006f $X=4.035 $Y=0.915
+ $X2=0 $Y2=0
cc_541 N_A_634_159#_c_714_n N_A_466_413#_c_799_n 0.00500472f $X=3.38 $Y=0.93
+ $X2=0 $Y2=0
cc_542 N_A_634_159#_M1029_g N_A_466_413#_c_800_n 0.00465771f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_543 N_A_634_159#_c_710_n N_A_466_413#_c_800_n 0.0064477f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_544 N_A_634_159#_c_711_n N_A_466_413#_c_800_n 2.46982e-19 $X=3.49 $Y=0.93
+ $X2=0 $Y2=0
cc_545 N_A_634_159#_c_712_n N_A_466_413#_c_800_n 0.00212952f $X=4.035 $Y=0.915
+ $X2=0 $Y2=0
cc_546 N_A_634_159#_c_713_n N_A_466_413#_c_800_n 0.00312426f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_547 N_A_634_159#_c_714_n N_A_466_413#_c_800_n 0.0049948f $X=3.38 $Y=0.93
+ $X2=0 $Y2=0
cc_548 N_A_634_159#_M1029_g N_A_466_413#_c_801_n 0.0173911f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_549 N_A_634_159#_c_710_n N_A_466_413#_c_801_n 0.00455719f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_550 N_A_634_159#_c_714_n N_A_466_413#_c_801_n 5.95332e-19 $X=3.38 $Y=0.93
+ $X2=0 $Y2=0
cc_551 N_A_634_159#_c_713_n N_A_466_413#_c_802_n 0.00562808f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_552 N_A_634_159#_M1029_g N_A_466_413#_c_818_n 0.0102787f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_553 N_A_634_159#_M1026_g N_A_466_413#_c_824_n 0.00143041f $X=3.38 $Y=0.445
+ $X2=0 $Y2=0
cc_554 N_A_634_159#_M1026_g N_A_466_413#_c_803_n 0.00406017f $X=3.38 $Y=0.445
+ $X2=0 $Y2=0
cc_555 N_A_634_159#_c_711_n N_A_466_413#_c_803_n 0.0222621f $X=3.49 $Y=0.93
+ $X2=0 $Y2=0
cc_556 N_A_634_159#_c_714_n N_A_466_413#_c_803_n 0.00601957f $X=3.38 $Y=0.93
+ $X2=0 $Y2=0
cc_557 N_A_634_159#_M1029_g N_A_466_413#_c_808_n 0.0108535f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_558 N_A_634_159#_M1029_g N_A_466_413#_c_810_n 0.0153425f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_559 N_A_634_159#_c_713_n N_A_466_413#_c_810_n 0.00722041f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_560 N_A_634_159#_M1029_g N_A_466_413#_c_804_n 0.00658437f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_561 N_A_634_159#_c_710_n N_A_466_413#_c_804_n 0.0189518f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_562 N_A_634_159#_c_711_n N_A_466_413#_c_804_n 0.0129752f $X=3.49 $Y=0.93
+ $X2=0 $Y2=0
cc_563 N_A_634_159#_c_713_n N_A_466_413#_c_804_n 0.0235594f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_564 N_A_634_159#_c_714_n N_A_466_413#_c_804_n 0.0020325f $X=3.38 $Y=0.93
+ $X2=0 $Y2=0
cc_565 N_A_634_159#_c_723_n N_A_891_413#_c_1076_n 0.0109209f $X=4.115 $Y=2.3
+ $X2=0 $Y2=0
cc_566 N_A_634_159#_M1029_g N_VPWR_c_1227_n 0.0057281f $X=3.245 $Y=2.275 $X2=0
+ $Y2=0
cc_567 N_A_634_159#_c_713_n N_VPWR_c_1227_n 0.0237f $X=4.075 $Y=2.135 $X2=0
+ $Y2=0
cc_568 N_A_634_159#_M1029_g N_VPWR_c_1234_n 0.00378797f $X=3.245 $Y=2.275 $X2=0
+ $Y2=0
cc_569 N_A_634_159#_c_723_n N_VPWR_c_1236_n 0.015079f $X=4.115 $Y=2.3 $X2=0
+ $Y2=0
cc_570 N_A_634_159#_M1008_d N_VPWR_c_1224_n 0.00285154f $X=3.98 $Y=1.735 $X2=0
+ $Y2=0
cc_571 N_A_634_159#_M1029_g N_VPWR_c_1224_n 0.00604354f $X=3.245 $Y=2.275 $X2=0
+ $Y2=0
cc_572 N_A_634_159#_c_723_n N_VPWR_c_1224_n 0.00439826f $X=4.115 $Y=2.3 $X2=0
+ $Y2=0
cc_573 N_A_634_159#_c_710_n N_VGND_M1026_d 0.00278876f $X=3.95 $Y=0.915 $X2=0
+ $Y2=0
cc_574 N_A_634_159#_M1026_g N_VGND_c_1485_n 0.0129352f $X=3.38 $Y=0.445 $X2=0
+ $Y2=0
cc_575 N_A_634_159#_c_733_n N_VGND_c_1485_n 0.00357337f $X=4.035 $Y=0.765 $X2=0
+ $Y2=0
cc_576 N_A_634_159#_c_711_n N_VGND_c_1485_n 0.0262751f $X=3.49 $Y=0.93 $X2=0
+ $Y2=0
cc_577 N_A_634_159#_c_750_p N_VGND_c_1485_n 0.0128408f $X=4.19 $Y=0.45 $X2=0
+ $Y2=0
cc_578 N_A_634_159#_c_714_n N_VGND_c_1485_n 4.63364e-19 $X=3.38 $Y=0.93 $X2=0
+ $Y2=0
cc_579 N_A_634_159#_c_750_p N_VGND_c_1492_n 0.0139094f $X=4.19 $Y=0.45 $X2=0
+ $Y2=0
cc_580 N_A_634_159#_M1026_g N_VGND_c_1500_n 0.00368966f $X=3.38 $Y=0.445 $X2=0
+ $Y2=0
cc_581 N_A_634_159#_M1013_d N_VGND_c_1507_n 0.00472956f $X=4.05 $Y=0.235 $X2=0
+ $Y2=0
cc_582 N_A_634_159#_M1026_g N_VGND_c_1507_n 0.0036978f $X=3.38 $Y=0.445 $X2=0
+ $Y2=0
cc_583 N_A_634_159#_c_710_n N_VGND_c_1507_n 0.00660235f $X=3.95 $Y=0.915 $X2=0
+ $Y2=0
cc_584 N_A_634_159#_c_711_n N_VGND_c_1507_n 0.00500137f $X=3.49 $Y=0.93 $X2=0
+ $Y2=0
cc_585 N_A_634_159#_c_750_p N_VGND_c_1507_n 0.0135555f $X=4.19 $Y=0.45 $X2=0
+ $Y2=0
cc_586 N_A_634_159#_c_714_n N_VGND_c_1507_n 0.00313291f $X=3.38 $Y=0.93 $X2=0
+ $Y2=0
cc_587 N_A_466_413#_c_818_n N_VPWR_M1029_d 0.00236303f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_588 N_A_466_413#_c_810_n N_VPWR_M1029_d 0.00412006f $X=3.355 $Y=2.19 $X2=0
+ $Y2=0
cc_589 N_A_466_413#_M1008_g N_VPWR_c_1227_n 0.00314007f $X=3.905 $Y=2.11 $X2=0
+ $Y2=0
cc_590 N_A_466_413#_c_801_n N_VPWR_c_1227_n 9.53331e-19 $X=3.83 $Y=1.41 $X2=0
+ $Y2=0
cc_591 N_A_466_413#_c_818_n N_VPWR_c_1227_n 0.0138309f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_592 N_A_466_413#_c_810_n N_VPWR_c_1227_n 0.0253561f $X=3.355 $Y=2.19 $X2=0
+ $Y2=0
cc_593 N_A_466_413#_c_804_n N_VPWR_c_1227_n 0.00781216f $X=3.355 $Y=1.41 $X2=0
+ $Y2=0
cc_594 N_A_466_413#_c_818_n N_VPWR_c_1234_n 0.0373829f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_595 N_A_466_413#_M1008_g N_VPWR_c_1236_n 0.00541359f $X=3.905 $Y=2.11 $X2=0
+ $Y2=0
cc_596 N_A_466_413#_M1012_d N_VPWR_c_1224_n 0.00227638f $X=2.33 $Y=2.065 $X2=0
+ $Y2=0
cc_597 N_A_466_413#_M1008_g N_VPWR_c_1224_n 0.00665748f $X=3.905 $Y=2.11 $X2=0
+ $Y2=0
cc_598 N_A_466_413#_c_818_n N_VPWR_c_1224_n 0.0167486f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_599 N_A_466_413#_c_824_n N_A_381_47#_c_1387_n 0.0125066f $X=2.91 $Y=0.45
+ $X2=0 $Y2=0
cc_600 N_A_466_413#_c_818_n A_561_413# 0.00531349f $X=3.27 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_601 N_A_466_413#_c_799_n N_VGND_c_1485_n 0.00803085f $X=3.94 $Y=0.95 $X2=0
+ $Y2=0
cc_602 N_A_466_413#_c_824_n N_VGND_c_1485_n 0.00869847f $X=2.91 $Y=0.45 $X2=0
+ $Y2=0
cc_603 N_A_466_413#_c_803_n N_VGND_c_1485_n 0.00226819f $X=2.995 $Y=1.315 $X2=0
+ $Y2=0
cc_604 N_A_466_413#_c_799_n N_VGND_c_1492_n 0.00448335f $X=3.94 $Y=0.95 $X2=0
+ $Y2=0
cc_605 N_A_466_413#_c_824_n N_VGND_c_1500_n 0.0225252f $X=2.91 $Y=0.45 $X2=0
+ $Y2=0
cc_606 N_A_466_413#_M1009_d N_VGND_c_1507_n 0.00293225f $X=2.465 $Y=0.235 $X2=0
+ $Y2=0
cc_607 N_A_466_413#_c_799_n N_VGND_c_1507_n 0.00626226f $X=3.94 $Y=0.95 $X2=0
+ $Y2=0
cc_608 N_A_466_413#_c_824_n N_VGND_c_1507_n 0.0226537f $X=2.91 $Y=0.45 $X2=0
+ $Y2=0
cc_609 N_A_466_413#_c_824_n A_592_47# 0.00271159f $X=2.91 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_610 N_A_466_413#_c_803_n A_592_47# 0.00138779f $X=2.995 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_611 N_A_1059_315#_M1014_g N_A_891_413#_M1025_g 0.0225645f $X=6.845 $Y=1.985
+ $X2=0 $Y2=0
cc_612 N_A_1059_315#_c_943_n N_A_891_413#_M1025_g 0.00606984f $X=6.205 $Y=2.34
+ $X2=0 $Y2=0
cc_613 N_A_1059_315#_c_944_n N_A_891_413#_M1025_g 0.0063384f $X=6.285 $Y=1.53
+ $X2=0 $Y2=0
cc_614 N_A_1059_315#_c_946_n N_A_891_413#_M1025_g 0.00459024f $X=6.205 $Y=1.63
+ $X2=0 $Y2=0
cc_615 N_A_1059_315#_c_919_n N_A_891_413#_c_1065_n 0.0221845f $X=6.855 $Y=0.995
+ $X2=0 $Y2=0
cc_616 N_A_1059_315#_c_927_n N_A_891_413#_c_1065_n 0.00404044f $X=6.225 $Y=0.385
+ $X2=0 $Y2=0
cc_617 N_A_1059_315#_c_928_n N_A_891_413#_c_1065_n 0.00496831f $X=6.29 $Y=0.995
+ $X2=0 $Y2=0
cc_618 N_A_1059_315#_c_930_n N_A_891_413#_c_1065_n 0.00262595f $X=6.225 $Y=0.825
+ $X2=0 $Y2=0
cc_619 N_A_1059_315#_M1011_g N_A_891_413#_c_1066_n 0.0181721f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_620 N_A_1059_315#_c_941_n N_A_891_413#_c_1066_n 0.00569718f $X=6.04 $Y=1.717
+ $X2=0 $Y2=0
cc_621 N_A_1059_315#_c_946_n N_A_891_413#_c_1066_n 0.00641947f $X=6.205 $Y=1.63
+ $X2=0 $Y2=0
cc_622 N_A_1059_315#_c_930_n N_A_891_413#_c_1066_n 0.00551597f $X=6.225 $Y=0.825
+ $X2=0 $Y2=0
cc_623 N_A_1059_315#_c_964_p N_A_891_413#_c_1066_n 0.0172129f $X=6.29 $Y=1.16
+ $X2=0 $Y2=0
cc_624 N_A_1059_315#_c_922_n N_A_891_413#_c_1067_n 0.0216197f $X=7.35 $Y=1.16
+ $X2=0 $Y2=0
cc_625 N_A_1059_315#_c_929_n N_A_891_413#_c_1067_n 0.0179674f $X=6.855 $Y=1.16
+ $X2=0 $Y2=0
cc_626 N_A_1059_315#_c_964_p N_A_891_413#_c_1067_n 0.00199985f $X=6.29 $Y=1.16
+ $X2=0 $Y2=0
cc_627 N_A_1059_315#_M1007_g N_A_891_413#_c_1076_n 0.00464573f $X=5.37 $Y=2.275
+ $X2=0 $Y2=0
cc_628 N_A_1059_315#_M1011_g N_A_891_413#_c_1079_n 0.00166852f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_629 N_A_1059_315#_M1011_g N_A_891_413#_c_1068_n 0.00941184f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_630 N_A_1059_315#_M1007_g N_A_891_413#_c_1074_n 0.0120276f $X=5.37 $Y=2.275
+ $X2=0 $Y2=0
cc_631 N_A_1059_315#_M1011_g N_A_891_413#_c_1074_n 0.00751613f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_632 N_A_1059_315#_c_941_n N_A_891_413#_c_1074_n 0.0282204f $X=6.04 $Y=1.717
+ $X2=0 $Y2=0
cc_633 N_A_1059_315#_c_942_n N_A_891_413#_c_1074_n 0.0079118f $X=5.565 $Y=1.74
+ $X2=0 $Y2=0
cc_634 N_A_1059_315#_M1011_g N_A_891_413#_c_1069_n 0.0232255f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_635 N_A_1059_315#_c_941_n N_A_891_413#_c_1069_n 0.0382059f $X=6.04 $Y=1.717
+ $X2=0 $Y2=0
cc_636 N_A_1059_315#_c_942_n N_A_891_413#_c_1069_n 0.00495398f $X=5.565 $Y=1.74
+ $X2=0 $Y2=0
cc_637 N_A_1059_315#_c_964_p N_A_891_413#_c_1069_n 0.0277655f $X=6.29 $Y=1.16
+ $X2=0 $Y2=0
cc_638 N_A_1059_315#_c_923_n N_A_1589_47#_c_1147_n 0.00368095f $X=8.235 $Y=0.995
+ $X2=0 $Y2=0
cc_639 N_A_1059_315#_c_924_n N_A_1589_47#_c_1147_n 0.0134165f $X=8.257 $Y=0.73
+ $X2=0 $Y2=0
cc_640 N_A_1059_315#_c_939_n N_A_1589_47#_M1027_g 0.0049186f $X=8.257 $Y=1.515
+ $X2=0 $Y2=0
cc_641 N_A_1059_315#_c_940_n N_A_1589_47#_M1027_g 0.0185375f $X=8.257 $Y=1.665
+ $X2=0 $Y2=0
cc_642 N_A_1059_315#_c_921_n N_A_1589_47#_c_1155_n 0.0020767f $X=8.16 $Y=1.16
+ $X2=0 $Y2=0
cc_643 N_A_1059_315#_M1010_g N_A_1589_47#_c_1155_n 0.00442235f $X=8.28 $Y=2.165
+ $X2=0 $Y2=0
cc_644 N_A_1059_315#_M1010_g N_A_1589_47#_c_1156_n 0.00647197f $X=8.28 $Y=2.165
+ $X2=0 $Y2=0
cc_645 N_A_1059_315#_c_920_n N_A_1589_47#_c_1149_n 0.0061678f $X=7.275 $Y=0.995
+ $X2=0 $Y2=0
cc_646 N_A_1059_315#_c_923_n N_A_1589_47#_c_1149_n 0.00509387f $X=8.235 $Y=0.995
+ $X2=0 $Y2=0
cc_647 N_A_1059_315#_c_924_n N_A_1589_47#_c_1149_n 0.00172506f $X=8.257 $Y=0.73
+ $X2=0 $Y2=0
cc_648 N_A_1059_315#_c_925_n N_A_1589_47#_c_1149_n 0.00370254f $X=8.257 $Y=0.85
+ $X2=0 $Y2=0
cc_649 N_A_1059_315#_c_925_n N_A_1589_47#_c_1150_n 0.00139755f $X=8.257 $Y=0.85
+ $X2=0 $Y2=0
cc_650 N_A_1059_315#_c_926_n N_A_1589_47#_c_1150_n 0.0123637f $X=8.235 $Y=1.16
+ $X2=0 $Y2=0
cc_651 N_A_1059_315#_c_940_n N_A_1589_47#_c_1150_n 0.00131663f $X=8.257 $Y=1.665
+ $X2=0 $Y2=0
cc_652 N_A_1059_315#_c_921_n N_A_1589_47#_c_1151_n 0.00186938f $X=8.16 $Y=1.16
+ $X2=0 $Y2=0
cc_653 N_A_1059_315#_M1019_g N_A_1589_47#_c_1158_n 0.00642633f $X=7.265 $Y=1.985
+ $X2=0 $Y2=0
cc_654 N_A_1059_315#_M1010_g N_A_1589_47#_c_1158_n 0.00145003f $X=8.28 $Y=2.165
+ $X2=0 $Y2=0
cc_655 N_A_1059_315#_c_939_n N_A_1589_47#_c_1158_n 0.00761479f $X=8.257 $Y=1.515
+ $X2=0 $Y2=0
cc_656 N_A_1059_315#_c_940_n N_A_1589_47#_c_1158_n 0.00617157f $X=8.257 $Y=1.665
+ $X2=0 $Y2=0
cc_657 N_A_1059_315#_c_921_n N_A_1589_47#_c_1179_n 0.0211857f $X=8.16 $Y=1.16
+ $X2=0 $Y2=0
cc_658 N_A_1059_315#_c_926_n N_A_1589_47#_c_1179_n 0.00575075f $X=8.235 $Y=1.16
+ $X2=0 $Y2=0
cc_659 N_A_1059_315#_c_926_n N_A_1589_47#_c_1152_n 0.0216214f $X=8.235 $Y=1.16
+ $X2=0 $Y2=0
cc_660 N_A_1059_315#_M1007_g N_VPWR_c_1228_n 0.00460353f $X=5.37 $Y=2.275 $X2=0
+ $Y2=0
cc_661 N_A_1059_315#_c_941_n N_VPWR_c_1228_n 0.0197488f $X=6.04 $Y=1.717 $X2=0
+ $Y2=0
cc_662 N_A_1059_315#_c_942_n N_VPWR_c_1228_n 0.00491995f $X=5.565 $Y=1.74 $X2=0
+ $Y2=0
cc_663 N_A_1059_315#_c_943_n N_VPWR_c_1228_n 0.0218928f $X=6.205 $Y=2.34 $X2=0
+ $Y2=0
cc_664 N_A_1059_315#_M1014_g N_VPWR_c_1229_n 0.00191466f $X=6.845 $Y=1.985 $X2=0
+ $Y2=0
cc_665 N_A_1059_315#_c_929_n N_VPWR_c_1229_n 0.00933114f $X=6.855 $Y=1.16 $X2=0
+ $Y2=0
cc_666 N_A_1059_315#_M1019_g N_VPWR_c_1230_n 0.00440592f $X=7.265 $Y=1.985 $X2=0
+ $Y2=0
cc_667 N_A_1059_315#_c_921_n N_VPWR_c_1230_n 0.00472325f $X=8.16 $Y=1.16 $X2=0
+ $Y2=0
cc_668 N_A_1059_315#_M1010_g N_VPWR_c_1230_n 0.00348891f $X=8.28 $Y=2.165 $X2=0
+ $Y2=0
cc_669 N_A_1059_315#_c_940_n N_VPWR_c_1231_n 0.011094f $X=8.257 $Y=1.665 $X2=0
+ $Y2=0
cc_670 N_A_1059_315#_M1007_g N_VPWR_c_1236_n 0.00565184f $X=5.37 $Y=2.275 $X2=0
+ $Y2=0
cc_671 N_A_1059_315#_c_943_n N_VPWR_c_1238_n 0.0217414f $X=6.205 $Y=2.34 $X2=0
+ $Y2=0
cc_672 N_A_1059_315#_M1014_g N_VPWR_c_1240_n 0.00543148f $X=6.845 $Y=1.985 $X2=0
+ $Y2=0
cc_673 N_A_1059_315#_M1019_g N_VPWR_c_1240_n 0.00543148f $X=7.265 $Y=1.985 $X2=0
+ $Y2=0
cc_674 N_A_1059_315#_M1010_g N_VPWR_c_1244_n 0.00542163f $X=8.28 $Y=2.165 $X2=0
+ $Y2=0
cc_675 N_A_1059_315#_M1025_s N_VPWR_c_1224_n 0.00217517f $X=6.08 $Y=1.485 $X2=0
+ $Y2=0
cc_676 N_A_1059_315#_M1007_g N_VPWR_c_1224_n 0.0117476f $X=5.37 $Y=2.275 $X2=0
+ $Y2=0
cc_677 N_A_1059_315#_M1014_g N_VPWR_c_1224_n 0.00960872f $X=6.845 $Y=1.985 $X2=0
+ $Y2=0
cc_678 N_A_1059_315#_M1019_g N_VPWR_c_1224_n 0.0109575f $X=7.265 $Y=1.985 $X2=0
+ $Y2=0
cc_679 N_A_1059_315#_M1010_g N_VPWR_c_1224_n 0.0111401f $X=8.28 $Y=2.165 $X2=0
+ $Y2=0
cc_680 N_A_1059_315#_c_941_n N_VPWR_c_1224_n 0.0104129f $X=6.04 $Y=1.717 $X2=0
+ $Y2=0
cc_681 N_A_1059_315#_c_942_n N_VPWR_c_1224_n 0.00115082f $X=5.565 $Y=1.74 $X2=0
+ $Y2=0
cc_682 N_A_1059_315#_c_943_n N_VPWR_c_1224_n 0.0128119f $X=6.205 $Y=2.34 $X2=0
+ $Y2=0
cc_683 N_A_1059_315#_M1014_g N_Q_c_1427_n 0.00943952f $X=6.845 $Y=1.985 $X2=0
+ $Y2=0
cc_684 N_A_1059_315#_M1019_g N_Q_c_1427_n 0.0142922f $X=7.265 $Y=1.985 $X2=0
+ $Y2=0
cc_685 N_A_1059_315#_c_946_n N_Q_c_1427_n 0.00160682f $X=6.205 $Y=1.63 $X2=0
+ $Y2=0
cc_686 N_A_1059_315#_M1014_g N_Q_c_1425_n 0.00535654f $X=6.845 $Y=1.985 $X2=0
+ $Y2=0
cc_687 N_A_1059_315#_c_919_n N_Q_c_1425_n 0.00261585f $X=6.855 $Y=0.995 $X2=0
+ $Y2=0
cc_688 N_A_1059_315#_M1019_g N_Q_c_1425_n 0.0119523f $X=7.265 $Y=1.985 $X2=0
+ $Y2=0
cc_689 N_A_1059_315#_c_920_n N_Q_c_1425_n 0.00411499f $X=7.275 $Y=0.995 $X2=0
+ $Y2=0
cc_690 N_A_1059_315#_c_922_n N_Q_c_1425_n 0.0225134f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_691 N_A_1059_315#_c_944_n N_Q_c_1425_n 0.00103347f $X=6.285 $Y=1.53 $X2=0
+ $Y2=0
cc_692 N_A_1059_315#_c_929_n N_Q_c_1425_n 0.0282849f $X=6.855 $Y=1.16 $X2=0
+ $Y2=0
cc_693 N_A_1059_315#_c_946_n N_Q_c_1425_n 0.00148631f $X=6.205 $Y=1.63 $X2=0
+ $Y2=0
cc_694 N_A_1059_315#_c_919_n N_Q_c_1438_n 0.00188476f $X=6.855 $Y=0.995 $X2=0
+ $Y2=0
cc_695 N_A_1059_315#_c_920_n N_Q_c_1438_n 0.00522811f $X=7.275 $Y=0.995 $X2=0
+ $Y2=0
cc_696 N_A_1059_315#_c_922_n N_Q_c_1438_n 0.00273743f $X=7.35 $Y=1.16 $X2=0
+ $Y2=0
cc_697 N_A_1059_315#_c_928_n N_Q_c_1438_n 9.78692e-19 $X=6.29 $Y=0.995 $X2=0
+ $Y2=0
cc_698 N_A_1059_315#_c_929_n N_Q_c_1438_n 0.00268244f $X=6.855 $Y=1.16 $X2=0
+ $Y2=0
cc_699 N_A_1059_315#_c_930_n N_Q_c_1438_n 0.00264475f $X=6.225 $Y=0.825 $X2=0
+ $Y2=0
cc_700 N_A_1059_315#_c_919_n N_Q_c_1444_n 0.00513559f $X=6.855 $Y=0.995 $X2=0
+ $Y2=0
cc_701 N_A_1059_315#_c_920_n N_Q_c_1444_n 0.00931238f $X=7.275 $Y=0.995 $X2=0
+ $Y2=0
cc_702 N_A_1059_315#_c_930_n N_Q_c_1444_n 0.00136135f $X=6.225 $Y=0.825 $X2=0
+ $Y2=0
cc_703 N_A_1059_315#_M1011_g N_VGND_c_1486_n 0.00502953f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_704 N_A_1059_315#_c_927_n N_VGND_c_1486_n 0.0181463f $X=6.225 $Y=0.385 $X2=0
+ $Y2=0
cc_705 N_A_1059_315#_c_919_n N_VGND_c_1487_n 0.00187348f $X=6.855 $Y=0.995 $X2=0
+ $Y2=0
cc_706 N_A_1059_315#_c_929_n N_VGND_c_1487_n 0.00929281f $X=6.855 $Y=1.16 $X2=0
+ $Y2=0
cc_707 N_A_1059_315#_c_920_n N_VGND_c_1488_n 0.00324666f $X=7.275 $Y=0.995 $X2=0
+ $Y2=0
cc_708 N_A_1059_315#_c_921_n N_VGND_c_1488_n 0.0044893f $X=8.16 $Y=1.16 $X2=0
+ $Y2=0
cc_709 N_A_1059_315#_c_924_n N_VGND_c_1488_n 0.00397682f $X=8.257 $Y=0.73 $X2=0
+ $Y2=0
cc_710 N_A_1059_315#_c_924_n N_VGND_c_1489_n 0.0068429f $X=8.257 $Y=0.73 $X2=0
+ $Y2=0
cc_711 N_A_1059_315#_M1011_g N_VGND_c_1492_n 0.00585385f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_712 N_A_1059_315#_c_927_n N_VGND_c_1494_n 0.016209f $X=6.225 $Y=0.385 $X2=0
+ $Y2=0
cc_713 N_A_1059_315#_c_919_n N_VGND_c_1496_n 0.00543342f $X=6.855 $Y=0.995 $X2=0
+ $Y2=0
cc_714 N_A_1059_315#_c_920_n N_VGND_c_1496_n 0.00475376f $X=7.275 $Y=0.995 $X2=0
+ $Y2=0
cc_715 N_A_1059_315#_c_924_n N_VGND_c_1501_n 0.00585385f $X=8.257 $Y=0.73 $X2=0
+ $Y2=0
cc_716 N_A_1059_315#_c_925_n N_VGND_c_1501_n 8.48802e-19 $X=8.257 $Y=0.85 $X2=0
+ $Y2=0
cc_717 N_A_1059_315#_M1015_s N_VGND_c_1507_n 0.00212021f $X=6.1 $Y=0.235 $X2=0
+ $Y2=0
cc_718 N_A_1059_315#_M1011_g N_VGND_c_1507_n 0.0121657f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_719 N_A_1059_315#_c_919_n N_VGND_c_1507_n 0.00960932f $X=6.855 $Y=0.995 $X2=0
+ $Y2=0
cc_720 N_A_1059_315#_c_920_n N_VGND_c_1507_n 0.00868278f $X=7.275 $Y=0.995 $X2=0
+ $Y2=0
cc_721 N_A_1059_315#_c_924_n N_VGND_c_1507_n 0.0122138f $X=8.257 $Y=0.73 $X2=0
+ $Y2=0
cc_722 N_A_1059_315#_c_925_n N_VGND_c_1507_n 0.00111161f $X=8.257 $Y=0.85 $X2=0
+ $Y2=0
cc_723 N_A_1059_315#_c_927_n N_VGND_c_1507_n 0.012105f $X=6.225 $Y=0.385 $X2=0
+ $Y2=0
cc_724 N_A_891_413#_M1025_g N_VPWR_c_1228_n 0.00213308f $X=6.425 $Y=1.985 $X2=0
+ $Y2=0
cc_725 N_A_891_413#_M1025_g N_VPWR_c_1229_n 0.00313741f $X=6.425 $Y=1.985 $X2=0
+ $Y2=0
cc_726 N_A_891_413#_c_1076_n N_VPWR_c_1236_n 0.0273429f $X=5.14 $Y=2.25 $X2=0
+ $Y2=0
cc_727 N_A_891_413#_M1025_g N_VPWR_c_1238_n 0.00541359f $X=6.425 $Y=1.985 $X2=0
+ $Y2=0
cc_728 N_A_891_413#_M1024_d N_VPWR_c_1224_n 0.00219484f $X=4.455 $Y=2.065 $X2=0
+ $Y2=0
cc_729 N_A_891_413#_M1025_g N_VPWR_c_1224_n 0.0109315f $X=6.425 $Y=1.985 $X2=0
+ $Y2=0
cc_730 N_A_891_413#_c_1076_n N_VPWR_c_1224_n 0.0275904f $X=5.14 $Y=2.25 $X2=0
+ $Y2=0
cc_731 N_A_891_413#_c_1076_n A_975_413# 0.00900936f $X=5.14 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_732 N_A_891_413#_c_1074_n A_975_413# 0.00123507f $X=5.225 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_733 N_A_891_413#_M1025_g N_Q_c_1427_n 3.15835e-19 $X=6.425 $Y=1.985 $X2=0
+ $Y2=0
cc_734 N_A_891_413#_M1025_g N_Q_c_1425_n 2.34774e-19 $X=6.425 $Y=1.985 $X2=0
+ $Y2=0
cc_735 N_A_891_413#_c_1065_n N_Q_c_1438_n 2.4955e-19 $X=6.435 $Y=0.995 $X2=0
+ $Y2=0
cc_736 N_A_891_413#_c_1065_n N_VGND_c_1486_n 0.00253884f $X=6.435 $Y=0.995 $X2=0
+ $Y2=0
cc_737 N_A_891_413#_c_1069_n N_VGND_c_1486_n 0.00938141f $X=5.935 $Y=1.16 $X2=0
+ $Y2=0
cc_738 N_A_891_413#_c_1065_n N_VGND_c_1487_n 0.00309623f $X=6.435 $Y=0.995 $X2=0
+ $Y2=0
cc_739 N_A_891_413#_c_1079_n N_VGND_c_1492_n 0.0268923f $X=5.14 $Y=0.45 $X2=0
+ $Y2=0
cc_740 N_A_891_413#_c_1065_n N_VGND_c_1494_n 0.00543148f $X=6.435 $Y=0.995 $X2=0
+ $Y2=0
cc_741 N_A_891_413#_M1031_d N_VGND_c_1507_n 0.00322972f $X=4.555 $Y=0.235 $X2=0
+ $Y2=0
cc_742 N_A_891_413#_c_1065_n N_VGND_c_1507_n 0.0109348f $X=6.435 $Y=0.995 $X2=0
+ $Y2=0
cc_743 N_A_891_413#_c_1079_n N_VGND_c_1507_n 0.0266007f $X=5.14 $Y=0.45 $X2=0
+ $Y2=0
cc_744 N_A_891_413#_c_1079_n A_1017_47# 0.00423935f $X=5.14 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_745 N_A_891_413#_c_1068_n A_1017_47# 0.00152168f $X=5.225 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_746 N_A_1589_47#_c_1155_n N_VPWR_c_1230_n 0.0345488f $X=8.07 $Y=1.88 $X2=0
+ $Y2=0
cc_747 N_A_1589_47#_M1027_g N_VPWR_c_1231_n 0.00159535f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_748 N_A_1589_47#_c_1150_n N_VPWR_c_1231_n 0.0177138f $X=8.675 $Y=1.16 $X2=0
+ $Y2=0
cc_749 N_A_1589_47#_c_1158_n N_VPWR_c_1231_n 0.0656425f $X=8.07 $Y=1.715 $X2=0
+ $Y2=0
cc_750 N_A_1589_47#_c_1152_n N_VPWR_c_1231_n 0.0027539f $X=9.185 $Y=1.16 $X2=0
+ $Y2=0
cc_751 N_A_1589_47#_M1030_g N_VPWR_c_1233_n 0.00318595f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_752 N_A_1589_47#_c_1156_n N_VPWR_c_1244_n 0.0186592f $X=8.07 $Y=2 $X2=0 $Y2=0
cc_753 N_A_1589_47#_M1027_g N_VPWR_c_1245_n 0.00541359f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_754 N_A_1589_47#_M1030_g N_VPWR_c_1245_n 0.00533769f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_755 N_A_1589_47#_M1010_s N_VPWR_c_1224_n 0.00210124f $X=7.945 $Y=1.845 $X2=0
+ $Y2=0
cc_756 N_A_1589_47#_M1027_g N_VPWR_c_1224_n 0.00968038f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_757 N_A_1589_47#_M1030_g N_VPWR_c_1224_n 0.0102881f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_758 N_A_1589_47#_c_1156_n N_VPWR_c_1224_n 0.0123045f $X=8.07 $Y=2 $X2=0 $Y2=0
cc_759 N_A_1589_47#_c_1149_n N_Q_c_1425_n 0.00333053f $X=8.065 $Y=0.995 $X2=0
+ $Y2=0
cc_760 N_A_1589_47#_c_1158_n N_Q_c_1425_n 0.00674652f $X=8.07 $Y=1.715 $X2=0
+ $Y2=0
cc_761 N_A_1589_47#_c_1179_n N_Q_c_1425_n 0.00808048f $X=8.1 $Y=1.16 $X2=0 $Y2=0
cc_762 N_A_1589_47#_c_1149_n N_Q_c_1438_n 0.00337456f $X=8.065 $Y=0.995 $X2=0
+ $Y2=0
cc_763 N_A_1589_47#_c_1151_n N_Q_c_1444_n 4.06938e-19 $X=8.07 $Y=0.51 $X2=0
+ $Y2=0
cc_764 N_A_1589_47#_c_1148_n N_Q_N_c_1466_n 0.00685312f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_765 N_A_1589_47#_c_1148_n N_Q_N_c_1463_n 0.00249693f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_766 N_A_1589_47#_M1027_g Q_N 0.0119052f $X=8.765 $Y=1.985 $X2=0 $Y2=0
cc_767 N_A_1589_47#_M1030_g Q_N 0.011267f $X=9.185 $Y=1.985 $X2=0 $Y2=0
cc_768 N_A_1589_47#_c_1147_n N_Q_N_c_1464_n 0.00258993f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_769 N_A_1589_47#_M1027_g N_Q_N_c_1464_n 0.00397766f $X=8.765 $Y=1.985 $X2=0
+ $Y2=0
cc_770 N_A_1589_47#_c_1148_n N_Q_N_c_1464_n 0.00482599f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_771 N_A_1589_47#_M1030_g N_Q_N_c_1464_n 0.00833812f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_772 N_A_1589_47#_c_1150_n N_Q_N_c_1464_n 0.0253962f $X=8.675 $Y=1.16 $X2=0
+ $Y2=0
cc_773 N_A_1589_47#_c_1152_n N_Q_N_c_1464_n 0.0282677f $X=9.185 $Y=1.16 $X2=0
+ $Y2=0
cc_774 N_A_1589_47#_c_1151_n N_VGND_c_1488_n 0.0120291f $X=8.07 $Y=0.51 $X2=0
+ $Y2=0
cc_775 N_A_1589_47#_c_1147_n N_VGND_c_1489_n 0.0106876f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_776 N_A_1589_47#_c_1148_n N_VGND_c_1489_n 7.94611e-19 $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_777 N_A_1589_47#_c_1149_n N_VGND_c_1489_n 0.0107592f $X=8.065 $Y=0.995 $X2=0
+ $Y2=0
cc_778 N_A_1589_47#_c_1150_n N_VGND_c_1489_n 0.0250055f $X=8.675 $Y=1.16 $X2=0
+ $Y2=0
cc_779 N_A_1589_47#_c_1152_n N_VGND_c_1489_n 0.00378658f $X=9.185 $Y=1.16 $X2=0
+ $Y2=0
cc_780 N_A_1589_47#_c_1148_n N_VGND_c_1491_n 0.00353346f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_781 N_A_1589_47#_c_1151_n N_VGND_c_1501_n 0.0109932f $X=8.07 $Y=0.51 $X2=0
+ $Y2=0
cc_782 N_A_1589_47#_c_1147_n N_VGND_c_1502_n 0.0046653f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_783 N_A_1589_47#_c_1148_n N_VGND_c_1502_n 0.00534242f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_784 N_A_1589_47#_M1002_s N_VGND_c_1507_n 0.00261104f $X=7.945 $Y=0.235 $X2=0
+ $Y2=0
cc_785 N_A_1589_47#_c_1147_n N_VGND_c_1507_n 0.00796766f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_786 N_A_1589_47#_c_1148_n N_VGND_c_1507_n 0.0103275f $X=9.185 $Y=0.995 $X2=0
+ $Y2=0
cc_787 N_A_1589_47#_c_1151_n N_VGND_c_1507_n 0.00940719f $X=8.07 $Y=0.51 $X2=0
+ $Y2=0
cc_788 N_VPWR_c_1224_n N_A_381_47#_M1023_d 0.00223112f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_789 N_VPWR_c_1234_n N_A_381_47#_c_1373_n 0.0151865f $X=3.61 $Y=2.72 $X2=0
+ $Y2=0
cc_790 N_VPWR_c_1224_n N_A_381_47#_c_1373_n 0.00442027f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_791 N_VPWR_c_1234_n N_A_381_47#_c_1375_n 8.77274e-19 $X=3.61 $Y=2.72 $X2=0
+ $Y2=0
cc_792 N_VPWR_c_1224_n N_A_381_47#_c_1375_n 6.01352e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_793 N_VPWR_c_1224_n A_561_413# 0.00247673f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_794 N_VPWR_c_1224_n A_975_413# 0.00364366f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_795 N_VPWR_c_1224_n N_Q_M1014_s 0.00217997f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_796 N_VPWR_c_1240_n N_Q_c_1427_n 0.0147046f $X=7.39 $Y=2.72 $X2=0 $Y2=0
cc_797 N_VPWR_c_1224_n N_Q_c_1427_n 0.0119354f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_798 N_VPWR_c_1224_n N_Q_N_M1027_s 0.00215201f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_799 N_VPWR_c_1245_n Q_N 0.0192448f $X=9.315 $Y=2.72 $X2=0 $Y2=0
cc_800 N_VPWR_c_1224_n Q_N 0.0123914f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_801 N_VPWR_c_1233_n N_VGND_c_1491_n 0.00931063f $X=9.4 $Y=1.66 $X2=0 $Y2=0
cc_802 N_A_381_47#_c_1371_n N_VGND_c_1500_n 8.86929e-19 $X=1.932 $Y=0.805 $X2=0
+ $Y2=0
cc_803 N_A_381_47#_c_1387_n N_VGND_c_1500_n 0.0115184f $X=2.045 $Y=0.45 $X2=0
+ $Y2=0
cc_804 N_A_381_47#_M1006_d N_VGND_c_1507_n 0.00412945f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_805 N_A_381_47#_c_1371_n N_VGND_c_1507_n 0.00130006f $X=1.932 $Y=0.805 $X2=0
+ $Y2=0
cc_806 N_A_381_47#_c_1387_n N_VGND_c_1507_n 0.0114633f $X=2.045 $Y=0.45 $X2=0
+ $Y2=0
cc_807 N_Q_c_1438_n N_VGND_c_1496_n 0.00100112f $X=7.065 $Y=0.74 $X2=0 $Y2=0
cc_808 N_Q_c_1444_n N_VGND_c_1496_n 0.0142147f $X=7.065 $Y=0.395 $X2=0 $Y2=0
cc_809 N_Q_M1021_s N_VGND_c_1507_n 0.00218509f $X=6.93 $Y=0.235 $X2=0 $Y2=0
cc_810 N_Q_c_1438_n N_VGND_c_1507_n 0.00158918f $X=7.065 $Y=0.74 $X2=0 $Y2=0
cc_811 N_Q_c_1444_n N_VGND_c_1507_n 0.0118437f $X=7.065 $Y=0.395 $X2=0 $Y2=0
cc_812 N_Q_N_c_1466_n N_VGND_c_1491_n 0.0237522f $X=8.975 $Y=0.57 $X2=0 $Y2=0
cc_813 N_Q_N_c_1466_n N_VGND_c_1502_n 0.0145794f $X=8.975 $Y=0.57 $X2=0 $Y2=0
cc_814 N_Q_N_M1003_s N_VGND_c_1507_n 0.0039413f $X=8.84 $Y=0.235 $X2=0 $Y2=0
cc_815 N_Q_N_c_1466_n N_VGND_c_1507_n 0.00953716f $X=8.975 $Y=0.57 $X2=0 $Y2=0
cc_816 N_VGND_c_1507_n A_592_47# 0.00749713f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_817 N_VGND_c_1507_n A_1017_47# 0.00618566f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24

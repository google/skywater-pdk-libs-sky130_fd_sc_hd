* NGSPICE file created from sky130_fd_sc_hd__a311o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_75_199# C1 a_544_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=4.15e+11p ps=2.83e+06u
M1001 VGND B1 a_75_199# VNB nshort w=650000u l=150000u
+  ad=4.94e+11p pd=4.12e+06u as=3.8025e+11p ps=3.77e+06u
M1002 VPWR A2 a_201_297# VPB phighvt w=1e+06u l=150000u
+  ad=8.95e+11p pd=5.79e+06u as=6.55e+11p ps=5.31e+06u
M1003 a_544_297# B1 a_201_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_75_199# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1005 a_315_47# A2 a_208_47# VNB nshort w=650000u l=150000u
+  ad=3.38e+11p pd=2.34e+06u as=2.5025e+11p ps=2.07e+06u
M1006 a_201_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_201_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_75_199# A1 a_315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_208_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_75_199# C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_75_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.765000 1.950000 1.015000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.039500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.040000 0.255000 6.460000 0.545000 ;
        RECT 6.040000 1.835000 7.300000 2.005000 ;
        RECT 6.040000 2.005000 6.370000 2.455000 ;
        RECT 6.290000 0.545000 6.460000 0.715000 ;
        RECT 6.290000 0.715000 7.300000 0.885000 ;
        RECT 6.585000 1.785000 7.300000 1.835000 ;
        RECT 6.750000 0.885000 7.300000 1.785000 ;
        RECT 6.970000 0.255000 7.300000 0.715000 ;
        RECT 6.970000 2.005000 7.300000 2.465000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.230000 1.055000 5.740000 1.325000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.090000 1.075000 0.380000 1.120000 ;
        RECT 0.090000 1.120000 5.460000 1.260000 ;
        RECT 0.090000 1.260000 0.380000 1.305000 ;
        RECT 5.170000 1.075000 5.460000 1.120000 ;
        RECT 5.170000 1.260000 5.460000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.450000  0.085000 1.785000 0.465000 ;
        RECT 3.315000  0.085000 3.650000 0.530000 ;
        RECT 4.295000  0.085000 4.580000 0.715000 ;
        RECT 5.590000  0.085000 5.870000 0.545000 ;
        RECT 6.630000  0.085000 6.800000 0.545000 ;
        RECT 7.470000  0.085000 7.735000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.450000 2.195000 1.815000 2.635000 ;
        RECT 3.335000 2.175000 3.695000 2.635000 ;
        RECT 4.295000 2.010000 4.580000 2.635000 ;
        RECT 5.575000 1.835000 5.840000 2.635000 ;
        RECT 6.540000 2.175000 6.800000 2.635000 ;
        RECT 7.470000 1.485000 7.735000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.345000 0.345000 0.635000 ;
      RECT 0.085000 0.635000 0.780000 0.805000 ;
      RECT 0.085000 1.795000 0.780000 1.965000 ;
      RECT 0.085000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.780000 1.070000 ;
      RECT 0.610000 1.070000 0.840000 1.400000 ;
      RECT 0.610000 1.400000 0.780000 1.795000 ;
      RECT 1.015000 0.345000 1.280000 1.355000 ;
      RECT 1.015000 1.355000 2.335000 1.585000 ;
      RECT 1.015000 1.585000 1.240000 2.465000 ;
      RECT 1.525000 1.785000 1.695000 1.855000 ;
      RECT 1.525000 1.855000 2.845000 1.905000 ;
      RECT 1.525000 1.905000 2.735000 2.025000 ;
      RECT 2.045000 1.585000 2.335000 1.685000 ;
      RECT 2.290000 0.705000 2.735000 1.035000 ;
      RECT 2.415000 0.365000 3.075000 0.535000 ;
      RECT 2.475000 2.195000 3.165000 2.425000 ;
      RECT 2.505000 1.575000 2.845000 1.855000 ;
      RECT 2.565000 1.035000 2.735000 1.575000 ;
      RECT 2.905000 0.535000 3.075000 0.995000 ;
      RECT 2.905000 0.995000 3.775000 1.165000 ;
      RECT 2.915000 2.060000 3.185000 2.090000 ;
      RECT 2.915000 2.090000 3.180000 2.105000 ;
      RECT 2.915000 2.105000 3.165000 2.195000 ;
      RECT 2.980000 2.015000 3.185000 2.060000 ;
      RECT 3.015000 1.165000 3.775000 1.325000 ;
      RECT 3.015000 1.325000 3.185000 2.015000 ;
      RECT 3.355000 1.535000 4.115000 1.865000 ;
      RECT 3.895000 0.415000 4.115000 0.745000 ;
      RECT 3.895000 1.865000 4.115000 2.435000 ;
      RECT 3.945000 0.745000 4.115000 0.995000 ;
      RECT 3.945000 0.995000 4.720000 1.325000 ;
      RECT 3.945000 1.325000 4.115000 1.535000 ;
      RECT 4.750000 0.290000 5.060000 0.715000 ;
      RECT 4.750000 0.715000 6.120000 0.825000 ;
      RECT 4.750000 1.495000 6.140000 1.665000 ;
      RECT 4.750000 1.665000 5.035000 2.465000 ;
      RECT 4.890000 0.825000 6.120000 0.885000 ;
      RECT 4.890000 0.885000 5.060000 1.495000 ;
      RECT 5.910000 0.885000 6.120000 1.055000 ;
      RECT 5.910000 1.055000 6.580000 1.290000 ;
      RECT 5.910000 1.290000 6.140000 1.495000 ;
    LAYER mcon ;
      RECT 0.610000 1.785000 0.780000 1.955000 ;
      RECT 1.525000 1.785000 1.695000 1.955000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 1.755000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.465000 1.755000 1.755000 1.800000 ;
      RECT 1.465000 1.940000 1.755000 1.985000 ;
  END
END sky130_fd_sc_hd__dlclkp_4
END LIBRARY

* File: sky130_fd_sc_hd__buf_12.pxi.spice
* Created: Tue Sep  1 18:58:54 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_12%A N_A_M1012_g N_A_M1004_g N_A_M1015_g N_A_M1008_g
+ N_A_M1018_g N_A_M1019_g N_A_c_138_n N_A_M1029_g N_A_M1027_g A A A A
+ PM_SKY130_FD_SC_HD__BUF_12%A
x_PM_SKY130_FD_SC_HD__BUF_12%A_109_47# N_A_109_47#_M1012_s N_A_109_47#_M1018_s
+ N_A_109_47#_M1004_d N_A_109_47#_M1019_d N_A_109_47#_M1000_g
+ N_A_109_47#_M1001_g N_A_109_47#_M1005_g N_A_109_47#_M1002_g
+ N_A_109_47#_M1007_g N_A_109_47#_M1003_g N_A_109_47#_M1016_g
+ N_A_109_47#_M1006_g N_A_109_47#_M1020_g N_A_109_47#_M1009_g
+ N_A_109_47#_M1021_g N_A_109_47#_M1010_g N_A_109_47#_M1023_g
+ N_A_109_47#_M1011_g N_A_109_47#_M1024_g N_A_109_47#_M1013_g
+ N_A_109_47#_M1025_g N_A_109_47#_M1014_g N_A_109_47#_M1026_g
+ N_A_109_47#_M1017_g N_A_109_47#_M1030_g N_A_109_47#_M1022_g
+ N_A_109_47#_M1031_g N_A_109_47#_M1028_g N_A_109_47#_c_266_n
+ N_A_109_47#_c_459_p N_A_109_47#_c_239_n N_A_109_47#_c_240_n
+ N_A_109_47#_c_260_n N_A_109_47#_c_261_n N_A_109_47#_c_284_n
+ N_A_109_47#_c_453_p N_A_109_47#_c_241_n N_A_109_47#_c_242_n
+ N_A_109_47#_c_243_n N_A_109_47#_c_244_n N_A_109_47#_c_263_n
+ N_A_109_47#_c_245_n N_A_109_47#_c_246_n N_A_109_47#_c_247_n
+ PM_SKY130_FD_SC_HD__BUF_12%A_109_47#
x_PM_SKY130_FD_SC_HD__BUF_12%VPWR N_VPWR_M1004_s N_VPWR_M1008_s N_VPWR_M1027_s
+ N_VPWR_M1002_s N_VPWR_M1006_s N_VPWR_M1010_s N_VPWR_M1013_s N_VPWR_M1017_s
+ N_VPWR_M1028_s N_VPWR_c_486_n N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n
+ N_VPWR_c_505_n VPWR VPWR N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_485_n
+ PM_SKY130_FD_SC_HD__BUF_12%VPWR
x_PM_SKY130_FD_SC_HD__BUF_12%X N_X_M1000_s N_X_M1007_s N_X_M1020_s N_X_M1023_s
+ N_X_M1025_s N_X_M1030_s N_X_M1001_d N_X_M1003_d N_X_M1009_d N_X_M1011_d
+ N_X_M1014_d N_X_M1022_d N_X_c_730_p N_X_c_695_n N_X_c_615_n N_X_c_616_n
+ N_X_c_622_n N_X_c_623_n N_X_c_733_p N_X_c_699_n N_X_c_617_n N_X_c_624_n
+ N_X_c_725_p N_X_c_703_n N_X_c_653_n N_X_c_654_n N_X_c_655_n N_X_c_656_n
+ N_X_c_657_n N_X_c_618_n N_X_c_625_n N_X_c_619_n N_X_c_626_n X N_X_c_672_n
+ N_X_c_621_n PM_SKY130_FD_SC_HD__BUF_12%X
x_PM_SKY130_FD_SC_HD__BUF_12%VGND N_VGND_M1012_d N_VGND_M1015_d N_VGND_M1029_d
+ N_VGND_M1005_d N_VGND_M1016_d N_VGND_M1021_d N_VGND_M1024_d N_VGND_M1026_d
+ N_VGND_M1031_d N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n
+ N_VGND_c_762_n N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n
+ N_VGND_c_767_n N_VGND_c_768_n N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n
+ N_VGND_c_772_n N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n VGND VGND
+ N_VGND_c_776_n VGND N_VGND_c_777_n N_VGND_c_778_n N_VGND_c_779_n
+ N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n N_VGND_c_784_n
+ VGND PM_SKY130_FD_SC_HD__BUF_12%VGND
cc_1 VNB N_A_M1012_g 0.0226823f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1015_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_A_M1008_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_4 VNB N_A_M1018_g 0.0170552f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_5 VNB N_A_M1019_g 4.49778e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_6 VNB N_A_c_138_n 0.0850733f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.025
cc_7 VNB N_A_M1029_g 0.0172396f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_A_M1027_g 4.62826e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=1.105
cc_10 VNB N_A_109_47#_M1000_g 0.0174794f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_11 VNB N_A_109_47#_M1001_g 4.62903e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_12 VNB N_A_109_47#_M1005_g 0.0170561f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_13 VNB N_A_109_47#_M1002_g 4.49847e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_14 VNB N_A_109_47#_M1007_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_15 VNB N_A_109_47#_M1003_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.105
cc_16 VNB N_A_109_47#_M1016_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_109_47#_M1006_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_18 VNB N_A_109_47#_M1020_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=1.405 $Y2=1.16
cc_19 VNB N_A_109_47#_M1009_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.175
cc_20 VNB N_A_109_47#_M1021_g 0.0170726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_109_47#_M1010_g 4.49522e-19 $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=1.175
cc_22 VNB N_A_109_47#_M1023_g 0.0165752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_109_47#_M1011_g 4.12504e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_109_47#_M1024_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_109_47#_M1013_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_109_47#_M1025_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_109_47#_M1014_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_109_47#_M1026_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_109_47#_M1017_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_109_47#_M1030_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_109_47#_M1022_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_109_47#_M1031_g 0.0233973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_109_47#_M1028_g 7.17859e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_109_47#_c_239_n 0.00308383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_109_47#_c_240_n 0.00149343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_109_47#_c_241_n 0.00104171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_109_47#_c_242_n 0.00305801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_109_47#_c_243_n 0.00102395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_109_47#_c_244_n 0.00274061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_109_47#_c_245_n 0.00127298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_109_47#_c_246_n 0.00134032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_109_47#_c_247_n 0.20655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VPWR_c_485_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_X_c_615_n 0.00308383f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_45 VNB N_X_c_616_n 0.00141134f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_46 VNB N_X_c_617_n 0.00308383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_X_c_618_n 0.00127314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_619_n 0.00127314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB X 0.00307662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_X_c_621_n 0.00160194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_758_n 0.0103086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_759_n 0.016957f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_53 VNB N_VGND_c_760_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.105
cc_54 VNB N_VGND_c_761_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_762_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_56 VNB N_VGND_c_763_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_57 VNB N_VGND_c_764_n 0.0112357f $X=-0.19 $Y=-0.24 $X2=1.405 $Y2=1.16
cc_58 VNB N_VGND_c_765_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_766_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.175
cc_60 VNB N_VGND_c_767_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_768_n 0.0141639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_769_n 0.00668519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_770_n 0.0112511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_771_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_772_n 0.0118636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_773_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_774_n 0.0112357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_775_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_776_n 0.0118636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_777_n 0.0112443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_778_n 0.0112541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_779_n 0.01186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_780_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_781_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_782_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_783_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_784_n 0.352987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VPB N_A_M1004_g 0.0274016f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_79 VPB N_A_M1008_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_80 VPB N_A_M1019_g 0.0191647f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_81 VPB N_A_c_138_n 0.00981082f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_82 VPB N_A_M1027_g 0.0194261f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_83 VPB N_A_109_47#_M1001_g 0.0198358f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_84 VPB N_A_109_47#_M1002_g 0.0189386f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_85 VPB N_A_109_47#_M1003_g 0.0189613f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.105
cc_86 VPB N_A_109_47#_M1006_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_87 VPB N_A_109_47#_M1009_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.175
cc_88 VPB N_A_109_47#_M1010_g 0.0189544f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.175
cc_89 VPB N_A_109_47#_M1011_g 0.0183706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_109_47#_M1013_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_109_47#_M1014_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_109_47#_M1017_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_109_47#_M1022_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_109_47#_M1028_g 0.0266676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_109_47#_c_260_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_109_47#_c_261_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_109_47#_c_243_n 0.00306481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_109_47#_c_263_n 0.00345546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_486_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_487_n 0.00416524f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_101 VPB N_VPWR_c_488_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.105
cc_102 VPB N_VPWR_c_489_n 0.00354062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_490_n 3.15634e-19 $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_104 VPB N_VPWR_c_491_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_105 VPB N_VPWR_c_492_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.16
cc_106 VPB N_VPWR_c_493_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_494_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.175
cc_108 VPB N_VPWR_c_495_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_496_n 0.014138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_497_n 0.00668519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_498_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_499_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_500_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_501_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_502_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_503_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_504_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_505_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_506_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_507_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_508_n 0.0124787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_509_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_510_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_511_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_485_n 0.0469734f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_X_c_622_n 0.00326551f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.16
cc_127 VPB N_X_c_623_n 0.00168851f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.16
cc_128 VPB N_X_c_624_n 0.00326551f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.175
cc_129 VPB N_X_c_625_n 0.00137166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_X_c_626_n 0.00137166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB X 0.00317321f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_X_c_621_n 0.00193594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 N_A_M1029_g N_A_109_47#_M1000_g 0.0213484f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_M1027_g N_A_109_47#_M1001_g 0.0213484f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1004_g N_A_109_47#_c_266_n 0.0167471f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1008_g N_A_109_47#_c_266_n 0.0106215f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1019_g N_A_109_47#_c_266_n 7.66249e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1015_g N_A_109_47#_c_239_n 0.0111101f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_M1018_g N_A_109_47#_c_239_n 0.0114493f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_c_138_n N_A_109_47#_c_239_n 0.00205431f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_141 A N_A_109_47#_c_239_n 0.0473018f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_142 N_A_M1012_g N_A_109_47#_c_240_n 0.00114299f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A_c_138_n N_A_109_47#_c_240_n 0.00213429f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_144 A N_A_109_47#_c_240_n 0.0138109f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_M1008_g N_A_109_47#_c_260_n 0.0107189f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1019_g N_A_109_47#_c_260_n 0.0107189f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_c_138_n N_A_109_47#_c_260_n 0.00198252f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_148 A N_A_109_47#_c_260_n 0.0578998f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A_M1004_g N_A_109_47#_c_261_n 0.00896105f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1008_g N_A_109_47#_c_261_n 0.00135419f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_c_138_n N_A_109_47#_c_261_n 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_152 A N_A_109_47#_c_261_n 0.026643f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A_M1008_g N_A_109_47#_c_284_n 7.67038e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_M1019_g N_A_109_47#_c_284_n 0.0107272f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1027_g N_A_109_47#_c_284_n 0.0109954f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1029_g N_A_109_47#_c_241_n 0.0126765f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_157 A N_A_109_47#_c_241_n 0.00392548f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A_M1029_g N_A_109_47#_c_242_n 0.00420813f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A_c_138_n N_A_109_47#_c_243_n 0.00448196f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_160 A N_A_109_47#_c_243_n 0.00218678f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A_M1019_g N_A_109_47#_c_263_n 0.00139111f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_c_138_n N_A_109_47#_c_263_n 0.00198252f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_163 N_A_M1027_g N_A_109_47#_c_263_n 0.0133819f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_c_138_n N_A_109_47#_c_245_n 0.00213376f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_165 A N_A_109_47#_c_245_n 0.0138019f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A_c_138_n N_A_109_47#_c_246_n 0.00177712f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_167 A N_A_109_47#_c_246_n 0.0144236f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A_c_138_n N_A_109_47#_c_247_n 0.0213484f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_169 N_A_M1004_g N_VPWR_c_487_n 0.00316354f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_c_138_n N_VPWR_c_487_n 0.00301634f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_171 A N_VPWR_c_487_n 0.00517703f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A_M1008_g N_VPWR_c_488_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_M1019_g N_VPWR_c_488_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_M1027_g N_VPWR_c_489_n 0.00146448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_M1004_g N_VPWR_c_498_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_M1008_g N_VPWR_c_498_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_M1019_g N_VPWR_c_500_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_M1027_g N_VPWR_c_500_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_M1004_g N_VPWR_c_485_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_M1008_g N_VPWR_c_485_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_M1019_g N_VPWR_c_485_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1027_g N_VPWR_c_485_n 0.00952874f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1012_g N_VGND_c_759_n 0.00913095f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_M1015_g N_VGND_c_759_n 5.77787e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_c_138_n N_VGND_c_759_n 0.00477275f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_186 A N_VGND_c_759_n 0.00857385f $X=1.49 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A_M1012_g N_VGND_c_760_n 5.77787e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A_M1015_g N_VGND_c_760_n 0.00769005f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A_M1018_g N_VGND_c_760_n 0.00772492f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A_M1029_g N_VGND_c_760_n 5.9099e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_M1018_g N_VGND_c_761_n 5.9099e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A_M1029_g N_VGND_c_761_n 0.00769102f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_M1018_g N_VGND_c_770_n 0.00350562f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A_M1029_g N_VGND_c_770_n 0.00350562f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A_M1012_g N_VGND_c_776_n 0.0046653f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_196 N_A_M1015_g N_VGND_c_776_n 0.00350562f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A_M1012_g N_VGND_c_784_n 0.00796766f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_M1015_g N_VGND_c_784_n 0.00418574f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_M1018_g N_VGND_c_784_n 0.00418574f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_M1029_g N_VGND_c_784_n 0.00418574f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_109_47#_c_260_n N_VPWR_M1008_s 0.00185611f $X=1.355 $Y=1.53 $X2=0
+ $Y2=0
cc_202 N_A_109_47#_c_263_n N_VPWR_M1027_s 0.00332925f $X=1.927 $Y=1.53 $X2=0
+ $Y2=0
cc_203 N_A_109_47#_c_260_n N_VPWR_c_488_n 0.0104788f $X=1.355 $Y=1.53 $X2=0
+ $Y2=0
cc_204 N_A_109_47#_M1001_g N_VPWR_c_489_n 0.00137415f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_109_47#_c_263_n N_VPWR_c_489_n 0.0102773f $X=1.927 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_109_47#_M1001_g N_VPWR_c_490_n 7.05049e-19 $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_109_47#_M1002_g N_VPWR_c_490_n 0.0112732f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_109_47#_M1003_g N_VPWR_c_490_n 0.0110878f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_109_47#_M1006_g N_VPWR_c_490_n 6.72101e-19 $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_109_47#_M1003_g N_VPWR_c_491_n 6.72101e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_109_47#_M1006_g N_VPWR_c_491_n 0.0110878f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_109_47#_M1009_g N_VPWR_c_491_n 0.0110878f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_109_47#_M1010_g N_VPWR_c_491_n 6.72101e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_109_47#_M1009_g N_VPWR_c_492_n 0.0046653f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_109_47#_M1010_g N_VPWR_c_492_n 0.0046653f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_109_47#_M1009_g N_VPWR_c_493_n 6.72101e-19 $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_109_47#_M1010_g N_VPWR_c_493_n 0.0110878f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_109_47#_M1011_g N_VPWR_c_493_n 0.0110878f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_109_47#_M1013_g N_VPWR_c_493_n 6.72101e-19 $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_109_47#_M1011_g N_VPWR_c_494_n 6.72101e-19 $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_109_47#_M1013_g N_VPWR_c_494_n 0.0110878f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_109_47#_M1014_g N_VPWR_c_494_n 0.0110878f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_109_47#_M1017_g N_VPWR_c_494_n 6.72101e-19 $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_109_47#_c_247_n N_VPWR_c_494_n 3.70191e-19 $X=6.77 $Y=1.16 $X2=0
+ $Y2=0
cc_225 N_A_109_47#_M1014_g N_VPWR_c_495_n 6.72101e-19 $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_109_47#_M1017_g N_VPWR_c_495_n 0.0110878f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_109_47#_M1022_g N_VPWR_c_495_n 0.0110878f $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_109_47#_M1028_g N_VPWR_c_495_n 6.72101e-19 $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_109_47#_c_247_n N_VPWR_c_495_n 3.70191e-19 $X=6.77 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_109_47#_M1022_g N_VPWR_c_497_n 8.11858e-19 $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_109_47#_M1028_g N_VPWR_c_497_n 0.0161769f $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_109_47#_c_266_n N_VPWR_c_498_n 0.0189039f $X=0.68 $Y=1.63 $X2=0 $Y2=0
cc_233 N_A_109_47#_c_284_n N_VPWR_c_500_n 0.0189039f $X=1.52 $Y=1.63 $X2=0 $Y2=0
cc_234 N_A_109_47#_M1001_g N_VPWR_c_502_n 0.00585385f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_109_47#_M1002_g N_VPWR_c_502_n 0.0046653f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_109_47#_M1003_g N_VPWR_c_504_n 0.0046653f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_109_47#_M1006_g N_VPWR_c_504_n 0.0046653f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_109_47#_M1011_g N_VPWR_c_506_n 0.0046653f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A_109_47#_M1013_g N_VPWR_c_506_n 0.0046653f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_109_47#_M1014_g N_VPWR_c_507_n 0.0046653f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_109_47#_M1017_g N_VPWR_c_507_n 0.0046653f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_109_47#_M1022_g N_VPWR_c_508_n 0.0046653f $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_109_47#_M1028_g N_VPWR_c_508_n 0.0046653f $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_A_109_47#_M1004_d N_VPWR_c_485_n 0.00215201f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_245 N_A_109_47#_M1019_d N_VPWR_c_485_n 0.00215201f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_246 N_A_109_47#_M1001_g N_VPWR_c_485_n 0.0106402f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_109_47#_M1002_g N_VPWR_c_485_n 0.00796766f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_248 N_A_109_47#_M1003_g N_VPWR_c_485_n 0.00796766f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_249 N_A_109_47#_M1006_g N_VPWR_c_485_n 0.00796766f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_250 N_A_109_47#_M1009_g N_VPWR_c_485_n 0.00796766f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_251 N_A_109_47#_M1010_g N_VPWR_c_485_n 0.00796766f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_252 N_A_109_47#_M1011_g N_VPWR_c_485_n 0.00796766f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_253 N_A_109_47#_M1013_g N_VPWR_c_485_n 0.00796766f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_A_109_47#_M1014_g N_VPWR_c_485_n 0.00796766f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_A_109_47#_M1017_g N_VPWR_c_485_n 0.00796766f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_109_47#_M1022_g N_VPWR_c_485_n 0.00796766f $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_A_109_47#_M1028_g N_VPWR_c_485_n 0.00796766f $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A_109_47#_c_266_n N_VPWR_c_485_n 0.0122217f $X=0.68 $Y=1.63 $X2=0 $Y2=0
cc_259 N_A_109_47#_c_284_n N_VPWR_c_485_n 0.0122217f $X=1.52 $Y=1.63 $X2=0 $Y2=0
cc_260 N_A_109_47#_M1005_g N_X_c_615_n 0.0111101f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_109_47#_M1007_g N_X_c_615_n 0.0114884f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_109_47#_c_244_n N_X_c_615_n 0.0467269f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_109_47#_c_247_n N_X_c_615_n 0.00205431f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_109_47#_M1000_g N_X_c_616_n 7.27465e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_265 N_A_109_47#_c_241_n N_X_c_616_n 0.00628034f $X=1.84 $Y=0.82 $X2=0 $Y2=0
cc_266 N_A_109_47#_c_244_n N_X_c_616_n 0.0136643f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_109_47#_c_247_n N_X_c_616_n 0.00213429f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_109_47#_M1002_g N_X_c_622_n 0.013304f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_109_47#_M1003_g N_X_c_622_n 0.0135832f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_109_47#_c_244_n N_X_c_622_n 0.0412229f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_109_47#_c_247_n N_X_c_622_n 0.00201555f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_109_47#_M1001_g N_X_c_623_n 7.19058e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_109_47#_c_244_n N_X_c_623_n 0.0121473f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_109_47#_c_263_n N_X_c_623_n 0.00690855f $X=1.927 $Y=1.53 $X2=0 $Y2=0
cc_275 N_A_109_47#_c_247_n N_X_c_623_n 0.00211055f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_109_47#_M1016_g N_X_c_617_n 0.0115326f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A_109_47#_M1020_g N_X_c_617_n 0.0115326f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A_109_47#_c_244_n N_X_c_617_n 0.0467269f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_109_47#_c_247_n N_X_c_617_n 0.00205431f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_109_47#_M1006_g N_X_c_624_n 0.0136273f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_109_47#_M1009_g N_X_c_624_n 0.0136273f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A_109_47#_c_244_n N_X_c_624_n 0.0412229f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A_109_47#_c_247_n N_X_c_624_n 0.00201555f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_109_47#_c_247_n N_X_c_653_n 3.16187e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_109_47#_c_247_n N_X_c_654_n 3.16187e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_109_47#_c_247_n N_X_c_655_n 2.95142e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A_109_47#_c_247_n N_X_c_656_n 3.16187e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_109_47#_c_247_n N_X_c_657_n 2.95142e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A_109_47#_c_244_n N_X_c_618_n 0.0136643f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_109_47#_c_247_n N_X_c_618_n 0.00213429f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A_109_47#_c_244_n N_X_c_625_n 0.0121473f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_109_47#_c_247_n N_X_c_625_n 0.00211055f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A_109_47#_c_244_n N_X_c_619_n 0.0136643f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_109_47#_c_247_n N_X_c_619_n 0.00213429f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A_109_47#_c_244_n N_X_c_626_n 0.0121473f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_109_47#_c_247_n N_X_c_626_n 0.00211055f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_109_47#_M1021_g X 0.0115326f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A_109_47#_M1010_g X 0.0136273f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_109_47#_M1023_g X 0.00915248f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_300 N_A_109_47#_M1011_g X 0.0108218f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A_109_47#_c_244_n X 0.0446492f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_109_47#_c_247_n X 0.00438115f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_109_47#_c_247_n N_X_c_672_n 2.95142e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A_109_47#_M1021_g N_X_c_621_n 3.46149e-19 $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A_109_47#_M1010_g N_X_c_621_n 4.94498e-19 $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A_109_47#_M1023_g N_X_c_621_n 0.00613332f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_109_47#_M1011_g N_X_c_621_n 0.00758103f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_109_47#_M1024_g N_X_c_621_n 0.0139761f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A_109_47#_M1013_g N_X_c_621_n 0.0179335f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_109_47#_M1025_g N_X_c_621_n 0.0139761f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A_109_47#_M1014_g N_X_c_621_n 0.0179335f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A_109_47#_M1026_g N_X_c_621_n 0.0139004f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A_109_47#_M1017_g N_X_c_621_n 0.0178499f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A_109_47#_M1030_g N_X_c_621_n 0.0132046f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A_109_47#_M1022_g N_X_c_621_n 0.0171762f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_109_47#_M1031_g N_X_c_621_n 0.00494338f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A_109_47#_M1028_g N_X_c_621_n 0.00630163f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A_109_47#_c_244_n N_X_c_621_n 0.0105888f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_109_47#_c_247_n N_X_c_621_n 0.0879788f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_109_47#_c_239_n N_VGND_M1015_d 0.00162006f $X=1.435 $Y=0.82 $X2=0
+ $Y2=0
cc_321 N_A_109_47#_c_241_n N_VGND_M1029_d 0.00337318f $X=1.84 $Y=0.82 $X2=0
+ $Y2=0
cc_322 N_A_109_47#_c_239_n N_VGND_c_760_n 0.016419f $X=1.435 $Y=0.82 $X2=0 $Y2=0
cc_323 N_A_109_47#_M1000_g N_VGND_c_761_n 0.00799556f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_324 N_A_109_47#_M1005_g N_VGND_c_761_n 5.77787e-19 $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_325 N_A_109_47#_c_241_n N_VGND_c_761_n 0.0153948f $X=1.84 $Y=0.82 $X2=0 $Y2=0
cc_326 N_A_109_47#_c_244_n N_VGND_c_761_n 0.00197677f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_109_47#_M1000_g N_VGND_c_762_n 5.77787e-19 $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_328 N_A_109_47#_M1005_g N_VGND_c_762_n 0.00769005f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_329 N_A_109_47#_M1007_g N_VGND_c_762_n 0.00769005f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_330 N_A_109_47#_M1016_g N_VGND_c_762_n 5.77787e-19 $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_331 N_A_109_47#_M1007_g N_VGND_c_763_n 5.77787e-19 $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_332 N_A_109_47#_M1016_g N_VGND_c_763_n 0.00769005f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_333 N_A_109_47#_M1020_g N_VGND_c_763_n 0.00769005f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_334 N_A_109_47#_M1021_g N_VGND_c_763_n 5.77787e-19 $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_335 N_A_109_47#_M1020_g N_VGND_c_764_n 0.00350562f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_336 N_A_109_47#_M1021_g N_VGND_c_764_n 0.00350562f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_337 N_A_109_47#_M1020_g N_VGND_c_765_n 5.77787e-19 $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_338 N_A_109_47#_M1021_g N_VGND_c_765_n 0.00769005f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_339 N_A_109_47#_M1023_g N_VGND_c_765_n 0.00769005f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_340 N_A_109_47#_M1024_g N_VGND_c_765_n 5.77787e-19 $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_341 N_A_109_47#_M1023_g N_VGND_c_766_n 5.77787e-19 $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_342 N_A_109_47#_M1024_g N_VGND_c_766_n 0.00769005f $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_343 N_A_109_47#_M1025_g N_VGND_c_766_n 0.00769005f $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_A_109_47#_M1026_g N_VGND_c_766_n 5.77787e-19 $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_345 N_A_109_47#_c_247_n N_VGND_c_766_n 3.77859e-19 $X=6.77 $Y=1.16 $X2=0
+ $Y2=0
cc_346 N_A_109_47#_M1025_g N_VGND_c_767_n 5.77787e-19 $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_347 N_A_109_47#_M1026_g N_VGND_c_767_n 0.00769005f $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_348 N_A_109_47#_M1030_g N_VGND_c_767_n 0.00769005f $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_349 N_A_109_47#_M1031_g N_VGND_c_767_n 5.77787e-19 $X=6.77 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_109_47#_c_247_n N_VGND_c_767_n 3.77859e-19 $X=6.77 $Y=1.16 $X2=0
+ $Y2=0
cc_351 N_A_109_47#_M1030_g N_VGND_c_769_n 7.33828e-19 $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_352 N_A_109_47#_M1031_g N_VGND_c_769_n 0.0125262f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A_109_47#_c_239_n N_VGND_c_770_n 0.00193763f $X=1.435 $Y=0.82 $X2=0
+ $Y2=0
cc_354 N_A_109_47#_c_453_p N_VGND_c_770_n 0.0110017f $X=1.52 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A_109_47#_c_241_n N_VGND_c_770_n 0.00193763f $X=1.84 $Y=0.82 $X2=0
+ $Y2=0
cc_356 N_A_109_47#_M1000_g N_VGND_c_772_n 0.0046653f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_109_47#_M1005_g N_VGND_c_772_n 0.00350562f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_358 N_A_109_47#_M1007_g N_VGND_c_774_n 0.00350562f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_359 N_A_109_47#_M1016_g N_VGND_c_774_n 0.00350562f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_109_47#_c_459_p N_VGND_c_776_n 0.0113595f $X=0.68 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_109_47#_c_239_n N_VGND_c_776_n 0.00193763f $X=1.435 $Y=0.82 $X2=0
+ $Y2=0
cc_362 N_A_109_47#_M1023_g N_VGND_c_777_n 0.0035053f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_109_47#_M1024_g N_VGND_c_777_n 0.00350562f $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_364 N_A_109_47#_M1025_g N_VGND_c_778_n 0.00350562f $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_109_47#_M1026_g N_VGND_c_778_n 0.00350562f $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_366 N_A_109_47#_M1030_g N_VGND_c_779_n 0.00350562f $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_367 N_A_109_47#_M1031_g N_VGND_c_779_n 0.0046653f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_109_47#_M1012_s N_VGND_c_784_n 0.00418657f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_369 N_A_109_47#_M1018_s N_VGND_c_784_n 0.00266498f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_370 N_A_109_47#_M1000_g N_VGND_c_784_n 0.00796766f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_371 N_A_109_47#_M1005_g N_VGND_c_784_n 0.00418574f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_372 N_A_109_47#_M1007_g N_VGND_c_784_n 0.00418574f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_373 N_A_109_47#_M1016_g N_VGND_c_784_n 0.00418574f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_374 N_A_109_47#_M1020_g N_VGND_c_784_n 0.00418574f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_375 N_A_109_47#_M1021_g N_VGND_c_784_n 0.00418574f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_376 N_A_109_47#_M1023_g N_VGND_c_784_n 0.00418516f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_377 N_A_109_47#_M1024_g N_VGND_c_784_n 0.00418574f $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_378 N_A_109_47#_M1025_g N_VGND_c_784_n 0.00418574f $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_379 N_A_109_47#_M1026_g N_VGND_c_784_n 0.00418574f $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_380 N_A_109_47#_M1030_g N_VGND_c_784_n 0.00418574f $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_381 N_A_109_47#_M1031_g N_VGND_c_784_n 0.00796766f $X=6.77 $Y=0.56 $X2=0
+ $Y2=0
cc_382 N_A_109_47#_c_459_p N_VGND_c_784_n 0.0064623f $X=0.68 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A_109_47#_c_239_n N_VGND_c_784_n 0.00895872f $X=1.435 $Y=0.82 $X2=0
+ $Y2=0
cc_384 N_A_109_47#_c_453_p N_VGND_c_784_n 0.00644569f $X=1.52 $Y=0.56 $X2=0
+ $Y2=0
cc_385 N_A_109_47#_c_241_n N_VGND_c_784_n 0.00485047f $X=1.84 $Y=0.82 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_485_n N_X_M1001_d 0.00570907f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_485_n N_X_M1003_d 0.00570907f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_c_485_n N_X_M1009_d 0.00570907f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_485_n N_X_M1011_d 0.00570907f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_485_n N_X_M1014_d 0.00570907f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_485_n N_X_M1022_d 0.00570907f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_502_n N_X_c_695_n 0.0113958f $X=2.615 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_485_n N_X_c_695_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_M1002_s N_X_c_622_n 0.00185611f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_395 N_VPWR_c_490_n N_X_c_622_n 0.0140015f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_396 N_VPWR_c_504_n N_X_c_699_n 0.0113958f $X=3.455 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_485_n N_X_c_699_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_M1006_s N_X_c_624_n 0.00185611f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_399 N_VPWR_c_491_n N_X_c_624_n 0.0140015f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_400 N_VPWR_c_492_n N_X_c_703_n 0.0113958f $X=4.295 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_485_n N_X_c_703_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_507_n N_X_c_655_n 0.0113958f $X=5.975 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_c_485_n N_X_c_655_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_508_n N_X_c_657_n 0.0113958f $X=6.815 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_c_485_n N_X_c_657_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_M1010_s X 0.00185611f $X=4.325 $Y=1.485 $X2=0 $Y2=0
cc_407 N_VPWR_c_493_n X 0.0140015f $X=4.46 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_c_506_n N_X_c_672_n 0.0113958f $X=5.135 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_485_n N_X_c_672_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_M1013_s N_X_c_621_n 0.00193841f $X=5.165 $Y=1.485 $X2=0 $Y2=0
cc_411 N_VPWR_M1017_s N_X_c_621_n 0.00193841f $X=6.005 $Y=1.485 $X2=0 $Y2=0
cc_412 N_VPWR_c_494_n N_X_c_621_n 0.0154647f $X=5.3 $Y=2 $X2=0 $Y2=0
cc_413 N_VPWR_c_495_n N_X_c_621_n 0.0154647f $X=6.14 $Y=2 $X2=0 $Y2=0
cc_414 N_VPWR_c_497_n N_VGND_c_769_n 0.00927817f $X=6.98 $Y=1.66 $X2=0 $Y2=0
cc_415 N_X_c_615_n N_VGND_M1005_d 0.00162006f $X=3.115 $Y=0.82 $X2=0 $Y2=0
cc_416 N_X_c_617_n N_VGND_M1016_d 0.00162006f $X=3.955 $Y=0.82 $X2=0 $Y2=0
cc_417 X N_VGND_M1021_d 0.00162006f $X=4.71 $Y=0.765 $X2=0 $Y2=0
cc_418 N_X_c_621_n N_VGND_M1024_d 0.00169066f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_419 N_X_c_621_n N_VGND_M1026_d 0.00169066f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_420 N_X_c_615_n N_VGND_c_762_n 0.016419f $X=3.115 $Y=0.82 $X2=0 $Y2=0
cc_421 N_X_c_617_n N_VGND_c_763_n 0.016419f $X=3.955 $Y=0.82 $X2=0 $Y2=0
cc_422 N_X_c_617_n N_VGND_c_764_n 0.00193763f $X=3.955 $Y=0.82 $X2=0 $Y2=0
cc_423 N_X_c_725_p N_VGND_c_764_n 0.0113595f $X=4.04 $Y=0.56 $X2=0 $Y2=0
cc_424 X N_VGND_c_764_n 0.00193763f $X=4.71 $Y=0.765 $X2=0 $Y2=0
cc_425 X N_VGND_c_765_n 0.016419f $X=4.71 $Y=0.765 $X2=0 $Y2=0
cc_426 N_X_c_621_n N_VGND_c_766_n 0.0180722f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_427 N_X_c_621_n N_VGND_c_767_n 0.0180722f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_428 N_X_c_730_p N_VGND_c_772_n 0.0113595f $X=2.36 $Y=0.56 $X2=0 $Y2=0
cc_429 N_X_c_615_n N_VGND_c_772_n 0.00193763f $X=3.115 $Y=0.82 $X2=0 $Y2=0
cc_430 N_X_c_615_n N_VGND_c_774_n 0.00193763f $X=3.115 $Y=0.82 $X2=0 $Y2=0
cc_431 N_X_c_733_p N_VGND_c_774_n 0.0113595f $X=3.2 $Y=0.56 $X2=0 $Y2=0
cc_432 N_X_c_617_n N_VGND_c_774_n 0.00193763f $X=3.955 $Y=0.82 $X2=0 $Y2=0
cc_433 N_X_c_653_n N_VGND_c_777_n 0.0111222f $X=4.88 $Y=0.56 $X2=0 $Y2=0
cc_434 X N_VGND_c_777_n 0.0011009f $X=4.71 $Y=0.765 $X2=0 $Y2=0
cc_435 N_X_c_621_n N_VGND_c_777_n 0.0029871f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_436 N_X_c_654_n N_VGND_c_778_n 0.0111222f $X=5.72 $Y=0.56 $X2=0 $Y2=0
cc_437 N_X_c_621_n N_VGND_c_778_n 0.0042033f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_438 N_X_c_656_n N_VGND_c_779_n 0.0111222f $X=6.56 $Y=0.56 $X2=0 $Y2=0
cc_439 N_X_c_621_n N_VGND_c_779_n 0.00210921f $X=6.56 $Y=1.175 $X2=0 $Y2=0
cc_440 N_X_M1000_s N_VGND_c_784_n 0.00418657f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_441 N_X_M1007_s N_VGND_c_784_n 0.00266406f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_442 N_X_M1020_s N_VGND_c_784_n 0.00266406f $X=3.905 $Y=0.235 $X2=0 $Y2=0
cc_443 N_X_M1023_s N_VGND_c_784_n 0.00267647f $X=4.745 $Y=0.235 $X2=0 $Y2=0
cc_444 N_X_M1025_s N_VGND_c_784_n 0.00269036f $X=5.585 $Y=0.235 $X2=0 $Y2=0
cc_445 N_X_M1030_s N_VGND_c_784_n 0.00415697f $X=6.425 $Y=0.235 $X2=0 $Y2=0
cc_446 N_X_c_730_p N_VGND_c_784_n 0.0064623f $X=2.36 $Y=0.56 $X2=0 $Y2=0
cc_447 N_X_c_615_n N_VGND_c_784_n 0.00895872f $X=3.115 $Y=0.82 $X2=0 $Y2=0
cc_448 N_X_c_733_p N_VGND_c_784_n 0.0064623f $X=3.2 $Y=0.56 $X2=0 $Y2=0
cc_449 N_X_c_617_n N_VGND_c_784_n 0.00895872f $X=3.955 $Y=0.82 $X2=0 $Y2=0
cc_450 N_X_c_725_p N_VGND_c_784_n 0.0064623f $X=4.04 $Y=0.56 $X2=0 $Y2=0
cc_451 N_X_c_653_n N_VGND_c_784_n 0.00641247f $X=4.88 $Y=0.56 $X2=0 $Y2=0
cc_452 N_X_c_654_n N_VGND_c_784_n 0.00641247f $X=5.72 $Y=0.56 $X2=0 $Y2=0
cc_453 N_X_c_656_n N_VGND_c_784_n 0.00641247f $X=6.56 $Y=0.56 $X2=0 $Y2=0
cc_454 X N_VGND_c_784_n 0.00691507f $X=4.71 $Y=0.765 $X2=0 $Y2=0
cc_455 N_X_c_621_n N_VGND_c_784_n 0.0217141f $X=6.56 $Y=1.175 $X2=0 $Y2=0

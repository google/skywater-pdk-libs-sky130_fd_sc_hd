* File: sky130_fd_sc_hd__nand2b_2.pxi.spice
* Created: Tue Sep  1 19:15:50 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2B_2%A_N N_A_N_M1009_g N_A_N_M1004_g A_N N_A_N_c_62_n
+ N_A_N_c_63_n PM_SKY130_FD_SC_HD__NAND2B_2%A_N
x_PM_SKY130_FD_SC_HD__NAND2B_2%A_27_93# N_A_27_93#_M1009_s N_A_27_93#_M1004_s
+ N_A_27_93#_M1001_g N_A_27_93#_M1006_g N_A_27_93#_M1002_g N_A_27_93#_M1005_g
+ N_A_27_93#_c_94_n N_A_27_93#_c_95_n N_A_27_93#_c_96_n N_A_27_93#_c_97_n
+ N_A_27_93#_c_110_n N_A_27_93#_c_102_n N_A_27_93#_c_98_n N_A_27_93#_c_103_n
+ PM_SKY130_FD_SC_HD__NAND2B_2%A_27_93#
x_PM_SKY130_FD_SC_HD__NAND2B_2%B N_B_M1000_g N_B_M1007_g N_B_M1003_g N_B_M1008_g
+ N_B_c_159_n B B B B N_B_c_163_n PM_SKY130_FD_SC_HD__NAND2B_2%B
x_PM_SKY130_FD_SC_HD__NAND2B_2%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1003_d
+ N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n VPWR N_VPWR_c_218_n
+ N_VPWR_c_219_n N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_214_n
+ PM_SKY130_FD_SC_HD__NAND2B_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND2B_2%Y N_Y_M1002_d N_Y_M1001_s N_Y_M1000_s N_Y_c_263_n
+ N_Y_c_264_n N_Y_c_278_n N_Y_c_281_n Y Y Y Y N_Y_c_260_n N_Y_c_301_n Y
+ PM_SKY130_FD_SC_HD__NAND2B_2%Y
x_PM_SKY130_FD_SC_HD__NAND2B_2%VGND N_VGND_M1009_d N_VGND_M1007_s N_VGND_c_308_n
+ N_VGND_c_309_n VGND N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n
+ N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n PM_SKY130_FD_SC_HD__NAND2B_2%VGND
x_PM_SKY130_FD_SC_HD__NAND2B_2%A_229_47# N_A_229_47#_M1002_s N_A_229_47#_M1005_s
+ N_A_229_47#_M1008_d N_A_229_47#_c_354_n N_A_229_47#_c_355_n
+ N_A_229_47#_c_364_n N_A_229_47#_c_367_n N_A_229_47#_c_356_n
+ N_A_229_47#_c_357_n N_A_229_47#_c_358_n PM_SKY130_FD_SC_HD__NAND2B_2%A_229_47#
cc_1 VNB A_N 0.00359475f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_2 VNB N_A_N_c_62_n 0.0231987f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_3 VNB N_A_N_c_63_n 0.0248851f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_4 VNB N_A_27_93#_M1001_g 4.26041e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_93#_M1006_g 5.73676e-19 $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_6 VNB N_A_27_93#_M1002_g 0.0227844f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_7 VNB N_A_27_93#_M1005_g 0.0176595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_93#_c_94_n 0.0171521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_93#_c_95_n 0.0230853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_93#_c_96_n 0.0401444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_93#_c_97_n 0.0213871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_93#_c_98_n 0.0123578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B_M1000_g 5.55993e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.675
cc_14 VNB N_B_M1007_g 0.0175567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B_M1008_g 0.0230765f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_16 VNB N_B_c_159_n 0.0280668f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_17 VNB B 0.00330317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB B 4.63871e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB B 0.00843946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_c_163_n 0.0268135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_214_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB Y 0.00126848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_260_n 5.45942e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_308_n 0.00863002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_309_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_26 VNB N_VGND_c_310_n 0.0172029f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_27 VNB N_VGND_c_311_n 0.0385811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_312_n 0.0173168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_313_n 0.19665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_314_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_315_n 0.00323511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_229_47#_c_354_n 0.00289512f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_33 VNB N_A_229_47#_c_355_n 0.0068998f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_34 VNB N_A_229_47#_c_356_n 0.00198362f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_35 VNB N_A_229_47#_c_357_n 0.0131994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_229_47#_c_358_n 0.0178665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_A_N_M1004_g 0.0255631f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_38 VPB A_N 0.00128469f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_39 VPB N_A_N_c_62_n 0.00439182f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_40 VPB N_A_27_93#_M1001_g 0.0228832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_93#_M1006_g 0.0238428f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=0.995
cc_42 VPB N_A_27_93#_c_97_n 0.00892971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_93#_c_102_n 0.00109431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_93#_c_103_n 0.0153447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B_M1000_g 0.0231962f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.675
cc_46 VPB N_B_M1003_g 0.0275749f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_47 VPB N_B_c_159_n 0.00305706f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_48 VPB B 0.0032262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_B_c_163_n 0.00721154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_215_n 0.0234672f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_51 VPB N_VPWR_c_216_n 0.0112306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_217_n 0.0469363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_218_n 0.0206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_219_n 0.0178481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_220_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_221_n 0.0183948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_222_n 0.0180355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_214_n 0.0592593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB Y 0.00238104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_A_N_M1004_g N_A_27_93#_M1001_g 0.0201227f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_61 A_N N_A_27_93#_M1002_g 6.79284e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_62 A_N N_A_27_93#_c_94_n 0.00339492f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_N_c_62_n N_A_27_93#_c_94_n 0.019421f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_64 A_N N_A_27_93#_c_97_n 0.024314f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_N_c_63_n N_A_27_93#_c_97_n 0.0189022f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_66 N_A_N_M1004_g N_A_27_93#_c_110_n 0.0130416f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_67 A_N N_A_27_93#_c_110_n 0.0237f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_N_c_62_n N_A_27_93#_c_110_n 0.00278962f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_N_M1004_g N_A_27_93#_c_102_n 7.74842e-19 $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_70 A_N N_A_27_93#_c_102_n 0.0158062f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_N_c_62_n N_A_27_93#_c_102_n 2.04341e-19 $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_N_M1004_g N_A_27_93#_c_103_n 0.00487393f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_73 N_A_N_M1004_g N_VPWR_c_215_n 0.0038843f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_74 N_A_N_M1004_g N_VPWR_c_218_n 0.00327927f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_75 N_A_N_M1004_g N_VPWR_c_214_n 0.00417489f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_76 A_N N_VGND_c_308_n 0.0212865f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_N_c_62_n N_VGND_c_308_n 0.00285475f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_N_c_63_n N_VGND_c_308_n 0.0159737f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_N_c_63_n N_VGND_c_310_n 0.00407165f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_N_c_63_n N_VGND_c_313_n 0.00413741f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_N_c_63_n N_A_229_47#_c_354_n 5.59778e-19 $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_N_c_63_n N_A_229_47#_c_355_n 0.00202997f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_27_93#_M1006_g N_B_M1000_g 0.0119603f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_27_93#_M1005_g N_B_M1007_g 0.0133281f $X=1.9 $Y=0.56 $X2=0 $Y2=0
cc_85 N_A_27_93#_c_96_n N_B_c_159_n 0.0183428f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_27_93#_c_96_n B 0.00190141f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_27_93#_c_110_n N_VPWR_M1004_d 0.00493585f $X=1.03 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_27_93#_M1001_g N_VPWR_c_215_n 0.00450113f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_27_93#_c_110_n N_VPWR_c_215_n 0.018387f $X=1.03 $Y=1.58 $X2=0 $Y2=0
cc_90 N_A_27_93#_M1001_g N_VPWR_c_221_n 0.00585385f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_27_93#_M1006_g N_VPWR_c_221_n 0.00436487f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_27_93#_M1006_g N_VPWR_c_222_n 0.00378613f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_27_93#_M1001_g N_VPWR_c_214_n 0.0120141f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_27_93#_M1006_g N_VPWR_c_214_n 0.00666539f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_27_93#_c_110_n N_Y_M1001_s 0.00321459f $X=1.03 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_27_93#_c_96_n N_Y_c_263_n 0.00465809f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_27_93#_M1006_g N_Y_c_264_n 0.0160948f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_27_93#_c_95_n N_Y_c_264_n 4.86978e-19 $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_27_93#_c_96_n N_Y_c_264_n 5.86337e-19 $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_27_93#_c_110_n N_Y_c_264_n 0.0173714f $X=1.03 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_27_93#_M1006_g Y 0.00563356f $X=1.44 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_27_93#_M1002_g Y 0.00613986f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_27_93#_M1005_g Y 0.00326985f $X=1.9 $Y=0.56 $X2=0 $Y2=0
cc_104 N_A_27_93#_c_96_n Y 0.0234185f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_27_93#_c_102_n Y 0.0318379f $X=1.195 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_27_93#_M1002_g N_Y_c_260_n 0.00380069f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A_27_93#_M1005_g N_Y_c_260_n 0.00473764f $X=1.9 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A_27_93#_M1002_g N_VGND_c_308_n 0.00208931f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_27_93#_c_110_n N_VGND_c_308_n 0.00106304f $X=1.03 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_27_93#_c_98_n N_VGND_c_310_n 0.00593412f $X=0.26 $Y=0.675 $X2=0 $Y2=0
cc_111 N_A_27_93#_M1002_g N_VGND_c_311_n 0.00357877f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_27_93#_M1005_g N_VGND_c_311_n 0.00357877f $X=1.9 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_27_93#_M1002_g N_VGND_c_313_n 0.00655123f $X=1.48 $Y=0.56 $X2=0 $Y2=0
cc_114 N_A_27_93#_M1005_g N_VGND_c_313_n 0.00525237f $X=1.9 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A_27_93#_c_98_n N_VGND_c_313_n 0.00761143f $X=0.26 $Y=0.675 $X2=0 $Y2=0
cc_116 N_A_27_93#_M1002_g N_A_229_47#_c_355_n 4.46102e-19 $X=1.48 $Y=0.56 $X2=0
+ $Y2=0
cc_117 N_A_27_93#_c_95_n N_A_229_47#_c_355_n 0.00709894f $X=1.365 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_A_27_93#_c_102_n N_A_229_47#_c_355_n 0.0240041f $X=1.195 $Y=1.16 $X2=0
+ $Y2=0
cc_119 N_A_27_93#_M1002_g N_A_229_47#_c_364_n 0.0124155f $X=1.48 $Y=0.56 $X2=0
+ $Y2=0
cc_120 N_A_27_93#_M1005_g N_A_229_47#_c_364_n 0.0124155f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_121 N_A_27_93#_c_96_n N_A_229_47#_c_364_n 2.87379e-19 $X=1.9 $Y=1.16 $X2=0
+ $Y2=0
cc_122 B N_VPWR_M1006_d 0.00447714f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_123 N_B_M1003_g N_VPWR_c_217_n 0.00457701f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B_c_159_n N_VPWR_c_217_n 0.0070915f $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_125 B N_VPWR_c_217_n 0.0214767f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B_M1000_g N_VPWR_c_219_n 0.00409104f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VPWR_c_219_n 0.00541359f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B_M1000_g N_VPWR_c_222_n 0.00484942f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B_M1000_g N_VPWR_c_214_n 0.00635193f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_130 N_B_M1003_g N_VPWR_c_214_n 0.0105165f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B_M1000_g N_Y_c_263_n 0.00972867f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_132 B N_Y_c_263_n 0.0105423f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_133 B N_Y_c_263_n 0.00250163f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B_M1003_g N_Y_c_278_n 0.00419276f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B_c_159_n N_Y_c_278_n 0.00229501f $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_136 B N_Y_c_278_n 0.0144864f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_137 N_B_M1000_g N_Y_c_281_n 0.014297f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B_M1003_g N_Y_c_281_n 0.00716293f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_139 B N_Y_c_281_n 0.00188606f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_140 N_B_M1000_g Y 0.00235751f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B_c_159_n Y 4.17935e-19 $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_142 B Y 0.0159738f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_143 B Y 0.0281888f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_144 N_B_M1007_g N_VGND_c_309_n 0.00268723f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_145 N_B_M1008_g N_VGND_c_309_n 0.00268723f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_146 N_B_M1007_g N_VGND_c_311_n 0.00418507f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_147 N_B_M1008_g N_VGND_c_312_n 0.00420025f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_148 N_B_M1007_g N_VGND_c_313_n 0.00569347f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_149 N_B_M1008_g N_VGND_c_313_n 0.00662088f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_150 N_B_M1007_g N_A_229_47#_c_367_n 0.00244813f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_151 N_B_M1007_g N_A_229_47#_c_356_n 0.00473177f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_152 N_B_M1008_g N_A_229_47#_c_356_n 4.52257e-19 $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_153 N_B_c_159_n N_A_229_47#_c_356_n 0.0017301f $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_154 B N_A_229_47#_c_356_n 0.0143035f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_155 B N_A_229_47#_c_356_n 0.00756265f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_156 N_B_M1007_g N_A_229_47#_c_357_n 0.00930481f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_157 N_B_M1008_g N_A_229_47#_c_357_n 0.0106332f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_158 N_B_c_159_n N_A_229_47#_c_357_n 0.00237212f $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_159 B N_A_229_47#_c_357_n 0.0648863f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_160 N_B_c_163_n N_A_229_47#_c_357_n 0.00728275f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B_M1007_g N_A_229_47#_c_358_n 5.13071e-19 $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_162 N_B_M1008_g N_A_229_47#_c_358_n 0.00599685f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_163 N_VPWR_c_214_n N_Y_M1001_s 0.0026338f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_164 N_VPWR_c_214_n N_Y_M1000_s 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_165 N_VPWR_M1006_d N_Y_c_263_n 0.00996823f $X=1.515 $Y=1.485 $X2=0 $Y2=0
cc_166 N_VPWR_c_219_n N_Y_c_263_n 0.00200535f $X=2.805 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_214_n N_Y_c_263_n 0.0040108f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_M1006_d N_Y_c_264_n 0.00417566f $X=1.515 $Y=1.485 $X2=0 $Y2=0
cc_169 N_VPWR_c_221_n N_Y_c_264_n 0.00221336f $X=1.535 $Y=2.49 $X2=0 $Y2=0
cc_170 N_VPWR_c_222_n N_Y_c_264_n 0.0417172f $X=2.11 $Y=2.49 $X2=0 $Y2=0
cc_171 N_VPWR_c_214_n N_Y_c_264_n 0.00591612f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_172 N_VPWR_c_219_n N_Y_c_281_n 0.0205884f $X=2.805 $Y=2.72 $X2=0 $Y2=0
cc_173 N_VPWR_c_222_n N_Y_c_281_n 0.0236692f $X=2.11 $Y=2.49 $X2=0 $Y2=0
cc_174 N_VPWR_c_214_n N_Y_c_281_n 0.0130643f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_175 N_VPWR_M1006_d Y 0.00819515f $X=1.515 $Y=1.485 $X2=0 $Y2=0
cc_176 N_VPWR_c_221_n N_Y_c_301_n 0.0187393f $X=1.535 $Y=2.49 $X2=0 $Y2=0
cc_177 N_VPWR_c_214_n N_Y_c_301_n 0.0125064f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_178 N_Y_M1002_d N_VGND_c_313_n 0.00216833f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_179 N_Y_c_260_n N_A_229_47#_c_355_n 0.00443415f $X=1.67 $Y=0.905 $X2=0 $Y2=0
cc_180 N_Y_M1002_d N_A_229_47#_c_364_n 0.00305226f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_181 N_Y_c_260_n N_A_229_47#_c_364_n 0.016295f $X=1.67 $Y=0.905 $X2=0 $Y2=0
cc_182 N_Y_c_260_n N_A_229_47#_c_356_n 0.00884302f $X=1.67 $Y=0.905 $X2=0 $Y2=0
cc_183 N_VGND_c_313_n N_A_229_47#_M1002_s 0.00209324f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_184 N_VGND_c_313_n N_A_229_47#_M1005_s 0.00215206f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_185 N_VGND_c_313_n N_A_229_47#_M1008_d 0.00209319f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_308_n N_A_229_47#_c_354_n 0.0144584f $X=0.745 $Y=0.38 $X2=0
+ $Y2=0
cc_187 N_VGND_c_311_n N_A_229_47#_c_354_n 0.0191208f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_c_313_n N_A_229_47#_c_354_n 0.0105783f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_c_308_n N_A_229_47#_c_355_n 0.0229678f $X=0.745 $Y=0.38 $X2=0
+ $Y2=0
cc_190 N_VGND_c_311_n N_A_229_47#_c_364_n 0.0362386f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_313_n N_A_229_47#_c_364_n 0.023553f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_311_n N_A_229_47#_c_367_n 0.0152108f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_313_n N_A_229_47#_c_367_n 0.00940698f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_M1007_s N_A_229_47#_c_357_n 0.00162194f $X=2.395 $Y=0.235 $X2=0
+ $Y2=0
cc_195 N_VGND_c_309_n N_A_229_47#_c_357_n 0.0122822f $X=2.53 $Y=0.36 $X2=0 $Y2=0
cc_196 N_VGND_c_311_n N_A_229_47#_c_357_n 0.00214238f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_312_n N_A_229_47#_c_357_n 0.00214238f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_313_n N_A_229_47#_c_357_n 0.0086619f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_312_n N_A_229_47#_c_358_n 0.0224042f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_313_n N_A_229_47#_c_358_n 0.0131812f $X=2.99 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__and4b_4.pxi.spice
* Created: Tue Sep  1 18:58:30 2020
* 
x_PM_SKY130_FD_SC_HD__AND4B_4%A_N N_A_N_M1016_g N_A_N_M1009_g A_N A_N A_N
+ N_A_N_c_84_n PM_SKY130_FD_SC_HD__AND4B_4%A_N
x_PM_SKY130_FD_SC_HD__AND4B_4%A_174_21# N_A_174_21#_M1005_d N_A_174_21#_M1012_d
+ N_A_174_21#_M1006_d N_A_174_21#_c_116_n N_A_174_21#_M1002_g
+ N_A_174_21#_M1001_g N_A_174_21#_c_117_n N_A_174_21#_M1004_g
+ N_A_174_21#_M1003_g N_A_174_21#_c_118_n N_A_174_21#_M1007_g
+ N_A_174_21#_M1013_g N_A_174_21#_c_119_n N_A_174_21#_M1017_g
+ N_A_174_21#_M1014_g N_A_174_21#_c_179_p N_A_174_21#_c_120_n
+ N_A_174_21#_c_121_n N_A_174_21#_c_122_n N_A_174_21#_c_141_p
+ N_A_174_21#_c_227_p N_A_174_21#_c_181_p N_A_174_21#_c_137_p
+ N_A_174_21#_c_154_p N_A_174_21#_c_123_n N_A_174_21#_c_156_p
+ N_A_174_21#_c_124_n PM_SKY130_FD_SC_HD__AND4B_4%A_174_21#
x_PM_SKY130_FD_SC_HD__AND4B_4%D N_D_M1011_g N_D_M1012_g D N_D_c_262_n
+ N_D_c_263_n PM_SKY130_FD_SC_HD__AND4B_4%D
x_PM_SKY130_FD_SC_HD__AND4B_4%C N_C_c_303_n N_C_M1008_g N_C_M1010_g C C
+ N_C_c_305_n PM_SKY130_FD_SC_HD__AND4B_4%C
x_PM_SKY130_FD_SC_HD__AND4B_4%B N_B_M1015_g N_B_M1006_g B B N_B_c_339_n
+ N_B_c_340_n PM_SKY130_FD_SC_HD__AND4B_4%B
x_PM_SKY130_FD_SC_HD__AND4B_4%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1009_s
+ N_A_27_47#_c_374_n N_A_27_47#_M1005_g N_A_27_47#_M1000_g N_A_27_47#_c_375_n
+ N_A_27_47#_c_381_n N_A_27_47#_c_382_n N_A_27_47#_c_376_n N_A_27_47#_c_377_n
+ N_A_27_47#_c_378_n N_A_27_47#_c_385_n PM_SKY130_FD_SC_HD__AND4B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4B_4%VPWR N_VPWR_M1009_d N_VPWR_M1003_d N_VPWR_M1014_d
+ N_VPWR_M1010_d N_VPWR_M1000_d N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n
+ VPWR N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n
+ N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_450_n
+ PM_SKY130_FD_SC_HD__AND4B_4%VPWR
x_PM_SKY130_FD_SC_HD__AND4B_4%X N_X_M1002_d N_X_M1007_d N_X_M1001_s N_X_M1013_s
+ N_X_c_564_p N_X_c_537_n N_X_c_541_n N_X_c_568_p X X X N_X_c_533_n X X
+ PM_SKY130_FD_SC_HD__AND4B_4%X
x_PM_SKY130_FD_SC_HD__AND4B_4%VGND N_VGND_M1016_d N_VGND_M1004_s N_VGND_M1017_s
+ N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n VGND N_VGND_c_578_n
+ N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n N_VGND_c_582_n N_VGND_c_583_n
+ N_VGND_c_584_n N_VGND_c_585_n PM_SKY130_FD_SC_HD__AND4B_4%VGND
cc_1 VNB N_A_N_M1016_g 0.0321441f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.00358216f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_3 VNB N_A_N_c_84_n 0.0227704f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_4 VNB N_A_174_21#_c_116_n 0.0159577f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_5 VNB N_A_174_21#_c_117_n 0.0157453f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_6 VNB N_A_174_21#_c_118_n 0.0157694f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.19
cc_7 VNB N_A_174_21#_c_119_n 0.0187605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_174_21#_c_120_n 0.0744831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_174_21#_c_121_n 0.00288958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_174_21#_c_122_n 4.58244e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_174_21#_c_123_n 0.022212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_174_21#_c_124_n 0.00135351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB D 0.00218032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_D_c_262_n 0.0219146f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_15 VNB N_D_c_263_n 0.0191016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_C_c_303_n 0.0164313f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_17 VNB C 0.00199419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_C_c_305_n 0.0244306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB B 0.00444113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_c_339_n 0.0239968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B_c_340_n 0.0178215f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_22 VNB N_A_27_47#_c_374_n 0.0236022f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_23 VNB N_A_27_47#_c_375_n 0.03336f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_24 VNB N_A_27_47#_c_376_n 0.00162108f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.19
cc_25 VNB N_A_27_47#_c_377_n 0.0448012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_378_n 0.0128993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_450_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB X 0.00104729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_575_n 0.00271064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_576_n 3.08095e-19 $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_31 VNB N_VGND_c_577_n 0.00494838f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.85
cc_32 VNB N_VGND_c_578_n 0.0178546f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.19
cc_33 VNB N_VGND_c_579_n 0.011348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_580_n 0.0138593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_581_n 0.0604534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_582_n 0.257164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_583_n 0.00507198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_584_n 0.00436184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_585_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_A_N_M1009_g 0.0549481f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_41 VPB A_N 0.00194922f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_42 VPB N_A_N_c_84_n 0.00469075f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_43 VPB N_A_174_21#_M1001_g 0.0186856f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_44 VPB N_A_174_21#_M1003_g 0.0182315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_174_21#_M1013_g 0.0182665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_174_21#_M1014_g 0.0214566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_174_21#_c_120_n 0.0163199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_174_21#_c_122_n 0.00346941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_D_M1012_g 0.0223425f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_50 VPB N_D_c_262_n 0.00420406f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_51 VPB N_C_M1010_g 0.0204101f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_52 VPB C 5.95777e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_C_c_305_n 0.00453286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_B_M1006_g 0.0223915f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_55 VPB B 0.00197506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_B_c_339_n 0.0045624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_M1000_g 0.0230296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_375_n 0.029221f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_59 VPB N_A_27_47#_c_381_n 0.0147617f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_60 VPB N_A_27_47#_c_382_n 0.00224522f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.85
cc_61 VPB N_A_27_47#_c_376_n 0.00695368f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.19
cc_62 VPB N_A_27_47#_c_377_n 0.0119156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_385_n 0.0110158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_451_n 0.00215067f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=0.995
cc_65 VPB N_VPWR_c_452_n 3.11529e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_453_n 0.00272466f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.53
cc_67 VPB N_VPWR_c_454_n 0.00281836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_455_n 0.010303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_456_n 0.0131478f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_457_n 0.0234027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_458_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_459_n 0.014294f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_460_n 0.0143676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_461_n 0.011815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_462_n 0.021623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_463_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_464_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_465_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_450_n 0.0437233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB X 0.00152769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 N_A_N_M1016_g N_A_174_21#_c_116_n 0.019384f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_82 A_N N_A_174_21#_c_116_n 0.00690255f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A_N_M1009_g N_A_174_21#_M1001_g 0.0348904f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_84 N_A_N_c_84_n N_A_174_21#_c_120_n 0.0216014f $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_N_M1016_g N_A_27_47#_c_375_n 0.0104714f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_N_M1009_g N_A_27_47#_c_375_n 0.0161698f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_87 A_N N_A_27_47#_c_375_n 0.0629743f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_N_c_84_n N_A_27_47#_c_375_n 0.00749129f $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_N_M1009_g N_A_27_47#_c_382_n 0.0150223f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_90 A_N N_A_27_47#_c_382_n 0.0192865f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_91 N_A_N_c_84_n N_A_27_47#_c_382_n 5.33633e-19 $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_92 A_N N_VPWR_M1009_d 0.00411499f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_93 N_A_N_M1009_g N_VPWR_c_451_n 0.00832549f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_94 N_A_N_M1009_g N_VPWR_c_459_n 0.00339367f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_95 N_A_N_M1009_g N_VPWR_c_450_n 0.00489827f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_96 N_A_N_M1016_g X 6.02166e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_97 A_N X 0.00417494f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A_N_M1009_g N_X_c_533_n 4.58489e-19 $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_99 A_N N_X_c_533_n 0.00683172f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_100 A_N X 0.0520765f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_101 N_A_N_c_84_n X 2.76793e-19 $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_102 A_N N_VGND_M1016_d 0.00356045f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_103 N_A_N_M1016_g N_VGND_c_575_n 0.00310635f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_104 A_N N_VGND_c_575_n 0.010711f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A_N_c_84_n N_VGND_c_575_n 3.38996e-19 $X=0.525 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_N_M1016_g N_VGND_c_578_n 0.00585385f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_N_M1016_g N_VGND_c_582_n 0.00841565f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_108 A_N N_VGND_c_582_n 0.00573938f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_109 N_A_174_21#_M1014_g N_D_M1012_g 0.0163059f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_174_21#_c_122_n N_D_M1012_g 0.00404479f $X=2.465 $Y=1.545 $X2=0 $Y2=0
cc_111 N_A_174_21#_c_137_p N_D_M1012_g 0.010157f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_112 N_A_174_21#_c_120_n D 3.44722e-19 $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_174_21#_c_121_n D 0.0036248f $X=2.465 $Y=1.075 $X2=0 $Y2=0
cc_114 N_A_174_21#_c_122_n D 0.0036248f $X=2.465 $Y=1.545 $X2=0 $Y2=0
cc_115 N_A_174_21#_c_141_p D 0.00466771f $X=2.795 $Y=0.7 $X2=0 $Y2=0
cc_116 N_A_174_21#_c_137_p D 0.0112164f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_117 N_A_174_21#_c_123_n D 0.00339299f $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_118 N_A_174_21#_c_124_n D 0.00885165f $X=2.465 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_174_21#_c_120_n N_D_c_262_n 0.0099699f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_174_21#_c_121_n N_D_c_262_n 5.86652e-19 $X=2.465 $Y=1.075 $X2=0 $Y2=0
cc_121 N_A_174_21#_c_122_n N_D_c_262_n 5.86652e-19 $X=2.465 $Y=1.545 $X2=0 $Y2=0
cc_122 N_A_174_21#_c_141_p N_D_c_262_n 0.00342681f $X=2.795 $Y=0.7 $X2=0 $Y2=0
cc_123 N_A_174_21#_c_137_p N_D_c_262_n 0.0031544f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_124 N_A_174_21#_c_124_n N_D_c_262_n 0.00144066f $X=2.465 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_174_21#_c_119_n N_D_c_263_n 0.00856086f $X=2.205 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_174_21#_c_121_n N_D_c_263_n 0.0038601f $X=2.465 $Y=1.075 $X2=0 $Y2=0
cc_127 N_A_174_21#_c_141_p N_D_c_263_n 0.00698434f $X=2.795 $Y=0.7 $X2=0 $Y2=0
cc_128 N_A_174_21#_c_154_p N_D_c_263_n 0.00439001f $X=2.88 $Y=0.615 $X2=0 $Y2=0
cc_129 N_A_174_21#_c_123_n N_D_c_263_n 0.00807289f $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_130 N_A_174_21#_c_156_p N_D_c_263_n 0.00306115f $X=2.965 $Y=0.385 $X2=0 $Y2=0
cc_131 N_A_174_21#_c_141_p N_C_c_303_n 7.19629e-19 $X=2.795 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A_174_21#_c_154_p N_C_c_303_n 7.17948e-19 $X=2.88 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_174_21#_c_123_n N_C_c_303_n 0.0112299f $X=4.39 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_174_21#_c_137_p N_C_M1010_g 0.00956284f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_135 N_A_174_21#_c_137_p C 0.0110571f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_136 N_A_174_21#_c_123_n C 0.00663419f $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_137 N_A_174_21#_c_137_p N_C_c_305_n 0.00128696f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_138 N_A_174_21#_c_123_n N_C_c_305_n 9.36849e-19 $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_139 N_A_174_21#_c_137_p N_B_M1006_g 0.0123442f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_140 N_A_174_21#_c_137_p B 0.0175693f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_141 N_A_174_21#_c_123_n B 0.0152421f $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_142 N_A_174_21#_c_137_p N_B_c_339_n 0.00213304f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_143 N_A_174_21#_c_123_n N_B_c_339_n 0.00149287f $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_144 N_A_174_21#_c_123_n N_B_c_340_n 0.0182249f $X=4.39 $Y=0.385 $X2=0 $Y2=0
cc_145 N_A_174_21#_c_123_n N_A_27_47#_c_374_n 0.0215854f $X=4.39 $Y=0.385 $X2=0
+ $Y2=0
cc_146 N_A_174_21#_c_137_p N_A_27_47#_M1000_g 0.00363421f $X=4.38 $Y=1.63 $X2=0
+ $Y2=0
cc_147 N_A_174_21#_M1012_d N_A_27_47#_c_382_n 0.00446851f $X=3.085 $Y=1.485
+ $X2=0 $Y2=0
cc_148 N_A_174_21#_M1006_d N_A_27_47#_c_382_n 0.0100877f $X=4.075 $Y=1.485 $X2=0
+ $Y2=0
cc_149 N_A_174_21#_M1001_g N_A_27_47#_c_382_n 0.0154059f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_174_21#_M1003_g N_A_27_47#_c_382_n 0.0116333f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_174_21#_M1013_g N_A_27_47#_c_382_n 0.0116333f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_174_21#_M1014_g N_A_27_47#_c_382_n 0.0147431f $X=2.205 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_174_21#_c_179_p N_A_27_47#_c_382_n 0.00420617f $X=2.38 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_174_21#_c_120_n N_A_27_47#_c_382_n 0.00197266f $X=2.285 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_174_21#_c_181_p N_A_27_47#_c_382_n 0.0121736f $X=2.55 $Y=1.63 $X2=0
+ $Y2=0
cc_156 N_A_174_21#_c_137_p N_A_27_47#_c_382_n 0.100306f $X=4.38 $Y=1.63 $X2=0
+ $Y2=0
cc_157 N_A_174_21#_c_137_p N_A_27_47#_c_376_n 0.0123627f $X=4.38 $Y=1.63 $X2=0
+ $Y2=0
cc_158 N_A_174_21#_c_123_n N_A_27_47#_c_376_n 0.0134493f $X=4.39 $Y=0.385 $X2=0
+ $Y2=0
cc_159 N_A_174_21#_c_123_n N_A_27_47#_c_377_n 0.00492599f $X=4.39 $Y=0.385 $X2=0
+ $Y2=0
cc_160 N_A_174_21#_c_122_n N_VPWR_M1014_d 0.00184028f $X=2.465 $Y=1.545 $X2=0
+ $Y2=0
cc_161 N_A_174_21#_c_181_p N_VPWR_M1014_d 0.00518332f $X=2.55 $Y=1.63 $X2=0
+ $Y2=0
cc_162 N_A_174_21#_c_137_p N_VPWR_M1014_d 0.0164292f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_163 N_A_174_21#_c_137_p N_VPWR_M1010_d 0.0142491f $X=4.38 $Y=1.63 $X2=0 $Y2=0
cc_164 N_A_174_21#_M1001_g N_VPWR_c_451_n 0.0016047f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_174_21#_M1001_g N_VPWR_c_452_n 0.00114039f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_174_21#_M1003_g N_VPWR_c_452_n 0.00842528f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_174_21#_M1013_g N_VPWR_c_452_n 0.00810864f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_174_21#_M1014_g N_VPWR_c_452_n 0.00110281f $X=2.205 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_174_21#_M1013_g N_VPWR_c_453_n 0.00110281f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_174_21#_M1014_g N_VPWR_c_453_n 0.00873606f $X=2.205 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_174_21#_M1001_g N_VPWR_c_460_n 0.00425094f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_174_21#_M1003_g N_VPWR_c_460_n 0.00339367f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_174_21#_M1013_g N_VPWR_c_461_n 0.00339367f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_174_21#_M1014_g N_VPWR_c_461_n 0.00339367f $X=2.205 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_174_21#_M1012_d N_VPWR_c_450_n 0.00315309f $X=3.085 $Y=1.485 $X2=0
+ $Y2=0
cc_176 N_A_174_21#_M1006_d N_VPWR_c_450_n 0.00515182f $X=4.075 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A_174_21#_M1001_g N_VPWR_c_450_n 0.00580516f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_174_21#_M1003_g N_VPWR_c_450_n 0.00398704f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_174_21#_M1013_g N_VPWR_c_450_n 0.00398704f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_174_21#_M1014_g N_VPWR_c_450_n 0.00398704f $X=2.205 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_174_21#_c_117_n N_X_c_537_n 0.0160528f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_174_21#_c_118_n N_X_c_537_n 0.0115365f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_174_21#_c_179_p N_X_c_537_n 0.0286246f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_174_21#_c_120_n N_X_c_537_n 0.00427833f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_174_21#_M1003_g N_X_c_541_n 0.0131115f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_174_21#_M1013_g N_X_c_541_n 0.00929518f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_174_21#_M1014_g N_X_c_541_n 0.00304053f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_174_21#_c_179_p N_X_c_541_n 0.0267852f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_174_21#_c_120_n N_X_c_541_n 0.00404946f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_174_21#_c_181_p N_X_c_541_n 0.0120185f $X=2.55 $Y=1.63 $X2=0 $Y2=0
cc_191 N_A_174_21#_c_116_n X 0.00604018f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_174_21#_M1001_g N_X_c_533_n 0.00338f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_174_21#_c_116_n X 0.00360971f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_174_21#_M1001_g X 0.00399679f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_174_21#_c_117_n X 0.0032178f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_174_21#_M1003_g X 0.0042867f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_174_21#_c_179_p X 0.0126559f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_174_21#_c_120_n X 0.0253785f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_174_21#_c_121_n N_VGND_M1017_s 0.00270979f $X=2.465 $Y=1.075 $X2=0
+ $Y2=0
cc_200 N_A_174_21#_c_141_p N_VGND_M1017_s 0.0165267f $X=2.795 $Y=0.7 $X2=0 $Y2=0
cc_201 N_A_174_21#_c_227_p N_VGND_M1017_s 0.00521187f $X=2.55 $Y=0.7 $X2=0 $Y2=0
cc_202 N_A_174_21#_c_154_p N_VGND_M1017_s 0.0022319f $X=2.88 $Y=0.615 $X2=0
+ $Y2=0
cc_203 N_A_174_21#_c_156_p N_VGND_M1017_s 0.0028145f $X=2.965 $Y=0.385 $X2=0
+ $Y2=0
cc_204 N_A_174_21#_c_116_n N_VGND_c_575_n 0.00769236f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_174_21#_c_117_n N_VGND_c_575_n 5.10275e-19 $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_174_21#_c_116_n N_VGND_c_576_n 5.10275e-19 $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_174_21#_c_117_n N_VGND_c_576_n 0.00670862f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_174_21#_c_118_n N_VGND_c_576_n 0.00679166f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_A_174_21#_c_119_n N_VGND_c_576_n 5.249e-19 $X=2.205 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_174_21#_c_119_n N_VGND_c_577_n 0.00212296f $X=2.205 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_174_21#_c_179_p N_VGND_c_577_n 0.00175693f $X=2.38 $Y=1.16 $X2=0
+ $Y2=0
cc_212 N_A_174_21#_c_120_n N_VGND_c_577_n 0.00173549f $X=2.285 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_174_21#_c_141_p N_VGND_c_577_n 0.00481916f $X=2.795 $Y=0.7 $X2=0
+ $Y2=0
cc_214 N_A_174_21#_c_227_p N_VGND_c_577_n 0.0142335f $X=2.55 $Y=0.7 $X2=0 $Y2=0
cc_215 N_A_174_21#_c_156_p N_VGND_c_577_n 0.0118319f $X=2.965 $Y=0.385 $X2=0
+ $Y2=0
cc_216 N_A_174_21#_c_116_n N_VGND_c_579_n 0.00424334f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_174_21#_c_117_n N_VGND_c_579_n 0.00341112f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_174_21#_c_118_n N_VGND_c_580_n 0.00341112f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_174_21#_c_119_n N_VGND_c_580_n 0.00585385f $X=2.205 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_174_21#_c_141_p N_VGND_c_581_n 0.00327636f $X=2.795 $Y=0.7 $X2=0
+ $Y2=0
cc_221 N_A_174_21#_c_123_n N_VGND_c_581_n 0.0909063f $X=4.39 $Y=0.385 $X2=0
+ $Y2=0
cc_222 N_A_174_21#_c_156_p N_VGND_c_581_n 0.00755799f $X=2.965 $Y=0.385 $X2=0
+ $Y2=0
cc_223 N_A_174_21#_M1005_d N_VGND_c_582_n 0.00212021f $X=4.665 $Y=0.235 $X2=0
+ $Y2=0
cc_224 N_A_174_21#_c_116_n N_VGND_c_582_n 0.0066176f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_174_21#_c_117_n N_VGND_c_582_n 0.00397316f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_174_21#_c_118_n N_VGND_c_582_n 0.00397316f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_174_21#_c_119_n N_VGND_c_582_n 0.0111361f $X=2.205 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_174_21#_c_141_p N_VGND_c_582_n 0.00550808f $X=2.795 $Y=0.7 $X2=0
+ $Y2=0
cc_229 N_A_174_21#_c_227_p N_VGND_c_582_n 8.89004e-19 $X=2.55 $Y=0.7 $X2=0 $Y2=0
cc_230 N_A_174_21#_c_123_n N_VGND_c_582_n 0.0702723f $X=4.39 $Y=0.385 $X2=0
+ $Y2=0
cc_231 N_A_174_21#_c_156_p N_VGND_c_582_n 0.00619596f $X=2.965 $Y=0.385 $X2=0
+ $Y2=0
cc_232 N_A_174_21#_c_123_n A_617_47# 0.00745008f $X=4.39 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_174_21#_c_123_n A_701_47# 0.0139731f $X=4.39 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_234 N_A_174_21#_c_123_n A_815_47# 0.021069f $X=4.39 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_235 N_D_c_263_n N_C_c_303_n 0.0420833f $X=2.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_236 N_D_M1012_g N_C_M1010_g 0.0477337f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_237 D C 0.0164762f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_238 N_D_c_262_n C 3.87016e-19 $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_239 N_D_c_263_n C 0.00245204f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_240 D N_C_c_305_n 0.00114946f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_241 N_D_c_262_n N_C_c_305_n 0.0204558f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_242 N_D_M1012_g N_A_27_47#_c_382_n 0.0133167f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_243 N_D_M1012_g N_VPWR_c_453_n 0.00674465f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_244 N_D_M1012_g N_VPWR_c_454_n 0.00217739f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_245 N_D_M1012_g N_VPWR_c_457_n 0.00425094f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_246 N_D_M1012_g N_VPWR_c_450_n 0.00664448f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_247 N_D_c_263_n N_VGND_c_577_n 0.0038505f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_248 N_D_c_263_n N_VGND_c_581_n 0.00367079f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_249 N_D_c_263_n N_VGND_c_582_n 0.00604949f $X=2.95 $Y=0.995 $X2=0 $Y2=0
cc_250 N_C_M1010_g N_B_M1006_g 0.0335271f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_251 N_C_c_303_n B 0.00131718f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_252 C B 0.0288138f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_253 N_C_c_305_n B 0.0024156f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_254 C N_B_c_339_n 3.57638e-19 $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_255 N_C_c_305_n N_B_c_339_n 0.0100722f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_256 N_C_c_303_n N_B_c_340_n 0.026681f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_257 C N_B_c_340_n 4.25482e-19 $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_258 N_C_M1010_g N_A_27_47#_c_382_n 0.0123f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_259 N_C_M1010_g N_VPWR_c_454_n 0.00975985f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_260 N_C_M1010_g N_VPWR_c_457_n 0.00339367f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_261 N_C_M1010_g N_VPWR_c_450_n 0.00401529f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_262 N_C_c_303_n N_VGND_c_581_n 0.00367119f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_263 N_C_c_303_n N_VGND_c_582_n 0.00567582f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_264 B N_A_27_47#_c_374_n 0.0038936f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_265 N_B_c_340_n N_A_27_47#_c_374_n 0.0218381f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_266 N_B_M1006_g N_A_27_47#_M1000_g 0.0317126f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_267 N_B_M1006_g N_A_27_47#_c_382_n 0.0134303f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_268 B N_A_27_47#_c_376_n 0.00849438f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_269 N_B_c_339_n N_A_27_47#_c_376_n 9.44974e-19 $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_270 B N_A_27_47#_c_377_n 0.00139934f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_271 N_B_c_339_n N_A_27_47#_c_377_n 0.0129363f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B_M1006_g N_VPWR_c_454_n 0.00874184f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B_M1006_g N_VPWR_c_456_n 0.00186865f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B_M1006_g N_VPWR_c_462_n 0.00425094f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B_M1006_g N_VPWR_c_450_n 0.00664632f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B_c_340_n N_VGND_c_581_n 0.00367119f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B_c_340_n N_VGND_c_582_n 0.00605146f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_278 B A_701_47# 0.00235594f $X=3.83 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_279 B A_815_47# 0.0020738f $X=3.83 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_280 N_A_27_47#_c_382_n N_VPWR_M1009_d 0.00527527f $X=4.73 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_281 N_A_27_47#_c_382_n N_VPWR_M1003_d 0.00328325f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_382_n N_VPWR_M1014_d 0.0167112f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_382_n N_VPWR_M1010_d 0.00759276f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_382_n N_VPWR_M1000_d 0.0101627f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_376_n N_VPWR_M1000_d 0.0233341f $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_382_n N_VPWR_c_451_n 0.0181288f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_382_n N_VPWR_c_452_n 0.0159625f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_382_n N_VPWR_c_453_n 0.020494f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_382_n N_VPWR_c_454_n 0.020494f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_290 N_A_27_47#_M1000_g N_VPWR_c_456_n 0.0112146f $X=4.59 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_382_n N_VPWR_c_456_n 0.016853f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_382_n N_VPWR_c_457_n 0.0140184f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_381_n N_VPWR_c_459_n 0.0179169f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_382_n N_VPWR_c_459_n 0.00244309f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_382_n N_VPWR_c_460_n 0.00848923f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_382_n N_VPWR_c_461_n 0.0077537f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_297 N_A_27_47#_M1000_g N_VPWR_c_462_n 0.00339367f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_382_n N_VPWR_c_462_n 0.0128806f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_299 N_A_27_47#_M1009_s N_VPWR_c_450_n 0.00226392f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1000_g N_VPWR_c_450_n 0.00439092f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_381_n N_VPWR_c_450_n 0.00991829f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_382_n N_VPWR_c_450_n 0.0855204f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_382_n N_X_M1001_s 0.00440505f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_382_n N_X_M1013_s 0.00440866f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_382_n N_X_c_541_n 0.0396402f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_382_n N_X_c_533_n 0.0138435f $X=4.73 $Y=2 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_378_n N_VGND_c_578_n 0.0177247f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_374_n N_VGND_c_581_n 0.00366918f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1016_s N_VGND_c_582_n 0.00382897f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_374_n N_VGND_c_582_n 0.00660056f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_378_n N_VGND_c_582_n 0.00987844f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_312 N_VPWR_c_450_n N_X_M1001_s 0.00315309f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_313 N_VPWR_c_450_n N_X_M1013_s 0.00315309f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_M1003_d N_X_c_541_n 0.00366235f $X=1.44 $Y=1.485 $X2=0 $Y2=0
cc_315 N_X_c_537_n N_VGND_M1004_s 0.00336712f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_316 N_X_c_537_n N_VGND_c_576_n 0.0152323f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_317 N_X_c_564_p N_VGND_c_579_n 0.0113958f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_318 N_X_c_537_n N_VGND_c_579_n 0.00216966f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_319 X N_VGND_c_579_n 0.00116615f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_320 N_X_c_537_n N_VGND_c_580_n 0.00235782f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_321 N_X_c_568_p N_VGND_c_580_n 0.0112485f $X=1.995 $Y=0.42 $X2=0 $Y2=0
cc_322 N_X_M1002_d N_VGND_c_582_n 0.00251375f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_323 N_X_M1007_d N_VGND_c_582_n 0.00406917f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_324 N_X_c_564_p N_VGND_c_582_n 0.00646998f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_325 N_X_c_537_n N_VGND_c_582_n 0.009166f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_326 N_X_c_568_p N_VGND_c_582_n 0.0064389f $X=1.995 $Y=0.42 $X2=0 $Y2=0
cc_327 X N_VGND_c_582_n 0.00302698f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_328 N_VGND_c_582_n A_617_47# 0.00219724f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_329 N_VGND_c_582_n A_701_47# 0.00342801f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_330 N_VGND_c_582_n A_815_47# 0.00358554f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24

* NGSPICE file created from sky130_fd_sc_hd__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u
M1001 Y A a_113_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_113_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1003 VPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__nand2b_4.spice
* Created: Thu Aug 27 14:29:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand2b_4.spice.pex"
.subckt sky130_fd_sc_hd__nand2b_4  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_A_N_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_215_47#_M1002_d N_A_27_47#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1003 N_A_215_47#_M1003_d N_A_27_47#_M1003_g N_Y_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1007 N_A_215_47#_M1003_d N_A_27_47#_M1007_g N_Y_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1010 N_A_215_47#_M1010_d N_A_27_47#_M1010_g N_Y_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.092625 AS=0.08775 PD=0.935 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75002 A=0.0975 P=1.6 MULT=1
MM1004 N_A_215_47#_M1010_d N_B_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.08775 PD=0.935 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_215_47#_M1008_d N_B_M1008_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_215_47#_M1008_d N_B_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_A_215_47#_M1013_d N_B_M1013_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2535 AS=0.08775 PD=2.08 PS=0.92 NRD=19.38 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_N_M1014_g N_A_27_47#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_27_47#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.3 A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1000_d N_A_27_47#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1015_d N_A_27_47#_M1015_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1016 N_Y_M1015_d N_A_27_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1425 PD=1.27 PS=1.285 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75001.4
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.1425 PD=1.27 PS=1.285 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75001.6
+ A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1001_d N_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75001.2
+ A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1009 N_Y_M1006_d N_B_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.39 PD=1.27 PS=2.78 NRD=0 NRS=20.685 M=1 R=6.66667 SA=75003.1 SB=75000.3
+ A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hd__nand2b_4.spice.SKY130_FD_SC_HD__NAND2B_4.pxi"
*
.ends
*
*

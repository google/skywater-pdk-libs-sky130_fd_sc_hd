# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__a31oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__a31oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 0.995000 5.420000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 3.550000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 1.735000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.670000 0.995000 6.855000 1.630000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.443500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.635000 7.585000 0.805000 ;
        RECT 6.075000 1.915000 7.245000 2.085000 ;
        RECT 6.575000 0.255000 6.745000 0.635000 ;
        RECT 7.045000 0.805000 7.245000 1.915000 ;
        RECT 7.415000 0.255000 7.585000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.355000  0.085000 1.685000 0.465000 ;
        RECT 6.075000  0.085000 6.405000 0.465000 ;
        RECT 6.915000  0.085000 7.245000 0.465000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.515000 1.915000 0.845000 2.635000 ;
        RECT 1.355000 1.915000 1.685000 2.635000 ;
        RECT 2.195000 1.915000 2.525000 2.635000 ;
        RECT 3.035000 1.915000 3.365000 2.635000 ;
        RECT 3.895000 1.915000 4.225000 2.635000 ;
        RECT 4.735000 2.255000 5.065000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.255000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 3.785000 0.805000 ;
      RECT 0.175000 1.495000 5.405000 1.665000 ;
      RECT 0.175000 1.665000 0.345000 2.465000 ;
      RECT 1.015000 0.255000 1.185000 0.635000 ;
      RECT 1.015000 1.665000 1.185000 2.465000 ;
      RECT 1.855000 0.255000 2.025000 0.635000 ;
      RECT 1.855000 1.665000 2.025000 2.465000 ;
      RECT 2.195000 0.295000 5.565000 0.465000 ;
      RECT 2.695000 1.665000 2.865000 2.465000 ;
      RECT 3.535000 1.665000 3.705000 2.465000 ;
      RECT 4.395000 1.665000 4.565000 2.465000 ;
      RECT 5.235000 1.665000 5.405000 2.255000 ;
      RECT 5.235000 2.255000 7.665000 2.425000 ;
      RECT 5.235000 2.425000 5.405000 2.465000 ;
      RECT 7.415000 1.495000 7.665000 2.255000 ;
  END
END sky130_fd_sc_hd__a31oi_4

* File: sky130_fd_sc_hd__mux2_2.pex.spice
* Created: Tue Sep  1 19:14:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2_2%A_79_21# 1 2 7 9 12 14 16 19 24 25 26 27 28
+ 30 32 33 35 37 39 42 43 44
r121 46 48 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r122 43 48 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.94 $Y=1.16 $X2=0.89
+ $Y2=1.16
r123 42 45 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.16
+ $X2=1.01 $Y2=1.325
r124 42 44 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.16
+ $X2=1.01 $Y2=0.995
r125 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r126 37 39 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=1.655 $Y=2.34
+ $X2=2.63 $Y2=2.34
r127 33 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.605 $Y=0.38
+ $X2=2.565 $Y2=0.38
r128 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=2.255
+ $X2=1.655 $Y2=2.34
r129 31 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.57 $Y=2.005
+ $X2=1.57 $Y2=2.255
r130 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.52 $Y=0.465
+ $X2=1.605 $Y2=0.38
r131 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.52 $Y=0.465
+ $X2=1.52 $Y2=0.635
r132 27 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=1.92
+ $X2=1.57 $Y2=2.005
r133 27 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.485 $Y=1.92
+ $X2=1.165 $Y2=1.92
r134 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=1.52 $Y2=0.635
r135 25 26 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=1.165 $Y2=0.72
r136 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.08 $Y=1.835
+ $X2=1.165 $Y2=1.92
r137 24 45 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.08 $Y=1.835
+ $X2=1.08 $Y2=1.325
r138 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.08 $Y=0.805
+ $X2=1.165 $Y2=0.72
r139 21 44 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.08 $Y=0.805
+ $X2=1.08 $Y2=0.995
r140 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r141 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r142 14 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r143 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r144 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r145 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r146 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r147 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r148 2 39 600 $w=1.7e-07 $l=6.01124e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.845 $X2=2.63 $Y2=2.34
r149 1 35 91 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.235 $X2=2.565 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%A_257_199# 1 2 9 13 17 18 20 21 23 24 25 30
+ 33
c91 25 0 1.28281e-19 $X=1.995 $Y=1.92
c92 13 0 3.54659e-20 $X=1.455 $Y=2.165
r93 28 33 2.86771 $w=3.32e-07 $l=8.6487e-08 $layer=LI1_cond $X=3.885 $Y=1.835
+ $X2=3.882 $Y2=1.92
r94 28 30 49.4154 $w=3.28e-07 $l=1.415e-06 $layer=LI1_cond $X=3.885 $Y=1.835
+ $X2=3.885 $Y2=0.42
r95 24 33 3.83825 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.715 $Y=1.92
+ $X2=3.882 $Y2=1.92
r96 24 25 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=3.715 $Y=1.92
+ $X2=1.995 $Y2=1.92
r97 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.91 $Y=1.835
+ $X2=1.995 $Y2=1.92
r98 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.91 $Y=1.665
+ $X2=1.91 $Y2=1.835
r99 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.825 $Y=1.58
+ $X2=1.91 $Y2=1.665
r100 20 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.825 $Y=1.58
+ $X2=1.505 $Y2=1.58
r101 18 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=1.42 $Y2=1.325
r102 18 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=1.42 $Y2=0.995
r103 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.16 $X2=1.42 $Y2=1.16
r104 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=1.495
+ $X2=1.505 $Y2=1.58
r105 15 17 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.42 $Y=1.495
+ $X2=1.42 $Y2=1.16
r106 13 36 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.455 $Y=2.165
+ $X2=1.455 $Y2=1.325
r107 9 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.365 $Y=0.445
+ $X2=1.365 $Y2=0.995
r108 2 33 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=3.735
+ $Y=1.845 $X2=3.88 $Y2=2
r109 1 30 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.235 $X2=3.88 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%A0 3 6 8 9 10 11 17 19 25
c51 25 0 1.53841e-19 $X=2.88 $Y=1.42
c52 9 0 1.50818e-19 $X=2.075 $Y=1.19
r53 22 25 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.79 $Y=1.42 $X2=2.88
+ $Y2=1.42
r54 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.42 $X2=2.79 $Y2=1.42
r55 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=0.93 $X2=1.9
+ $Y2=0.765
r56 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9
+ $Y=0.93 $X2=1.9 $Y2=0.93
r57 11 23 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=2.995 $Y=1.47
+ $X2=2.79 $Y2=1.47
r58 10 23 9.47977 $w=3.08e-07 $l=2.55e-07 $layer=LI1_cond $X=2.535 $Y=1.47
+ $X2=2.79 $Y2=1.47
r59 10 27 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=2.535 $Y=1.47 $X2=2.445
+ $Y2=1.47
r60 9 27 7.6764 $w=4.45e-07 $l=4.32926e-07 $layer=LI1_cond $X=2.13 $Y=1.19
+ $X2=2.445 $Y2=1.47
r61 9 18 7.12809 $w=4.45e-07 $l=2.6e-07 $layer=LI1_cond $X=2.13 $Y=1.19 $X2=2.13
+ $Y2=0.93
r62 8 18 2.19326 $w=4.45e-07 $l=8e-08 $layer=LI1_cond $X=2.13 $Y=0.85 $X2=2.13
+ $Y2=0.93
r63 4 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.88 $Y=1.555
+ $X2=2.88 $Y2=1.42
r64 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.88 $Y=1.555 $X2=2.88
+ $Y2=2.165
r65 3 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.84 $Y=0.445
+ $X2=1.84 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%A1 3 5 6 9 11 12 16
c53 9 0 1.50818e-19 $X=2.815 $Y=0.445
r54 16 19 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.79 $Y=0.94 $X2=2.79
+ $Y2=1
r55 16 18 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.79 $Y=0.94
+ $X2=2.79 $Y2=0.805
r56 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=0.94 $X2=2.79 $Y2=0.94
r57 12 17 8.14658 $w=2.88e-07 $l=2.05e-07 $layer=LI1_cond $X=2.995 $Y=0.88
+ $X2=2.79 $Y2=0.88
r58 12 21 3.21194 $w=1.9e-07 $l=1.45e-07 $layer=LI1_cond $X=2.995 $Y=0.88
+ $X2=2.995 $Y2=0.735
r59 11 21 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=2.995 $Y=0.51
+ $X2=2.995 $Y2=0.735
r60 9 18 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.815 $Y=0.445
+ $X2=2.815 $Y2=0.805
r61 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1 $X2=2.79
+ $Y2=1
r62 5 6 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.625 $Y=1 $X2=2.395
+ $Y2=1
r63 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.32 $Y=1.075
+ $X2=2.395 $Y2=1
r64 1 3 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=2.32 $Y=1.075
+ $X2=2.32 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%S 3 7 11 15 17 18 19 28
c45 17 0 1.53841e-19 $X=3.455 $Y=0.85
r46 26 28 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.455 $Y=1.16
+ $X2=3.66 $Y2=1.16
r47 23 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.24 $Y=1.16
+ $X2=3.455 $Y2=1.16
r48 18 19 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.455 $Y2=1.53
r49 18 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.455
+ $Y=1.16 $X2=3.455 $Y2=1.16
r50 17 18 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=3.455 $Y=0.85
+ $X2=3.455 $Y2=1.16
r51 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.325
+ $X2=3.66 $Y2=1.16
r52 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.66 $Y=1.325
+ $X2=3.66 $Y2=2.165
r53 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=0.995
+ $X2=3.66 $Y2=1.16
r54 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.66 $Y=0.995
+ $X2=3.66 $Y2=0.445
r55 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.325
+ $X2=3.24 $Y2=1.16
r56 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.24 $Y=1.325 $X2=3.24
+ $Y2=2.165
r57 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=0.995
+ $X2=3.24 $Y2=1.16
r58 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.24 $Y=0.995 $X2=3.24
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%VPWR 1 2 3 10 12 18 22 24 26 31 41 42 48 51
r61 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 39 51 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.545 $Y=2.72
+ $X2=3.435 $Y2=2.72
r66 39 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.545 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 32 48 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.315 $Y=2.72
+ $X2=1.17 $Y2=2.72
r74 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.315 $Y=2.72
+ $X2=1.61 $Y2=2.72
r75 31 51 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.435 $Y2=2.72
r76 31 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 30 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 27 45 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r80 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 26 48 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=1.17 $Y2=2.72
r82 26 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r84 24 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 20 51 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.435 $Y=2.635
+ $X2=3.435 $Y2=2.72
r86 20 22 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.435 $Y=2.635
+ $X2=3.435 $Y2=2.34
r87 16 48 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=2.635
+ $X2=1.17 $Y2=2.72
r88 16 18 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.17 $Y=2.635
+ $X2=1.17 $Y2=2.34
r89 12 15 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r90 10 45 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r91 10 15 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r92 3 22 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.845 $X2=3.45 $Y2=2.34
r93 2 18 600 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.15 $Y2=2.34
r94 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r95 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%X 1 2 9 13 14 15 16 17
c27 14 0 3.54659e-20 $X=0.67 $Y=1.75
r28 17 23 9.29389 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=0.67 $Y=2.21
+ $X2=0.67 $Y2=1.96
r29 16 23 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=0.67 $Y=1.87 $X2=0.67
+ $Y2=1.96
r30 14 16 4.46107 $w=3.08e-07 $l=1.2e-07 $layer=LI1_cond $X=0.67 $Y=1.75
+ $X2=0.67 $Y2=1.87
r31 14 15 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.67 $Y=1.75
+ $X2=0.67 $Y2=1.595
r32 13 15 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.6 $Y=0.75 $X2=0.6
+ $Y2=1.595
r33 7 13 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.64 $Y=0.625
+ $X2=0.64 $Y2=0.75
r34 7 9 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.64 $Y=0.625
+ $X2=0.64 $Y2=0.42
r35 2 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
r36 1 9 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r61 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r62 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 40 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r64 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r65 37 49 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.45
+ $Y2=0
r66 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.91
+ $Y2=0
r67 36 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r68 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r69 33 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r70 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r71 32 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r72 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r73 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r74 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r75 29 49 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.45
+ $Y2=0
r76 29 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=2.99
+ $Y2=0
r77 28 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r78 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r79 25 43 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r80 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r81 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r82 24 27 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r83 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r84 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r85 18 49 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=0.085 $X2=3.45
+ $Y2=0
r86 18 20 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.45 $Y=0.085
+ $X2=3.45 $Y2=0.42
r87 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r88 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r89 10 43 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r90 10 12 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.38
r91 3 20 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.315
+ $Y=0.235 $X2=3.45 $Y2=0.42
r92 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r93 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


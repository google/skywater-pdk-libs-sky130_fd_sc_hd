* File: sky130_fd_sc_hd__and2_0.spice
* Created: Thu Aug 27 14:06:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and2_0.pex.spice"
.subckt sky130_fd_sc_hd__and2_0  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_123_47# N_A_M1001_g N_A_40_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g A_123_47# VNB NSHORT L=0.15 W=0.42 AD=0.0966
+ AS=0.0441 PD=0.88 PS=0.63 NRD=18.564 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_40_47#_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0966 PD=1.37 PS=0.88 NRD=0 NRS=32.856 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_40_47#_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0609 AS=0.1113 PD=0.71 PS=1.37 NRD=4.6886 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_40_47#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.145891 AS=0.0609 PD=0.998491 PS=0.71 NRD=78.5636 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_40_47#_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.222309 PD=1.81 PS=1.52151 NRD=0 NRS=1.5366 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__and2_0.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a2bb2oi_1.pxi.spice
* Created: Tue Sep  1 18:54:09 2020
* 
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%A1_N N_A1_N_M1008_g N_A1_N_M1007_g A1_N A1_N
+ N_A1_N_c_58_n N_A1_N_c_59_n N_A1_N_c_60_n PM_SKY130_FD_SC_HD__A2BB2OI_1%A1_N
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%A2_N N_A2_N_M1005_g N_A2_N_c_85_n N_A2_N_M1006_g
+ A2_N N_A2_N_c_87_n A2_N PM_SKY130_FD_SC_HD__A2BB2OI_1%A2_N
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%A_109_47# N_A_109_47#_M1008_d
+ N_A_109_47#_M1005_d N_A_109_47#_c_119_n N_A_109_47#_M1002_g
+ N_A_109_47#_M1003_g N_A_109_47#_c_120_n N_A_109_47#_c_121_n
+ N_A_109_47#_c_180_p N_A_109_47#_c_135_n N_A_109_47#_c_138_n
+ N_A_109_47#_c_126_n N_A_109_47#_c_127_n N_A_109_47#_c_128_n
+ N_A_109_47#_c_122_n PM_SKY130_FD_SC_HD__A2BB2OI_1%A_109_47#
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%B2 N_B2_c_189_n N_B2_M1001_g N_B2_M1000_g B2 B2
+ B2 B2 N_B2_c_192_n B2 PM_SKY130_FD_SC_HD__A2BB2OI_1%B2
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%B1 N_B1_M1004_g N_B1_M1009_g B1 N_B1_c_236_n
+ N_B1_c_237_n PM_SKY130_FD_SC_HD__A2BB2OI_1%B1
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%VPWR N_VPWR_M1007_s N_VPWR_M1000_d
+ N_VPWR_c_265_n VPWR VPWR N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_264_n
+ N_VPWR_c_270_n N_VPWR_c_271_n PM_SKY130_FD_SC_HD__A2BB2OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%Y N_Y_M1002_d N_Y_M1003_s N_Y_c_308_n Y Y Y
+ PM_SKY130_FD_SC_HD__A2BB2OI_1%Y
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%A_397_297# N_A_397_297#_M1003_d
+ N_A_397_297#_M1009_d N_A_397_297#_c_343_n N_A_397_297#_c_347_n
+ N_A_397_297#_c_344_n N_A_397_297#_c_341_n N_A_397_297#_c_342_n
+ N_A_397_297#_c_345_n PM_SKY130_FD_SC_HD__A2BB2OI_1%A_397_297#
x_PM_SKY130_FD_SC_HD__A2BB2OI_1%VGND N_VGND_M1008_s N_VGND_M1006_d
+ N_VGND_M1004_d N_VGND_c_369_n N_VGND_c_370_n VGND VGND N_VGND_c_372_n
+ N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_1%VGND
cc_1 VNB N_A1_N_c_58_n 0.0262988f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_2 VNB N_A1_N_c_59_n 0.0139994f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_3 VNB N_A1_N_c_60_n 0.0213312f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_4 VNB N_A2_N_c_85_n 0.0191856f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_5 VNB A2_N 0.00892467f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A2_N_c_87_n 0.0203614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_109_47#_c_119_n 0.0201685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_109_47#_c_120_n 0.0397473f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_9 VNB N_A_109_47#_c_121_n 0.0101847f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_10 VNB N_A_109_47#_c_122_n 0.00206149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B2_c_189_n 0.0164433f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_12 VNB B2 0.00190399f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_13 VNB B2 0.0028337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B2_c_192_n 0.021448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB B2 7.44967e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB B1 0.0120009f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_17 VNB N_B1_c_236_n 0.0288746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_c_237_n 0.0212964f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_19 VNB N_VPWR_c_264_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_308_n 0.00105946f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_VGND_c_369_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_370_n 0.0271113f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_23 VNB VGND 0.0103361f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_24 VNB N_VGND_c_372_n 0.0314288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_373_n 0.0117584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_374_n 0.0162605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_375_n 0.179928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_376_n 0.027016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A1_N_M1007_g 0.0217215f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_30 VPB N_A1_N_c_58_n 0.00490856f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_31 VPB N_A1_N_c_59_n 0.00680297f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_32 VPB N_A2_N_M1005_g 0.022574f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_33 VPB N_A2_N_c_87_n 0.00427188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_109_47#_M1003_g 0.0233145f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_35 VPB N_A_109_47#_c_120_n 0.0150371f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_36 VPB N_A_109_47#_c_121_n 6.57079e-19 $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_37 VPB N_A_109_47#_c_126_n 0.00921317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_109_47#_c_127_n 0.0119914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_109_47#_c_128_n 0.00274243f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_109_47#_c_122_n 0.00231195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B2_M1000_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_42 VPB N_B2_c_192_n 0.00459565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB B2 0.00228415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_B1_M1009_g 0.0230255f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB B1 0.00660854f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_46 VPB N_B1_c_236_n 0.00659506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_265_n 0.00231024f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_48 VPB VPWR 0.0103102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_267_n 0.0535368f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.325
cc_50 VPB N_VPWR_c_268_n 0.0151047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_264_n 0.0536626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_270_n 0.00353634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_271_n 0.0306083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_Y_c_308_n 0.00154032f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_55 VPB Y 0.00833523f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_397_297#_c_341_n 0.00899863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_397_297#_c_342_n 0.0195283f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_58 N_A1_N_M1007_g N_A2_N_M1005_g 0.048214f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A1_N_c_60_n N_A2_N_c_85_n 0.0235077f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A1_N_c_58_n A2_N 0.00162517f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A1_N_c_59_n A2_N 0.0189845f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A1_N_c_58_n N_A2_N_c_87_n 0.048214f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A1_N_c_59_n N_A2_N_c_87_n 0.00202629f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A1_N_M1007_g N_A_109_47#_c_126_n 0.00276518f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_65 N_A1_N_M1007_g N_A_109_47#_c_128_n 4.37046e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_66 N_A1_N_c_59_n N_A_109_47#_c_128_n 0.0075813f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A1_N_c_59_n N_VPWR_M1007_s 0.00800252f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A1_N_M1007_g N_VPWR_c_267_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A1_N_M1007_g N_VPWR_c_264_n 0.00783311f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A1_N_M1007_g N_VPWR_c_271_n 0.0173908f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A1_N_c_58_n N_VPWR_c_271_n 4.03133e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A1_N_c_59_n N_VPWR_c_271_n 0.0175924f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A1_N_c_60_n N_VGND_c_373_n 0.0046653f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A1_N_c_60_n N_VGND_c_374_n 5.71175e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_75 N_A1_N_c_60_n N_VGND_c_375_n 0.00799591f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A1_N_c_58_n N_VGND_c_376_n 7.77033e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A1_N_c_59_n N_VGND_c_376_n 0.0215627f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A1_N_c_60_n N_VGND_c_376_n 0.0114888f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_79 A2_N N_A_109_47#_c_120_n 0.00240279f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A2_N_c_87_n N_A_109_47#_c_120_n 0.0123653f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A2_N_c_85_n N_A_109_47#_c_135_n 0.0122302f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_82 A2_N N_A_109_47#_c_135_n 0.0297714f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A2_N_c_87_n N_A_109_47#_c_135_n 0.00122718f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_84 A2_N N_A_109_47#_c_138_n 0.00289746f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A2_N_c_87_n N_A_109_47#_c_138_n 2.52487e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A2_N_M1005_g N_A_109_47#_c_126_n 0.0141945f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_87 A2_N N_A_109_47#_c_127_n 0.00268974f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_88 N_A2_N_M1005_g N_A_109_47#_c_128_n 0.00380164f $X=0.83 $Y=1.985 $X2=0
+ $Y2=0
cc_89 A2_N N_A_109_47#_c_128_n 0.0280044f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A2_N_c_87_n N_A_109_47#_c_128_n 0.00321967f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A2_N_M1005_g N_A_109_47#_c_122_n 0.00286789f $X=0.83 $Y=1.985 $X2=0
+ $Y2=0
cc_92 N_A2_N_c_85_n N_A_109_47#_c_122_n 0.0042018f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_93 A2_N N_A_109_47#_c_122_n 0.0207162f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A2_N_c_87_n N_A_109_47#_c_122_n 6.15083e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A2_N_M1005_g N_VPWR_c_267_n 0.00541359f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A2_N_M1005_g N_VPWR_c_264_n 0.0108917f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A2_N_M1005_g N_VPWR_c_271_n 0.00303228f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A2_N_c_85_n N_VGND_c_373_n 0.00342263f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A2_N_c_85_n N_VGND_c_374_n 0.0084862f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A2_N_c_85_n N_VGND_c_375_n 0.00404827f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A2_N_c_85_n N_VGND_c_376_n 6.85747e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_109_47#_c_119_n N_B2_c_189_n 0.0224527f $X=1.91 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_109_47#_M1003_g N_B2_M1000_g 0.041627f $X=1.91 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_109_47#_c_121_n B2 0.00123007f $X=1.91 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_109_47#_c_121_n N_B2_c_192_n 0.0211836f $X=1.91 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_109_47#_M1003_g B2 0.00137155f $X=1.91 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_109_47#_M1003_g N_VPWR_c_267_n 0.00539883f $X=1.91 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_109_47#_c_126_n N_VPWR_c_267_n 0.0210382f $X=1.04 $Y=1.64 $X2=0 $Y2=0
cc_109 N_A_109_47#_M1005_d N_VPWR_c_264_n 0.00209319f $X=0.905 $Y=1.485 $X2=0
+ $Y2=0
cc_110 N_A_109_47#_M1003_g N_VPWR_c_264_n 0.00768248f $X=1.91 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_109_47#_c_126_n N_VPWR_c_264_n 0.0124268f $X=1.04 $Y=1.64 $X2=0 $Y2=0
cc_112 N_A_109_47#_c_126_n N_VPWR_c_271_n 0.0225012f $X=1.04 $Y=1.64 $X2=0 $Y2=0
cc_113 N_A_109_47#_c_127_n N_Y_M1003_s 0.00269266f $X=1.41 $Y=1.53 $X2=0 $Y2=0
cc_114 N_A_109_47#_c_119_n N_Y_c_308_n 0.00628353f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_109_47#_M1003_g N_Y_c_308_n 0.0163786f $X=1.91 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_109_47#_c_120_n N_Y_c_308_n 0.00945143f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_109_47#_c_121_n N_Y_c_308_n 0.00613012f $X=1.91 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_109_47#_c_126_n N_Y_c_308_n 0.00552823f $X=1.04 $Y=1.64 $X2=0 $Y2=0
cc_119 N_A_109_47#_c_127_n N_Y_c_308_n 0.0126507f $X=1.41 $Y=1.53 $X2=0 $Y2=0
cc_120 N_A_109_47#_c_122_n N_Y_c_308_n 0.0393066f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_109_47#_M1003_g Y 0.00543326f $X=1.91 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_109_47#_c_120_n Y 0.0070244f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_109_47#_c_126_n Y 0.0489281f $X=1.04 $Y=1.64 $X2=0 $Y2=0
cc_124 N_A_109_47#_c_127_n Y 0.014691f $X=1.41 $Y=1.53 $X2=0 $Y2=0
cc_125 N_A_109_47#_c_119_n Y 0.0215976f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_109_47#_c_135_n Y 0.0132607f $X=1.41 $Y=0.745 $X2=0 $Y2=0
cc_127 N_A_109_47#_M1003_g N_A_397_297#_c_343_n 0.00179375f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_128 N_A_109_47#_M1003_g N_A_397_297#_c_344_n 0.0011544f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_129 N_A_109_47#_M1003_g N_A_397_297#_c_345_n 0.00408878f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_130 N_A_109_47#_c_135_n N_VGND_M1006_d 0.0164521f $X=1.41 $Y=0.745 $X2=0
+ $Y2=0
cc_131 N_A_109_47#_c_122_n N_VGND_M1006_d 0.00128389f $X=1.495 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_109_47#_c_119_n N_VGND_c_372_n 0.00357668f $X=1.91 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_109_47#_c_180_p N_VGND_c_373_n 0.0112623f $X=0.68 $Y=0.66 $X2=0 $Y2=0
cc_134 N_A_109_47#_c_135_n N_VGND_c_373_n 0.00229693f $X=1.41 $Y=0.745 $X2=0
+ $Y2=0
cc_135 N_A_109_47#_c_119_n N_VGND_c_374_n 0.00577023f $X=1.91 $Y=0.995 $X2=0
+ $Y2=0
cc_136 N_A_109_47#_c_120_n N_VGND_c_374_n 0.00151821f $X=1.835 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_109_47#_c_135_n N_VGND_c_374_n 0.046106f $X=1.41 $Y=0.745 $X2=0 $Y2=0
cc_138 N_A_109_47#_M1008_d N_VGND_c_375_n 0.00413109f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_139 N_A_109_47#_c_119_n N_VGND_c_375_n 0.00666921f $X=1.91 $Y=0.995 $X2=0
+ $Y2=0
cc_140 N_A_109_47#_c_180_p N_VGND_c_375_n 0.0064418f $X=0.68 $Y=0.66 $X2=0 $Y2=0
cc_141 N_A_109_47#_c_135_n N_VGND_c_375_n 0.00694049f $X=1.41 $Y=0.745 $X2=0
+ $Y2=0
cc_142 N_B2_M1000_g N_B1_M1009_g 0.0445273f $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_143 B2 N_B1_M1009_g 0.00372559f $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_144 N_B2_M1000_g B1 2.26215e-19 $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_145 B2 B1 0.0488063f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_146 N_B2_c_192_n B1 2.68837e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_147 B2 N_B1_c_236_n 0.00372559f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_148 N_B2_c_192_n N_B1_c_236_n 0.0203393f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B2_c_189_n N_B1_c_237_n 0.0360034f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_150 B2 N_B1_c_237_n 0.00372559f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_151 B2 N_VPWR_M1000_d 0.00278837f $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_152 N_B2_M1000_g N_VPWR_c_265_n 0.00291989f $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B2_M1000_g N_VPWR_c_267_n 0.00539883f $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B2_M1000_g N_VPWR_c_264_n 0.00584993f $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B2_c_189_n N_Y_c_308_n 5.83845e-19 $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B2_M1000_g N_Y_c_308_n 0.00134166f $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_157 B2 N_Y_c_308_n 0.00430323f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_158 B2 N_Y_c_308_n 0.0258081f $X=2.44 $Y=1.105 $X2=0 $Y2=0
cc_159 N_B2_c_192_n N_Y_c_308_n 0.00108576f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B2_c_192_n Y 2.51049e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B2_M1000_g N_A_397_297#_c_343_n 0.00573833f $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_B2_M1000_g N_A_397_297#_c_347_n 0.00801436f $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_163 B2 N_A_397_297#_c_347_n 0.0209961f $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_164 N_B2_M1000_g N_A_397_297#_c_344_n 0.00207117f $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_B2_c_192_n N_A_397_297#_c_344_n 8.09007e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_166 B2 N_A_397_297#_c_344_n 0.00244706f $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_167 N_B2_M1000_g N_A_397_297#_c_345_n 0.00272627f $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_B2_c_189_n N_VGND_c_370_n 0.00178306f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_169 B2 N_VGND_c_370_n 0.0276664f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_170 N_B2_c_189_n N_VGND_c_372_n 0.00585385f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_171 B2 N_VGND_c_372_n 0.00525379f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_172 N_B2_c_189_n N_VGND_c_375_n 0.0108681f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_173 B2 N_VGND_c_375_n 0.00586314f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_174 B2 A_481_47# 0.0091941f $X=2.44 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_175 N_B1_M1009_g N_VPWR_c_265_n 0.00957278f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B1_M1009_g N_VPWR_c_268_n 0.0046653f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B1_M1009_g N_VPWR_c_264_n 0.00515525f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_178 B1 N_A_397_297#_M1009_d 0.00772628f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_179 N_B1_M1009_g N_A_397_297#_c_343_n 5.9207e-19 $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1009_g N_A_397_297#_c_347_n 0.0125389f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_181 B1 N_A_397_297#_c_347_n 0.00335055f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_182 B1 N_A_397_297#_c_341_n 0.0167568f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_183 N_B1_c_236_n N_A_397_297#_c_341_n 5.13239e-19 $X=2.865 $Y=1.16 $X2=0
+ $Y2=0
cc_184 B1 N_VGND_c_370_n 0.0213054f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_185 N_B1_c_236_n N_VGND_c_370_n 0.00390305f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_186 N_B1_c_237_n N_VGND_c_370_n 0.0142495f $X=2.837 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_237_n N_VGND_c_372_n 0.0046653f $X=2.837 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_237_n N_VGND_c_375_n 0.00799591f $X=2.837 $Y=0.995 $X2=0 $Y2=0
cc_189 N_VPWR_c_264_n A_109_297# 0.00897657f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_190 N_VPWR_c_264_n N_Y_M1003_s 0.00303476f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_267_n Y 0.0254566f $X=2.455 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_264_n Y 0.0198308f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_264_n N_A_397_297#_M1003_d 0.00215227f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_194 N_VPWR_c_264_n N_A_397_297#_M1009_d 0.00235804f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_195 N_VPWR_M1000_d N_A_397_297#_c_347_n 0.00353814f $X=2.405 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_265_n N_A_397_297#_c_347_n 0.0137794f $X=2.54 $Y=2.36 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_264_n N_A_397_297#_c_347_n 0.0115157f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_268_n N_A_397_297#_c_342_n 0.0176426f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_264_n N_A_397_297#_c_342_n 0.00974347f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_267_n N_A_397_297#_c_345_n 0.0178243f $X=2.455 $Y=2.72 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_264_n N_A_397_297#_c_345_n 0.0119575f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_202 Y N_A_397_297#_c_344_n 0.0145809f $X=1.52 $Y=2.125 $X2=0 $Y2=0
cc_203 N_Y_c_308_n N_VGND_M1006_d 6.2131e-19 $X=1.86 $Y=1.785 $X2=0 $Y2=0
cc_204 Y N_VGND_M1006_d 0.0117713f $X=1.98 $Y=0.425 $X2=0 $Y2=0
cc_205 Y N_VGND_c_372_n 0.0253507f $X=1.98 $Y=0.425 $X2=0 $Y2=0
cc_206 Y N_VGND_c_374_n 0.0202845f $X=1.98 $Y=0.425 $X2=0 $Y2=0
cc_207 N_Y_M1002_d N_VGND_c_375_n 0.00393857f $X=1.985 $Y=0.235 $X2=0 $Y2=0
cc_208 Y N_VGND_c_375_n 0.015741f $X=1.98 $Y=0.425 $X2=0 $Y2=0
cc_209 N_VGND_c_375_n A_481_47# 0.00587338f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o311a_1.spice
* Created: Thu Aug 27 14:38:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o311a_1.pex.spice"
.subckt sky130_fd_sc_hd__o311a_1  VNB VPB A1 A2 A3 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_81_21#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.203125 AS=0.169 PD=1.275 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1003 N_A_266_47#_M1003_d N_A1_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.203125 PD=1.01 PS=1.275 NRD=7.38 NRS=1.836 M=1 R=4.33333
+ SA=75001 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_266_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1365 AS=0.117 PD=1.07 PS=1.01 NRD=12.912 NRS=7.38 M=1 R=4.33333
+ SA=75001.5 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_266_47#_M1008_d N_A3_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.1365 PD=1.015 PS=1.07 NRD=8.304 NRS=12.912 M=1 R=4.33333
+ SA=75002 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 A_585_47# N_B1_M1009_g N_A_266_47#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.118625 PD=0.86 PS=1.015 NRD=9.228 NRS=7.38 M=1 R=4.33333
+ SA=75002.6 SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1010 N_A_81_21#_M1010_d N_C1_M1010_g A_585_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.06825 PD=1.82 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_81_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3125 AS=0.26 PD=1.625 PS=2.52 NRD=25.5903 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1002 A_266_297# N_A1_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.18
+ AS=0.3125 PD=1.36 PS=1.625 NRD=24.6053 NRS=42.3353 M=1 R=6.66667 SA=75001
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1004 A_368_297# N_A2_M1004_g A_266_297# VPB PHIGHVT L=0.15 W=1 AD=0.21 AS=0.18
+ PD=1.42 PS=1.36 NRD=30.5153 NRS=24.6053 M=1 R=6.66667 SA=75001.5 SB=75001.6
+ A=0.15 P=2.3 MULT=1
MM1011 N_A_81_21#_M1011_d N_A3_M1011_g A_368_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.21 PD=1.275 PS=1.42 NRD=0 NRS=30.5153 M=1 R=6.66667 SA=75002
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_81_21#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.1375 PD=1.3 PS=1.275 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75002.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_81_21#_M1000_d N_C1_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.15 PD=2.52 PS=1.3 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75002.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__o311a_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o21bai_2.pxi.spice
* Created: Thu Aug 27 14:36:32 2020
* 
x_PM_SKY130_FD_SC_HD__O21BAI_2%B1_N N_B1_N_M1005_g N_B1_N_M1006_g B1_N
+ N_B1_N_c_74_n N_B1_N_c_75_n N_B1_N_c_76_n PM_SKY130_FD_SC_HD__O21BAI_2%B1_N
x_PM_SKY130_FD_SC_HD__O21BAI_2%A_28_297# N_A_28_297#_M1005_d N_A_28_297#_M1006_s
+ N_A_28_297#_M1008_g N_A_28_297#_M1011_g N_A_28_297#_c_104_n
+ N_A_28_297#_M1007_g N_A_28_297#_c_105_n N_A_28_297#_M1009_g
+ N_A_28_297#_c_118_n N_A_28_297#_c_106_n N_A_28_297#_c_107_n
+ N_A_28_297#_c_108_n N_A_28_297#_c_115_n N_A_28_297#_c_109_n
+ N_A_28_297#_c_110_n N_A_28_297#_c_111_n PM_SKY130_FD_SC_HD__O21BAI_2%A_28_297#
x_PM_SKY130_FD_SC_HD__O21BAI_2%A2 N_A2_c_178_n N_A2_M1012_g N_A2_M1003_g
+ N_A2_c_179_n N_A2_M1013_g N_A2_M1004_g A2 N_A2_c_181_n
+ PM_SKY130_FD_SC_HD__O21BAI_2%A2
x_PM_SKY130_FD_SC_HD__O21BAI_2%A1 N_A1_c_230_n N_A1_M1001_g N_A1_M1000_g
+ N_A1_c_231_n N_A1_M1002_g N_A1_M1010_g A1 N_A1_c_233_n
+ PM_SKY130_FD_SC_HD__O21BAI_2%A1
x_PM_SKY130_FD_SC_HD__O21BAI_2%VPWR N_VPWR_M1006_d N_VPWR_M1011_d N_VPWR_M1000_d
+ N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n VPWR N_VPWR_c_272_n
+ N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_268_n N_VPWR_c_277_n
+ N_VPWR_c_278_n N_VPWR_c_279_n PM_SKY130_FD_SC_HD__O21BAI_2%VPWR
x_PM_SKY130_FD_SC_HD__O21BAI_2%Y N_Y_M1007_d N_Y_M1008_s N_Y_M1003_s N_Y_c_357_n
+ N_Y_c_331_n N_Y_c_364_p N_Y_c_332_n N_Y_c_329_n Y
+ PM_SKY130_FD_SC_HD__O21BAI_2%Y
x_PM_SKY130_FD_SC_HD__O21BAI_2%A_397_297# N_A_397_297#_M1003_d
+ N_A_397_297#_M1004_d N_A_397_297#_M1010_s N_A_397_297#_c_372_n
+ N_A_397_297#_c_378_n N_A_397_297#_c_373_n N_A_397_297#_c_374_n
+ N_A_397_297#_c_397_n N_A_397_297#_c_375_n N_A_397_297#_c_376_n
+ N_A_397_297#_c_377_n PM_SKY130_FD_SC_HD__O21BAI_2%A_397_297#
x_PM_SKY130_FD_SC_HD__O21BAI_2%VGND N_VGND_M1005_s N_VGND_M1012_s N_VGND_M1001_s
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n
+ N_VGND_c_415_n VGND N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n
+ N_VGND_c_419_n PM_SKY130_FD_SC_HD__O21BAI_2%VGND
x_PM_SKY130_FD_SC_HD__O21BAI_2%A_229_47# N_A_229_47#_M1007_s N_A_229_47#_M1009_s
+ N_A_229_47#_M1013_d N_A_229_47#_M1002_d N_A_229_47#_c_469_n
+ N_A_229_47#_c_470_n N_A_229_47#_c_483_n N_A_229_47#_c_487_n
+ N_A_229_47#_c_471_n N_A_229_47#_c_472_n N_A_229_47#_c_495_n
+ N_A_229_47#_c_473_n N_A_229_47#_c_474_n N_A_229_47#_c_475_n
+ PM_SKY130_FD_SC_HD__O21BAI_2%A_229_47#
cc_1 VNB N_B1_N_c_74_n 0.0347541f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_2 VNB N_B1_N_c_75_n 0.0152894f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_3 VNB N_B1_N_c_76_n 0.0218216f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.995
cc_4 VNB N_A_28_297#_c_104_n 0.0193714f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_5 VNB N_A_28_297#_c_105_n 0.0161165f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_6 VNB N_A_28_297#_c_106_n 0.0043177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_28_297#_c_107_n 9.05065e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_28_297#_c_108_n 9.61753e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_28_297#_c_109_n 0.00679699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_28_297#_c_110_n 0.00101775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_28_297#_c_111_n 0.0678428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_178_n 0.0160068f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_13 VNB N_A2_c_179_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_14 VNB A2 0.0115907f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_15 VNB N_A2_c_181_n 0.0302945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_230_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_17 VNB N_A1_c_231_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB A1 0.0209839f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_19 VNB N_A1_c_233_n 0.0372217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_268_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_329_n 5.95106e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB Y 8.47613e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_410_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=1.16
cc_24 VNB N_VGND_c_411_n 0.0184161f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_25 VNB N_VGND_c_412_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_413_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_414_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_415_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_416_n 0.0526102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_417_n 0.0200444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_418_n 0.243353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_419_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_229_47#_c_469_n 0.00628458f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.995
cc_34 VNB N_A_229_47#_c_470_n 0.00632785f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_35 VNB N_A_229_47#_c_471_n 0.00218403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_229_47#_c_472_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_229_47#_c_473_n 0.0130716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_229_47#_c_474_n 0.0183327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_229_47#_c_475_n 0.00252847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_B1_N_M1006_g 0.0292612f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.695
cc_41 VPB N_B1_N_c_74_n 0.00733828f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_42 VPB N_B1_N_c_75_n 0.00408805f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_43 VPB N_A_28_297#_M1008_g 0.0208772f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_28_297#_M1011_g 0.0219282f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.995
cc_45 VPB N_A_28_297#_c_107_n 0.0034884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_28_297#_c_115_n 0.00361181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_28_297#_c_111_n 0.0192246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A2_M1003_g 0.0226707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.695
cc_49 VPB N_A2_M1004_g 0.0188152f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.995
cc_50 VPB N_A2_c_181_n 0.00410911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A1_M1000_g 0.0182767f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.695
cc_52 VPB N_A1_M1010_g 0.0250431f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.995
cc_53 VPB N_A1_c_233_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_269_n 0.0214531f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_55 VPB N_VPWR_c_270_n 0.0103161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_271_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_272_n 0.0207592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_273_n 0.0149703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_274_n 0.0357219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_275_n 0.0177805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_268_n 0.0686865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_277_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_278_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_279_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_Y_c_331_n 0.0137573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_Y_c_332_n 0.00167421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB Y 0.00656124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_397_297#_c_372_n 0.004784f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_69 VPB N_A_397_297#_c_373_n 0.00178643f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_70 VPB N_A_397_297#_c_374_n 0.00185317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_397_297#_c_375_n 0.00330345f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_72 VPB N_A_397_297#_c_376_n 0.0116415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_397_297#_c_377_n 0.0307403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_B1_N_M1006_g N_A_28_297#_M1008_g 0.0141662f $X=0.475 $Y=1.695 $X2=0
+ $Y2=0
cc_75 N_B1_N_M1006_g N_A_28_297#_c_118_n 0.0137464f $X=0.475 $Y=1.695 $X2=0
+ $Y2=0
cc_76 N_B1_N_c_75_n N_A_28_297#_c_118_n 0.0108027f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B1_N_c_75_n N_A_28_297#_c_106_n 0.00606206f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_N_c_76_n N_A_28_297#_c_106_n 0.00604363f $X=0.362 $Y=0.995 $X2=0
+ $Y2=0
cc_79 N_B1_N_c_74_n N_A_28_297#_c_107_n 0.00430707f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B1_N_c_75_n N_A_28_297#_c_107_n 0.00606206f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B1_N_M1006_g N_A_28_297#_c_115_n 2.26469e-19 $X=0.475 $Y=1.695 $X2=0
+ $Y2=0
cc_82 N_B1_N_c_74_n N_A_28_297#_c_115_n 0.00383828f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B1_N_c_75_n N_A_28_297#_c_115_n 0.0131028f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B1_N_c_76_n N_A_28_297#_c_109_n 4.45628e-19 $X=0.362 $Y=0.995 $X2=0
+ $Y2=0
cc_85 N_B1_N_c_74_n N_A_28_297#_c_110_n 0.00139007f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B1_N_c_75_n N_A_28_297#_c_110_n 0.0146232f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_N_c_74_n N_A_28_297#_c_111_n 0.0141662f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B1_N_c_75_n N_A_28_297#_c_111_n 2.09592e-19 $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B1_N_M1006_g N_VPWR_c_269_n 0.00366987f $X=0.475 $Y=1.695 $X2=0 $Y2=0
cc_90 N_B1_N_M1006_g N_VPWR_c_272_n 0.00327927f $X=0.475 $Y=1.695 $X2=0 $Y2=0
cc_91 N_B1_N_M1006_g N_VPWR_c_268_n 0.00417489f $X=0.475 $Y=1.695 $X2=0 $Y2=0
cc_92 N_B1_N_c_74_n N_VGND_c_411_n 0.00389539f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B1_N_c_75_n N_VGND_c_411_n 0.0136043f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_N_c_76_n N_VGND_c_411_n 0.00476913f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B1_N_c_76_n N_VGND_c_416_n 0.00510437f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B1_N_c_76_n N_VGND_c_418_n 0.00512902f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B1_N_c_76_n N_A_229_47#_c_469_n 0.00320334f $X=0.362 $Y=0.995 $X2=0
+ $Y2=0
cc_98 N_A_28_297#_c_105_n N_A2_c_178_n 0.0146384f $X=1.9 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_28_297#_c_111_n A2 0.00647538f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_28_297#_c_111_n N_A2_c_181_n 0.0146384f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_28_297#_c_118_n N_VPWR_M1006_d 0.00528106f $X=0.695 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A_28_297#_M1008_g N_VPWR_c_269_n 0.0122482f $X=0.96 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_28_297#_M1011_g N_VPWR_c_269_n 6.39542e-19 $X=1.38 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_28_297#_c_118_n N_VPWR_c_269_n 0.0162855f $X=0.695 $Y=1.58 $X2=0
+ $Y2=0
cc_105 N_A_28_297#_c_108_n N_VPWR_c_269_n 0.00101503f $X=1.17 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_A_28_297#_c_115_n N_VPWR_c_269_n 5.6836e-19 $X=0.265 $Y=1.58 $X2=0
+ $Y2=0
cc_107 N_A_28_297#_M1011_g N_VPWR_c_270_n 0.00329978f $X=1.38 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_28_297#_c_111_n N_VPWR_c_270_n 8.56004e-19 $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_28_297#_M1008_g N_VPWR_c_273_n 0.0046653f $X=0.96 $Y=1.985 $X2=0
+ $Y2=0
cc_110 N_A_28_297#_M1011_g N_VPWR_c_273_n 0.00585385f $X=1.38 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_28_297#_M1008_g N_VPWR_c_268_n 0.00789179f $X=0.96 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_28_297#_M1011_g N_VPWR_c_268_n 0.0117754f $X=1.38 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_28_297#_c_115_n N_VPWR_c_268_n 0.00647432f $X=0.265 $Y=1.58 $X2=0
+ $Y2=0
cc_114 N_A_28_297#_c_111_n N_Y_c_331_n 0.00729082f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_28_297#_M1008_g N_Y_c_332_n 3.5749e-19 $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_28_297#_c_107_n N_Y_c_332_n 0.00274402f $X=0.78 $Y=1.495 $X2=0 $Y2=0
cc_117 N_A_28_297#_c_108_n N_Y_c_332_n 0.0121469f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_28_297#_c_111_n N_Y_c_332_n 0.00227631f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_28_297#_c_104_n N_Y_c_329_n 0.00347361f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_28_297#_c_105_n N_Y_c_329_n 0.00396956f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_28_297#_M1011_g Y 0.0218847f $X=1.38 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_28_297#_c_104_n Y 0.00276455f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_28_297#_c_105_n Y 0.00231234f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_28_297#_c_106_n Y 0.00439456f $X=0.78 $Y=1.075 $X2=0 $Y2=0
cc_125 N_A_28_297#_c_107_n Y 0.00558599f $X=0.78 $Y=1.495 $X2=0 $Y2=0
cc_126 N_A_28_297#_c_108_n Y 0.0168964f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_28_297#_c_111_n Y 0.0294218f $X=1.9 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_28_297#_c_109_n N_VGND_c_411_n 0.00107392f $X=0.78 $Y=0.635 $X2=0
+ $Y2=0
cc_129 N_A_28_297#_c_104_n N_VGND_c_416_n 0.00357877f $X=1.48 $Y=0.995 $X2=0
+ $Y2=0
cc_130 N_A_28_297#_c_105_n N_VGND_c_416_n 0.00357877f $X=1.9 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_28_297#_c_109_n N_VGND_c_416_n 0.00818069f $X=0.78 $Y=0.635 $X2=0
+ $Y2=0
cc_132 N_A_28_297#_c_104_n N_VGND_c_418_n 0.00655123f $X=1.48 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_28_297#_c_105_n N_VGND_c_418_n 0.00525237f $X=1.9 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_28_297#_c_109_n N_VGND_c_418_n 0.00891815f $X=0.78 $Y=0.635 $X2=0
+ $Y2=0
cc_135 N_A_28_297#_c_109_n N_A_229_47#_c_469_n 0.00218471f $X=0.78 $Y=0.635
+ $X2=0 $Y2=0
cc_136 N_A_28_297#_c_104_n N_A_229_47#_c_470_n 4.45069e-19 $X=1.48 $Y=0.995
+ $X2=0 $Y2=0
cc_137 N_A_28_297#_c_106_n N_A_229_47#_c_470_n 0.00539924f $X=0.78 $Y=1.075
+ $X2=0 $Y2=0
cc_138 N_A_28_297#_c_108_n N_A_229_47#_c_470_n 0.020813f $X=1.17 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_28_297#_c_109_n N_A_229_47#_c_470_n 0.0244038f $X=0.78 $Y=0.635 $X2=0
+ $Y2=0
cc_140 N_A_28_297#_c_111_n N_A_229_47#_c_470_n 0.00803853f $X=1.9 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_28_297#_c_104_n N_A_229_47#_c_483_n 0.0127333f $X=1.48 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_A_28_297#_c_105_n N_A_229_47#_c_483_n 0.0123199f $X=1.9 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_28_297#_c_111_n N_A_229_47#_c_483_n 3.07604e-19 $X=1.9 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A2_c_179_n N_A1_c_230_n 0.0150406f $X=2.74 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_145 N_A2_M1004_g N_A1_M1000_g 0.0150406f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_146 A2 A1 0.01677f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_147 A2 N_A1_c_233_n 0.00529309f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A2_c_181_n N_A1_c_233_n 0.0150406f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A2_M1003_g N_VPWR_c_270_n 0.00216742f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A2_M1004_g N_VPWR_c_271_n 0.00110007f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_M1003_g N_VPWR_c_274_n 0.00357877f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A2_M1004_g N_VPWR_c_274_n 0.00357877f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A2_M1003_g N_VPWR_c_268_n 0.00655123f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A2_M1004_g N_VPWR_c_268_n 0.00525237f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A2_M1003_g N_Y_c_331_n 0.0154024f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A2_M1004_g N_Y_c_331_n 6.14663e-19 $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_157 A2 N_Y_c_331_n 0.0535594f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A2_c_181_n N_Y_c_331_n 0.00222181f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_M1003_g Y 0.00313515f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_160 A2 Y 0.0155988f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A2_c_181_n Y 7.70674e-19 $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A2_M1003_g N_A_397_297#_c_378_n 0.0121306f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_M1004_g N_A_397_297#_c_378_n 0.0121306f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_M1004_g N_A_397_297#_c_374_n 2.63361e-19 $X=2.74 $Y=1.985 $X2=0
+ $Y2=0
cc_165 A2 N_A_397_297#_c_374_n 0.0140069f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_166 A2 N_A_397_297#_c_375_n 0.00396848f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A2_c_178_n N_VGND_c_412_n 0.00268723f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_179_n N_VGND_c_412_n 0.00146448f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A2_c_179_n N_VGND_c_414_n 0.00423334f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A2_c_178_n N_VGND_c_416_n 0.00421816f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_c_178_n N_VGND_c_418_n 0.00575258f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_179_n N_VGND_c_418_n 0.0057435f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_173 A2 N_A_229_47#_c_483_n 0.00138616f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A2_c_178_n N_A_229_47#_c_487_n 0.00255288f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A2_c_178_n N_A_229_47#_c_471_n 0.00485712f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A2_c_179_n N_A_229_47#_c_471_n 4.58193e-19 $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_177 A2 N_A_229_47#_c_471_n 0.0211267f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A2_c_178_n N_A_229_47#_c_472_n 0.00869873f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A2_c_179_n N_A_229_47#_c_472_n 0.00865195f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_180 A2 N_A_229_47#_c_472_n 0.0363039f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A2_c_181_n N_A_229_47#_c_472_n 0.00222006f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A2_c_178_n N_A_229_47#_c_495_n 5.22228e-19 $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_179_n N_A_229_47#_c_495_n 0.00630972f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_179_n N_A_229_47#_c_475_n 0.00112659f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_185 A2 N_A_229_47#_c_475_n 0.025711f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A1_M1000_g N_VPWR_c_271_n 0.0122146f $X=3.16 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A1_M1010_g N_VPWR_c_271_n 0.0129691f $X=3.58 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A1_M1000_g N_VPWR_c_274_n 0.0046653f $X=3.16 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A1_M1010_g N_VPWR_c_275_n 0.0046653f $X=3.58 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A1_M1000_g N_VPWR_c_268_n 0.007919f $X=3.16 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A1_M1010_g N_VPWR_c_268_n 0.00892182f $X=3.58 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A1_M1000_g N_A_397_297#_c_375_n 0.0152539f $X=3.16 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A1_M1010_g N_A_397_297#_c_375_n 0.013814f $X=3.58 $Y=1.985 $X2=0 $Y2=0
cc_194 A1 N_A_397_297#_c_375_n 0.0310409f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_195 N_A1_c_233_n N_A_397_297#_c_375_n 0.00213668f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_196 A1 N_A_397_297#_c_376_n 0.0226583f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A1_c_230_n N_VGND_c_413_n 0.00146448f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_231_n N_VGND_c_413_n 0.00268723f $X=3.58 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_230_n N_VGND_c_414_n 0.00423334f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_231_n N_VGND_c_417_n 0.00423737f $X=3.58 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_230_n N_VGND_c_418_n 0.0057435f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A1_c_231_n N_VGND_c_418_n 0.00674672f $X=3.58 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_230_n N_A_229_47#_c_495_n 0.00630972f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_231_n N_A_229_47#_c_495_n 5.22228e-19 $X=3.58 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A1_c_230_n N_A_229_47#_c_473_n 0.0101811f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A1_c_231_n N_A_229_47#_c_473_n 0.0099997f $X=3.58 $Y=0.995 $X2=0 $Y2=0
cc_207 A1 N_A_229_47#_c_473_n 0.0561868f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A1_c_233_n N_A_229_47#_c_473_n 0.00222006f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A1_c_230_n N_A_229_47#_c_474_n 5.18879e-19 $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_231_n N_A_229_47#_c_474_n 0.00621819f $X=3.58 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A1_c_230_n N_A_229_47#_c_475_n 0.0014009f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_212 N_VPWR_c_268_n N_Y_M1008_s 0.00562358f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_268_n N_Y_M1003_s 0.00216833f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_273_n N_Y_c_357_n 0.0113958f $X=1.47 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_c_268_n N_Y_c_357_n 0.00646998f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_M1011_d Y 0.00264121f $X=1.455 $Y=1.485 $X2=0 $Y2=0
cc_217 N_VPWR_c_270_n Y 0.0177477f $X=1.59 $Y=1.96 $X2=0 $Y2=0
cc_218 N_VPWR_c_268_n N_A_397_297#_M1003_d 0.0020932f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_219 N_VPWR_c_268_n N_A_397_297#_M1004_d 0.00385313f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_268_n N_A_397_297#_M1010_s 0.00399293f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_270_n N_A_397_297#_c_372_n 0.0320877f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_274_n N_A_397_297#_c_378_n 0.0344282f $X=3.205 $Y=2.72 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_268_n N_A_397_297#_c_378_n 0.0219525f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_270_n N_A_397_297#_c_373_n 0.0117482f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_274_n N_A_397_297#_c_373_n 0.0180757f $X=3.205 $Y=2.72 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_268_n N_A_397_297#_c_373_n 0.0107791f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_274_n N_A_397_297#_c_397_n 0.0114668f $X=3.205 $Y=2.72 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_268_n N_A_397_297#_c_397_n 0.006547f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_M1000_d N_A_397_297#_c_375_n 0.00166915f $X=3.235 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_271_n N_A_397_297#_c_375_n 0.0172742f $X=3.37 $Y=2 $X2=0 $Y2=0
cc_231 N_VPWR_c_275_n N_A_397_297#_c_377_n 0.019049f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_268_n N_A_397_297#_c_377_n 0.0105137f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_Y_c_331_n N_A_397_297#_M1003_d 0.00278154f $X=2.405 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_234 N_Y_c_331_n N_A_397_297#_c_372_n 0.0181545f $X=2.405 $Y=1.53 $X2=0 $Y2=0
cc_235 N_Y_M1003_s N_A_397_297#_c_378_n 0.00312348f $X=2.395 $Y=1.485 $X2=0
+ $Y2=0
cc_236 N_Y_c_364_p N_A_397_297#_c_378_n 0.0118865f $X=2.53 $Y=1.62 $X2=0 $Y2=0
cc_237 N_Y_c_331_n N_A_397_297#_c_374_n 0.00229817f $X=2.405 $Y=1.53 $X2=0 $Y2=0
cc_238 N_Y_M1007_d N_VGND_c_418_n 0.00216833f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_329_n N_A_229_47#_c_470_n 0.0105269f $X=1.69 $Y=0.73 $X2=0 $Y2=0
cc_240 Y N_A_229_47#_c_470_n 6.39493e-19 $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_241 N_Y_M1007_d N_A_229_47#_c_483_n 0.00304656f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_242 N_Y_c_329_n N_A_229_47#_c_483_n 0.016271f $X=1.69 $Y=0.73 $X2=0 $Y2=0
cc_243 N_Y_c_329_n N_A_229_47#_c_471_n 0.00767188f $X=1.69 $Y=0.73 $X2=0 $Y2=0
cc_244 N_A_397_297#_c_375_n N_A_229_47#_c_473_n 0.00403925f $X=3.705 $Y=1.56
+ $X2=0 $Y2=0
cc_245 N_A_397_297#_c_375_n N_A_229_47#_c_475_n 7.61366e-19 $X=3.705 $Y=1.56
+ $X2=0 $Y2=0
cc_246 N_VGND_c_418_n N_A_229_47#_M1007_s 0.00209324f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_247 N_VGND_c_418_n N_A_229_47#_M1009_s 0.00215206f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_418_n N_A_229_47#_M1013_d 0.00215201f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_418_n N_A_229_47#_M1002_d 0.00226063f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_c_416_n N_A_229_47#_c_469_n 0.0194781f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_251 N_VGND_c_418_n N_A_229_47#_c_469_n 0.0107706f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_416_n N_A_229_47#_c_483_n 0.0363282f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_418_n N_A_229_47#_c_483_n 0.023578f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_416_n N_A_229_47#_c_487_n 0.0152108f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_418_n N_A_229_47#_c_487_n 0.00940698f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_M1012_s N_A_229_47#_c_472_n 0.00162089f $X=2.395 $Y=0.235 $X2=0
+ $Y2=0
cc_257 N_VGND_c_412_n N_A_229_47#_c_472_n 0.0122559f $X=2.53 $Y=0.39 $X2=0 $Y2=0
cc_258 N_VGND_c_414_n N_A_229_47#_c_472_n 0.00198695f $X=3.285 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_c_416_n N_A_229_47#_c_472_n 0.00198695f $X=2.445 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_418_n N_A_229_47#_c_472_n 0.00835832f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_414_n N_A_229_47#_c_495_n 0.0188551f $X=3.285 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_418_n N_A_229_47#_c_495_n 0.0122069f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_M1001_s N_A_229_47#_c_473_n 0.00162089f $X=3.235 $Y=0.235 $X2=0
+ $Y2=0
cc_264 N_VGND_c_413_n N_A_229_47#_c_473_n 0.0122559f $X=3.37 $Y=0.39 $X2=0 $Y2=0
cc_265 N_VGND_c_414_n N_A_229_47#_c_473_n 0.00198695f $X=3.285 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_417_n N_A_229_47#_c_473_n 0.00198695f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_267 N_VGND_c_418_n N_A_229_47#_c_473_n 0.00835832f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_417_n N_A_229_47#_c_474_n 0.0213509f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_418_n N_A_229_47#_c_474_n 0.0133027f $X=3.91 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkbuf_1.pxi.spice
* Created: Thu Aug 27 14:10:48 2020
* 
x_PM_SKY130_FD_SC_HD__CLKBUF_1%A_75_212# N_A_75_212#_M1001_d N_A_75_212#_M1002_d
+ N_A_75_212#_M1003_g N_A_75_212#_M1000_g N_A_75_212#_c_41_n N_A_75_212#_c_36_n
+ N_A_75_212#_c_63_p N_A_75_212#_c_42_n N_A_75_212#_c_65_p N_A_75_212#_c_97_p
+ N_A_75_212#_c_83_p N_A_75_212#_c_37_n N_A_75_212#_c_38_n N_A_75_212#_c_39_n
+ PM_SKY130_FD_SC_HD__CLKBUF_1%A_75_212#
x_PM_SKY130_FD_SC_HD__CLKBUF_1%A N_A_c_101_n N_A_M1001_g N_A_M1002_g N_A_c_102_n
+ N_A_c_105_n N_A_c_106_n A PM_SKY130_FD_SC_HD__CLKBUF_1%A
x_PM_SKY130_FD_SC_HD__CLKBUF_1%X N_X_M1003_s N_X_M1000_s N_X_c_131_n N_X_c_134_n
+ N_X_c_132_n X X X PM_SKY130_FD_SC_HD__CLKBUF_1%X
x_PM_SKY130_FD_SC_HD__CLKBUF_1%VPWR N_VPWR_M1000_d N_VPWR_c_156_n VPWR
+ N_VPWR_c_158_n N_VPWR_c_159_n N_VPWR_c_160_n PM_SKY130_FD_SC_HD__CLKBUF_1%VPWR
x_PM_SKY130_FD_SC_HD__CLKBUF_1%VGND N_VGND_M1003_d N_VGND_c_179_n VGND
+ N_VGND_c_181_n N_VGND_c_182_n N_VGND_c_183_n PM_SKY130_FD_SC_HD__CLKBUF_1%VGND
cc_1 VNB N_A_75_212#_M1003_g 0.0289893f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_2 VNB N_A_75_212#_c_36_n 0.00771329f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=0.72
cc_3 VNB N_A_75_212#_c_37_n 0.00163395f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.225
cc_4 VNB N_A_75_212#_c_38_n 0.0191693f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.225
cc_5 VNB N_A_75_212#_c_39_n 0.0021693f $X=-0.19 $Y=-0.24 $X2=0.567 $Y2=1.06
cc_6 VNB N_A_c_101_n 0.0179813f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=0.235
cc_7 VNB N_A_c_102_n 0.048966f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.06
cc_8 VNB A 0.0163436f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.39
cc_9 VNB N_X_c_131_n 0.00847523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_X_c_132_n 0.0254822f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.09
cc_11 VNB X 0.0145716f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.09
cc_12 VNB VPWR 0.0609879f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_13 VNB N_VGND_c_179_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB VGND 0.10585f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_15 VNB N_VGND_c_181_n 0.0153759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_182_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.39
cc_17 VNB N_VGND_c_183_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.62
cc_18 VPB N_A_75_212#_M1000_g 0.0288945f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.09
cc_19 VPB N_A_75_212#_c_41_n 0.00135348f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.535
cc_20 VPB N_A_75_212#_c_42_n 0.0120187f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.62
cc_21 VPB N_A_75_212#_c_37_n 6.91362e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.225
cc_22 VPB N_A_75_212#_c_38_n 0.00918419f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.225
cc_23 VPB N_A_c_102_n 0.00829456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.06
cc_24 VPB N_A_c_105_n 0.0136585f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.495
cc_25 VPB N_A_c_106_n 0.0273733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB A 0.00627368f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.39
cc_27 VPB N_X_c_134_n 0.0110375f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.39
cc_28 VPB N_X_c_132_n 0.0119115f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.09
cc_29 VPB X 0.0297138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_156_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB VPWR 0.0448622f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.495
cc_32 VPB N_VPWR_c_158_n 0.0152818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_159_n 0.0162226f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.39
cc_34 VPB N_VPWR_c_160_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.62
cc_35 N_A_75_212#_M1003_g N_A_c_101_n 0.0209393f $X=0.47 $Y=0.495 $X2=-0.19
+ $Y2=-0.24
cc_36 N_A_75_212#_c_36_n N_A_c_101_n 0.015302f $X=1.035 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_37 N_A_75_212#_c_39_n N_A_c_101_n 0.00318324f $X=0.567 $Y=1.06 $X2=-0.19
+ $Y2=-0.24
cc_38 N_A_75_212#_M1003_g N_A_c_102_n 0.003841f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_39 N_A_75_212#_c_36_n N_A_c_102_n 0.00234783f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_40 N_A_75_212#_c_42_n N_A_c_102_n 0.00154723f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_41 N_A_75_212#_c_38_n N_A_c_102_n 0.0193066f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_42 N_A_75_212#_c_39_n N_A_c_102_n 0.00324151f $X=0.567 $Y=1.06 $X2=0 $Y2=0
cc_43 N_A_75_212#_M1000_g N_A_c_105_n 0.00368068f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_44 N_A_75_212#_c_37_n N_A_c_105_n 0.00324151f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_45 N_A_75_212#_M1000_g N_A_c_106_n 0.0166651f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_46 N_A_75_212#_c_41_n N_A_c_106_n 7.5643e-19 $X=0.625 $Y=1.535 $X2=0 $Y2=0
cc_47 N_A_75_212#_c_42_n N_A_c_106_n 0.0192508f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_48 N_A_75_212#_c_36_n A 0.0207534f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_49 N_A_75_212#_c_42_n A 0.0208772f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_50 N_A_75_212#_c_38_n A 2.94551e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_51 N_A_75_212#_c_39_n A 0.0224427f $X=0.567 $Y=1.06 $X2=0 $Y2=0
cc_52 N_A_75_212#_M1003_g N_X_c_131_n 0.00222896f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_53 N_A_75_212#_c_63_p N_X_c_131_n 0.00484499f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_54 N_A_75_212#_M1000_g N_X_c_134_n 0.00347811f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_55 N_A_75_212#_c_65_p N_X_c_134_n 0.0108006f $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_56 N_A_75_212#_M1003_g N_X_c_132_n 0.00632981f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_57 N_A_75_212#_M1000_g N_X_c_132_n 0.00357773f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_58 N_A_75_212#_c_41_n N_X_c_132_n 0.0070136f $X=0.625 $Y=1.535 $X2=0 $Y2=0
cc_59 N_A_75_212#_c_63_p N_X_c_132_n 0.00240564f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_60 N_A_75_212#_c_65_p N_X_c_132_n 0.00132477f $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_61 N_A_75_212#_c_37_n N_X_c_132_n 0.0245251f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_62 N_A_75_212#_c_38_n N_X_c_132_n 0.00753248f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_63 N_A_75_212#_c_39_n N_X_c_132_n 0.0123683f $X=0.567 $Y=1.06 $X2=0 $Y2=0
cc_64 N_A_75_212#_c_42_n N_VPWR_M1000_d 7.12223e-19 $X=1.035 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_75_212#_c_65_p N_VPWR_M1000_d 0.00119515f $X=0.71 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_75_212#_M1000_g N_VPWR_c_156_n 0.0118404f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_67 N_A_75_212#_c_42_n N_VPWR_c_156_n 0.00690111f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_68 N_A_75_212#_c_65_p N_VPWR_c_156_n 0.0100761f $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_69 N_A_75_212#_c_37_n N_VPWR_c_156_n 4.75835e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_70 N_A_75_212#_c_38_n N_VPWR_c_156_n 3.07082e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_71 N_A_75_212#_M1002_d VPWR 0.00525232f $X=0.985 $Y=1.695 $X2=0 $Y2=0
cc_72 N_A_75_212#_M1000_g VPWR 0.00946027f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_73 N_A_75_212#_c_83_p VPWR 0.00646998f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_74 N_A_75_212#_M1000_g N_VPWR_c_158_n 0.00505556f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_75 N_A_75_212#_c_83_p N_VPWR_c_159_n 0.0116048f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_76 N_A_75_212#_c_36_n N_VGND_M1003_d 6.85198e-19 $X=1.035 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_75_212#_c_63_p N_VGND_M1003_d 0.00114971f $X=0.71 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_75_212#_M1003_g N_VGND_c_179_n 0.00801602f $X=0.47 $Y=0.495 $X2=0
+ $Y2=0
cc_79 N_A_75_212#_c_36_n N_VGND_c_179_n 0.00647139f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_80 N_A_75_212#_c_63_p N_VGND_c_179_n 0.00945604f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_81 N_A_75_212#_c_37_n N_VGND_c_179_n 3.89729e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_82 N_A_75_212#_c_38_n N_VGND_c_179_n 2.51407e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_83 N_A_75_212#_M1001_d VGND 0.00369894f $X=0.985 $Y=0.235 $X2=0 $Y2=0
cc_84 N_A_75_212#_M1003_g VGND 0.00957284f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A_75_212#_c_36_n VGND 0.0050992f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_86 N_A_75_212#_c_63_p VGND 8.54935e-19 $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_87 N_A_75_212#_c_97_p VGND 0.00643448f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_75_212#_M1003_g N_VGND_c_181_n 0.00505556f $X=0.47 $Y=0.495 $X2=0
+ $Y2=0
cc_89 N_A_75_212#_c_36_n N_VGND_c_182_n 0.00260015f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_90 N_A_75_212#_c_97_p N_VGND_c_182_n 0.01143f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_c_106_n N_VPWR_c_156_n 0.0118915f $X=0.925 $Y=1.62 $X2=0 $Y2=0
cc_92 N_A_c_106_n VPWR 0.00946027f $X=0.925 $Y=1.62 $X2=0 $Y2=0
cc_93 N_A_c_106_n N_VPWR_c_159_n 0.00505556f $X=0.925 $Y=1.62 $X2=0 $Y2=0
cc_94 N_A_c_101_n N_VGND_c_179_n 0.00787353f $X=0.91 $Y=0.83 $X2=0 $Y2=0
cc_95 N_A_c_101_n VGND 0.00526324f $X=0.91 $Y=0.83 $X2=0 $Y2=0
cc_96 N_A_c_101_n N_VGND_c_182_n 0.00367706f $X=0.91 $Y=0.83 $X2=0 $Y2=0
cc_97 N_X_M1000_s VPWR 0.00348182f $X=0.135 $Y=1.695 $X2=0 $Y2=0
cc_98 X VPWR 0.0103212f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_99 X N_VPWR_c_158_n 0.0183559f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_100 N_X_M1003_s VGND 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_101 X VGND 0.00990988f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_102 X N_VGND_c_181_n 0.0178762f $X=0.145 $Y=0.425 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o311ai_0.spice
* Created: Thu Aug 27 14:39:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o311ai_0.spice.pex"
.subckt sky130_fd_sc_hd__o311ai_0  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_138_47#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_138_47#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_138_47#_M1004_d N_A3_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1281 AS=0.0567 PD=1.03 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1007 A_458_47# N_B1_M1007_g N_A_138_47#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1281 PD=0.63 PS=1.03 NRD=14.28 NRS=95.712 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_C1_M1006_g A_458_47# VNB NSHORT L=0.15 W=0.42 AD=0.1176
+ AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1008 A_138_369# N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1792 PD=0.91 PS=1.84 NRD=24.625 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1001 A_222_369# N_A2_M1001_g A_138_369# VPB PHIGHVT L=0.15 W=0.64 AD=0.0864
+ AS=0.0864 PD=0.91 PS=0.91 NRD=24.625 NRS=24.625 M=1 R=4.26667 SA=75000.6
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1009 N_Y_M1009_d N_A3_M1009_g A_222_369# VPB PHIGHVT L=0.15 W=0.64 AD=0.144
+ AS=0.0864 PD=1.09 PS=0.91 NRD=26.1616 NRS=24.625 M=1 R=4.26667 SA=75001
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_Y_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1184 AS=0.144 PD=1.01 PS=1.09 NRD=13.8491 NRS=26.1616 M=1 R=4.26667
+ SA=75001.6 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1984 AS=0.1184 PD=1.9 PS=1.01 NRD=7.683 NRS=13.8491 M=1 R=4.26667
+ SA=75002.2 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o311ai_0.spice.SKY130_FD_SC_HD__O311AI_0.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_2.pxi.spice
* Created: Tue Sep  1 19:10:44 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%A N_A_M1001_g N_A_M1002_g N_A_c_39_n
+ N_A_c_40_n A N_A_c_42_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%A_27_47# N_A_27_47#_M1001_s
+ N_A_27_47#_M1002_s N_A_27_47#_c_72_n N_A_27_47#_M1003_g N_A_27_47#_c_77_n
+ N_A_27_47#_M1000_g N_A_27_47#_c_73_n N_A_27_47#_M1004_g N_A_27_47#_c_78_n
+ N_A_27_47#_M1005_g N_A_27_47#_c_74_n N_A_27_47#_c_80_n N_A_27_47#_c_81_n
+ N_A_27_47#_c_93_n N_A_27_47#_c_75_n N_A_27_47#_c_76_n N_A_27_47#_c_83_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%A_27_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%KAPWR N_KAPWR_M1002_d N_KAPWR_M1005_s
+ N_KAPWR_c_144_n N_KAPWR_c_145_n N_KAPWR_c_156_n N_KAPWR_c_146_n KAPWR
+ N_KAPWR_c_148_n KAPWR PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%X N_X_M1003_d N_X_M1000_d N_X_c_179_n
+ N_X_c_188_n N_X_c_182_n X X X X PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%X
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%VGND N_VGND_M1001_d N_VGND_M1004_s
+ N_VGND_c_222_n N_VGND_c_223_n N_VGND_c_224_n VGND N_VGND_c_225_n
+ N_VGND_c_226_n N_VGND_c_227_n N_VGND_c_228_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%VPWR VPWR N_VPWR_c_253_n
+ N_VPWR_c_252_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%VPWR
cc_1 VNB N_A_M1001_g 0.0270129f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_c_39_n 0.0169866f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.06
cc_3 VNB N_A_c_40_n 0.00513444f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.395
cc_4 VNB A 0.00679649f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_5 VNB N_A_c_42_n 0.0116517f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.065
cc_6 VNB N_A_27_47#_c_72_n 0.0156271f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_7 VNB N_A_27_47#_c_73_n 0.0174297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_74_n 0.0331156f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.065
cc_9 VNB N_A_27_47#_c_75_n 0.0625076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_76_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_X_c_179_n 3.57995e-19 $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=0.9
cc_12 VNB X 0.0126029f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.065
cc_13 VNB X 0.0204789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_222_n 0.00468168f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=0.9
cc_15 VNB N_VGND_c_223_n 0.0102408f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.395
cc_16 VNB N_VGND_c_224_n 0.013519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_225_n 0.0168654f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.85
cc_18 VNB N_VGND_c_226_n 0.014857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_227_n 0.0052624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_228_n 0.122794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_252_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=0.9
cc_22 VPB N_A_c_40_n 0.0294846f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.395
cc_23 VPB N_A_27_47#_c_77_n 0.014798f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.235
cc_24 VPB N_A_27_47#_c_78_n 0.018678f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.065
cc_25 VPB N_A_27_47#_c_74_n 0.00504729f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.065
cc_26 VPB N_A_27_47#_c_80_n 0.0282758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_27_47#_c_81_n 0.00572179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_c_75_n 0.0121119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_27_47#_c_83_n 0.0112463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_KAPWR_c_144_n 0.0122621f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_31 VPB N_KAPWR_c_145_n 0.00876329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_KAPWR_c_146_n 0.00846083f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.85
cc_33 VPB N_X_c_182_n 0.00920858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB X 0.0175394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_253_n 0.0518026f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.06
cc_36 VPB N_VPWR_c_252_n 0.0419517f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.9
cc_37 N_A_M1001_g N_A_27_47#_c_72_n 0.0164192f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_38 N_A_c_40_n N_A_27_47#_c_77_n 0.0193489f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_39 N_A_M1001_g N_A_27_47#_c_74_n 0.00813844f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_40 N_A_c_39_n N_A_27_47#_c_74_n 0.0146119f $X=0.505 $Y=1.06 $X2=0 $Y2=0
cc_41 N_A_c_40_n N_A_27_47#_c_74_n 4.92465e-19 $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_42 A N_A_27_47#_c_74_n 0.0373345f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_43 N_A_c_40_n N_A_27_47#_c_80_n 0.00287179f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_44 N_A_c_40_n N_A_27_47#_c_81_n 0.0190503f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_45 A N_A_27_47#_c_81_n 0.0279518f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_46 N_A_c_39_n N_A_27_47#_c_93_n 2.12331e-19 $X=0.505 $Y=1.06 $X2=0 $Y2=0
cc_47 N_A_c_40_n N_A_27_47#_c_93_n 8.99015e-19 $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_48 A N_A_27_47#_c_93_n 0.0183358f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_49 N_A_c_39_n N_A_27_47#_c_75_n 0.0325342f $X=0.505 $Y=1.06 $X2=0 $Y2=0
cc_50 A N_A_27_47#_c_75_n 0.0050302f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_51 N_A_c_40_n N_A_27_47#_c_83_n 5.49807e-19 $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_52 N_A_c_40_n N_KAPWR_c_145_n 0.00257081f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_53 N_A_c_40_n N_KAPWR_c_148_n 0.00735225f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_54 A X 0.00492153f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_55 A X 0.00519615f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_56 N_A_M1001_g N_VGND_c_222_n 0.00317144f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_57 N_A_c_39_n N_VGND_c_222_n 4.71188e-19 $X=0.505 $Y=1.06 $X2=0 $Y2=0
cc_58 A N_VGND_c_222_n 0.0166012f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VGND_c_225_n 0.00465542f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_60 A N_VGND_c_225_n 0.00178819f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_VGND_c_228_n 0.00771383f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_62 A N_VGND_c_228_n 0.0038034f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_40_n N_VPWR_c_253_n 0.0054895f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_64 N_A_c_40_n N_VPWR_c_252_n 0.00630403f $X=0.505 $Y=1.395 $X2=0 $Y2=0
cc_65 N_A_27_47#_c_81_n N_KAPWR_M1002_d 0.00270677f $X=0.965 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_27_47#_c_77_n N_KAPWR_c_144_n 0.00310566f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_67 N_A_27_47#_c_78_n N_KAPWR_c_144_n 0.00282671f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_68 N_A_27_47#_c_81_n N_KAPWR_c_144_n 0.00597432f $X=0.965 $Y=1.495 $X2=0
+ $Y2=0
cc_69 N_A_27_47#_M1002_s N_KAPWR_c_145_n 7.68319e-19 $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_70 N_A_27_47#_c_80_n N_KAPWR_c_145_n 0.028294f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_71 N_A_27_47#_c_81_n N_KAPWR_c_145_n 0.00468787f $X=0.965 $Y=1.495 $X2=0
+ $Y2=0
cc_72 N_A_27_47#_c_80_n N_KAPWR_c_156_n 4.3931e-19 $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_73 N_A_27_47#_c_81_n N_KAPWR_c_156_n 0.00137056f $X=0.965 $Y=1.495 $X2=0
+ $Y2=0
cc_74 N_A_27_47#_c_78_n N_KAPWR_c_146_n 0.00341733f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_80_n N_KAPWR_c_148_n 0.0243626f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_81_n N_KAPWR_c_148_n 0.0119975f $X=0.965 $Y=1.495 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_81_n N_X_M1000_d 0.00224161f $X=0.965 $Y=1.495 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_75_n N_X_c_179_n 6.13678e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_77_n N_X_c_188_n 7.45291e-19 $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_78_n N_X_c_188_n 6.74448e-19 $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_78_n N_X_c_182_n 0.0169371f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_81_n N_X_c_182_n 0.010554f $X=0.965 $Y=1.495 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_75_n N_X_c_182_n 4.12318e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_72_n X 0.00291318f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_73_n X 0.00702038f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_93_n X 0.0130886f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_75_n X 0.0170488f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_77_n X 0.00104199f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_78_n X 0.0130361f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_81_n X 0.0141986f $X=0.965 $Y=1.495 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_93_n X 0.0305477f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_75_n X 0.0244793f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_72_n N_VGND_c_222_n 0.00152531f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_72_n N_VGND_c_224_n 5.45981e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_73_n N_VGND_c_224_n 0.00813915f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_76_n N_VGND_c_225_n 0.017242f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_72_n N_VGND_c_226_n 0.00585385f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_73_n N_VGND_c_226_n 0.00341689f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1001_s N_VGND_c_228_n 0.00400903f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_72_n N_VGND_c_228_n 0.0106812f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_73_n N_VGND_c_228_n 0.0039829f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_76_n N_VGND_c_228_n 0.00981906f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_77_n N_VPWR_c_253_n 0.00585385f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_78_n N_VPWR_c_253_n 0.00425061f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_80_n N_VPWR_c_253_n 0.015543f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1002_s N_VPWR_c_252_n 0.00128591f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_77_n N_VPWR_c_252_n 0.00539971f $X=0.95 $Y=1.395 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_78_n N_VPWR_c_252_n 0.00581205f $X=1.37 $Y=1.395 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_80_n N_VPWR_c_252_n 0.00254601f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_110 N_KAPWR_c_144_n N_X_M1000_d 0.00121495f $X=1.435 $Y=2.24 $X2=0 $Y2=0
cc_111 N_KAPWR_c_144_n N_X_c_188_n 0.0145148f $X=1.435 $Y=2.24 $X2=0 $Y2=0
cc_112 N_KAPWR_c_156_n N_X_c_188_n 4.29016e-19 $X=0.84 $Y=2.21 $X2=0 $Y2=0
cc_113 N_KAPWR_c_146_n N_X_c_188_n 0.0136354f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_114 N_KAPWR_c_148_n N_X_c_188_n 0.00593488f $X=0.69 $Y=1.94 $X2=0 $Y2=0
cc_115 N_KAPWR_M1005_s N_X_c_182_n 0.00350959f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_116 N_KAPWR_c_144_n N_X_c_182_n 0.0148019f $X=1.435 $Y=2.24 $X2=0 $Y2=0
cc_117 N_KAPWR_c_146_n N_X_c_182_n 0.0173761f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_118 N_KAPWR_M1005_s X 0.00175457f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_119 N_KAPWR_c_144_n N_VPWR_c_253_n 0.00200978f $X=1.435 $Y=2.24 $X2=0 $Y2=0
cc_120 N_KAPWR_c_145_n N_VPWR_c_253_n 0.00137036f $X=0.55 $Y=2.21 $X2=0 $Y2=0
cc_121 N_KAPWR_c_146_n N_VPWR_c_253_n 0.0203984f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_122 N_KAPWR_c_148_n N_VPWR_c_253_n 0.0196112f $X=0.69 $Y=1.94 $X2=0 $Y2=0
cc_123 N_KAPWR_M1002_d N_VPWR_c_252_n 0.00141094f $X=0.55 $Y=1.485 $X2=0 $Y2=0
cc_124 N_KAPWR_M1005_s N_VPWR_c_252_n 0.0010704f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_125 N_KAPWR_c_145_n N_VPWR_c_252_n 0.174842f $X=0.55 $Y=2.21 $X2=0 $Y2=0
cc_126 N_KAPWR_c_146_n N_VPWR_c_252_n 0.00281098f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_127 N_KAPWR_c_148_n N_VPWR_c_252_n 0.00297304f $X=0.69 $Y=1.94 $X2=0 $Y2=0
cc_128 X N_VGND_c_224_n 0.0214173f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_129 N_X_c_179_n N_VGND_c_226_n 0.0122263f $X=1.16 $Y=0.42 $X2=0 $Y2=0
cc_130 X N_VGND_c_226_n 0.00275256f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_131 N_X_M1003_d N_VGND_c_228_n 0.0028269f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_132 N_X_c_179_n N_VGND_c_228_n 0.00771386f $X=1.16 $Y=0.42 $X2=0 $Y2=0
cc_133 X N_VGND_c_228_n 0.00550683f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_134 N_X_c_188_n N_VPWR_c_253_n 0.00976296f $X=1.16 $Y=2.27 $X2=0 $Y2=0
cc_135 N_X_c_182_n N_VPWR_c_253_n 0.00173573f $X=1.555 $Y=1.75 $X2=0 $Y2=0
cc_136 N_X_M1000_d N_VPWR_c_252_n 0.0013312f $X=1.025 $Y=1.485 $X2=0 $Y2=0
cc_137 N_X_c_188_n N_VPWR_c_252_n 0.00166426f $X=1.16 $Y=2.27 $X2=0 $Y2=0
cc_138 N_X_c_182_n N_VPWR_c_252_n 2.49894e-19 $X=1.555 $Y=1.75 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__tapvgnd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ends


* File: sky130_fd_sc_hd__dlrtp_2.pex.spice
* Created: Thu Aug 27 14:17:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRTP_2%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39414e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.21 $Y=1.19
+ $X2=0.21 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%A_27_47# 1 2 9 13 17 19 20 23 27 30 34 35 36
+ 41 44 46 49 50 53 56 57 60 64
c151 57 0 7.21753e-20 $X=2.535 $Y=1.53
c152 19 0 1.56925e-19 $X=3.135 $Y=1.325
c153 13 0 2.69707e-20 $X=0.89 $Y=2.135
c154 9 0 2.69707e-20 $X=0.89 $Y=0.445
r155 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r156 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.53
+ $X2=2.535 $Y2=1.53
r157 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r158 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r159 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.39 $Y=1.53
+ $X2=2.535 $Y2=1.53
r160 49 50 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.39 $Y=1.53
+ $X2=0.84 $Y2=1.53
r161 48 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r162 47 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r163 45 64 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r164 44 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r165 44 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r166 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r167 38 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r168 37 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r169 36 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r170 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r171 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r172 34 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r173 28 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r174 28 30 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r175 26 60 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r176 26 27 40.8463 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r177 25 60 26.6608 $w=2.7e-07 $l=1.2e-07 $layer=POLY_cond $X=2.67 $Y=1.4
+ $X2=2.67 $Y2=1.52
r178 21 23 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=3.21 $Y=1.25
+ $X2=3.21 $Y2=0.415
r179 20 25 72.6412 $w=8.6e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.325
+ $X2=2.67 $Y2=1.4
r180 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.135 $Y=1.325
+ $X2=3.21 $Y2=1.25
r181 19 20 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.135 $Y=1.325
+ $X2=2.805 $Y2=1.325
r182 17 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.725 $Y=2.275
+ $X2=2.725 $Y2=1.685
r183 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r184 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r185 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r186 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r187 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r188 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%D 3 7 9 13 15
c39 13 0 1.05996e-19 $X=1.605 $Y=1.04
r40 12 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.605 $Y=1.04
+ $X2=1.83 $Y2=1.04
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.04 $X2=1.605 $Y2=1.04
r42 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.605 $Y=1.19
+ $X2=1.605 $Y2=1.04
r43 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r44 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r45 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r46 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%A_299_47# 1 2 7 9 12 16 18 20 21 24 27 34
c85 34 0 1.28593e-19 $X=2.25 $Y=0.93
c86 20 0 4.79766e-21 $X=2.035 $Y=1.095
r87 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=0.93 $X2=2.25 $Y2=0.93
r88 27 29 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=1.61 $Y=0.51
+ $X2=1.61 $Y2=0.7
r89 21 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=1.495
+ $X2=2.035 $Y2=1.58
r90 20 33 8.95737 $w=3.17e-07 $l=2.11849e-07 $layer=LI1_cond $X=2.035 $Y=1.095
+ $X2=2.142 $Y2=0.93
r91 20 21 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.035 $Y=1.095
+ $X2=2.035 $Y2=1.495
r92 19 29 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7 $X2=1.61
+ $Y2=0.7
r93 18 33 8.85174 $w=3.17e-07 $l=3.11545e-07 $layer=LI1_cond $X=1.95 $Y=0.7
+ $X2=2.142 $Y2=0.93
r94 18 19 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.95 $Y=0.7
+ $X2=1.705 $Y2=0.7
r95 14 24 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.61 $Y=1.58
+ $X2=2.035 $Y2=1.58
r96 14 16 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.61 $Y=1.665
+ $X2=1.61 $Y2=1.99
r97 10 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.095
+ $X2=2.25 $Y2=0.93
r98 10 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=1.095
+ $X2=2.25 $Y2=2.165
r99 7 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.765
+ $X2=2.25 $Y2=0.93
r100 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.765
+ $X2=2.25 $Y2=0.445
r101 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r102 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%A_193_47# 1 2 9 13 17 19 22 25 26 28 29 32
+ 35 42 43
c127 43 0 1.73085e-19 $X=3.18 $Y=1.745
c128 42 0 7.21753e-20 $X=3.18 $Y=1.745
c129 25 0 2.48451e-19 $X=3.015 $Y=1.57
c130 22 0 3.79282e-19 $X=2.76 $Y=0.905
c131 19 0 1.56925e-19 $X=2.93 $Y=0.887
c132 9 0 4.79766e-21 $X=2.725 $Y=0.415
r133 42 45 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.745
+ $X2=3.18 $Y2=1.88
r134 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.745 $X2=3.18 $Y2=1.745
r135 35 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.01 $Y=1.87
+ $X2=3.01 $Y2=1.87
r136 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r137 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r138 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.865 $Y=1.87
+ $X2=3.01 $Y2=1.87
r139 28 29 1.93688 $w=1.4e-07 $l=1.565e-06 $layer=MET1_cond $X=2.865 $Y=1.87
+ $X2=1.3 $Y2=1.87
r140 26 32 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r141 26 27 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r142 25 43 9.32846 $w=3.29e-07 $l=2.07063e-07 $layer=LI1_cond $X=3.015 $Y=1.57
+ $X2=3.085 $Y2=1.745
r143 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.015 $Y=1.04
+ $X2=3.015 $Y2=1.57
r144 22 39 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=0.905
+ $X2=2.76 $Y2=0.77
r145 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=0.905 $X2=2.76 $Y2=0.905
r146 19 24 7.55824 $w=3.05e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.93 $Y=0.887
+ $X2=3.015 $Y2=1.04
r147 19 21 6.42345 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=2.93 $Y=0.887
+ $X2=2.76 $Y2=0.887
r148 17 27 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r149 13 45 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.145 $Y=2.275
+ $X2=3.145 $Y2=1.88
r150 9 39 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=2.725 $Y=0.415
+ $X2=2.725 $Y2=0.77
r151 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r152 1 17 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%A_711_307# 1 2 9 13 17 19 21 22 24 27 29 32
+ 36 39 42 44 46 48 49 51 52 53 67
c146 67 0 2.66825e-20 $X=5.97 $Y=1.16
c147 32 0 1.67596e-19 $X=3.86 $Y=1.7
c148 13 0 8.08555e-20 $X=3.685 $Y=0.445
c149 9 0 1.73085e-19 $X=3.63 $Y=2.275
r150 66 67 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.55 $Y=1.16
+ $X2=5.97 $Y2=1.16
r151 58 60 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.63 $Y=1.7
+ $X2=3.685 $Y2=1.7
r152 57 66 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.53 $Y=1.16 $X2=5.55
+ $Y2=1.16
r153 57 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.53 $Y=1.16
+ $X2=5.515 $Y2=1.16
r154 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.16 $X2=5.53 $Y2=1.16
r155 54 56 25.0595 $w=1.85e-07 $l=3.8e-07 $layer=LI1_cond $X=5.515 $Y=0.78
+ $X2=5.515 $Y2=1.16
r156 52 53 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=4.955 $Y=0.76
+ $X2=5.095 $Y2=0.76
r157 48 56 10.9829 $w=1.85e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.5 $Y=1.325
+ $X2=5.515 $Y2=1.16
r158 48 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.5 $Y=1.325
+ $X2=5.5 $Y2=1.535
r159 46 54 1.22693 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.415 $Y=0.78
+ $X2=5.515 $Y2=0.78
r160 46 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.415 $Y=0.78
+ $X2=5.095 $Y2=0.78
r161 45 51 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.97 $Y=1.62
+ $X2=4.885 $Y2=1.7
r162 44 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=1.62
+ $X2=5.5 $Y2=1.535
r163 44 45 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.415 $Y=1.62
+ $X2=4.97 $Y2=1.62
r164 40 51 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=1.865
+ $X2=4.885 $Y2=1.7
r165 40 42 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.885 $Y=1.865
+ $X2=4.885 $Y2=2.27
r166 39 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.58 $Y=0.74
+ $X2=4.955 $Y2=0.74
r167 34 39 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.41 $Y=0.655
+ $X2=4.58 $Y2=0.74
r168 34 36 8.64332 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=4.41 $Y=0.655
+ $X2=4.41 $Y2=0.4
r169 32 60 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.86 $Y=1.7
+ $X2=3.685 $Y2=1.7
r170 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.86
+ $Y=1.7 $X2=3.86 $Y2=1.7
r171 29 51 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=1.7 $X2=4.885
+ $Y2=1.7
r172 29 31 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=4.8 $Y=1.7 $X2=3.86
+ $Y2=1.7
r173 25 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.325
+ $X2=5.97 $Y2=1.16
r174 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.97 $Y=1.325
+ $X2=5.97 $Y2=1.985
r175 22 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=1.16
r176 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=0.56
r177 19 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.55 $Y=0.995
+ $X2=5.55 $Y2=1.16
r178 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.55 $Y=0.995
+ $X2=5.55 $Y2=0.56
r179 15 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.515 $Y=1.325
+ $X2=5.515 $Y2=1.16
r180 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.515 $Y=1.325
+ $X2=5.515 $Y2=1.985
r181 11 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=1.535
+ $X2=3.685 $Y2=1.7
r182 11 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.685 $Y=1.535
+ $X2=3.685 $Y2=0.445
r183 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=1.7
r184 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=2.275
r185 2 51 600 $w=1.7e-07 $l=3.505e-07 $layer=licon1_PDIFF $count=1 $X=4.7
+ $Y=1.485 $X2=4.885 $Y2=1.755
r186 2 42 600 $w=1.7e-07 $l=8.72611e-07 $layer=licon1_PDIFF $count=1 $X=4.7
+ $Y=1.485 $X2=4.885 $Y2=2.27
r187 1 36 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.29
+ $Y=0.235 $X2=4.415 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%A_560_47# 1 2 9 13 15 16 17 21 26 28 30 31
+ 33
c95 33 0 1.02902e-19 $X=4.135 $Y=1.16
c96 31 0 3.14158e-20 $X=3.605 $Y=1.16
c97 26 0 1.66981e-19 $X=3.357 $Y=0.995
r98 36 38 5.69237 $w=3.28e-07 $l=1.63e-07 $layer=LI1_cond $X=3.357 $Y=1.16
+ $X2=3.52 $Y2=1.16
r99 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.16 $X2=4.135 $Y2=1.16
r100 31 38 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=3.52 $Y2=1.16
r101 31 33 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=4.135 $Y2=1.16
r102 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.16
r103 29 30 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.985
r104 27 30 6.32124 $w=1.93e-07 $l=1.11803e-07 $layer=LI1_cond $X=3.495 $Y=2.085
+ $X2=3.52 $Y2=1.985
r105 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.495 $Y=2.085
+ $X2=3.495 $Y2=2.255
r106 26 36 4.47052 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=3.357 $Y=0.995
+ $X2=3.357 $Y2=1.16
r107 25 26 29.1532 $w=1.73e-07 $l=4.6e-07 $layer=LI1_cond $X=3.357 $Y=0.535
+ $X2=3.357 $Y2=0.995
r108 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=2.34
+ $X2=3.495 $Y2=2.255
r109 21 23 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.41 $Y=2.34
+ $X2=2.935 $Y2=2.34
r110 17 25 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.27 $Y=0.45
+ $X2=3.357 $Y2=0.535
r111 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.27 $Y=0.45
+ $X2=2.935 $Y2=0.45
r112 15 34 92.2021 $w=2.7e-07 $l=4.15e-07 $layer=POLY_cond $X=4.55 $Y=1.16
+ $X2=4.135 $Y2=1.16
r113 15 16 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.55 $Y=1.16
+ $X2=4.625 $Y2=1.16
r114 11 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.625 $Y=1.295
+ $X2=4.625 $Y2=1.16
r115 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.625 $Y=1.295
+ $X2=4.625 $Y2=1.985
r116 7 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.625 $Y=1.025
+ $X2=4.625 $Y2=1.16
r117 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.625 $Y=1.025
+ $X2=4.625 $Y2=0.56
r118 2 23 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=2.065 $X2=2.935 $Y2=2.34
r119 1 19 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.935 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%RESET_B 3 6 8 12 13 14 16 18
c47 12 0 1.02902e-19 $X=5.05 $Y=1.16
r48 16 18 1.58958 $w=2.88e-07 $l=4e-08 $layer=LI1_cond $X=4.815 $Y=1.18
+ $X2=4.855 $Y2=1.18
r49 12 15 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=5.047 $Y=1.16
+ $X2=5.047 $Y2=1.325
r50 12 14 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=5.047 $Y=1.16
+ $X2=5.047 $Y2=0.995
r51 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.16 $X2=5.05 $Y2=1.16
r52 8 16 1.06065 $w=3.3e-07 $l=2.3e-08 $layer=LI1_cond $X=4.792 $Y=1.18
+ $X2=4.815 $Y2=1.18
r53 8 13 6.87492 $w=2.88e-07 $l=1.73e-07 $layer=LI1_cond $X=4.877 $Y=1.18
+ $X2=5.05 $Y2=1.18
r54 8 18 0.874267 $w=2.88e-07 $l=2.2e-08 $layer=LI1_cond $X=4.877 $Y=1.18
+ $X2=4.855 $Y2=1.18
r55 6 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.095 $Y=1.985
+ $X2=5.095 $Y2=1.325
r56 3 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.095 $Y=0.56
+ $X2=5.095 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%VPWR 1 2 3 4 5 6 21 25 29 31 35 39 41 43 45
+ 47 52 57 65 70 76 79 82 85 88 92
r107 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r108 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r109 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r110 83 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r111 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r112 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r113 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 74 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 74 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r116 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r117 71 88 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.312 $Y2=2.72
r118 71 73 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.75 $Y2=2.72
r119 70 91 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.267 $Y2=2.72
r120 70 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r121 69 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r122 69 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r123 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r124 66 85 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.56 $Y=2.72 $X2=4.42
+ $Y2=2.72
r125 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.56 $Y=2.72
+ $X2=4.83 $Y2=2.72
r126 65 88 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.14 $Y=2.72
+ $X2=5.312 $Y2=2.72
r127 65 68 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.14 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r130 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r131 61 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 58 79 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.102 $Y2=2.72
r135 58 60 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 57 82 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.75 $Y=2.72
+ $X2=3.92 $Y2=2.72
r137 57 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.75 $Y=2.72 $X2=3.45
+ $Y2=2.72
r138 56 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r139 56 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r140 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r141 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r142 53 55 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r143 52 79 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.102 $Y2=2.72
r144 52 55 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r145 47 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r146 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 45 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 45 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r149 41 91 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.225 $Y=2.635
+ $X2=6.267 $Y2=2.72
r150 41 43 35.4598 $w=2.58e-07 $l=8e-07 $layer=LI1_cond $X=6.225 $Y=2.635
+ $X2=6.225 $Y2=1.835
r151 37 88 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.312 $Y=2.635
+ $X2=5.312 $Y2=2.72
r152 37 39 20.5435 $w=3.43e-07 $l=6.15e-07 $layer=LI1_cond $X=5.312 $Y=2.635
+ $X2=5.312 $Y2=2.02
r153 33 85 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.635
+ $X2=4.42 $Y2=2.72
r154 33 35 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.42 $Y=2.635
+ $X2=4.42 $Y2=2.34
r155 32 82 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.09 $Y=2.72
+ $X2=3.92 $Y2=2.72
r156 31 85 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.28 $Y=2.72 $X2=4.42
+ $Y2=2.72
r157 31 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.28 $Y=2.72
+ $X2=4.09 $Y2=2.72
r158 27 82 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.72
r159 27 29 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.34
r160 23 79 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.102 $Y=2.635
+ $X2=2.102 $Y2=2.72
r161 23 25 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=2.102 $Y=2.635
+ $X2=2.102 $Y2=2
r162 19 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r163 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r164 6 43 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=1.835
r165 5 39 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.17
+ $Y=1.485 $X2=5.305 $Y2=2.02
r166 4 35 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.485 $X2=4.405 $Y2=2.34
r167 3 29 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=2.065 $X2=3.84 $Y2=2.34
r168 2 25 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r169 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%Q 1 2 8 14 16 17 18 19 20 21 31 37
r47 31 37 0.81742 $w=5.97e-07 $l=4.69042e-08 $layer=LI1_cond $X=6.07 $Y=0.89
+ $X2=6.055 $Y2=0.85
r48 20 37 0.470017 $w=5.97e-07 $l=2.3e-08 $layer=LI1_cond $X=6.055 $Y=0.827
+ $X2=6.055 $Y2=0.85
r49 20 21 5.83351 $w=5.68e-07 $l=2.78e-07 $layer=LI1_cond $X=6.07 $Y=0.912
+ $X2=6.07 $Y2=1.19
r50 20 31 0.461644 $w=5.68e-07 $l=2.2e-08 $layer=LI1_cond $X=6.07 $Y=0.912
+ $X2=6.07 $Y2=0.89
r51 19 29 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=5.79 $Y=2.21 $X2=5.79
+ $Y2=2.3
r52 18 21 4.09185 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.07 $Y=1.385
+ $X2=6.07 $Y2=1.19
r53 16 19 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=5.79 $Y=2.01 $X2=5.79
+ $Y2=2.21
r54 16 17 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.79 $Y=2.01
+ $X2=5.79 $Y2=1.875
r55 12 14 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=5.76 $Y=0.37 $X2=5.84
+ $Y2=0.37
r56 9 18 2.36195 $w=5.94e-07 $l=2.81691e-07 $layer=LI1_cond $X=5.84 $Y=1.5
+ $X2=6.07 $Y2=1.385
r57 9 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.84 $Y=1.5 $X2=5.84
+ $Y2=1.875
r58 8 20 8.23439 $w=5.97e-07 $l=2.44039e-07 $layer=LI1_cond $X=5.84 $Y=0.765
+ $X2=6.055 $Y2=0.827
r59 7 14 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.84 $Y=0.485
+ $X2=5.84 $Y2=0.37
r60 7 8 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.84 $Y=0.485 $X2=5.84
+ $Y2=0.765
r61 2 29 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.59
+ $Y=1.485 $X2=5.74 $Y2=2.3
r62 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.76 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_2%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 56 61 67 70 73 76 80
c107 80 0 2.71124e-20 $X=6.21 $Y=0
c108 48 0 1.80885e-19 $X=3.72 $Y=0
c109 30 0 2.66825e-20 $X=5.34 $Y=0.36
c110 22 0 2.25971e-20 $X=2.04 $Y=0.36
r111 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r112 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r113 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r114 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r115 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 65 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r117 65 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r118 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r119 62 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0 $X2=5.34
+ $Y2=0
r120 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.425 $Y=0
+ $X2=5.75 $Y2=0
r121 61 79 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.267 $Y2=0
r122 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.75
+ $Y2=0
r123 60 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r124 60 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r125 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r126 57 73 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.06 $Y=0 $X2=3.89
+ $Y2=0
r127 57 59 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.06 $Y=0 $X2=4.37
+ $Y2=0
r128 56 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.255 $Y=0 $X2=5.34
+ $Y2=0
r129 56 59 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=5.255 $Y=0 $X2=4.37
+ $Y2=0
r130 55 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r131 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r132 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r133 52 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r134 51 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r135 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r136 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r137 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r138 48 73 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.89
+ $Y2=0
r139 48 54 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.45
+ $Y2=0
r140 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r141 47 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r142 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r143 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r144 44 46 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r145 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r146 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r147 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r148 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r149 36 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r150 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r151 32 79 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.267 $Y2=0
r152 32 34 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0.38
r153 28 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0
r154 28 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0.36
r155 24 73 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=0.085
+ $X2=3.89 $Y2=0
r156 24 26 12.2023 $w=3.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.89 $Y=0.085
+ $X2=3.89 $Y2=0.445
r157 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r158 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r159 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r160 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r161 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.38
r162 4 30 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=5.17
+ $Y=0.235 $X2=5.34 $Y2=0.36
r163 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.235 $X2=3.895 $Y2=0.445
r164 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r165 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o211ai_1.pxi.spice
* Created: Tue Sep  1 19:20:47 2020
* 
x_PM_SKY130_FD_SC_HD__O211AI_1%A1 N_A1_M1002_g N_A1_M1003_g A1 N_A1_c_46_n
+ N_A1_c_47_n PM_SKY130_FD_SC_HD__O211AI_1%A1
x_PM_SKY130_FD_SC_HD__O211AI_1%A2 N_A2_M1001_g N_A2_M1004_g N_A2_c_71_n
+ N_A2_c_72_n A2 N_A2_c_73_n PM_SKY130_FD_SC_HD__O211AI_1%A2
x_PM_SKY130_FD_SC_HD__O211AI_1%B1 N_B1_M1005_g N_B1_M1006_g B1 B1 N_B1_c_109_n
+ N_B1_c_110_n PM_SKY130_FD_SC_HD__O211AI_1%B1
x_PM_SKY130_FD_SC_HD__O211AI_1%C1 N_C1_c_141_n N_C1_M1007_g N_C1_M1000_g C1
+ N_C1_c_142_n N_C1_c_143_n PM_SKY130_FD_SC_HD__O211AI_1%C1
x_PM_SKY130_FD_SC_HD__O211AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_c_171_n
+ N_VPWR_c_172_n N_VPWR_c_173_n VPWR N_VPWR_c_174_n N_VPWR_c_175_n
+ N_VPWR_c_170_n N_VPWR_c_177_n PM_SKY130_FD_SC_HD__O211AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O211AI_1%Y N_Y_M1007_d N_Y_M1001_d N_Y_M1000_d N_Y_c_211_n
+ N_Y_c_215_n N_Y_c_237_n N_Y_c_218_n N_Y_c_214_n Y N_Y_c_212_n
+ PM_SKY130_FD_SC_HD__O211AI_1%Y
x_PM_SKY130_FD_SC_HD__O211AI_1%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1004_d
+ N_A_27_47#_c_250_n N_A_27_47#_c_253_n N_A_27_47#_c_251_n N_A_27_47#_c_261_n
+ N_A_27_47#_c_268_p PM_SKY130_FD_SC_HD__O211AI_1%A_27_47#
x_PM_SKY130_FD_SC_HD__O211AI_1%VGND N_VGND_M1002_d N_VGND_c_274_n VGND
+ N_VGND_c_275_n N_VGND_c_276_n N_VGND_c_277_n N_VGND_c_278_n
+ PM_SKY130_FD_SC_HD__O211AI_1%VGND
cc_1 VNB A1 0.0125518f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_2 VNB N_A1_c_46_n 0.0317275f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_3 VNB N_A1_c_47_n 0.0232607f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.995
cc_4 VNB N_A2_c_71_n 0.00337049f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_5 VNB N_A2_c_72_n 0.0237978f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.995
cc_6 VNB N_A2_c_73_n 0.0185641f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB B1 0.0135722f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_B1_c_109_n 0.0222936f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.995
cc_9 VNB N_B1_c_110_n 0.0169284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_C1_c_141_n 0.0195269f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_11 VNB N_C1_c_142_n 0.034594f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.995
cc_12 VNB N_C1_c_143_n 0.00244002f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=1.325
cc_13 VNB N_VPWR_c_170_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_211_n 0.0232932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Y_c_212_n 0.0266214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_250_n 0.0141804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_251_n 0.00921527f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_18 VNB N_VGND_c_274_n 0.0055721f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_19 VNB N_VGND_c_275_n 0.0170734f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=1.16
cc_20 VNB N_VGND_c_276_n 0.0497381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_277_n 0.162421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_278_n 0.00630985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VPB N_A1_M1003_g 0.0246947f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_24 VPB A1 0.00195821f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_25 VPB N_A1_c_46_n 0.00737518f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_26 VPB N_A2_M1001_g 0.0186932f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_27 VPB N_A2_c_71_n 5.58377e-19 $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_28 VPB N_A2_c_72_n 0.00711074f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.995
cc_29 VPB A2 0.0018837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_B1_M1005_g 0.0194538f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_31 VPB B1 0.00246253f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_B1_c_109_n 0.00832628f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.995
cc_33 VPB N_C1_M1000_g 0.0243129f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_34 VPB N_C1_c_142_n 0.0098219f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.995
cc_35 VPB N_C1_c_143_n 0.00167263f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=1.325
cc_36 VPB N_VPWR_c_171_n 0.0103398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_172_n 0.0383737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_173_n 0.00295613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_174_n 0.0255781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_175_n 0.0259849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_170_n 0.0437029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_177_n 0.00521838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_Y_c_211_n 0.0212792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_Y_c_214_n 0.0281471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 N_A1_M1003_g N_A2_M1001_g 0.0484957f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_46 A1 N_A2_c_71_n 0.0224666f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A1_c_46_n N_A2_c_71_n 0.00263499f $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_48 A1 N_A2_c_72_n 2.50948e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A1_c_46_n N_A2_c_72_n 0.0484957f $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_50 N_A1_M1003_g A2 0.00613049f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_51 N_A1_c_47_n N_A2_c_73_n 0.0223869f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A1_M1003_g N_VPWR_c_172_n 0.017933f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_53 A1 N_VPWR_c_172_n 0.0170103f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A1_c_46_n N_VPWR_c_172_n 0.00480561f $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A1_M1003_g N_VPWR_c_174_n 0.00486043f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_56 N_A1_M1003_g N_VPWR_c_170_n 0.00814024f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A1_c_47_n N_A_27_47#_c_250_n 0.00551286f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_58 N_A1_c_47_n N_A_27_47#_c_253_n 0.013941f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_59 A1 N_A_27_47#_c_251_n 0.0225513f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_60 N_A1_c_46_n N_A_27_47#_c_251_n 0.00504127f $X=0.31 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A1_c_47_n N_A_27_47#_c_251_n 0.00164474f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A1_c_47_n N_VGND_c_274_n 0.00427574f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A1_c_47_n N_VGND_c_275_n 0.0041289f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A1_c_47_n N_VGND_c_277_n 0.00681546f $X=0.362 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A2_c_71_n B1 0.015545f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A2_c_72_n B1 0.0012505f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A2_M1001_g N_B1_c_109_n 0.0200969f $X=0.835 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A2_c_71_n N_B1_c_109_n 3.52567e-19 $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A2_c_72_n N_B1_c_109_n 0.020758f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_70 A2 N_B1_c_109_n 0.00103545f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_71 N_A2_c_73_n N_B1_c_110_n 0.0169403f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A2_M1001_g N_VPWR_c_172_n 0.00239535f $X=0.835 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A2_M1001_g N_VPWR_c_173_n 0.00105516f $X=0.835 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A2_M1001_g N_VPWR_c_174_n 0.00567951f $X=0.835 $Y=1.985 $X2=0 $Y2=0
cc_75 A2 N_VPWR_c_174_n 0.00406515f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_76 N_A2_M1001_g N_VPWR_c_170_n 0.0104874f $X=0.835 $Y=1.985 $X2=0 $Y2=0
cc_77 A2 N_VPWR_c_170_n 0.00561063f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_78 A2 A_110_297# 0.0014015f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_79 N_A2_c_71_n N_Y_c_215_n 0.00129848f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A2_c_72_n N_Y_c_215_n 0.0055705f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A2_c_73_n N_A_27_47#_c_250_n 5.60696e-19 $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A2_c_71_n N_A_27_47#_c_253_n 0.0264545f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A2_c_72_n N_A_27_47#_c_253_n 0.00451511f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A2_c_73_n N_A_27_47#_c_253_n 0.0175094f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A2_c_73_n N_VGND_c_274_n 0.00326685f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A2_c_73_n N_VGND_c_276_n 0.00422112f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A2_c_73_n N_VGND_c_277_n 0.0061748f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B1_c_110_n N_C1_c_141_n 0.0382142f $X=1.465 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_89 N_B1_M1005_g N_C1_M1000_g 0.0299692f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_90 B1 N_C1_c_142_n 0.00537356f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_91 N_B1_c_109_n N_C1_c_142_n 0.0382142f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_92 B1 N_C1_c_143_n 0.0372336f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B1_c_109_n N_C1_c_143_n 2.11598e-19 $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_94 B1 N_VPWR_M1005_d 0.0044971f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B1_M1005_g N_VPWR_c_173_n 0.00654544f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_96 N_B1_M1005_g N_VPWR_c_174_n 0.00415785f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B1_M1005_g N_VPWR_c_170_n 0.00504548f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_98 B1 N_Y_c_211_n 0.00248917f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B1_M1005_g N_Y_c_218_n 0.013783f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_100 B1 N_Y_c_218_n 0.0250963f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B1_c_109_n N_Y_c_218_n 5.79761e-19 $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B1_M1005_g N_Y_c_214_n 7.78793e-19 $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_c_110_n N_Y_c_212_n 0.0016788f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_104 B1 N_A_27_47#_c_261_n 0.0112784f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_105 N_B1_c_109_n N_A_27_47#_c_261_n 0.00109624f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B1_c_110_n N_VGND_c_276_n 0.00585385f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_c_110_n N_VGND_c_277_n 0.0108951f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_108 N_C1_M1000_g N_VPWR_c_173_n 0.00521722f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_109 N_C1_M1000_g N_VPWR_c_175_n 0.00423594f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_110 N_C1_M1000_g N_VPWR_c_170_n 0.00741047f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_111 N_C1_c_143_n N_Y_M1000_d 0.00517677f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C1_c_141_n N_Y_c_211_n 0.00329063f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_113 N_C1_M1000_g N_Y_c_211_n 0.00612419f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_114 N_C1_c_142_n N_Y_c_211_n 0.00386675f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C1_c_143_n N_Y_c_211_n 0.0430183f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C1_M1000_g N_Y_c_218_n 0.015453f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_117 N_C1_c_143_n N_Y_c_218_n 0.020954f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C1_M1000_g N_Y_c_214_n 0.00763549f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_119 N_C1_c_142_n N_Y_c_214_n 0.00107603f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C1_c_141_n N_Y_c_212_n 0.0107379f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_121 N_C1_c_142_n N_Y_c_212_n 0.00667683f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C1_c_143_n N_Y_c_212_n 0.0200206f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_123 N_C1_c_141_n N_VGND_c_276_n 0.00547467f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_124 N_C1_c_141_n N_VGND_c_277_n 0.0110397f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_125 N_VPWR_c_170_n A_110_297# 0.00385482f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_126 N_VPWR_c_170_n N_Y_M1001_d 0.0044771f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_127 N_VPWR_c_170_n N_Y_M1000_d 0.00516805f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_128 N_VPWR_c_174_n N_Y_c_237_n 0.018848f $X=1.445 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_170_n N_Y_c_237_n 0.0125105f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_130 N_VPWR_M1005_d N_Y_c_218_n 0.00667527f $X=1.45 $Y=1.485 $X2=0 $Y2=0
cc_131 N_VPWR_c_173_n N_Y_c_218_n 0.0162136f $X=1.61 $Y=2.36 $X2=0 $Y2=0
cc_132 N_VPWR_c_174_n N_Y_c_218_n 0.00241332f $X=1.445 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_175_n N_Y_c_218_n 0.00267427f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_134 N_VPWR_c_170_n N_Y_c_218_n 0.0104913f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_c_173_n N_Y_c_214_n 0.0137599f $X=1.61 $Y=2.36 $X2=0 $Y2=0
cc_136 N_VPWR_c_175_n N_Y_c_214_n 0.0467484f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_137 N_VPWR_c_170_n N_Y_c_214_n 0.0267653f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_138 N_Y_c_212_n N_VGND_c_276_n 0.0471777f $X=2.572 $Y=0.55 $X2=0 $Y2=0
cc_139 N_Y_M1007_d N_VGND_c_277_n 0.00492208f $X=1.99 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Y_c_212_n N_VGND_c_277_n 0.0270403f $X=2.572 $Y=0.55 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_253_n N_VGND_M1002_d 0.00583929f $X=1.125 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_142 N_A_27_47#_c_253_n N_VGND_c_274_n 0.0212122f $X=1.125 $Y=0.72 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_250_n N_VGND_c_275_n 0.0208048f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_253_n N_VGND_c_275_n 0.0026189f $X=1.125 $Y=0.72 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_253_n N_VGND_c_276_n 0.00311196f $X=1.125 $Y=0.72 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_268_p N_VGND_c_276_n 0.0210051f $X=1.29 $Y=0.38 $X2=0 $Y2=0
cc_147 N_A_27_47#_M1002_s N_VGND_c_277_n 0.00213418f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_M1004_d N_VGND_c_277_n 0.00410115f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_250_n N_VGND_c_277_n 0.0123922f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_253_n N_VGND_c_277_n 0.0108339f $X=1.125 $Y=0.72 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_268_p N_VGND_c_277_n 0.012574f $X=1.29 $Y=0.38 $X2=0 $Y2=0
cc_152 N_VGND_c_277_n A_326_47# 0.00897657f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

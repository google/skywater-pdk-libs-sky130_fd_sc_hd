* File: sky130_fd_sc_hd__dlrtn_1.pex.spice
* Created: Thu Aug 27 14:17:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRTN_1%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%A_27_47# 1 2 9 13 17 20 24 28 29 30 38 42 45
+ 47 52 54 56 57 60 63 64 68 71 75 79
c167 20 0 1.41946e-19 $X=3.335 $Y=2.275
c168 13 0 2.6965e-20 $X=0.89 $Y=2.135
c169 9 0 2.6965e-20 $X=0.89 $Y=0.445
r170 64 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.095 $Y=1.53
+ $X2=3.095 $Y2=1.415
r171 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.53
+ $X2=3.015 $Y2=1.53
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r173 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=3.015 $Y2=1.53
r175 56 57 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=0.84 $Y2=1.53
r176 52 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.87
+ $X2=2.8 $Y2=0.705
r177 51 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0.87
+ $X2=3.01 $Y2=0.87
r178 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=0.87 $X2=2.8 $Y2=0.87
r179 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r180 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r181 46 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r182 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r183 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r184 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r185 39 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.335 $Y2=1.74
r186 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r187 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.53
r188 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.74
r189 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=0.87
r190 34 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.415
r191 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r192 31 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r193 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r194 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r195 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r196 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r197 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r198 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r199 18 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=1.74
r200 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=2.275
r201 17 71 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.79 $Y=0.415
+ $X2=2.79 $Y2=0.705
r202 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r203 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r204 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r206 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 32 0 1.12109e-19 $X=2.255 $Y=0.93
c84 18 0 7.13094e-20 $X=1.97 $Y=0.7
r85 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r86 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r87 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r88 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r89 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r90 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r92 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r93 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r94 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r95 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r96 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r97 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r98 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r99 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r101 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c113 38 0 1.41946e-19 $X=2.67 $Y=1.52
r114 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r115 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.612 $Y=1.87
+ $X2=2.612 $Y2=1.52
r116 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.87
+ $X2=2.555 $Y2=1.87
r117 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r119 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=2.555 $Y2=1.87
r120 26 27 1.37376 $w=1.4e-07 $l=1.11e-06 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=1.3 $Y2=1.87
r121 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r122 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r123 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r124 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r125 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r126 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r127 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.22 $Y=1.245
+ $X2=3.22 $Y2=0.415
r128 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r129 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=3.22 $Y2=1.245
r130 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=2.805 $Y2=1.32
r131 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r132 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r133 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%A_724_21# 1 2 9 13 17 20 22 25 29 31 32 35
+ 37 42 43 45 51
r95 43 52 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=5.875 $Y=1.16
+ $X2=5.875 $Y2=1.325
r96 43 51 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=5.875 $Y=1.16
+ $X2=5.875 $Y2=0.995
r97 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.16 $X2=5.84 $Y2=1.16
r98 40 42 13.5052 $w=3.18e-07 $l=3.75e-07 $layer=LI1_cond $X=5.765 $Y=1.535
+ $X2=5.765 $Y2=1.16
r99 39 42 12.0646 $w=3.18e-07 $l=3.35e-07 $layer=LI1_cond $X=5.765 $Y=0.825
+ $X2=5.765 $Y2=1.16
r100 38 45 3.19459 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.94 $Y=1.7
+ $X2=4.845 $Y2=1.7
r101 37 40 6.81859 $w=3.3e-07 $l=2.31571e-07 $layer=LI1_cond $X=5.605 $Y=1.7
+ $X2=5.765 $Y2=1.535
r102 37 38 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=5.605 $Y=1.7
+ $X2=4.94 $Y2=1.7
r103 33 45 3.38787 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=1.865
+ $X2=4.845 $Y2=1.7
r104 33 35 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=4.845 $Y=1.865
+ $X2=4.845 $Y2=2.27
r105 31 39 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=5.605 $Y=0.74
+ $X2=5.765 $Y2=0.825
r106 31 32 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=5.605 $Y=0.74
+ $X2=4.59 $Y2=0.74
r107 27 32 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.415 $Y=0.655
+ $X2=4.59 $Y2=0.74
r108 27 29 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.415 $Y=0.655
+ $X2=4.415 $Y2=0.4
r109 25 46 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.695 $Y2=1.7
r110 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r111 22 45 3.19459 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.75 $Y=1.7
+ $X2=4.845 $Y2=1.7
r112 22 24 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.75 $Y=1.7
+ $X2=3.925 $Y2=1.7
r113 20 52 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.97 $Y=1.985
+ $X2=5.97 $Y2=1.325
r114 17 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.97 $Y=0.56
+ $X2=5.97 $Y2=0.995
r115 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=1.7
r116 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=2.275
r117 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=1.7
r118 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=0.445
r119 2 45 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.845 $Y2=1.755
r120 2 35 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.845 $Y2=2.27
r121 1 29 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.3
+ $Y=0.235 $X2=4.425 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%A_561_413# 1 2 9 13 15 16 17 21 26 28 29 31
c86 31 0 1.05716e-19 $X=4.145 $Y=1.16
c87 29 0 1.65126e-19 $X=3.65 $Y=1.175
r88 34 35 6.98473 $w=2.62e-07 $l=1.5e-07 $layer=LI1_cond $X=3.415 $Y=1.175
+ $X2=3.565 $Y2=1.175
r89 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=1.16 $X2=4.145 $Y2=1.16
r90 29 35 3.68445 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.175 $X2=3.565
+ $Y2=1.175
r91 29 31 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=3.65 $Y=1.175
+ $X2=4.145 $Y2=1.175
r92 27 35 3.26844 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.175
r93 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=2.255
r94 26 34 3.26844 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.415 $Y=1.025
+ $X2=3.415 $Y2=1.175
r95 25 26 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=1.025
r96 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.565 $Y2=2.255
r97 21 23 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.065 $Y2=2.34
r98 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r99 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.005 $Y2=0.45
r100 15 32 92.2021 $w=2.7e-07 $l=4.15e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.145 $Y2=1.16
r101 15 16 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.635 $Y2=1.16
r102 11 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.635 $Y=1.295
+ $X2=4.635 $Y2=1.16
r103 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.635 $Y=1.295
+ $X2=4.635 $Y2=1.985
r104 7 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.635 $Y=1.025
+ $X2=4.635 $Y2=1.16
r105 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.635 $Y=1.025
+ $X2=4.635 $Y2=0.56
r106 2 23 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=3.065 $Y2=2.34
r107 1 19 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3.005 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%RESET_B 3 6 8 9 13 15 22
c37 13 0 1.05716e-19 $X=5.065 $Y=1.16
r38 14 22 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.065 $Y=1.16
+ $X2=5.315 $Y2=1.16
r39 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.065 $Y=1.16
+ $X2=5.065 $Y2=1.325
r40 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.065 $Y=1.16
+ $X2=5.065 $Y2=0.995
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.065
+ $Y=1.16 $X2=5.065 $Y2=1.16
r42 9 22 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=5.335 $Y=1.16 $X2=5.315
+ $Y2=1.16
r43 8 14 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.875 $Y=1.16
+ $X2=5.065 $Y2=1.16
r44 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.055 $Y=1.985
+ $X2=5.055 $Y2=1.325
r45 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.055 $Y=0.56
+ $X2=5.055 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%VPWR 1 2 3 4 5 18 22 26 28 32 34 36 41 46 61
+ 62 65 68 71 74 79 82
r97 81 82 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=2.47
+ $X2=5.925 $Y2=2.47
r98 77 81 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=5.75 $Y=2.47 $X2=5.76
+ $Y2=2.47
r99 77 79 19.0914 $w=6.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.75 $Y=2.47
+ $X2=5.11 $Y2=2.47
r100 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r102 72 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r105 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r106 62 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r107 61 82 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=5.925 $Y2=2.72
r108 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r109 58 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 58 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r111 57 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.11 $Y2=2.72
r112 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r113 55 74 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.58 $Y=2.72 $X2=4.44
+ $Y2=2.72
r114 55 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.58 $Y=2.72
+ $X2=4.83 $Y2=2.72
r115 53 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r116 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r117 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 50 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 49 52 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r120 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r121 47 68 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r122 47 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r123 46 71 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=3.965 $Y2=2.72
r124 46 52 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=3.45 $Y2=2.72
r125 45 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 45 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r128 42 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r129 42 44 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r130 41 68 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r131 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r132 36 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r133 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r134 34 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 34 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r136 30 74 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=2.635
+ $X2=4.44 $Y2=2.72
r137 30 32 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.44 $Y=2.635
+ $X2=4.44 $Y2=2.34
r138 29 71 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=3.965 $Y2=2.72
r139 28 74 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.3 $Y=2.72 $X2=4.44
+ $Y2=2.72
r140 28 29 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.3 $Y=2.72
+ $X2=4.11 $Y2=2.72
r141 24 71 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=2.635
+ $X2=3.965 $Y2=2.72
r142 24 26 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.965 $Y=2.635
+ $X2=3.965 $Y2=2.3
r143 20 68 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r144 20 22 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r145 16 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r146 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r147 5 81 300 $w=1.7e-07 $l=1.1268e-06 $layer=licon1_PDIFF $count=2 $X=5.13
+ $Y=1.485 $X2=5.76 $Y2=2.34
r148 4 32 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.485 $X2=4.425 $Y2=2.34
r149 3 26 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=2.065 $X2=3.905 $Y2=2.3
r150 2 22 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r151 1 18 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%Q 1 2 7 8 9 10 11 12
r10 11 12 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=6.225 $Y=1.835
+ $X2=6.225 $Y2=2.21
r11 10 11 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=6.225 $Y=1.53
+ $X2=6.225 $Y2=1.835
r12 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=6.225 $Y=1.19
+ $X2=6.225 $Y2=1.53
r13 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=6.225 $Y=0.85
+ $X2=6.225 $Y2=1.19
r14 7 8 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=6.225 $Y=0.51
+ $X2=6.225 $Y2=0.85
r15 2 11 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=1.835
r16 1 7 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_1%VGND 1 2 3 4 15 19 23 25 27 32 37 52 53 56
+ 59 62 67 73
c97 53 0 2.71124e-20 $X=6.21 $Y=0
c98 2 0 7.13094e-20 $X=1.905 $Y=0.235
r99 72 73 10.0659 $w=5.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.755 $Y=0.2
+ $X2=5.925 $Y2=0.2
r100 69 72 0.104919 $w=5.68e-07 $l=5e-09 $layer=LI1_cond $X=5.75 $Y=0.2
+ $X2=5.755 $Y2=0.2
r101 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r102 66 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r103 65 69 9.65256 $w=5.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=0.2
+ $X2=5.75 $Y2=0.2
r104 65 67 10.5905 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.29 $Y=0.2
+ $X2=5.095 $Y2=0.2
r105 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r106 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r107 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r108 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r109 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r110 52 73 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=5.925 $Y2=0
r111 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r112 49 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r113 49 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r114 48 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=5.095 $Y2=0
r115 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r116 46 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.905
+ $Y2=0
r117 46 48 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.83
+ $Y2=0
r118 44 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r119 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r120 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r121 41 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r122 40 43 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r123 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r124 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r125 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r126 37 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.905
+ $Y2=0
r127 37 43 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.45
+ $Y2=0
r128 36 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r129 36 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r130 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r131 33 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r132 33 35 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r133 32 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r134 32 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r135 27 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r136 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r137 25 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r138 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r139 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r140 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0.445
r141 17 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r142 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r143 13 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r144 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r145 4 72 91 $w=1.7e-07 $l=6.93722e-07 $layer=licon1_NDIFF $count=2 $X=5.13
+ $Y=0.235 $X2=5.755 $Y2=0.38
r146 3 23 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.235 $X2=3.905 $Y2=0.445
r147 2 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r148 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__nor4bb_2.spice
* Created: Thu Aug 27 14:33:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor4bb_2.pex.spice"
.subckt sky130_fd_sc_hd__nor4bb_2  VNB VPB D_N C_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_D_N_M1003_g N_A_27_410#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_201_93#_M1016_d N_C_N_M1016_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_201_93#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.221 AS=0.08775 PD=1.98 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75000.3
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_201_93#_M1005_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1005_d N_A_27_410#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_27_410#_M1007_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.65 AD=0.182
+ AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.5
+ A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_B_M1017_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1017_d N_A_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_M1014_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.08775 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 N_VPWR_M1015_d N_D_N_M1015_g N_A_27_410#_M1015_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.122612 AS=0.1092 PD=1.32 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_201_93#_M1018_d N_C_N_M1018_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.122612 PD=1.36 PS=1.32 NRD=0 NRS=111.128 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_418_297#_M1001_d N_A_201_93#_M1001_g N_A_336_297#_M1001_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1019 N_A_418_297#_M1001_d N_A_201_93#_M1019_g N_A_336_297#_M1019_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001 A=0.15 P=2.3 MULT=1
MM1008 N_A_336_297#_M1019_s N_A_27_410#_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_A_336_297#_M1011_d N_A_27_410#_M1011_g N_Y_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_776_297#_M1009_d N_B_M1009_g N_A_418_297#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1013 N_A_776_297#_M1013_d N_B_M1013_g N_A_418_297#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_776_297#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1004_d N_A_M1012_g N_A_776_297#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__nor4bb_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a21oi_4.spice.pex
* Created: Thu Aug 27 14:01:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 34 35 43
+ 45
c73 22 0 5.96372e-20 $X=1.765 $Y=0.995
c74 6 0 2.99299e-20 $X=0.475 $Y=1.985
r75 44 45 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.765 $Y2=1.16
r76 42 44 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.265 $Y=1.16
+ $X2=1.335 $Y2=1.16
r77 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.265
+ $Y=1.16 $X2=1.265 $Y2=1.16
r78 40 42 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=0.905 $Y=1.16
+ $X2=1.265 $Y2=1.16
r79 39 40 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.905 $Y2=1.16
r80 35 43 3.33602 $w=3.78e-07 $l=1.1e-07 $layer=LI1_cond $X=1.155 $Y=1.225
+ $X2=1.265 $Y2=1.225
r81 34 35 22.8972 $w=3.78e-07 $l=7.55e-07 $layer=LI1_cond $X=0.4 $Y=1.225
+ $X2=1.155 $Y2=1.225
r82 32 39 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.475 $Y2=1.16
r83 31 34 4.3816 $w=4.18e-07 $l=1.55e-07 $layer=LI1_cond $X=0.245 $Y=1.205
+ $X2=0.4 $Y2=1.205
r84 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r85 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.325
+ $X2=1.765 $Y2=1.16
r86 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.325
+ $X2=1.765 $Y2=1.985
r87 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=0.995
+ $X2=1.765 $Y2=1.16
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.765 $Y=0.995
+ $X2=1.765 $Y2=0.56
r89 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.16
r90 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.985
r91 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=1.16
r92 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=0.56
r93 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r95 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r97 4 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.16
r98 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.985
r99 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%A2 3 7 8 10 13 15 17 20 22 24 27 31 32 35 36
+ 37 38 41 54 55
c128 35 0 3.12905e-20 $X=2.395 $Y=1.592
c129 32 0 3.88689e-19 $X=2.215 $Y=1.16
c130 8 0 6.41563e-20 $X=4.385 $Y=0.995
r131 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.305
+ $Y=1.16 $X2=5.305 $Y2=1.16
r132 52 54 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.245 $Y=1.16
+ $X2=5.305 $Y2=1.16
r133 50 52 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=4.965 $Y=1.16
+ $X2=5.245 $Y2=1.16
r134 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.965
+ $Y=1.16 $X2=4.965 $Y2=1.16
r135 48 50 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.815 $Y=1.16
+ $X2=4.965 $Y2=1.16
r136 47 51 6.45503 $w=6.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.625 $Y=1.39
+ $X2=4.965 $Y2=1.39
r137 46 48 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.625 $Y=1.16
+ $X2=4.815 $Y2=1.16
r138 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.625
+ $Y=1.16 $X2=4.625 $Y2=1.16
r139 43 46 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.385 $Y=1.16
+ $X2=4.625 $Y2=1.16
r140 38 55 0.189854 $w=6.28e-07 $l=1e-08 $layer=LI1_cond $X=5.295 $Y=1.39
+ $X2=5.305 $Y2=1.39
r141 38 51 6.26517 $w=6.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.295 $Y=1.39
+ $X2=4.965 $Y2=1.39
r142 36 47 1.61376 $w=6.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=1.39
+ $X2=4.625 $Y2=1.39
r143 36 37 11.207 $w=6.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.54 $Y=1.39
+ $X2=4.225 $Y2=1.39
r144 35 37 93.732 $w=2.23e-07 $l=1.83e-06 $layer=LI1_cond $X=2.395 $Y=1.592
+ $X2=4.225 $Y2=1.592
r145 32 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.215 $Y2=1.325
r146 32 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.215 $Y2=0.995
r147 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.215
+ $Y=1.16 $X2=2.215 $Y2=1.16
r148 29 35 7.21695 $w=2.25e-07 $l=2.22047e-07 $layer=LI1_cond $X=2.222 $Y=1.48
+ $X2=2.395 $Y2=1.592
r149 29 31 10.6893 $w=3.43e-07 $l=3.2e-07 $layer=LI1_cond $X=2.222 $Y=1.48
+ $X2=2.222 $Y2=1.16
r150 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.325
+ $X2=5.245 $Y2=1.16
r151 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.245 $Y=1.325
+ $X2=5.245 $Y2=1.985
r152 22 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=0.995
+ $X2=5.245 $Y2=1.16
r153 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.245 $Y=0.995
+ $X2=5.245 $Y2=0.56
r154 18 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.325
+ $X2=4.815 $Y2=1.16
r155 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.815 $Y=1.325
+ $X2=4.815 $Y2=1.985
r156 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=1.16
r157 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=0.56
r158 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=1.325
+ $X2=4.385 $Y2=1.16
r159 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.385 $Y=1.325
+ $X2=4.385 $Y2=1.985
r160 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=1.16
r161 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=0.56
r162 7 41 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.235 $Y=0.56
+ $X2=2.235 $Y2=0.995
r163 3 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.225 $Y=1.985
+ $X2=2.225 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29
r72 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.815
+ $Y=1.16 $X2=3.815 $Y2=1.16
r73 39 43 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.475 $Y=1.187
+ $X2=3.815 $Y2=1.187
r74 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.475
+ $Y=1.16 $X2=3.475 $Y2=1.16
r75 35 39 31.9862 $w=2.43e-07 $l=6.8e-07 $layer=LI1_cond $X=2.795 $Y=1.187
+ $X2=3.475 $Y2=1.187
r76 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.16 $X2=2.795 $Y2=1.16
r77 29 43 4.70385 $w=2.43e-07 $l=1e-07 $layer=LI1_cond $X=3.915 $Y=1.187
+ $X2=3.815 $Y2=1.187
r78 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.955 $Y=1.295
+ $X2=3.955 $Y2=1.985
r79 22 25 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=3.955 $Y=1.142
+ $X2=3.955 $Y2=1.295
r80 22 42 27.535 $w=3.05e-07 $l=1.4e-07 $layer=POLY_cond $X=3.955 $Y=1.142
+ $X2=3.815 $Y2=1.142
r81 22 24 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.955 $Y=0.99
+ $X2=3.955 $Y2=0.56
r82 18 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.525 $Y=1.295
+ $X2=3.525 $Y2=1.985
r83 15 42 57.0367 $w=3.05e-07 $l=2.9e-07 $layer=POLY_cond $X=3.525 $Y=1.142
+ $X2=3.815 $Y2=1.142
r84 15 18 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=3.525 $Y=1.142
+ $X2=3.525 $Y2=1.295
r85 15 38 9.83392 $w=3.05e-07 $l=5e-08 $layer=POLY_cond $X=3.525 $Y=1.142
+ $X2=3.475 $Y2=1.142
r86 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.525 $Y=0.99
+ $X2=3.525 $Y2=0.56
r87 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.095 $Y=1.295
+ $X2=3.095 $Y2=1.985
r88 8 38 74.7378 $w=3.05e-07 $l=3.8e-07 $layer=POLY_cond $X=3.095 $Y=1.142
+ $X2=3.475 $Y2=1.142
r89 8 11 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=3.095 $Y=1.142
+ $X2=3.095 $Y2=1.295
r90 8 34 59.0035 $w=3.05e-07 $l=3e-07 $layer=POLY_cond $X=3.095 $Y=1.142
+ $X2=2.795 $Y2=1.142
r91 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.095 $Y=0.99
+ $X2=3.095 $Y2=0.56
r92 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.665 $Y2=1.985
r93 1 34 25.5682 $w=3.05e-07 $l=1.3e-07 $layer=POLY_cond $X=2.665 $Y=1.142
+ $X2=2.795 $Y2=1.142
r94 1 4 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=2.665 $Y=1.142
+ $X2=2.665 $Y2=1.295
r95 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.665 $Y=0.99
+ $X2=2.665 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%A_28_297# 1 2 3 4 5 6 7 22 24 26 28 29 32 34
+ 38 40 44 46 48 50 59 61 62
c83 29 0 2.24772e-19 $X=2.115 $Y=1.99
c84 28 0 1.93847e-19 $X=2.785 $Y=1.99
r85 55 57 34.3608 $w=3.16e-07 $l=8.9e-07 $layer=LI1_cond $X=1.12 $Y=2.205
+ $X2=2.01 $Y2=2.205
r86 48 64 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=5.495 $Y=2.105
+ $X2=5.495 $Y2=1.99
r87 48 50 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=5.495 $Y=2.105
+ $X2=5.495 $Y2=2.3
r88 47 62 4.19361 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=4.685 $Y=1.99 $X2=4.595
+ $Y2=1.99
r89 46 64 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=1.99
+ $X2=5.495 $Y2=1.99
r90 46 47 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.365 $Y=1.99
+ $X2=4.685 $Y2=1.99
r91 42 62 2.23839 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=4.595 $Y=2.105
+ $X2=4.595 $Y2=1.99
r92 42 44 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=4.595 $Y=2.105
+ $X2=4.595 $Y2=2.3
r93 41 61 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.835 $Y=1.99
+ $X2=3.74 $Y2=1.99
r94 40 62 4.19361 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=4.505 $Y=1.99 $X2=4.595
+ $Y2=1.99
r95 40 41 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=4.505 $Y=1.99
+ $X2=3.835 $Y2=1.99
r96 36 61 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.74 $Y=2.105
+ $X2=3.74 $Y2=1.99
r97 36 38 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.74 $Y=2.105
+ $X2=3.74 $Y2=2.3
r98 35 59 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.975 $Y=1.99
+ $X2=2.88 $Y2=1.99
r99 34 61 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.645 $Y=1.99
+ $X2=3.74 $Y2=1.99
r100 34 35 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.645 $Y=1.99
+ $X2=2.975 $Y2=1.99
r101 30 59 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.88 $Y=2.105
+ $X2=2.88 $Y2=1.99
r102 30 32 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.88 $Y=2.105
+ $X2=2.88 $Y2=2.3
r103 29 57 4.97931 $w=3.16e-07 $l=2.62298e-07 $layer=LI1_cond $X=2.115 $Y=1.99
+ $X2=2.01 $Y2=2.205
r104 28 59 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.785 $Y=1.99
+ $X2=2.88 $Y2=1.99
r105 28 29 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.785 $Y=1.99
+ $X2=2.115 $Y2=1.99
r106 27 53 3.05549 $w=2.5e-07 $l=9.8e-08 $layer=LI1_cond $X=0.375 $Y=2.34
+ $X2=0.277 $Y2=2.34
r107 26 55 6.93673 $w=3.16e-07 $l=2.22486e-07 $layer=LI1_cond $X=0.955 $Y=2.34
+ $X2=1.12 $Y2=2.205
r108 26 27 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=0.955 $Y=2.34
+ $X2=0.375 $Y2=2.34
r109 22 53 3.89731 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=0.277 $Y=2.215
+ $X2=0.277 $Y2=2.34
r110 22 24 14.5035 $w=1.93e-07 $l=2.55e-07 $layer=LI1_cond $X=0.277 $Y=2.215
+ $X2=0.277 $Y2=1.96
r111 7 64 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=5.32
+ $Y=1.485 $X2=5.46 $Y2=1.96
r112 7 50 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=5.32
+ $Y=1.485 $X2=5.46 $Y2=2.3
r113 6 44 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.485 $X2=4.6 $Y2=2.3
r114 5 61 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.485 $X2=3.74 $Y2=1.96
r115 5 38 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.485 $X2=3.74 $Y2=2.3
r116 4 59 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=1.485 $X2=2.88 $Y2=1.96
r117 4 32 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=1.485 $X2=2.88 $Y2=2.3
r118 3 57 600 $w=1.7e-07 $l=8.95977e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.485 $X2=2.01 $Y2=2.3
r119 2 55 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=2.36
r120 1 53 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2.3
r121 1 24 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%Y 1 2 3 4 5 6 19 23 26 28 29 33 36 43 44 47
c75 33 0 6.41563e-20 $X=3.74 $Y=0.76
c76 29 0 3.98769e-19 $X=2.385 $Y=0.785
c77 28 0 1.1531e-19 $X=1.88 $Y=0.795
r78 44 47 2.80331 $w=4.5e-07 $l=1.4e-07 $layer=LI1_cond $X=1.74 $Y=1.81 $X2=1.6
+ $Y2=1.81
r79 44 47 1.32898 $w=4.48e-07 $l=5e-08 $layer=LI1_cond $X=1.55 $Y=1.81 $X2=1.6
+ $Y2=1.81
r80 44 49 22.8584 $w=4.48e-07 $l=8.6e-07 $layer=LI1_cond $X=1.55 $Y=1.81
+ $X2=0.69 $Y2=1.81
r81 31 33 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=2.88 $Y=0.785 $X2=3.74
+ $Y2=0.785
r82 29 43 5.8804 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=2.385 $Y=0.785
+ $X2=2.275 $Y2=0.785
r83 29 31 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=2.385 $Y=0.785
+ $X2=2.88 $Y2=0.785
r84 28 43 21.9045 $w=1.98e-07 $l=3.95e-07 $layer=LI1_cond $X=1.88 $Y=0.795
+ $X2=2.275 $Y2=0.795
r85 26 44 4.50532 $w=2.8e-07 $l=2.25e-07 $layer=LI1_cond $X=1.74 $Y=1.585
+ $X2=1.74 $Y2=1.81
r86 25 28 7.77084 $w=2.25e-07 $l=1.58745e-07 $layer=LI1_cond $X=1.74 $Y=0.755
+ $X2=1.88 $Y2=0.795
r87 25 41 10.3022 $w=2.25e-07 $l=1.9e-07 $layer=LI1_cond $X=1.74 $Y=0.755
+ $X2=1.55 $Y2=0.755
r88 25 26 28.3995 $w=2.78e-07 $l=6.9e-07 $layer=LI1_cond $X=1.74 $Y=0.895
+ $X2=1.74 $Y2=1.585
r89 21 41 1.72863 $w=1.9e-07 $l=1.4e-07 $layer=LI1_cond $X=1.55 $Y=0.615
+ $X2=1.55 $Y2=0.755
r90 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.55 $Y=0.615
+ $X2=1.55 $Y2=0.42
r91 20 36 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=0.69 $Y=0.74
+ $X2=0.69 $Y2=0.535
r92 19 41 4.78459 $w=2.5e-07 $l=1.02225e-07 $layer=LI1_cond $X=1.455 $Y=0.74
+ $X2=1.55 $Y2=0.755
r93 19 20 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=0.74
+ $X2=0.785 $Y2=0.74
r94 6 44 600 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=1.89
r95 5 49 600 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.85
r96 4 33 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.6
+ $Y=0.235 $X2=3.74 $Y2=0.76
r97 3 31 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=0.235 $X2=2.88 $Y2=0.76
r98 2 41 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.76
r99 2 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.42
r100 1 36 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
r103 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r104 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r105 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r107 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r109 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r110 51 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r111 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r112 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.45 $Y2=2.72
r113 48 50 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.99 $Y2=2.72
r114 47 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r115 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r116 42 46 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r117 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.45 $Y2=2.72
r118 40 46 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 38 47 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r120 38 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r121 36 56 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.865 $Y=2.72
+ $X2=4.83 $Y2=2.72
r122 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=2.72
+ $X2=5.03 $Y2=2.72
r123 35 59 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.195 $Y=2.72
+ $X2=5.75 $Y2=2.72
r124 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=2.72
+ $X2=5.03 $Y2=2.72
r125 33 53 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=3.91 $Y2=2.72
r126 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=4.17 $Y2=2.72
r127 32 56 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.335 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=2.72
+ $X2=4.17 $Y2=2.72
r129 30 50 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.145 $Y=2.72
+ $X2=2.99 $Y2=2.72
r130 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=2.72
+ $X2=3.31 $Y2=2.72
r131 29 53 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.91 $Y2=2.72
r132 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.31 $Y2=2.72
r133 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=2.635
+ $X2=5.03 $Y2=2.72
r134 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.03 $Y=2.635
+ $X2=5.03 $Y2=2.36
r135 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=2.635
+ $X2=4.17 $Y2=2.72
r136 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.17 $Y=2.635
+ $X2=4.17 $Y2=2.36
r137 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=2.635
+ $X2=3.31 $Y2=2.72
r138 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.31 $Y=2.635
+ $X2=3.31 $Y2=2.36
r139 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=2.635
+ $X2=2.45 $Y2=2.72
r140 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.45 $Y=2.635
+ $X2=2.45 $Y2=2.36
r141 4 27 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.485 $X2=5.03 $Y2=2.36
r142 3 23 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.485 $X2=4.17 $Y2=2.36
r143 2 19 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.17
+ $Y=1.485 $X2=3.31 $Y2=2.36
r144 1 15 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.485 $X2=2.45 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 49 62 63 69 72
c93 37 0 1.51849e-19 $X=4.505 $Y=0
r94 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r95 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r96 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r97 60 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r98 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r99 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r100 57 73 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=2.07
+ $Y2=0
r101 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r102 54 72 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.975
+ $Y2=0
r103 54 56 147.118 $w=1.68e-07 $l=2.255e-06 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=4.37 $Y2=0
r104 53 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r105 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r106 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r107 50 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r108 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.61 $Y2=0
r109 49 72 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.975
+ $Y2=0
r110 49 52 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=1.61 $Y2=0
r111 48 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r112 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r113 45 66 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r114 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r115 44 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r116 44 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.69 $Y2=0
r117 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r118 42 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r119 40 59 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.365 $Y=0 $X2=5.29
+ $Y2=0
r120 40 41 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=0 $X2=5.495
+ $Y2=0
r121 39 62 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.625 $Y=0
+ $X2=5.75 $Y2=0
r122 39 41 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.625 $Y=0 $X2=5.495
+ $Y2=0
r123 37 56 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=4.37 $Y2=0
r124 37 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.505 $Y=0 $X2=4.6
+ $Y2=0
r125 36 59 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=5.29 $Y2=0
r126 36 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.695 $Y=0 $X2=4.6
+ $Y2=0
r127 32 41 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=0.085
+ $X2=5.495 $Y2=0
r128 32 34 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.495 $Y=0.085
+ $X2=5.495 $Y2=0.38
r129 28 38 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.085
+ $X2=4.6 $Y2=0
r130 28 30 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=4.6 $Y=0.085
+ $X2=4.6 $Y2=0.4
r131 24 72 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0
r132 24 26 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0.36
r133 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r134 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r135 16 66 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r136 16 18 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r137 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.32
+ $Y=0.235 $X2=5.46 $Y2=0.38
r138 4 30 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.235 $X2=4.6 $Y2=0.4
r139 3 26 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=2.02 $Y2=0.36
r140 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.36
r141 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_4%A_462_47# 1 2 3 4 13 19 22 23 24 27
c45 1 0 1.87282e-19 $X=2.31 $Y=0.235
r46 25 27 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.03 $Y=0.735
+ $X2=5.03 $Y2=0.395
r47 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.865 $Y=0.82
+ $X2=5.03 $Y2=0.735
r48 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.865 $Y=0.82
+ $X2=4.335 $Y2=0.82
r49 20 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.205 $Y=0.735
+ $X2=4.335 $Y2=0.82
r50 20 22 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.205 $Y=0.735
+ $X2=4.205 $Y2=0.7
r51 19 30 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=4.205 $Y=0.505
+ $X2=4.205 $Y2=0.38
r52 19 22 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.205 $Y=0.505
+ $X2=4.205 $Y2=0.7
r53 15 18 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=2.45 $Y=0.38 $X2=3.31
+ $Y2=0.38
r54 13 30 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=4.075 $Y=0.38
+ $X2=4.205 $Y2=0.38
r55 13 18 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=4.075 $Y=0.38
+ $X2=3.31 $Y2=0.38
r56 4 27 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=4.89
+ $Y=0.235 $X2=5.03 $Y2=0.395
r57 3 30 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.235 $X2=4.17 $Y2=0.36
r58 3 22 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.235 $X2=4.17 $Y2=0.7
r59 2 18 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.31 $Y2=0.42
r60 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.235 $X2=2.45 $Y2=0.42
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__ebufn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.780000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.280000 1.425000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 1.445000 5.895000 1.725000 ;
        RECT 4.145000 0.615000 5.895000 0.855000 ;
        RECT 5.675000 0.855000 5.895000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.515000  0.085000 0.930000 0.595000 ;
        RECT 2.345000  0.085000 2.675000 0.485000 ;
        RECT 3.185000  0.085000 3.515000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.515000 1.845000 0.930000 2.635000 ;
        RECT 1.980000 2.275000 2.310000 2.635000 ;
        RECT 2.820000 2.275000 3.150000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.280000 0.345000 0.665000 ;
      RECT 0.085000 0.665000 0.320000 1.765000 ;
      RECT 0.085000 1.765000 0.345000 2.465000 ;
      RECT 1.100000 0.255000 1.725000 0.595000 ;
      RECT 1.100000 1.595000 1.725000 1.765000 ;
      RECT 1.100000 1.765000 1.355000 2.465000 ;
      RECT 1.450000 0.595000 1.725000 1.025000 ;
      RECT 1.450000 1.025000 3.810000 1.275000 ;
      RECT 1.450000 1.275000 1.725000 1.595000 ;
      RECT 1.565000 1.935000 5.895000 2.105000 ;
      RECT 1.565000 2.105000 1.810000 2.465000 ;
      RECT 1.895000 0.255000 2.175000 0.655000 ;
      RECT 1.895000 0.655000 3.975000 0.855000 ;
      RECT 1.895000 1.895000 5.895000 1.935000 ;
      RECT 2.480000 2.105000 2.650000 2.465000 ;
      RECT 2.845000 0.275000 3.015000 0.655000 ;
      RECT 3.320000 2.105000 5.895000 2.465000 ;
      RECT 3.685000 0.255000 5.735000 0.445000 ;
      RECT 3.685000 0.445000 3.975000 0.655000 ;
      RECT 3.980000 1.025000 5.505000 1.275000 ;
    LAYER mcon ;
      RECT 0.150000 1.105000 0.320000 1.275000 ;
      RECT 4.310000 1.105000 4.480000 1.275000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 4.540000 1.260000 ;
      RECT 0.085000 1.260000 0.380000 1.305000 ;
      RECT 4.250000 1.075000 4.540000 1.120000 ;
      RECT 4.250000 1.260000 4.540000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_4
END LIBRARY

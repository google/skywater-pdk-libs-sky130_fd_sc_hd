* File: sky130_fd_sc_hd__lpflow_isobufsrc_8.pxi.spice
* Created: Thu Aug 27 14:25:58 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A N_A_M1010_g N_A_c_131_n N_A_M1023_g
+ N_A_M1029_g N_A_c_132_n N_A_M1025_g A N_A_c_134_n A
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A_123_297# N_A_123_297#_M1023_d
+ N_A_123_297#_M1010_d N_A_123_297#_c_174_n N_A_123_297#_M1002_g
+ N_A_123_297#_M1000_g N_A_123_297#_c_175_n N_A_123_297#_M1003_g
+ N_A_123_297#_M1001_g N_A_123_297#_c_176_n N_A_123_297#_M1007_g
+ N_A_123_297#_M1014_g N_A_123_297#_c_177_n N_A_123_297#_M1008_g
+ N_A_123_297#_M1022_g N_A_123_297#_c_178_n N_A_123_297#_M1013_g
+ N_A_123_297#_M1024_g N_A_123_297#_c_179_n N_A_123_297#_M1028_g
+ N_A_123_297#_M1026_g N_A_123_297#_c_180_n N_A_123_297#_M1032_g
+ N_A_123_297#_M1027_g N_A_123_297#_c_181_n N_A_123_297#_M1035_g
+ N_A_123_297#_M1033_g N_A_123_297#_c_192_n N_A_123_297#_c_199_n
+ N_A_123_297#_c_201_n N_A_123_297#_c_182_n N_A_123_297#_c_193_n
+ N_A_123_297#_c_209_n N_A_123_297#_c_183_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A_123_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%SLEEP N_SLEEP_c_350_n N_SLEEP_M1005_g
+ N_SLEEP_M1004_g N_SLEEP_c_351_n N_SLEEP_M1006_g N_SLEEP_M1011_g
+ N_SLEEP_c_352_n N_SLEEP_M1009_g N_SLEEP_M1012_g N_SLEEP_c_353_n
+ N_SLEEP_M1015_g N_SLEEP_M1017_g N_SLEEP_c_354_n N_SLEEP_M1016_g
+ N_SLEEP_M1020_g N_SLEEP_c_355_n N_SLEEP_M1018_g N_SLEEP_M1030_g
+ N_SLEEP_c_356_n N_SLEEP_M1019_g N_SLEEP_M1031_g N_SLEEP_c_357_n
+ N_SLEEP_M1021_g N_SLEEP_M1034_g SLEEP N_SLEEP_c_370_n N_SLEEP_c_358_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%SLEEP
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%VPWR N_VPWR_M1010_s N_VPWR_M1029_s
+ N_VPWR_M1000_s N_VPWR_M1014_s N_VPWR_M1024_s N_VPWR_M1027_s N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n
+ N_VPWR_c_505_n N_VPWR_c_506_n VPWR N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_493_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A_321_297# N_A_321_297#_M1000_d
+ N_A_321_297#_M1001_d N_A_321_297#_M1022_d N_A_321_297#_M1026_d
+ N_A_321_297#_M1033_d N_A_321_297#_M1011_s N_A_321_297#_M1017_s
+ N_A_321_297#_M1030_s N_A_321_297#_M1034_s N_A_321_297#_c_617_n
+ N_A_321_297#_c_618_n N_A_321_297#_c_619_n N_A_321_297#_c_675_n
+ N_A_321_297#_c_620_n N_A_321_297#_c_679_n N_A_321_297#_c_621_n
+ N_A_321_297#_c_683_n N_A_321_297#_c_622_n N_A_321_297#_c_623_n
+ N_A_321_297#_c_687_n N_A_321_297#_c_652_n N_A_321_297#_c_710_p
+ N_A_321_297#_c_654_n N_A_321_297#_c_714_p N_A_321_297#_c_656_n
+ N_A_321_297#_c_717_p N_A_321_297#_c_658_n N_A_321_297#_c_720_p
+ N_A_321_297#_c_624_n N_A_321_297#_c_625_n N_A_321_297#_c_626_n
+ N_A_321_297#_c_697_n N_A_321_297#_c_699_n N_A_321_297#_c_701_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A_321_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%X N_X_M1002_d N_X_M1007_d N_X_M1013_d
+ N_X_M1032_d N_X_M1005_s N_X_M1009_s N_X_M1016_s N_X_M1019_s N_X_M1004_d
+ N_X_M1012_d N_X_M1020_d N_X_M1031_d N_X_c_744_n N_X_c_721_n N_X_c_722_n
+ N_X_c_755_n N_X_c_723_n N_X_c_763_n N_X_c_724_n N_X_c_771_n N_X_c_725_n
+ N_X_c_776_n N_X_c_868_n N_X_c_737_n N_X_c_738_n N_X_c_726_n N_X_c_806_n
+ N_X_c_872_n N_X_c_739_n N_X_c_727_n N_X_c_818_n N_X_c_875_n N_X_c_740_n
+ N_X_c_728_n N_X_c_830_n N_X_c_878_n N_X_c_729_n N_X_c_730_n N_X_c_731_n
+ N_X_c_732_n N_X_c_733_n N_X_c_741_n N_X_c_734_n N_X_c_742_n N_X_c_735_n X
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%X
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%VGND N_VGND_M1023_s N_VGND_M1025_s
+ N_VGND_M1003_s N_VGND_M1008_s N_VGND_M1028_s N_VGND_M1035_s N_VGND_M1006_d
+ N_VGND_M1015_d N_VGND_M1018_d N_VGND_M1021_d N_VGND_c_945_n N_VGND_c_946_n
+ N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n
+ N_VGND_c_952_n N_VGND_c_953_n N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n
+ N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n
+ N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n
+ N_VGND_c_967_n N_VGND_c_968_n N_VGND_c_969_n VGND N_VGND_c_970_n
+ N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n N_VGND_c_975_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%VGND
cc_1 VNB N_A_c_131_n 0.0192657f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.995
cc_2 VNB N_A_c_132_n 0.0182175f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.995
cc_3 VNB A 0.0507065f $X=-0.19 $Y=-0.24 $X2=0.185 $Y2=1.105
cc_4 VNB N_A_c_134_n 0.0755148f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=1.16
cc_5 VNB N_A_123_297#_c_174_n 0.0185904f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.56
cc_6 VNB N_A_123_297#_c_175_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.56
cc_7 VNB N_A_123_297#_c_176_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_8 VNB N_A_123_297#_c_177_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_123_297#_c_178_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_123_297#_c_179_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_123_297#_c_180_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_123_297#_c_181_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_123_297#_c_182_n 0.0237489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_123_297#_c_183_n 0.128815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_SLEEP_c_350_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.325
cc_16 VNB N_SLEEP_c_351_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.325
cc_17 VNB N_SLEEP_c_352_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_SLEEP_c_353_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_19 VNB N_SLEEP_c_354_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.175
cc_20 VNB N_SLEEP_c_355_n 0.0157999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SLEEP_c_356_n 0.0157944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_SLEEP_c_357_n 0.019415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_SLEEP_c_358_n 0.131227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_493_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_721_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_722_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_723_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_724_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_725_n 0.00414888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_726_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_727_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_728_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_729_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_730_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_731_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_732_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_733_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_734_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_735_n 0.0109568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB X 0.0181545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_945_n 0.0127748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_946_n 0.0107395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_947_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_948_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_949_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_950_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_951_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_952_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_953_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_954_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_955_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_956_n 0.0100749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_957_n 0.0174928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_958_n 0.0143113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_959_n 0.00422832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_960_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_961_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_962_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_963_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_964_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_965_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_966_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_967_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_968_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_969_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_970_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_971_n 0.0166671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_972_n 0.00980307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_973_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_974_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_975_n 0.41623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VPB N_A_M1010_g 0.0250347f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.985
cc_73 VPB N_A_M1029_g 0.024514f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.985
cc_74 VPB N_A_c_134_n 0.0229749f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=1.16
cc_75 VPB N_A_123_297#_M1000_g 0.0252703f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=0.995
cc_76 VPB N_A_123_297#_M1001_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_123_297#_M1014_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_78 VPB N_A_123_297#_M1022_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_123_297#_M1024_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_123_297#_M1026_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_123_297#_M1027_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_123_297#_M1033_g 0.0185038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_123_297#_c_192_n 0.00313685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_123_297#_c_193_n 0.00120802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_123_297#_c_183_n 0.0224782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_SLEEP_M1004_g 0.018815f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.56
cc_87 VPB N_SLEEP_M1011_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=0.56
cc_88 VPB N_SLEEP_M1012_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_89 VPB N_SLEEP_M1017_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=1.16
cc_90 VPB N_SLEEP_M1020_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.175 $Y2=1.175
cc_91 VPB N_SLEEP_M1030_g 0.0181374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_SLEEP_M1031_g 0.0181277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_SLEEP_M1034_g 0.022286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_SLEEP_c_358_n 0.0223627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_494_n 0.0126236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_495_n 0.0428287f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_97 VPB N_VPWR_c_496_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.16
cc_98 VPB N_VPWR_c_497_n 0.0155448f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.175
cc_99 VPB N_VPWR_c_498_n 0.0196975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_499_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_500_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_501_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_502_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_503_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_504_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_505_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_506_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_507_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_508_n 0.0921061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_493_n 0.0596462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_510_n 0.00468329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_511_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_512_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_321_297#_c_617_n 0.00520781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_321_297#_c_618_n 0.00821221f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.175
cc_116 VPB N_A_321_297#_c_619_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.175
cc_117 VPB N_A_321_297#_c_620_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_321_297#_c_621_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_321_297#_c_622_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_321_297#_c_623_n 0.00407886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_321_297#_c_624_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_321_297#_c_625_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_321_297#_c_626_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_X_c_737_n 0.00234891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_X_c_738_n 0.0023869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_X_c_739_n 0.00234891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_X_c_740_n 0.00234891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_X_c_741_n 0.00202537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_X_c_742_n 0.00202537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB X 0.0189514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 N_A_c_132_n N_A_123_297#_c_174_n 0.00572906f $X=1.2 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_M1010_g N_A_123_297#_c_192_n 0.0028315f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1029_g N_A_123_297#_c_192_n 0.00215259f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_c_134_n N_A_123_297#_c_192_n 0.00202121f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_M1010_g N_A_123_297#_c_199_n 0.00951962f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1029_g N_A_123_297#_c_199_n 0.00951962f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_c_131_n N_A_123_297#_c_201_n 0.0105637f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_132_n N_A_123_297#_c_201_n 0.01254f $X=1.2 $Y=0.995 $X2=0 $Y2=0
cc_139 A N_A_123_297#_c_201_n 0.00490807f $X=0.185 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A_c_134_n N_A_123_297#_c_201_n 0.00910258f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_c_134_n N_A_123_297#_c_182_n 0.0126f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_M1010_g N_A_123_297#_c_193_n 0.00278727f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1029_g N_A_123_297#_c_193_n 0.00610341f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_c_134_n N_A_123_297#_c_193_n 0.00508115f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_145 A N_A_123_297#_c_209_n 0.0179768f $X=0.185 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A_c_134_n N_A_123_297#_c_209_n 0.0250762f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_134_n N_A_123_297#_c_183_n 0.00572906f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_M1010_g N_VPWR_c_495_n 0.00386041f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_149 A N_VPWR_c_495_n 0.0182999f $X=0.185 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A_c_134_n N_VPWR_c_495_n 0.00532863f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_M1010_g N_VPWR_c_496_n 0.00541359f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1029_g N_VPWR_c_496_n 0.00541359f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_M1029_g N_VPWR_c_497_n 0.00387648f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_c_134_n N_VPWR_c_497_n 0.0053981f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_M1010_g N_VPWR_c_493_n 0.0105165f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1029_g N_VPWR_c_493_n 0.0108276f $X=0.96 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_c_131_n N_VGND_c_945_n 0.00341559f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_158 A N_VGND_c_945_n 0.0607701f $X=0.185 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A_c_134_n N_VGND_c_945_n 0.00701224f $X=1.2 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_132_n N_VGND_c_946_n 0.00228475f $X=1.2 $Y=0.995 $X2=0 $Y2=0
cc_161 A N_VGND_c_958_n 0.0127617f $X=0.185 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A_c_131_n N_VGND_c_970_n 0.00541359f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_132_n N_VGND_c_970_n 0.00541359f $X=1.2 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_131_n N_VGND_c_975_n 0.010649f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_132_n N_VGND_c_975_n 0.0101559f $X=1.2 $Y=0.995 $X2=0 $Y2=0
cc_166 A N_VGND_c_975_n 0.00685509f $X=0.185 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A_123_297#_c_181_n N_SLEEP_c_350_n 0.0196453f $X=4.9 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_123_297#_M1033_g N_SLEEP_M1004_g 0.0196453f $X=4.9 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_123_297#_c_182_n N_SLEEP_c_370_n 0.0124677f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_170 N_A_123_297#_c_183_n N_SLEEP_c_370_n 2.30564e-19 $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_171 N_A_123_297#_c_182_n N_SLEEP_c_358_n 0.00185127f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_123_297#_c_183_n N_SLEEP_c_358_n 0.0196453f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_173 N_A_123_297#_c_192_n N_VPWR_c_495_n 0.0389948f $X=0.75 $Y=1.62 $X2=0
+ $Y2=0
cc_174 N_A_123_297#_c_199_n N_VPWR_c_496_n 0.0189039f $X=0.75 $Y=2.3 $X2=0 $Y2=0
cc_175 N_A_123_297#_M1000_g N_VPWR_c_497_n 0.00366507f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_123_297#_c_192_n N_VPWR_c_497_n 0.0390134f $X=0.75 $Y=1.62 $X2=0
+ $Y2=0
cc_177 N_A_123_297#_c_182_n N_VPWR_c_497_n 0.0144088f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_A_123_297#_c_209_n N_VPWR_c_497_n 0.006109f $X=0.95 $Y=1.175 $X2=0
+ $Y2=0
cc_179 N_A_123_297#_M1000_g N_VPWR_c_498_n 0.00585385f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_123_297#_M1000_g N_VPWR_c_499_n 0.00302074f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_123_297#_M1001_g N_VPWR_c_499_n 0.00157837f $X=2.38 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_123_297#_M1014_g N_VPWR_c_500_n 0.00157837f $X=2.8 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_123_297#_M1022_g N_VPWR_c_500_n 0.00157837f $X=3.22 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_123_297#_M1024_g N_VPWR_c_501_n 0.00157837f $X=3.64 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_123_297#_M1026_g N_VPWR_c_501_n 0.00157837f $X=4.06 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_123_297#_M1027_g N_VPWR_c_502_n 0.00157837f $X=4.48 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_123_297#_M1033_g N_VPWR_c_502_n 0.00302074f $X=4.9 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_123_297#_M1022_g N_VPWR_c_503_n 0.00585385f $X=3.22 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_123_297#_M1024_g N_VPWR_c_503_n 0.00585385f $X=3.64 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_123_297#_M1026_g N_VPWR_c_505_n 0.00585385f $X=4.06 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_123_297#_M1027_g N_VPWR_c_505_n 0.00585385f $X=4.48 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_123_297#_M1001_g N_VPWR_c_507_n 0.00585385f $X=2.38 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_123_297#_M1014_g N_VPWR_c_507_n 0.00585385f $X=2.8 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_123_297#_M1033_g N_VPWR_c_508_n 0.00585385f $X=4.9 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_123_297#_M1010_d N_VPWR_c_493_n 0.00215201f $X=0.615 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_A_123_297#_M1000_g N_VPWR_c_493_n 0.0117628f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_123_297#_M1001_g N_VPWR_c_493_n 0.0104367f $X=2.38 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_123_297#_M1014_g N_VPWR_c_493_n 0.0104367f $X=2.8 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_123_297#_M1022_g N_VPWR_c_493_n 0.0104367f $X=3.22 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_123_297#_M1024_g N_VPWR_c_493_n 0.0104367f $X=3.64 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_123_297#_M1026_g N_VPWR_c_493_n 0.0104367f $X=4.06 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_A_123_297#_M1027_g N_VPWR_c_493_n 0.0104367f $X=4.48 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_123_297#_M1033_g N_VPWR_c_493_n 0.010464f $X=4.9 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_123_297#_c_199_n N_VPWR_c_493_n 0.0122217f $X=0.75 $Y=2.3 $X2=0 $Y2=0
cc_205 N_A_123_297#_c_182_n N_A_321_297#_c_617_n 0.0274221f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_206 N_A_123_297#_M1000_g N_A_321_297#_c_619_n 0.0147299f $X=1.96 $Y=1.985
+ $X2=0 $Y2=0
cc_207 N_A_123_297#_M1001_g N_A_321_297#_c_619_n 0.0144778f $X=2.38 $Y=1.985
+ $X2=0 $Y2=0
cc_208 N_A_123_297#_c_182_n N_A_321_297#_c_619_n 0.0423927f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_209 N_A_123_297#_c_183_n N_A_321_297#_c_619_n 0.00212577f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_210 N_A_123_297#_M1014_g N_A_321_297#_c_620_n 0.0144778f $X=2.8 $Y=1.985
+ $X2=0 $Y2=0
cc_211 N_A_123_297#_M1022_g N_A_321_297#_c_620_n 0.0144778f $X=3.22 $Y=1.985
+ $X2=0 $Y2=0
cc_212 N_A_123_297#_c_182_n N_A_321_297#_c_620_n 0.042354f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_123_297#_c_183_n N_A_321_297#_c_620_n 0.00212577f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_214 N_A_123_297#_M1024_g N_A_321_297#_c_621_n 0.0144778f $X=3.64 $Y=1.985
+ $X2=0 $Y2=0
cc_215 N_A_123_297#_M1026_g N_A_321_297#_c_621_n 0.0144778f $X=4.06 $Y=1.985
+ $X2=0 $Y2=0
cc_216 N_A_123_297#_c_182_n N_A_321_297#_c_621_n 0.042354f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_217 N_A_123_297#_c_183_n N_A_321_297#_c_621_n 0.00212577f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_218 N_A_123_297#_M1027_g N_A_321_297#_c_622_n 0.0144232f $X=4.48 $Y=1.985
+ $X2=0 $Y2=0
cc_219 N_A_123_297#_M1033_g N_A_321_297#_c_622_n 0.0144195f $X=4.9 $Y=1.985
+ $X2=0 $Y2=0
cc_220 N_A_123_297#_c_182_n N_A_321_297#_c_622_n 0.0423927f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_221 N_A_123_297#_c_183_n N_A_321_297#_c_622_n 0.00212577f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_222 N_A_123_297#_c_182_n N_A_321_297#_c_623_n 0.00128541f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_223 N_A_123_297#_c_182_n N_A_321_297#_c_624_n 0.0204549f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_224 N_A_123_297#_c_183_n N_A_321_297#_c_624_n 0.00220041f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_225 N_A_123_297#_c_182_n N_A_321_297#_c_625_n 0.0204549f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_226 N_A_123_297#_c_183_n N_A_321_297#_c_625_n 0.00220041f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_227 N_A_123_297#_c_182_n N_A_321_297#_c_626_n 0.0204549f $X=4.79 $Y=1.16
+ $X2=0 $Y2=0
cc_228 N_A_123_297#_c_183_n N_A_321_297#_c_626_n 0.00220041f $X=4.9 $Y=1.16
+ $X2=0 $Y2=0
cc_229 N_A_123_297#_c_174_n N_X_c_744_n 0.00539651f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_123_297#_c_175_n N_X_c_744_n 0.00630972f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_123_297#_c_176_n N_X_c_744_n 5.22228e-19 $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_123_297#_c_175_n N_X_c_721_n 0.00870364f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_123_297#_c_176_n N_X_c_721_n 0.00870364f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_123_297#_c_182_n N_X_c_721_n 0.0362443f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_123_297#_c_183_n N_X_c_721_n 0.00222133f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_123_297#_c_174_n N_X_c_722_n 0.00262807f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_123_297#_c_175_n N_X_c_722_n 0.00113286f $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_123_297#_c_182_n N_X_c_722_n 0.0266272f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_123_297#_c_183_n N_X_c_722_n 0.00230339f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_123_297#_c_175_n N_X_c_755_n 5.22228e-19 $X=2.38 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_123_297#_c_176_n N_X_c_755_n 0.00630972f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_123_297#_c_177_n N_X_c_755_n 0.00630972f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_123_297#_c_178_n N_X_c_755_n 5.22228e-19 $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_123_297#_c_177_n N_X_c_723_n 0.00870364f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_123_297#_c_178_n N_X_c_723_n 0.00870364f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_123_297#_c_182_n N_X_c_723_n 0.0362443f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_123_297#_c_183_n N_X_c_723_n 0.00222133f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_123_297#_c_177_n N_X_c_763_n 5.22228e-19 $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_123_297#_c_178_n N_X_c_763_n 0.00630972f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_123_297#_c_179_n N_X_c_763_n 0.00630972f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_123_297#_c_180_n N_X_c_763_n 5.22228e-19 $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_123_297#_c_179_n N_X_c_724_n 0.00870364f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_123_297#_c_180_n N_X_c_724_n 0.00870364f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_123_297#_c_182_n N_X_c_724_n 0.0362443f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_123_297#_c_183_n N_X_c_724_n 0.00222133f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_123_297#_c_179_n N_X_c_771_n 5.22228e-19 $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A_123_297#_c_180_n N_X_c_771_n 0.00630972f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A_123_297#_c_181_n N_X_c_771_n 0.00630972f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_123_297#_c_181_n N_X_c_725_n 0.00865686f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_123_297#_c_182_n N_X_c_725_n 0.0101912f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_123_297#_c_181_n N_X_c_776_n 5.22228e-19 $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_123_297#_c_176_n N_X_c_729_n 0.00113286f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_123_297#_c_177_n N_X_c_729_n 0.00113286f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_123_297#_c_182_n N_X_c_729_n 0.0266272f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_123_297#_c_183_n N_X_c_729_n 0.00230339f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_123_297#_c_178_n N_X_c_730_n 0.00113286f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_123_297#_c_179_n N_X_c_730_n 0.00113286f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_123_297#_c_182_n N_X_c_730_n 0.0266272f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_123_297#_c_183_n N_X_c_730_n 0.00230339f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_123_297#_c_180_n N_X_c_731_n 0.00113286f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_123_297#_c_181_n N_X_c_731_n 0.00113286f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_123_297#_c_182_n N_X_c_731_n 0.0266272f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_123_297#_c_183_n N_X_c_731_n 0.00230339f $X=4.9 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_123_297#_c_192_n N_VGND_c_945_n 0.00262006f $X=0.75 $Y=1.62 $X2=0
+ $Y2=0
cc_275 N_A_123_297#_c_201_n N_VGND_c_945_n 0.0243665f $X=0.99 $Y=0.39 $X2=0
+ $Y2=0
cc_276 N_A_123_297#_c_174_n N_VGND_c_946_n 0.00228438f $X=1.96 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_123_297#_c_201_n N_VGND_c_946_n 0.0252338f $X=0.99 $Y=0.39 $X2=0
+ $Y2=0
cc_278 N_A_123_297#_c_182_n N_VGND_c_946_n 0.0435327f $X=4.79 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_A_123_297#_c_174_n N_VGND_c_947_n 0.00541359f $X=1.96 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_123_297#_c_175_n N_VGND_c_947_n 0.00423334f $X=2.38 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_123_297#_c_175_n N_VGND_c_948_n 0.00146448f $X=2.38 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_123_297#_c_176_n N_VGND_c_948_n 0.00146448f $X=2.8 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_123_297#_c_177_n N_VGND_c_949_n 0.00146448f $X=3.22 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_123_297#_c_178_n N_VGND_c_949_n 0.00146448f $X=3.64 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A_123_297#_c_179_n N_VGND_c_950_n 0.00146448f $X=4.06 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_123_297#_c_180_n N_VGND_c_950_n 0.00146448f $X=4.48 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_123_297#_c_181_n N_VGND_c_951_n 0.00146448f $X=4.9 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_123_297#_c_176_n N_VGND_c_960_n 0.00423334f $X=2.8 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_A_123_297#_c_177_n N_VGND_c_960_n 0.00423334f $X=3.22 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_123_297#_c_178_n N_VGND_c_962_n 0.00423334f $X=3.64 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_123_297#_c_179_n N_VGND_c_962_n 0.00423334f $X=4.06 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_123_297#_c_180_n N_VGND_c_964_n 0.00423334f $X=4.48 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_123_297#_c_181_n N_VGND_c_964_n 0.00423334f $X=4.9 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_123_297#_c_201_n N_VGND_c_970_n 0.0189039f $X=0.99 $Y=0.39 $X2=0
+ $Y2=0
cc_295 N_A_123_297#_M1023_d N_VGND_c_975_n 0.00215201f $X=0.855 $Y=0.235 $X2=0
+ $Y2=0
cc_296 N_A_123_297#_c_174_n N_VGND_c_975_n 0.0101559f $X=1.96 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_123_297#_c_175_n N_VGND_c_975_n 0.0057163f $X=2.38 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_123_297#_c_176_n N_VGND_c_975_n 0.0057163f $X=2.8 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_A_123_297#_c_177_n N_VGND_c_975_n 0.0057163f $X=3.22 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_A_123_297#_c_178_n N_VGND_c_975_n 0.0057163f $X=3.64 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_A_123_297#_c_179_n N_VGND_c_975_n 0.0057163f $X=4.06 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_123_297#_c_180_n N_VGND_c_975_n 0.0057163f $X=4.48 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_123_297#_c_181_n N_VGND_c_975_n 0.0057435f $X=4.9 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_123_297#_c_201_n N_VGND_c_975_n 0.0122217f $X=0.99 $Y=0.39 $X2=0
+ $Y2=0
cc_305 N_SLEEP_M1004_g N_VPWR_c_508_n 0.00357877f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_306 N_SLEEP_M1011_g N_VPWR_c_508_n 0.00357877f $X=5.74 $Y=1.985 $X2=0 $Y2=0
cc_307 N_SLEEP_M1012_g N_VPWR_c_508_n 0.00357877f $X=6.16 $Y=1.985 $X2=0 $Y2=0
cc_308 N_SLEEP_M1017_g N_VPWR_c_508_n 0.00357877f $X=6.58 $Y=1.985 $X2=0 $Y2=0
cc_309 N_SLEEP_M1020_g N_VPWR_c_508_n 0.00357877f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_310 N_SLEEP_M1030_g N_VPWR_c_508_n 0.00357877f $X=7.42 $Y=1.985 $X2=0 $Y2=0
cc_311 N_SLEEP_M1031_g N_VPWR_c_508_n 0.00357877f $X=7.84 $Y=1.985 $X2=0 $Y2=0
cc_312 N_SLEEP_M1034_g N_VPWR_c_508_n 0.00357877f $X=8.26 $Y=1.985 $X2=0 $Y2=0
cc_313 N_SLEEP_M1004_g N_VPWR_c_493_n 0.00525237f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_314 N_SLEEP_M1011_g N_VPWR_c_493_n 0.00522516f $X=5.74 $Y=1.985 $X2=0 $Y2=0
cc_315 N_SLEEP_M1012_g N_VPWR_c_493_n 0.00522516f $X=6.16 $Y=1.985 $X2=0 $Y2=0
cc_316 N_SLEEP_M1017_g N_VPWR_c_493_n 0.00522516f $X=6.58 $Y=1.985 $X2=0 $Y2=0
cc_317 N_SLEEP_M1020_g N_VPWR_c_493_n 0.00522516f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_318 N_SLEEP_M1030_g N_VPWR_c_493_n 0.00522516f $X=7.42 $Y=1.985 $X2=0 $Y2=0
cc_319 N_SLEEP_M1031_g N_VPWR_c_493_n 0.00522516f $X=7.84 $Y=1.985 $X2=0 $Y2=0
cc_320 N_SLEEP_M1034_g N_VPWR_c_493_n 0.00618885f $X=8.26 $Y=1.985 $X2=0 $Y2=0
cc_321 N_SLEEP_M1004_g N_A_321_297#_c_623_n 2.57315e-19 $X=5.32 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_SLEEP_M1004_g N_A_321_297#_c_652_n 0.0121747f $X=5.32 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_SLEEP_M1011_g N_A_321_297#_c_652_n 0.0121306f $X=5.74 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_SLEEP_M1012_g N_A_321_297#_c_654_n 0.0121747f $X=6.16 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_SLEEP_M1017_g N_A_321_297#_c_654_n 0.0121747f $X=6.58 $Y=1.985 $X2=0
+ $Y2=0
cc_326 N_SLEEP_M1020_g N_A_321_297#_c_656_n 0.0121747f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_327 N_SLEEP_M1030_g N_A_321_297#_c_656_n 0.0121747f $X=7.42 $Y=1.985 $X2=0
+ $Y2=0
cc_328 N_SLEEP_M1031_g N_A_321_297#_c_658_n 0.0121306f $X=7.84 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_SLEEP_M1034_g N_A_321_297#_c_658_n 0.0121747f $X=8.26 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_SLEEP_c_350_n N_X_c_771_n 5.22228e-19 $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_331 N_SLEEP_c_350_n N_X_c_725_n 0.00942689f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_332 N_SLEEP_c_370_n N_X_c_725_n 0.00651491f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_333 N_SLEEP_c_350_n N_X_c_776_n 0.00630972f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_334 N_SLEEP_c_351_n N_X_c_776_n 0.00630972f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_335 N_SLEEP_c_352_n N_X_c_776_n 5.22228e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_336 N_SLEEP_M1011_g N_X_c_737_n 0.0133089f $X=5.74 $Y=1.985 $X2=0 $Y2=0
cc_337 N_SLEEP_M1012_g N_X_c_737_n 0.0133439f $X=6.16 $Y=1.985 $X2=0 $Y2=0
cc_338 N_SLEEP_c_370_n N_X_c_737_n 0.0415099f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_339 N_SLEEP_c_358_n N_X_c_737_n 0.00214031f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_340 N_SLEEP_M1004_g N_X_c_738_n 5.90444e-19 $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_341 N_SLEEP_c_370_n N_X_c_738_n 0.0203891f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_342 N_SLEEP_c_358_n N_X_c_738_n 0.00222344f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_343 N_SLEEP_c_351_n N_X_c_726_n 0.00870364f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_344 N_SLEEP_c_352_n N_X_c_726_n 0.00870364f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_345 N_SLEEP_c_370_n N_X_c_726_n 0.036111f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_346 N_SLEEP_c_358_n N_X_c_726_n 0.00222133f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_347 N_SLEEP_c_351_n N_X_c_806_n 5.22228e-19 $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_348 N_SLEEP_c_352_n N_X_c_806_n 0.00630972f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_349 N_SLEEP_c_353_n N_X_c_806_n 0.00630972f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_350 N_SLEEP_c_354_n N_X_c_806_n 5.22228e-19 $X=7 $Y=0.995 $X2=0 $Y2=0
cc_351 N_SLEEP_M1017_g N_X_c_739_n 0.0133881f $X=6.58 $Y=1.985 $X2=0 $Y2=0
cc_352 N_SLEEP_M1020_g N_X_c_739_n 0.0133881f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_353 N_SLEEP_c_370_n N_X_c_739_n 0.0415099f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_354 N_SLEEP_c_358_n N_X_c_739_n 0.00214031f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_355 N_SLEEP_c_353_n N_X_c_727_n 0.00870364f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_356 N_SLEEP_c_354_n N_X_c_727_n 0.00870364f $X=7 $Y=0.995 $X2=0 $Y2=0
cc_357 N_SLEEP_c_370_n N_X_c_727_n 0.036111f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_358 N_SLEEP_c_358_n N_X_c_727_n 0.00222133f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_359 N_SLEEP_c_353_n N_X_c_818_n 5.22228e-19 $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_360 N_SLEEP_c_354_n N_X_c_818_n 0.00630972f $X=7 $Y=0.995 $X2=0 $Y2=0
cc_361 N_SLEEP_c_355_n N_X_c_818_n 0.00630972f $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_362 N_SLEEP_c_356_n N_X_c_818_n 5.22228e-19 $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_363 N_SLEEP_M1030_g N_X_c_740_n 0.0133881f $X=7.42 $Y=1.985 $X2=0 $Y2=0
cc_364 N_SLEEP_M1031_g N_X_c_740_n 0.0133881f $X=7.84 $Y=1.985 $X2=0 $Y2=0
cc_365 N_SLEEP_c_370_n N_X_c_740_n 0.0415099f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_366 N_SLEEP_c_358_n N_X_c_740_n 0.00214031f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_367 N_SLEEP_c_355_n N_X_c_728_n 0.00870364f $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_368 N_SLEEP_c_356_n N_X_c_728_n 0.00870364f $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_369 N_SLEEP_c_370_n N_X_c_728_n 0.036111f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_370 N_SLEEP_c_358_n N_X_c_728_n 0.00222133f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_371 N_SLEEP_c_355_n N_X_c_830_n 5.22228e-19 $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_372 N_SLEEP_c_356_n N_X_c_830_n 0.00630972f $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_373 N_SLEEP_c_357_n N_X_c_830_n 0.0109314f $X=8.26 $Y=0.995 $X2=0 $Y2=0
cc_374 N_SLEEP_c_350_n N_X_c_732_n 0.00113286f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_375 N_SLEEP_c_351_n N_X_c_732_n 0.00113286f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_376 N_SLEEP_c_370_n N_X_c_732_n 0.0265405f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_377 N_SLEEP_c_358_n N_X_c_732_n 0.00230339f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_378 N_SLEEP_c_352_n N_X_c_733_n 0.00113286f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_379 N_SLEEP_c_353_n N_X_c_733_n 0.00113286f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_380 N_SLEEP_c_370_n N_X_c_733_n 0.0265405f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_381 N_SLEEP_c_358_n N_X_c_733_n 0.00230339f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_382 N_SLEEP_c_370_n N_X_c_741_n 0.0203891f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_383 N_SLEEP_c_358_n N_X_c_741_n 0.00222344f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_384 N_SLEEP_c_354_n N_X_c_734_n 0.00113286f $X=7 $Y=0.995 $X2=0 $Y2=0
cc_385 N_SLEEP_c_355_n N_X_c_734_n 0.00113286f $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_386 N_SLEEP_c_370_n N_X_c_734_n 0.0265405f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_387 N_SLEEP_c_358_n N_X_c_734_n 0.00230339f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_388 N_SLEEP_c_370_n N_X_c_742_n 0.0203891f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_389 N_SLEEP_c_358_n N_X_c_742_n 0.00222344f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_390 N_SLEEP_c_356_n N_X_c_735_n 0.00113286f $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_391 N_SLEEP_c_357_n N_X_c_735_n 0.00946293f $X=8.26 $Y=0.995 $X2=0 $Y2=0
cc_392 N_SLEEP_c_370_n N_X_c_735_n 0.0100214f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_393 N_SLEEP_c_358_n N_X_c_735_n 0.00281533f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_394 N_SLEEP_c_356_n X 8.984e-19 $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_395 N_SLEEP_M1031_g X 0.00157422f $X=7.84 $Y=1.985 $X2=0 $Y2=0
cc_396 N_SLEEP_c_357_n X 0.00371247f $X=8.26 $Y=0.995 $X2=0 $Y2=0
cc_397 N_SLEEP_M1034_g X 0.0188787f $X=8.26 $Y=1.985 $X2=0 $Y2=0
cc_398 N_SLEEP_c_370_n X 0.0231659f $X=7.825 $Y=1.16 $X2=0 $Y2=0
cc_399 N_SLEEP_c_358_n X 0.0236342f $X=8.26 $Y=1.16 $X2=0 $Y2=0
cc_400 N_SLEEP_c_350_n N_VGND_c_951_n 0.00146448f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_401 N_SLEEP_c_351_n N_VGND_c_952_n 0.00146448f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_402 N_SLEEP_c_352_n N_VGND_c_952_n 0.00146448f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_403 N_SLEEP_c_353_n N_VGND_c_953_n 0.00146448f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_404 N_SLEEP_c_354_n N_VGND_c_953_n 0.00146448f $X=7 $Y=0.995 $X2=0 $Y2=0
cc_405 N_SLEEP_c_354_n N_VGND_c_954_n 0.00423334f $X=7 $Y=0.995 $X2=0 $Y2=0
cc_406 N_SLEEP_c_355_n N_VGND_c_954_n 0.00423334f $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_407 N_SLEEP_c_355_n N_VGND_c_955_n 0.00146448f $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_408 N_SLEEP_c_356_n N_VGND_c_955_n 0.00146448f $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_409 N_SLEEP_c_357_n N_VGND_c_957_n 0.00322276f $X=8.26 $Y=0.995 $X2=0 $Y2=0
cc_410 N_SLEEP_c_350_n N_VGND_c_966_n 0.00423334f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_411 N_SLEEP_c_351_n N_VGND_c_966_n 0.00423334f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_412 N_SLEEP_c_352_n N_VGND_c_968_n 0.00423334f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_413 N_SLEEP_c_353_n N_VGND_c_968_n 0.00423334f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_414 N_SLEEP_c_356_n N_VGND_c_971_n 0.00423334f $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_415 N_SLEEP_c_357_n N_VGND_c_971_n 0.00423225f $X=8.26 $Y=0.995 $X2=0 $Y2=0
cc_416 N_SLEEP_c_350_n N_VGND_c_975_n 0.0057435f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_417 N_SLEEP_c_351_n N_VGND_c_975_n 0.0057163f $X=5.74 $Y=0.995 $X2=0 $Y2=0
cc_418 N_SLEEP_c_352_n N_VGND_c_975_n 0.0057163f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_419 N_SLEEP_c_353_n N_VGND_c_975_n 0.0057163f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_420 N_SLEEP_c_354_n N_VGND_c_975_n 0.0057163f $X=7 $Y=0.995 $X2=0 $Y2=0
cc_421 N_SLEEP_c_355_n N_VGND_c_975_n 0.0057163f $X=7.42 $Y=0.995 $X2=0 $Y2=0
cc_422 N_SLEEP_c_356_n N_VGND_c_975_n 0.0057163f $X=7.84 $Y=0.995 $X2=0 $Y2=0
cc_423 N_SLEEP_c_357_n N_VGND_c_975_n 0.00667801f $X=8.26 $Y=0.995 $X2=0 $Y2=0
cc_424 N_VPWR_c_493_n N_A_321_297#_M1000_d 0.00260431f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_425 N_VPWR_c_493_n N_A_321_297#_M1001_d 0.00284632f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_493_n N_A_321_297#_M1022_d 0.00284632f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_493_n N_A_321_297#_M1026_d 0.00284632f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_493_n N_A_321_297#_M1033_d 0.00246446f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_493_n N_A_321_297#_M1011_s 0.00215203f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_493_n N_A_321_297#_M1017_s 0.00215203f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_493_n N_A_321_297#_M1030_s 0.00215203f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_493_n N_A_321_297#_M1034_s 0.00252233f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_497_n N_A_321_297#_c_617_n 0.0149366f $X=1.17 $Y=1.64 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_497_n N_A_321_297#_c_618_n 0.0533927f $X=1.17 $Y=1.64 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_498_n N_A_321_297#_c_618_n 0.0208267f $X=2.045 $Y=2.72 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_493_n N_A_321_297#_c_618_n 0.0122467f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_437 N_VPWR_M1000_s N_A_321_297#_c_619_n 0.00166915f $X=2.035 $Y=1.485 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_499_n N_A_321_297#_c_619_n 0.0128751f $X=2.17 $Y=2 $X2=0 $Y2=0
cc_439 N_VPWR_c_507_n N_A_321_297#_c_675_n 0.0142343f $X=2.885 $Y=2.72 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_493_n N_A_321_297#_c_675_n 0.00955092f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_M1014_s N_A_321_297#_c_620_n 0.00166915f $X=2.875 $Y=1.485 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_500_n N_A_321_297#_c_620_n 0.0128751f $X=3.01 $Y=2 $X2=0 $Y2=0
cc_443 N_VPWR_c_503_n N_A_321_297#_c_679_n 0.0142343f $X=3.725 $Y=2.72 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_493_n N_A_321_297#_c_679_n 0.00955092f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_M1024_s N_A_321_297#_c_621_n 0.00166915f $X=3.715 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_501_n N_A_321_297#_c_621_n 0.0128751f $X=3.85 $Y=2 $X2=0 $Y2=0
cc_447 N_VPWR_c_505_n N_A_321_297#_c_683_n 0.0142343f $X=4.565 $Y=2.72 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_493_n N_A_321_297#_c_683_n 0.00955092f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_449 N_VPWR_M1027_s N_A_321_297#_c_622_n 0.00166915f $X=4.555 $Y=1.485 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_502_n N_A_321_297#_c_622_n 0.0128751f $X=4.69 $Y=2 $X2=0 $Y2=0
cc_451 N_VPWR_c_508_n N_A_321_297#_c_687_n 0.0143053f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_493_n N_A_321_297#_c_687_n 0.00962794f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_508_n N_A_321_297#_c_652_n 0.0330174f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_493_n N_A_321_297#_c_652_n 0.0204627f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_508_n N_A_321_297#_c_654_n 0.0330174f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_493_n N_A_321_297#_c_654_n 0.0204627f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_508_n N_A_321_297#_c_656_n 0.0330174f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_493_n N_A_321_297#_c_656_n 0.0204627f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_508_n N_A_321_297#_c_658_n 0.0489601f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_493_n N_A_321_297#_c_658_n 0.0300907f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_508_n N_A_321_297#_c_697_n 0.0143053f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_493_n N_A_321_297#_c_697_n 0.00962794f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_508_n N_A_321_297#_c_699_n 0.0143053f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_493_n N_A_321_297#_c_699_n 0.00962794f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_508_n N_A_321_297#_c_701_n 0.0143053f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_493_n N_A_321_297#_c_701_n 0.00962794f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_493_n N_X_M1004_d 0.00216833f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_468 N_VPWR_c_493_n N_X_M1012_d 0.00216833f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_469 N_VPWR_c_493_n N_X_M1020_d 0.00216833f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_470 N_VPWR_c_493_n N_X_M1031_d 0.00216833f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_471 N_A_321_297#_c_652_n N_X_M1004_d 0.00312348f $X=5.825 $Y=2.38 $X2=0 $Y2=0
cc_472 N_A_321_297#_c_654_n N_X_M1012_d 0.00312348f $X=6.665 $Y=2.38 $X2=0 $Y2=0
cc_473 N_A_321_297#_c_656_n N_X_M1020_d 0.00312348f $X=7.505 $Y=2.38 $X2=0 $Y2=0
cc_474 N_A_321_297#_c_658_n N_X_M1031_d 0.00312348f $X=8.345 $Y=2.38 $X2=0 $Y2=0
cc_475 N_A_321_297#_c_623_n N_X_c_725_n 0.0088033f $X=5.11 $Y=1.665 $X2=0 $Y2=0
cc_476 N_A_321_297#_c_652_n N_X_c_868_n 0.0118865f $X=5.825 $Y=2.38 $X2=0 $Y2=0
cc_477 N_A_321_297#_M1011_s N_X_c_737_n 0.00165831f $X=5.815 $Y=1.485 $X2=0
+ $Y2=0
cc_478 N_A_321_297#_c_710_p N_X_c_737_n 0.0126919f $X=5.95 $Y=1.96 $X2=0 $Y2=0
cc_479 N_A_321_297#_c_623_n N_X_c_738_n 0.00271526f $X=5.11 $Y=1.665 $X2=0 $Y2=0
cc_480 N_A_321_297#_c_654_n N_X_c_872_n 0.0118865f $X=6.665 $Y=2.38 $X2=0 $Y2=0
cc_481 N_A_321_297#_M1017_s N_X_c_739_n 0.00165831f $X=6.655 $Y=1.485 $X2=0
+ $Y2=0
cc_482 N_A_321_297#_c_714_p N_X_c_739_n 0.0126919f $X=6.79 $Y=1.96 $X2=0 $Y2=0
cc_483 N_A_321_297#_c_656_n N_X_c_875_n 0.0118865f $X=7.505 $Y=2.38 $X2=0 $Y2=0
cc_484 N_A_321_297#_M1030_s N_X_c_740_n 0.00165831f $X=7.495 $Y=1.485 $X2=0
+ $Y2=0
cc_485 N_A_321_297#_c_717_p N_X_c_740_n 0.0126919f $X=7.63 $Y=1.96 $X2=0 $Y2=0
cc_486 N_A_321_297#_c_658_n N_X_c_878_n 0.0118865f $X=8.345 $Y=2.38 $X2=0 $Y2=0
cc_487 N_A_321_297#_M1034_s X 0.0033792f $X=8.335 $Y=1.485 $X2=0 $Y2=0
cc_488 N_A_321_297#_c_720_p X 0.0182127f $X=8.47 $Y=1.96 $X2=0 $Y2=0
cc_489 N_X_c_721_n N_VGND_M1003_s 0.00162089f $X=2.845 $Y=0.815 $X2=0 $Y2=0
cc_490 N_X_c_723_n N_VGND_M1008_s 0.00162089f $X=3.685 $Y=0.815 $X2=0 $Y2=0
cc_491 N_X_c_724_n N_VGND_M1028_s 0.00162089f $X=4.525 $Y=0.815 $X2=0 $Y2=0
cc_492 N_X_c_725_n N_VGND_M1035_s 0.00162089f $X=5.365 $Y=0.815 $X2=0 $Y2=0
cc_493 N_X_c_726_n N_VGND_M1006_d 0.00162089f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_494 N_X_c_727_n N_VGND_M1015_d 0.00162089f $X=7.045 $Y=0.815 $X2=0 $Y2=0
cc_495 N_X_c_728_n N_VGND_M1018_d 0.00162089f $X=7.885 $Y=0.815 $X2=0 $Y2=0
cc_496 N_X_c_735_n N_VGND_M1021_d 0.00290026f $X=8.27 $Y=0.815 $X2=0 $Y2=0
cc_497 N_X_c_722_n N_VGND_c_946_n 0.00843013f $X=2.335 $Y=0.815 $X2=0 $Y2=0
cc_498 N_X_c_744_n N_VGND_c_947_n 0.0188551f $X=2.17 $Y=0.39 $X2=0 $Y2=0
cc_499 N_X_c_721_n N_VGND_c_947_n 0.00198695f $X=2.845 $Y=0.815 $X2=0 $Y2=0
cc_500 N_X_c_721_n N_VGND_c_948_n 0.0122559f $X=2.845 $Y=0.815 $X2=0 $Y2=0
cc_501 N_X_c_723_n N_VGND_c_949_n 0.0122559f $X=3.685 $Y=0.815 $X2=0 $Y2=0
cc_502 N_X_c_724_n N_VGND_c_950_n 0.0122559f $X=4.525 $Y=0.815 $X2=0 $Y2=0
cc_503 N_X_c_725_n N_VGND_c_951_n 0.0122559f $X=5.365 $Y=0.815 $X2=0 $Y2=0
cc_504 N_X_c_726_n N_VGND_c_952_n 0.0122559f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_505 N_X_c_727_n N_VGND_c_953_n 0.0122559f $X=7.045 $Y=0.815 $X2=0 $Y2=0
cc_506 N_X_c_727_n N_VGND_c_954_n 0.00198695f $X=7.045 $Y=0.815 $X2=0 $Y2=0
cc_507 N_X_c_818_n N_VGND_c_954_n 0.0188551f $X=7.21 $Y=0.39 $X2=0 $Y2=0
cc_508 N_X_c_728_n N_VGND_c_954_n 0.00198695f $X=7.885 $Y=0.815 $X2=0 $Y2=0
cc_509 N_X_c_728_n N_VGND_c_955_n 0.0122559f $X=7.885 $Y=0.815 $X2=0 $Y2=0
cc_510 N_X_c_735_n N_VGND_c_957_n 0.0228574f $X=8.27 $Y=0.815 $X2=0 $Y2=0
cc_511 N_X_c_721_n N_VGND_c_960_n 0.00198695f $X=2.845 $Y=0.815 $X2=0 $Y2=0
cc_512 N_X_c_755_n N_VGND_c_960_n 0.0188551f $X=3.01 $Y=0.39 $X2=0 $Y2=0
cc_513 N_X_c_723_n N_VGND_c_960_n 0.00198695f $X=3.685 $Y=0.815 $X2=0 $Y2=0
cc_514 N_X_c_723_n N_VGND_c_962_n 0.00198695f $X=3.685 $Y=0.815 $X2=0 $Y2=0
cc_515 N_X_c_763_n N_VGND_c_962_n 0.0188551f $X=3.85 $Y=0.39 $X2=0 $Y2=0
cc_516 N_X_c_724_n N_VGND_c_962_n 0.00198695f $X=4.525 $Y=0.815 $X2=0 $Y2=0
cc_517 N_X_c_724_n N_VGND_c_964_n 0.00198695f $X=4.525 $Y=0.815 $X2=0 $Y2=0
cc_518 N_X_c_771_n N_VGND_c_964_n 0.0188551f $X=4.69 $Y=0.39 $X2=0 $Y2=0
cc_519 N_X_c_725_n N_VGND_c_964_n 0.00198695f $X=5.365 $Y=0.815 $X2=0 $Y2=0
cc_520 N_X_c_725_n N_VGND_c_966_n 0.00198695f $X=5.365 $Y=0.815 $X2=0 $Y2=0
cc_521 N_X_c_776_n N_VGND_c_966_n 0.0188551f $X=5.53 $Y=0.39 $X2=0 $Y2=0
cc_522 N_X_c_726_n N_VGND_c_966_n 0.00198695f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_523 N_X_c_726_n N_VGND_c_968_n 0.00198695f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_524 N_X_c_806_n N_VGND_c_968_n 0.0188551f $X=6.37 $Y=0.39 $X2=0 $Y2=0
cc_525 N_X_c_727_n N_VGND_c_968_n 0.00198695f $X=7.045 $Y=0.815 $X2=0 $Y2=0
cc_526 N_X_c_728_n N_VGND_c_971_n 0.00198695f $X=7.885 $Y=0.815 $X2=0 $Y2=0
cc_527 N_X_c_830_n N_VGND_c_971_n 0.0188614f $X=8.05 $Y=0.39 $X2=0 $Y2=0
cc_528 N_X_c_735_n N_VGND_c_971_n 0.00215161f $X=8.27 $Y=0.815 $X2=0 $Y2=0
cc_529 N_X_M1002_d N_VGND_c_975_n 0.00215201f $X=2.035 $Y=0.235 $X2=0 $Y2=0
cc_530 N_X_M1007_d N_VGND_c_975_n 0.00215201f $X=2.875 $Y=0.235 $X2=0 $Y2=0
cc_531 N_X_M1013_d N_VGND_c_975_n 0.00215201f $X=3.715 $Y=0.235 $X2=0 $Y2=0
cc_532 N_X_M1032_d N_VGND_c_975_n 0.00215201f $X=4.555 $Y=0.235 $X2=0 $Y2=0
cc_533 N_X_M1005_s N_VGND_c_975_n 0.00215201f $X=5.395 $Y=0.235 $X2=0 $Y2=0
cc_534 N_X_M1009_s N_VGND_c_975_n 0.00215201f $X=6.235 $Y=0.235 $X2=0 $Y2=0
cc_535 N_X_M1016_s N_VGND_c_975_n 0.00215201f $X=7.075 $Y=0.235 $X2=0 $Y2=0
cc_536 N_X_M1019_s N_VGND_c_975_n 0.00215201f $X=7.915 $Y=0.235 $X2=0 $Y2=0
cc_537 N_X_c_744_n N_VGND_c_975_n 0.0122069f $X=2.17 $Y=0.39 $X2=0 $Y2=0
cc_538 N_X_c_721_n N_VGND_c_975_n 0.00835832f $X=2.845 $Y=0.815 $X2=0 $Y2=0
cc_539 N_X_c_755_n N_VGND_c_975_n 0.0122069f $X=3.01 $Y=0.39 $X2=0 $Y2=0
cc_540 N_X_c_723_n N_VGND_c_975_n 0.00835832f $X=3.685 $Y=0.815 $X2=0 $Y2=0
cc_541 N_X_c_763_n N_VGND_c_975_n 0.0122069f $X=3.85 $Y=0.39 $X2=0 $Y2=0
cc_542 N_X_c_724_n N_VGND_c_975_n 0.00835832f $X=4.525 $Y=0.815 $X2=0 $Y2=0
cc_543 N_X_c_771_n N_VGND_c_975_n 0.0122069f $X=4.69 $Y=0.39 $X2=0 $Y2=0
cc_544 N_X_c_725_n N_VGND_c_975_n 0.00835832f $X=5.365 $Y=0.815 $X2=0 $Y2=0
cc_545 N_X_c_776_n N_VGND_c_975_n 0.0122069f $X=5.53 $Y=0.39 $X2=0 $Y2=0
cc_546 N_X_c_726_n N_VGND_c_975_n 0.00835832f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_547 N_X_c_806_n N_VGND_c_975_n 0.0122069f $X=6.37 $Y=0.39 $X2=0 $Y2=0
cc_548 N_X_c_727_n N_VGND_c_975_n 0.00835832f $X=7.045 $Y=0.815 $X2=0 $Y2=0
cc_549 N_X_c_818_n N_VGND_c_975_n 0.0122069f $X=7.21 $Y=0.39 $X2=0 $Y2=0
cc_550 N_X_c_728_n N_VGND_c_975_n 0.00835832f $X=7.885 $Y=0.815 $X2=0 $Y2=0
cc_551 N_X_c_830_n N_VGND_c_975_n 0.0122084f $X=8.05 $Y=0.39 $X2=0 $Y2=0
cc_552 N_X_c_735_n N_VGND_c_975_n 0.00529045f $X=8.27 $Y=0.815 $X2=0 $Y2=0

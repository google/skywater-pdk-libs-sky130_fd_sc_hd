* File: sky130_fd_sc_hd__or4b_1.spice
* Created: Thu Aug 27 14:44:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4b_1.spice.pex"
.subckt sky130_fd_sc_hd__or4b_1  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1002 N_A_109_53#_M1002_d N_D_N_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_215_297#_M1005_d N_A_109_53#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.06405 AS=0.1092 PD=0.725 PS=1.36 NRD=7.14 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g N_A_215_297#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.06405 PD=0.69 PS=0.725 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1003 N_A_215_297#_M1003_d N_B_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_215_297#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_215_297#_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.123773 PD=1.85 PS=1.2028 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_109_53#_M1007_d N_D_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_297_297# N_A_109_53#_M1000_g N_A_215_297#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06825 AS=0.1092 PD=0.745 PS=1.36 NRD=50.4123 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1009 A_392_297# N_C_M1009_g A_297_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.04515
+ AS=0.06825 PD=0.635 PS=0.745 NRD=24.6053 NRS=50.4123 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1010 A_465_297# N_B_M1010_g A_392_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.06405
+ AS=0.04515 PD=0.725 PS=0.635 NRD=45.7237 NRS=24.6053 M=1 R=2.8 SA=75001
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g A_465_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.06405 PD=0.792676 PS=0.725 NRD=72.1217 NRS=45.7237 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_215_297#_M1001_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.208803 PD=2.55 PS=1.88732 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_73 VPB 0 1.14153e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__or4b_1.spice.SKY130_FD_SC_HD__OR4B_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__nand2_8.pex.spice
* Created: Tue Sep  1 19:15:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2_8%B 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 66 67 68 69 70 90 91
c169 90 0 1.93909e-19 $X=3.2 $Y=1.16
c170 59 0 8.09502e-20 $X=3.41 $Y=0.56
r171 89 91 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.2 $Y=1.16
+ $X2=3.41 $Y2=1.16
r172 89 90 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.2
+ $Y=1.16 $X2=3.2 $Y2=1.16
r173 87 89 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.2 $Y2=1.16
r174 86 87 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r175 85 86 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r176 84 85 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=2.15 $Y2=1.16
r177 83 84 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r178 82 83 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r179 80 82 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=0.675 $Y=1.16
+ $X2=0.89 $Y2=1.16
r180 77 80 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.675 $Y2=1.16
r181 70 90 10.7387 $w=2.18e-07 $l=2.05e-07 $layer=LI1_cond $X=2.995 $Y=1.185
+ $X2=3.2 $Y2=1.185
r182 69 70 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.185
+ $X2=2.995 $Y2=1.185
r183 68 69 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=2.075 $Y=1.185
+ $X2=2.535 $Y2=1.185
r184 67 68 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=1.615 $Y=1.185
+ $X2=2.075 $Y2=1.185
r185 66 67 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.185
+ $X2=1.615 $Y2=1.185
r186 65 66 25.1442 $w=2.18e-07 $l=4.8e-07 $layer=LI1_cond $X=0.675 $Y=1.185
+ $X2=1.155 $Y2=1.185
r187 65 80 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.675
+ $Y=1.16 $X2=0.675 $Y2=1.16
r188 61 91 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r189 61 63 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r190 57 91 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r191 57 59 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r192 53 87 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r193 53 55 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r194 49 87 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r195 49 51 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r196 45 86 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r197 45 47 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r198 41 86 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r199 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r200 37 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r201 37 39 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r202 33 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r203 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r204 29 84 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r205 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r206 25 84 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r207 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r208 21 83 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r209 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r210 17 83 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r211 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r212 13 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r213 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r214 9 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r215 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r216 5 77 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r217 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.985
r218 1 77 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r219 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 66 67 68 69 89
c138 89 0 1.93909e-19 $X=6.77 $Y=1.16
c139 3 0 1.56255e-19 $X=3.83 $Y=0.56
r140 88 89 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.35 $Y=1.16
+ $X2=6.77 $Y2=1.16
r141 86 88 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=6.14 $Y=1.16
+ $X2=6.35 $Y2=1.16
r142 84 86 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.93 $Y=1.16
+ $X2=6.14 $Y2=1.16
r143 83 84 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.93 $Y2=1.16
r144 82 83 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.51 $Y2=1.16
r145 81 82 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.67 $Y=1.16
+ $X2=5.09 $Y2=1.16
r146 79 81 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.67 $Y2=1.16
r147 77 79 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.46 $Y2=1.16
r148 75 77 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.83 $Y=1.16
+ $X2=4.25 $Y2=1.16
r149 69 86 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.14
+ $Y=1.16 $X2=6.14 $Y2=1.16
r150 68 69 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=5.755 $Y=1.175
+ $X2=6.14 $Y2=1.175
r151 67 68 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=5.295 $Y=1.175
+ $X2=5.755 $Y2=1.175
r152 66 67 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.835 $Y=1.175
+ $X2=5.295 $Y2=1.175
r153 65 66 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=4.835 $Y2=1.175
r154 65 79 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r155 61 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.16
r156 61 63 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.985
r157 57 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=1.16
r158 57 59 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=0.56
r159 53 88 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.16
r160 53 55 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.985
r161 49 88 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=1.16
r162 49 51 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=0.56
r163 45 84 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.16
r164 45 47 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.985
r165 41 84 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=1.16
r166 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=0.56
r167 37 83 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.16
r168 37 39 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.985
r169 33 83 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=1.16
r170 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=0.56
r171 29 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.16
r172 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.985
r173 25 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=1.16
r174 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=0.56
r175 21 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.16
r176 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.985
r177 17 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=1.16
r178 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=0.56
r179 13 77 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.16
r180 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.985
r181 9 77 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=1.16
r182 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
r183 5 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.16
r184 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.985
r185 1 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.16
r186 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_8%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 48 52
+ 54 58 62 64 66 71 72 74 75 77 78 80 81 82 83 85 86 87 109 117 121
r120 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r121 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r122 112 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r123 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r124 109 120 5.03279 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.915 $Y=2.72
+ $X2=7.137 $Y2=2.72
r125 109 111 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=2.72
+ $X2=6.67 $Y2=2.72
r126 108 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r127 108 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r129 105 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.3 $Y2=2.72
r130 105 107 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.75 $Y2=2.72
r131 104 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r132 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r134 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r135 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r136 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r137 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r138 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r139 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r141 89 114 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r142 89 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r143 87 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r144 87 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 85 107 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=5.75 $Y2=2.72
r146 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=6.14 $Y2=2.72
r147 84 111 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.225 $Y=2.72
+ $X2=6.67 $Y2=2.72
r148 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=2.72
+ $X2=6.14 $Y2=2.72
r149 82 103 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.37 $Y2=2.72
r150 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.46 $Y2=2.72
r151 80 100 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r152 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.62 $Y2=2.72
r153 79 103 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.705 $Y=2.72
+ $X2=4.37 $Y2=2.72
r154 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=2.72
+ $X2=3.62 $Y2=2.72
r155 77 97 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r156 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.78 $Y2=2.72
r157 76 100 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.45 $Y2=2.72
r158 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.78 $Y2=2.72
r159 74 94 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r160 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r161 73 97 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r162 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r163 71 91 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r164 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r165 70 94 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r166 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r167 66 69 22.075 $w=3.53e-07 $l=6.8e-07 $layer=LI1_cond $X=7.092 $Y=1.66
+ $X2=7.092 $Y2=2.34
r168 64 120 2.94713 $w=3.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=7.092 $Y=2.635
+ $X2=7.137 $Y2=2.72
r169 64 69 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=7.092 $Y=2.635
+ $X2=7.092 $Y2=2.34
r170 60 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=2.635
+ $X2=6.14 $Y2=2.72
r171 60 62 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.14 $Y=2.635
+ $X2=6.14 $Y2=2
r172 56 117 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r173 56 58 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2
r174 55 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.46 $Y2=2.72
r175 54 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=2.72
+ $X2=5.3 $Y2=2.72
r176 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.215 $Y=2.72
+ $X2=4.545 $Y2=2.72
r177 50 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2.72
r178 50 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2
r179 46 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r180 46 48 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2
r181 42 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r182 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r183 38 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r184 38 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r185 34 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r186 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r187 30 33 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r188 28 114 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r189 28 33 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r190 9 69 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=7.08 $Y2=2.34
r191 9 66 400 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=7.08 $Y2=1.66
r192 8 62 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.005
+ $Y=1.485 $X2=6.14 $Y2=2
r193 7 58 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2
r194 6 52 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2
r195 5 48 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2
r196 4 44 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r197 3 40 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r198 2 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r199 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r200 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 37 39 41 45 47
+ 51 53 57 59 61 62 63 65 67 73 77 79 83 85 89 91 92 96 98 100 104 106 108 111
+ 112
c189 61 0 8.09502e-20 $X=3.997 $Y=0.905
r190 119 121 2.2815 $w=5.08e-07 $l=9.5e-08 $layer=LI1_cond $X=3.922 $Y=1.565
+ $X2=3.922 $Y2=1.66
r191 112 119 0.840551 $w=5.08e-07 $l=3.5e-08 $layer=LI1_cond $X=3.922 $Y=1.53
+ $X2=3.922 $Y2=1.565
r192 111 112 8.16535 $w=5.08e-07 $l=3.4e-07 $layer=LI1_cond $X=3.922 $Y=1.19
+ $X2=3.922 $Y2=1.53
r193 92 108 3.75388 $w=2.9e-07 $l=1.18322e-07 $layer=LI1_cond $X=6.6 $Y=1.465
+ $X2=6.56 $Y2=1.565
r194 91 110 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.6 $Y=0.905
+ $X2=6.6 $Y2=0.78
r195 91 92 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=6.6 $Y=0.905
+ $X2=6.6 $Y2=1.465
r196 87 108 3.75388 $w=2.9e-07 $l=1e-07 $layer=LI1_cond $X=6.56 $Y=1.665
+ $X2=6.56 $Y2=1.565
r197 87 89 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.56 $Y=1.665
+ $X2=6.56 $Y2=2.34
r198 86 106 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.885 $Y=1.565
+ $X2=5.72 $Y2=1.565
r199 85 108 2.70891 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.565
+ $X2=6.56 $Y2=1.565
r200 85 86 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=6.395 $Y=1.565
+ $X2=5.885 $Y2=1.565
r201 81 106 0.381419 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=5.72 $Y=1.665
+ $X2=5.72 $Y2=1.565
r202 81 83 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.72 $Y=1.665
+ $X2=5.72 $Y2=2.34
r203 80 104 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=1.565
+ $X2=4.88 $Y2=1.565
r204 79 106 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.555 $Y=1.565
+ $X2=5.72 $Y2=1.565
r205 79 80 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=5.555 $Y=1.565
+ $X2=5.045 $Y2=1.565
r206 75 104 0.381419 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=4.88 $Y=1.665
+ $X2=4.88 $Y2=1.565
r207 75 77 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.88 $Y=1.665
+ $X2=4.88 $Y2=2.34
r208 74 119 6.24589 $w=2e-07 $l=2.83e-07 $layer=LI1_cond $X=4.205 $Y=1.565
+ $X2=3.922 $Y2=1.565
r209 73 104 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=1.565
+ $X2=4.88 $Y2=1.565
r210 73 74 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=4.715 $Y=1.565
+ $X2=4.205 $Y2=1.565
r211 70 72 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=4.88 $Y=0.78
+ $X2=5.72 $Y2=0.78
r212 68 102 3.38121 $w=2.5e-07 $l=1.23e-07 $layer=LI1_cond $X=4.12 $Y=0.78
+ $X2=3.997 $Y2=0.78
r213 68 70 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=4.12 $Y=0.78
+ $X2=4.88 $Y2=0.78
r214 67 110 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=0.78
+ $X2=6.6 $Y2=0.78
r215 67 72 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=6.475 $Y=0.78
+ $X2=5.72 $Y2=0.78
r216 63 121 1.61573 $w=5.08e-07 $l=1.20474e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=3.922 $Y2=1.66
r217 63 65 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=2.34
r218 62 111 6.04247 $w=5.08e-07 $l=1.47817e-07 $layer=LI1_cond $X=3.997 $Y=1.075
+ $X2=3.922 $Y2=1.19
r219 61 102 3.43619 $w=2.45e-07 $l=1.25e-07 $layer=LI1_cond $X=3.997 $Y=0.905
+ $X2=3.997 $Y2=0.78
r220 61 62 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=3.997 $Y=0.905
+ $X2=3.997 $Y2=1.075
r221 60 100 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=1.565
+ $X2=3.2 $Y2=1.565
r222 59 119 6.24589 $w=2e-07 $l=2.82e-07 $layer=LI1_cond $X=3.64 $Y=1.565
+ $X2=3.922 $Y2=1.565
r223 59 60 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.64 $Y=1.565
+ $X2=3.365 $Y2=1.565
r224 55 100 0.381419 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=3.2 $Y=1.665 $X2=3.2
+ $Y2=1.565
r225 55 57 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.2 $Y=1.665
+ $X2=3.2 $Y2=2.34
r226 54 98 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=1.565
+ $X2=2.36 $Y2=1.565
r227 53 100 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.565
+ $X2=3.2 $Y2=1.565
r228 53 54 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=3.035 $Y=1.565
+ $X2=2.525 $Y2=1.565
r229 49 98 0.381419 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=1.565
r230 49 51 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=2.34
r231 48 96 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.565
+ $X2=1.52 $Y2=1.565
r232 47 98 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=1.565
+ $X2=2.36 $Y2=1.565
r233 47 48 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=2.195 $Y=1.565
+ $X2=1.685 $Y2=1.565
r234 43 96 0.381419 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.565
r235 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r236 42 94 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.565
+ $X2=0.68 $Y2=1.565
r237 41 96 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.565
+ $X2=1.52 $Y2=1.565
r238 41 42 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.565
+ $X2=0.845 $Y2=1.565
r239 37 94 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=0.68 $Y=1.665 $X2=0.68
+ $Y2=1.565
r240 37 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r241 12 108 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.485 $X2=6.56 $Y2=1.66
r242 12 89 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.485 $X2=6.56 $Y2=2.34
r243 11 106 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=1.66
r244 11 83 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=2.34
r245 10 104 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.66
r246 10 77 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2.34
r247 9 121 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=1.66
r248 9 65 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=2.34
r249 8 100 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.66
r250 8 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.34
r251 7 98 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.66
r252 7 51 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.34
r253 6 96 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r254 6 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r255 5 94 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r256 5 39 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r257 4 110 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=6.425
+ $Y=0.235 $X2=6.56 $Y2=0.74
r258 3 72 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.74
r259 2 70 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.74
r260 1 102 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_8%A_27_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 52 53 54 62 64 66 67 68
c129 53 0 1.56255e-19 $X=3.58 $Y=0.735
r130 62 74 2.79446 $w=3.75e-07 $l=1.15e-07 $layer=LI1_cond $X=7.082 $Y=0.485
+ $X2=7.082 $Y2=0.37
r131 62 64 7.83661 $w=3.73e-07 $l=2.55e-07 $layer=LI1_cond $X=7.082 $Y=0.485
+ $X2=7.082 $Y2=0.74
r132 59 61 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=5.3 $Y=0.37
+ $X2=6.14 $Y2=0.37
r133 57 59 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=4.46 $Y=0.37
+ $X2=5.3 $Y2=0.37
r134 55 70 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.705 $Y=0.37
+ $X2=3.58 $Y2=0.37
r135 55 57 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=3.705 $Y=0.37
+ $X2=4.46 $Y2=0.37
r136 54 74 4.54403 $w=2.3e-07 $l=1.87e-07 $layer=LI1_cond $X=6.895 $Y=0.37
+ $X2=7.082 $Y2=0.37
r137 54 61 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=6.895 $Y=0.37
+ $X2=6.14 $Y2=0.37
r138 53 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=0.735
+ $X2=3.58 $Y2=0.82
r139 52 70 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=3.58 $Y=0.485
+ $X2=3.58 $Y2=0.37
r140 52 53 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.58 $Y=0.485
+ $X2=3.58 $Y2=0.735
r141 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0.82
+ $X2=2.78 $Y2=0.82
r142 50 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.455 $Y=0.82
+ $X2=3.58 $Y2=0.82
r143 50 51 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.455 $Y=0.82
+ $X2=2.945 $Y2=0.82
r144 46 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.82
r145 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.4
r146 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0.82
+ $X2=1.94 $Y2=0.82
r147 44 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0.82
+ $X2=2.78 $Y2=0.82
r148 44 45 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.615 $Y=0.82
+ $X2=2.105 $Y2=0.82
r149 40 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.82
r150 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.4
r151 39 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0.82
+ $X2=1.1 $Y2=0.82
r152 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0.82
+ $X2=1.94 $Y2=0.82
r153 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=0.82
+ $X2=1.265 $Y2=0.82
r154 34 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.735 $X2=1.1
+ $Y2=0.82
r155 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.4
r156 32 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=1.1 $Y2=0.82
r157 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=0.425 $Y2=0.82
r158 28 33 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r159 28 30 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.4
r160 9 74 182 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=1 $X=6.845
+ $Y=0.235 $X2=7.08 $Y2=0.4
r161 9 64 182 $w=1.7e-07 $l=6.1131e-07 $layer=licon1_NDIFF $count=1 $X=6.845
+ $Y=0.235 $X2=7.08 $Y2=0.74
r162 8 61 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.005
+ $Y=0.235 $X2=6.14 $Y2=0.4
r163 7 59 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.165
+ $Y=0.235 $X2=5.3 $Y2=0.4
r164 6 57 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.4
r165 5 72 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.74
r166 5 70 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.4
r167 4 48 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.4
r168 3 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.4
r169 2 36 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r170 1 30 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_8%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 39 40 41 60 61
r101 60 61 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r102 58 61 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=7.13
+ $Y2=0
r103 57 60 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=7.13
+ $Y2=0
r104 57 58 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r105 55 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r106 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r107 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r108 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r109 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r110 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r111 41 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r112 41 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r113 39 54 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=0
+ $X2=2.99 $Y2=0
r114 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.2
+ $Y2=0
r115 38 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.45 $Y2=0
r116 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.2
+ $Y2=0
r117 36 51 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.07 $Y2=0
r118 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.36
+ $Y2=0
r119 35 54 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.99 $Y2=0
r120 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.36
+ $Y2=0
r121 33 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.15 $Y2=0
r122 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.52
+ $Y2=0
r123 32 51 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=2.07 $Y2=0
r124 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.52
+ $Y2=0
r125 30 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r126 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r127 29 48 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=1.15 $Y2=0
r128 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r129 25 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.085 $X2=3.2
+ $Y2=0
r130 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0.4
r131 21 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r132 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.4
r133 17 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r134 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r135 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r136 13 15 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r137 4 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.4
r138 3 23 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.4
r139 2 19 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r140 1 15 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends


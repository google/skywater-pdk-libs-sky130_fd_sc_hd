* NGSPICE file created from sky130_fd_sc_hd__nand3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
M1000 VPWR B Y VPB phighvt w=1e+06u l=150000u
+  ad=5.9e+11p pd=5.18e+06u as=5.3e+11p ps=5.06e+06u
M1001 a_193_47# B a_109_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u
M1002 Y C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A a_193_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1004 a_109_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1005 Y A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__and3b_4.spice.pex
* Created: Thu Aug 27 14:08:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND3B_4%A_98_199# 1 2 9 12 15 16 17 18 20 24 26 31
c81 16 0 1.70701e-19 $X=4.165 $Y=1.99
c82 12 0 1.97561e-19 $X=0.685 $Y=1.985
r83 24 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.16
+ $X2=0.625 $Y2=1.325
r84 24 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.16
+ $X2=0.625 $Y2=0.995
r85 23 26 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.625 $Y=1.16
+ $X2=0.765 $Y2=1.16
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.16 $X2=0.625 $Y2=1.16
r87 18 29 3.11269 $w=2.8e-07 $l=1.15e-07 $layer=LI1_cond $X=4.305 $Y=1.875
+ $X2=4.305 $Y2=1.99
r88 18 20 52.8889 $w=2.78e-07 $l=1.285e-06 $layer=LI1_cond $X=4.305 $Y=1.875
+ $X2=4.305 $Y2=0.59
r89 16 29 3.78936 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=4.165 $Y=1.99
+ $X2=4.305 $Y2=1.99
r90 16 17 166.102 $w=2.28e-07 $l=3.315e-06 $layer=LI1_cond $X=4.165 $Y=1.99
+ $X2=0.85 $Y2=1.99
r91 15 17 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.765 $Y=1.875
+ $X2=0.85 $Y2=1.99
r92 14 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=1.325
+ $X2=0.765 $Y2=1.16
r93 14 15 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.765 $Y=1.325
+ $X2=0.765 $Y2=1.875
r94 12 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.685 $Y=1.985
+ $X2=0.685 $Y2=1.325
r95 9 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.685 $Y=0.56
+ $X2=0.685 $Y2=0.995
r96 2 29 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.725 $X2=4.18 $Y2=2.02
r97 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.465 $X2=4.25 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%B 3 6 8 9 13 15
c41 8 0 5.73368e-20 $X=1.065 $Y=0.765
c42 6 0 9.13552e-20 $X=1.21 $Y=1.985
r43 13 16 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=1.127 $Y=1.16
+ $X2=1.127 $Y2=1.325
r44 13 15 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=1.127 $Y=1.16
+ $X2=1.127 $Y2=0.995
r45 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.16 $X2=1.105 $Y2=1.16
r46 8 9 16.6166 $w=2.13e-07 $l=3.1e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.16
r47 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.21 $Y=1.985
+ $X2=1.21 $Y2=1.325
r48 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.21 $Y=0.56 $X2=1.21
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%C 3 6 8 11 13
c40 11 0 1.82625e-19 $X=1.63 $Y=1.16
c41 8 0 9.13552e-20 $X=1.61 $Y=1.19
c42 6 0 1.66082e-19 $X=1.66 $Y=1.985
r43 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=1.325
r44 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=0.995
r45 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.16 $X2=1.63 $Y2=1.16
r46 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.66 $Y=1.985
+ $X2=1.66 $Y2=1.325
r47 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.59 $Y=0.56 $X2=1.59
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%A_56_297# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 42 44 48 51 53 59 63 68 69 70 74 82
c146 82 0 1.70701e-19 $X=3.455 $Y=1.16
c147 51 0 1.82625e-19 $X=2 $Y=1.02
c148 48 0 8.37355e-20 $X=1.885 $Y=0.71
c149 44 0 1.55732e-19 $X=1.885 $Y=1.61
r150 81 82 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.025 $Y=1.16
+ $X2=3.455 $Y2=1.16
r151 78 79 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.605 $Y2=1.16
r152 70 72 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=1.51 $Y=0.45
+ $X2=1.51 $Y2=0.71
r153 68 69 7.01282 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.33 $Y=1.66
+ $X2=0.33 $Y2=1.495
r154 66 69 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=0.26 $Y=0.805
+ $X2=0.26 $Y2=1.495
r155 65 66 12.3665 $w=4.83e-07 $l=3.55e-07 $layer=LI1_cond $X=0.392 $Y=0.45
+ $X2=0.392 $Y2=0.805
r156 63 65 1.7263 $w=4.83e-07 $l=7e-08 $layer=LI1_cond $X=0.392 $Y=0.38
+ $X2=0.392 $Y2=0.45
r157 60 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.935 $Y=1.16
+ $X2=3.025 $Y2=1.16
r158 60 79 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.935 $Y=1.16
+ $X2=2.605 $Y2=1.16
r159 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.16 $X2=2.935 $Y2=1.16
r160 57 78 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.595 $Y2=1.16
r161 57 75 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.165 $Y2=1.16
r162 56 59 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=2.255 $Y=1.187
+ $X2=2.935 $Y2=1.187
r163 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=1.16 $X2=2.255 $Y2=1.16
r164 54 74 0.43014 $w=3.35e-07 $l=1.15e-07 $layer=LI1_cond $X=2.115 $Y=1.187
+ $X2=2 $Y2=1.187
r165 54 56 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=2.115 $Y=1.187
+ $X2=2.255 $Y2=1.187
r166 52 74 7.74634 $w=2e-07 $l=1.82384e-07 $layer=LI1_cond $X=1.97 $Y=1.355
+ $X2=2 $Y2=1.187
r167 52 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.97 $Y=1.355
+ $X2=1.97 $Y2=1.525
r168 51 74 7.74634 $w=2e-07 $l=1.67e-07 $layer=LI1_cond $X=2 $Y=1.02 $X2=2
+ $Y2=1.187
r169 50 51 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2 $Y=0.805 $X2=2
+ $Y2=1.02
r170 49 72 0.384081 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.6 $Y=0.71 $X2=1.51
+ $Y2=0.71
r171 48 50 6.89722 $w=1.9e-07 $l=1.55403e-07 $layer=LI1_cond $X=1.885 $Y=0.71
+ $X2=2 $Y2=0.805
r172 48 49 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=1.885 $Y=0.71
+ $X2=1.6 $Y2=0.71
r173 44 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.885 $Y=1.61
+ $X2=1.97 $Y2=1.525
r174 44 46 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.885 $Y=1.61
+ $X2=1.445 $Y2=1.61
r175 43 65 6.27638 $w=1.9e-07 $l=2.43e-07 $layer=LI1_cond $X=0.635 $Y=0.45
+ $X2=0.392 $Y2=0.45
r176 42 70 0.384081 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.42 $Y=0.45 $X2=1.51
+ $Y2=0.45
r177 42 43 45.823 $w=1.88e-07 $l=7.85e-07 $layer=LI1_cond $X=1.42 $Y=0.45
+ $X2=0.635 $Y2=0.45
r178 34 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.455 $Y=1.325
+ $X2=3.455 $Y2=1.16
r179 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.455 $Y=1.325
+ $X2=3.455 $Y2=1.985
r180 31 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=1.16
r181 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=0.56
r182 27 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.025 $Y=1.325
+ $X2=3.025 $Y2=1.16
r183 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.025 $Y=1.325
+ $X2=3.025 $Y2=1.985
r184 24 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.025 $Y=0.995
+ $X2=3.025 $Y2=1.16
r185 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.025 $Y=0.995
+ $X2=3.025 $Y2=0.56
r186 20 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.605 $Y=1.325
+ $X2=2.605 $Y2=1.16
r187 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.605 $Y=1.325
+ $X2=2.605 $Y2=1.985
r188 17 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.595 $Y=0.995
+ $X2=2.595 $Y2=1.16
r189 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.595 $Y=0.995
+ $X2=2.595 $Y2=0.56
r190 13 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=1.325
+ $X2=2.165 $Y2=1.16
r191 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.165 $Y=1.325
+ $X2=2.165 $Y2=1.985
r192 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=1.16
r193 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=0.56
r194 3 46 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=1.285
+ $Y=1.485 $X2=1.445 $Y2=1.61
r195 2 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=1.485 $X2=0.425 $Y2=1.66
r196 1 63 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=0.305
+ $Y=0.235 $X2=0.47 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%A_N 3 6 7 8 12 14 15
r31 12 15 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.902 $Y=1.16
+ $X2=3.902 $Y2=1.325
r32 12 14 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.902 $Y=1.16
+ $X2=3.902 $Y2=0.995
r33 7 8 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.855 $Y=1.16
+ $X2=3.855 $Y2=1.53
r34 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9 $Y=1.16
+ $X2=3.9 $Y2=1.16
r35 6 15 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.965 $Y=1.935
+ $X2=3.965 $Y2=1.325
r36 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.965 $Y=0.675
+ $X2=3.965 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%VPWR 1 2 3 4 15 19 23 26 29 33 34 36 37 39
+ 40 41 57 58
r72 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r74 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r75 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r76 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r79 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r80 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 41 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 39 54 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.67 $Y2=2.72
r84 38 57 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.835 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=2.72
+ $X2=3.67 $Y2=2.72
r86 36 51 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.645 $Y=2.72
+ $X2=2.53 $Y2=2.72
r87 36 37 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.645 $Y=2.72
+ $X2=2.812 $Y2=2.72
r88 35 54 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 35 37 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=2.812 $Y2=2.72
r90 33 48 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=1.61 $Y2=2.72
r91 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=1.91 $Y2=2.72
r92 32 51 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=2.53 $Y2=2.72
r93 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=1.91 $Y2=2.72
r94 30 48 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.18 $Y=2.72
+ $X2=1.61 $Y2=2.72
r95 29 44 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.73 $Y=2.72 $X2=0.69
+ $Y2=2.72
r96 28 30 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.18 $Y2=2.72
r97 28 29 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.73 $Y2=2.72
r98 26 28 9.56863 $w=4.48e-07 $l=3.6e-07 $layer=LI1_cond $X=0.955 $Y=2.36
+ $X2=0.955 $Y2=2.72
r99 21 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=2.635
+ $X2=3.67 $Y2=2.72
r100 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.67 $Y=2.635
+ $X2=3.67 $Y2=2.36
r101 17 37 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.812 $Y=2.635
+ $X2=2.812 $Y2=2.72
r102 17 19 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.812 $Y=2.635
+ $X2=2.812 $Y2=2.36
r103 13 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=2.635
+ $X2=1.91 $Y2=2.72
r104 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.91 $Y=2.635
+ $X2=1.91 $Y2=2.36
r105 4 23 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.485 $X2=3.67 $Y2=2.36
r106 3 19 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.815 $Y2=2.36
r107 2 15 600 $w=1.7e-07 $l=9.58514e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=1.485 $X2=1.91 $Y2=2.36
r108 1 26 600 $w=1.7e-07 $l=9.72111e-07 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=1.485 $X2=0.965 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%X 1 2 3 4 13 19 23 28 30 35
c45 13 0 1.50574e-19 $X=3.27 $Y=1.62
r46 33 35 0.217442 $w=2.63e-07 $l=5e-09 $layer=LI1_cond $X=3.402 $Y=0.845
+ $X2=3.402 $Y2=0.85
r47 30 33 5.21318 $w=2.27e-07 $l=1.42671e-07 $layer=LI1_cond $X=3.34 $Y=0.73
+ $X2=3.402 $Y2=0.845
r48 30 35 1.73954 $w=2.63e-07 $l=4e-08 $layer=LI1_cond $X=3.402 $Y=0.89
+ $X2=3.402 $Y2=0.85
r49 29 30 28.05 $w=2.63e-07 $l=6.45e-07 $layer=LI1_cond $X=3.402 $Y=1.535
+ $X2=3.402 $Y2=0.89
r50 26 28 4.38803 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=0.68
+ $X2=2.475 $Y2=0.68
r51 21 30 5.21318 $w=2.27e-07 $l=1.57242e-07 $layer=LI1_cond $X=3.24 $Y=0.615
+ $X2=3.34 $Y2=0.73
r52 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.24 $Y=0.615
+ $X2=3.24 $Y2=0.42
r53 19 30 1.30324 $w=2.3e-07 $l=1.95e-07 $layer=LI1_cond $X=3.145 $Y=0.73
+ $X2=3.34 $Y2=0.73
r54 19 28 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.145 $Y=0.73
+ $X2=2.475 $Y2=0.73
r55 15 18 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.39 $Y=1.62
+ $X2=3.24 $Y2=1.62
r56 13 29 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.27 $Y=1.62
+ $X2=3.402 $Y2=1.535
r57 13 18 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.27 $Y=1.62 $X2=3.24
+ $Y2=1.62
r58 4 18 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=1.485 $X2=3.24 $Y2=1.62
r59 3 15 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.485 $X2=2.39 $Y2=1.62
r60 2 30 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.1
+ $Y=0.235 $X2=3.24 $Y2=0.76
r61 2 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.1
+ $Y=0.235 $X2=3.24 $Y2=0.42
r62 1 26 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.38 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_4%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 47
+ 48
c74 26 0 8.37355e-20 $X=2.645 $Y=0
r75 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r76 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r77 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r78 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r79 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r80 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r81 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r82 34 38 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r83 31 39 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r84 31 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r85 29 44 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.45
+ $Y2=0
r86 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.67
+ $Y2=0
r87 28 47 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.835 $Y=0 $X2=4.37
+ $Y2=0
r88 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.67
+ $Y2=0
r89 26 41 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.53
+ $Y2=0
r90 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.81
+ $Y2=0
r91 25 44 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.45
+ $Y2=0
r92 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.81
+ $Y2=0
r93 23 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.61
+ $Y2=0
r94 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.945
+ $Y2=0
r95 22 41 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.53
+ $Y2=0
r96 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.945
+ $Y2=0
r97 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0.085
+ $X2=3.67 $Y2=0
r98 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.67 $Y=0.085
+ $X2=3.67 $Y2=0.36
r99 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.085
+ $X2=2.81 $Y2=0
r100 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.81 $Y=0.085
+ $X2=2.81 $Y2=0.36
r101 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=0.085
+ $X2=1.945 $Y2=0
r102 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.945 $Y=0.085
+ $X2=1.945 $Y2=0.36
r103 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.53
+ $Y=0.235 $X2=3.67 $Y2=0.36
r104 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.235 $X2=2.81 $Y2=0.36
r105 1 12 182 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.235 $X2=1.945 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__nor2_2.pxi.spice
* Created: Tue Sep  1 19:17:41 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2_2%A N_A_c_43_n N_A_M1002_g N_A_M1000_g N_A_c_44_n
+ N_A_M1004_g N_A_M1007_g A A N_A_c_46_n PM_SKY130_FD_SC_HD__NOR2_2%A
x_PM_SKY130_FD_SC_HD__NOR2_2%B N_B_c_81_n N_B_M1001_g N_B_M1005_g N_B_c_82_n
+ N_B_M1003_g N_B_M1006_g B B N_B_c_84_n PM_SKY130_FD_SC_HD__NOR2_2%B
x_PM_SKY130_FD_SC_HD__NOR2_2%A_27_297# N_A_27_297#_M1000_s N_A_27_297#_M1007_s
+ N_A_27_297#_M1006_d N_A_27_297#_c_128_n N_A_27_297#_c_129_n
+ N_A_27_297#_c_130_n N_A_27_297#_c_131_n N_A_27_297#_c_147_p
+ N_A_27_297#_c_132_n N_A_27_297#_c_133_n PM_SKY130_FD_SC_HD__NOR2_2%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR2_2%VPWR N_VPWR_M1000_d N_VPWR_c_164_n VPWR
+ N_VPWR_c_165_n N_VPWR_c_166_n N_VPWR_c_163_n N_VPWR_c_168_n
+ PM_SKY130_FD_SC_HD__NOR2_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR2_2%Y N_Y_M1002_s N_Y_M1001_d N_Y_M1005_s N_Y_c_199_n
+ N_Y_c_192_n N_Y_c_193_n N_Y_c_206_n N_Y_c_194_n N_Y_c_195_n N_Y_c_196_n
+ N_Y_c_198_n Y PM_SKY130_FD_SC_HD__NOR2_2%Y
x_PM_SKY130_FD_SC_HD__NOR2_2%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_M1003_s
+ N_VGND_c_251_n N_VGND_c_252_n N_VGND_c_253_n N_VGND_c_254_n N_VGND_c_255_n
+ N_VGND_c_256_n N_VGND_c_257_n VGND N_VGND_c_258_n N_VGND_c_259_n
+ PM_SKY130_FD_SC_HD__NOR2_2%VGND
cc_1 VNB N_A_c_43_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_44_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB A 0.0165272f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_A_c_46_n 0.0372851f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_5 VNB N_B_c_81_n 0.0160101f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_82_n 0.0191673f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_7 VNB B 0.00630293f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_B_c_84_n 0.033234f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_9 VNB N_VPWR_c_163_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_10 VNB N_Y_c_192_n 0.00248283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_193_n 0.00238181f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_Y_c_194_n 0.00897642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_Y_c_195_n 0.0195815f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_14 VNB N_Y_c_196_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_15 VNB N_VGND_c_251_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_16 VNB N_VGND_c_252_n 0.0329389f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_17 VNB N_VGND_c_253_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_18 VNB N_VGND_c_254_n 0.0120543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_255_n 0.019039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_256_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_21 VNB N_VGND_c_257_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_22 VNB N_VGND_c_258_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_259_n 0.143274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_A_M1000_g 0.0250431f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_25 VPB N_A_M1007_g 0.0182765f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_26 VPB N_A_c_46_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_27 VPB N_B_M1005_g 0.018627f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_28 VPB N_B_M1006_g 0.0219547f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_29 VPB N_B_c_84_n 0.0042141f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_30 VPB N_A_27_297#_c_128_n 0.0116274f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_31 VPB N_A_27_297#_c_129_n 0.0307403f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_32 VPB N_A_27_297#_c_130_n 0.00330266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_297#_c_131_n 0.00183229f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_34 VPB N_A_27_297#_c_132_n 0.00813676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_297#_c_133_n 0.0204518f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_36 VPB N_VPWR_c_164_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_37 VPB N_VPWR_c_165_n 0.015553f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_38 VPB N_VPWR_c_166_n 0.035774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_163_n 0.0455404f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_40 VPB N_VPWR_c_168_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_41 VPB N_Y_c_195_n 0.00755322f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_42 VPB N_Y_c_198_n 0.0139077f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.175
cc_43 N_A_c_44_n N_B_c_81_n 0.0195336f $X=0.91 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_44 N_A_M1007_g N_B_M1005_g 0.0195336f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_45 A B 0.0168341f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_46 N_A_c_46_n B 0.00538133f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A_c_46_n N_B_c_84_n 0.0195336f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_48 A N_A_27_297#_c_128_n 0.0225537f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_A_27_297#_c_130_n 0.0138201f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_M1007_g N_A_27_297#_c_130_n 0.0152986f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_51 A N_A_27_297#_c_130_n 0.0309573f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_52 N_A_c_46_n N_A_27_297#_c_130_n 0.00213789f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_M1000_g N_VPWR_c_164_n 0.0129691f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_54 N_A_M1007_g N_VPWR_c_164_n 0.0122146f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_55 N_A_M1000_g N_VPWR_c_165_n 0.0046653f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_56 N_A_M1007_g N_VPWR_c_166_n 0.0046653f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A_M1000_g N_VPWR_c_163_n 0.00886468f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A_M1007_g N_VPWR_c_163_n 0.007919f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_c_43_n N_Y_c_199_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A_c_44_n N_Y_c_199_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_61 N_A_c_44_n N_Y_c_192_n 0.0100722f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A_c_43_n N_Y_c_193_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A_c_44_n N_Y_c_193_n 0.00151671f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_64 A N_Y_c_193_n 0.0222065f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_c_46_n N_Y_c_193_n 0.00230339f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_44_n N_Y_c_206_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A_c_43_n N_VGND_c_252_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_68 A N_VGND_c_252_n 0.0233158f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_c_44_n N_VGND_c_253_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_c_43_n N_VGND_c_256_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_c_44_n N_VGND_c_256_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_c_43_n N_VGND_c_259_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_c_44_n N_VGND_c_259_n 0.0057435f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_74 B N_A_27_297#_c_130_n 0.00401644f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_75 N_B_M1005_g N_A_27_297#_c_131_n 2.36323e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_76 B N_A_27_297#_c_131_n 0.0139423f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_77 N_B_M1005_g N_A_27_297#_c_132_n 0.0112436f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B_M1006_g N_A_27_297#_c_132_n 0.00929492f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B_M1005_g N_VPWR_c_164_n 0.00110007f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_80 N_B_M1005_g N_VPWR_c_166_n 0.00357877f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_81 N_B_M1006_g N_VPWR_c_166_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_82 N_B_M1005_g N_VPWR_c_163_n 0.00525237f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_83 N_B_M1006_g N_VPWR_c_163_n 0.00624775f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_84 N_B_c_81_n N_Y_c_199_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B_c_81_n N_Y_c_192_n 0.00865686f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_86 B N_Y_c_192_n 0.0292573f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B_c_81_n N_Y_c_206_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B_c_82_n N_Y_c_206_n 0.0109314f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B_c_82_n N_Y_c_194_n 0.0108204f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_90 B N_Y_c_194_n 0.00305484f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_91 N_B_c_82_n N_Y_c_195_n 0.0193198f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_92 B N_Y_c_195_n 0.0160937f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B_c_81_n N_Y_c_196_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B_c_82_n N_Y_c_196_n 0.00158032f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_95 B N_Y_c_196_n 0.0265405f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B_c_84_n N_Y_c_196_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_M1005_g N_Y_c_198_n 0.00330354f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B_M1006_g N_Y_c_198_n 0.0143596f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_99 B N_Y_c_198_n 0.0273027f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_100 N_B_c_84_n N_Y_c_198_n 0.00215368f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B_M1005_g Y 0.00527894f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B_M1006_g Y 0.0111068f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B_c_81_n N_VGND_c_253_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B_c_82_n N_VGND_c_255_n 0.0032322f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_c_81_n N_VGND_c_258_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B_c_82_n N_VGND_c_258_n 0.00424416f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B_c_81_n N_VGND_c_259_n 0.0057435f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B_c_82_n N_VGND_c_259_n 0.00675866f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_27_297#_c_130_n N_VPWR_M1000_d 0.00166915f $X=1.035 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_110 N_A_27_297#_c_130_n N_VPWR_c_164_n 0.0172742f $X=1.035 $Y=1.56 $X2=0
+ $Y2=0
cc_111 N_A_27_297#_c_129_n N_VPWR_c_165_n 0.019049f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_112 N_A_27_297#_c_147_p N_VPWR_c_166_n 0.0114668f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_113 N_A_27_297#_c_132_n N_VPWR_c_166_n 0.0566987f $X=1.875 $Y=2.38 $X2=0
+ $Y2=0
cc_114 N_A_27_297#_M1000_s N_VPWR_c_163_n 0.00399293f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_115 N_A_27_297#_M1007_s N_VPWR_c_163_n 0.00385313f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_116 N_A_27_297#_M1006_d N_VPWR_c_163_n 0.00209324f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_117 N_A_27_297#_c_129_n N_VPWR_c_163_n 0.0105137f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_118 N_A_27_297#_c_147_p N_VPWR_c_163_n 0.00653655f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_119 N_A_27_297#_c_132_n N_VPWR_c_163_n 0.0349677f $X=1.875 $Y=2.38 $X2=0
+ $Y2=0
cc_120 N_A_27_297#_c_132_n N_Y_M1005_s 0.00312348f $X=1.875 $Y=2.38 $X2=0 $Y2=0
cc_121 N_A_27_297#_c_130_n N_Y_c_192_n 0.00302189f $X=1.035 $Y=1.56 $X2=0 $Y2=0
cc_122 N_A_27_297#_c_130_n N_Y_c_193_n 0.0018215f $X=1.035 $Y=1.56 $X2=0 $Y2=0
cc_123 N_A_27_297#_M1006_d N_Y_c_198_n 0.00296777f $X=1.825 $Y=1.485 $X2=0 $Y2=0
cc_124 N_A_27_297#_c_131_n N_Y_c_198_n 0.0102037f $X=1.12 $Y=1.665 $X2=0 $Y2=0
cc_125 N_A_27_297#_c_132_n N_Y_c_198_n 0.00282992f $X=1.875 $Y=2.38 $X2=0 $Y2=0
cc_126 N_A_27_297#_c_133_n N_Y_c_198_n 0.0209375f $X=1.96 $Y=2 $X2=0 $Y2=0
cc_127 N_A_27_297#_c_132_n Y 0.0154795f $X=1.875 $Y=2.38 $X2=0 $Y2=0
cc_128 N_VPWR_c_163_n N_Y_M1005_s 0.00216833f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_129 N_Y_c_192_n N_VGND_M1004_d 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_130 N_Y_c_194_n N_VGND_M1003_s 0.00287493f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_131 N_Y_c_193_n N_VGND_c_252_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_132 N_Y_c_192_n N_VGND_c_253_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_133 N_Y_c_194_n N_VGND_c_255_n 0.0207632f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_134 N_Y_c_199_n N_VGND_c_256_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_135 N_Y_c_192_n N_VGND_c_256_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_136 N_Y_c_192_n N_VGND_c_258_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_137 N_Y_c_206_n N_VGND_c_258_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_138 N_Y_c_194_n N_VGND_c_258_n 0.00193763f $X=1.92 $Y=0.82 $X2=0 $Y2=0
cc_139 N_Y_M1002_s N_VGND_c_259_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Y_M1001_d N_VGND_c_259_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_141 N_Y_c_199_n N_VGND_c_259_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_142 N_Y_c_192_n N_VGND_c_259_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_143 N_Y_c_206_n N_VGND_c_259_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_144 N_Y_c_194_n N_VGND_c_259_n 0.00492504f $X=1.92 $Y=0.82 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__fahcin_1.spice.pex
* Created: Thu Aug 27 14:21:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_67_199# 1 2 3 4 5 18 21 23 24 25 27 28 29
+ 32 33 37 42 47 51 54 55 56 57 60 64 66 67 70
c188 57 0 1.08163e-19 $X=2.8 $Y=1.87
c189 55 0 1.08972e-19 $X=2.11 $Y=1.87
c190 51 0 1.21052e-19 $X=2.1 $Y=0.36
c191 42 0 3.27481e-19 $X=0.51 $Y=1.16
r192 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.225 $Y=1.87
+ $X2=4.225 $Y2=1.87
r193 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.655 $Y=1.87
+ $X2=2.655 $Y2=1.87
r194 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.965 $Y=1.87
+ $X2=1.965 $Y2=1.87
r195 57 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.8 $Y=1.87
+ $X2=2.655 $Y2=1.87
r196 56 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.08 $Y=1.87
+ $X2=4.225 $Y2=1.87
r197 56 57 1.58416 $w=1.4e-07 $l=1.28e-06 $layer=MET1_cond $X=4.08 $Y=1.87
+ $X2=2.8 $Y2=1.87
r198 55 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.11 $Y=1.87
+ $X2=1.965 $Y2=1.87
r199 54 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.51 $Y=1.87
+ $X2=2.655 $Y2=1.87
r200 54 55 0.495049 $w=1.4e-07 $l=4e-07 $layer=MET1_cond $X=2.51 $Y=1.87
+ $X2=2.11 $Y2=1.87
r201 49 60 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.45 $Y=1.87
+ $X2=1.965 $Y2=1.87
r202 48 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=1.87
+ $X2=1.45 $Y2=1.87
r203 47 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.365 $Y=1.585
+ $X2=1.365 $Y2=1.87
r204 42 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.16
+ $X2=0.5 $Y2=1.325
r205 42 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.16
+ $X2=0.5 $Y2=0.995
r206 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r207 37 53 42.1222 $w=2.34e-07 $l=8.29036e-07 $layer=LI1_cond $X=2.515 $Y=0.34
+ $X2=3.305 $Y2=0.42
r208 37 51 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.515 $Y=0.34
+ $X2=2.1 $Y2=0.34
r209 34 44 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=0.36
+ $X2=1.16 $Y2=0.36
r210 34 36 29.5758 $w=2.08e-07 $l=5.6e-07 $layer=LI1_cond $X=1.325 $Y=0.36
+ $X2=1.885 $Y2=0.36
r211 33 51 5.98033 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=1.995 $Y=0.36
+ $X2=2.1 $Y2=0.36
r212 33 36 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=1.995 $Y=0.36
+ $X2=1.885 $Y2=0.36
r213 30 32 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.16 $Y=0.735
+ $X2=1.16 $Y2=0.72
r214 29 44 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.36
r215 29 32 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.72
r216 27 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.585
+ $X2=1.365 $Y2=1.585
r217 27 28 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.28 $Y=1.585
+ $X2=0.78 $Y2=1.585
r218 26 41 15.1941 $w=2.73e-07 $l=4.19667e-07 $layer=LI1_cond $X=0.78 $Y=0.82
+ $X2=0.602 $Y2=1.16
r219 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.995 $Y=0.82
+ $X2=1.16 $Y2=0.735
r220 25 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.995 $Y=0.82
+ $X2=0.78 $Y2=0.82
r221 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.695 $Y=1.5
+ $X2=0.78 $Y2=1.585
r222 23 41 9.1003 $w=2.73e-07 $l=2.06325e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.602 $Y2=1.16
r223 23 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.5
r224 21 71 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r225 18 70 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.475 $Y=0.555
+ $X2=0.475 $Y2=0.995
r226 5 67 600 $w=1.7e-07 $l=4.32262e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=1.61 $X2=4.28 $Y2=1.98
r227 4 64 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=1.485 $X2=2.73 $Y2=1.96
r228 3 47 600 $w=1.7e-07 $l=3.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.485 $X2=1.365 $Y2=1.665
r229 2 53 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.235 $X2=3.305 $Y2=0.42
r230 1 44 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.16 $Y2=0.38
r231 1 36 182 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.885 $Y2=0.38
r232 1 32 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.16 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A 1 3 6 8 14
c42 8 0 1.76755e-19 $X=1.15 $Y=1.19
c43 1 0 5.07203e-20 $X=0.95 $Y=0.995
r44 12 14 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=1.175 $Y2=1.16
r45 10 12 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.975 $Y2=1.16
r46 8 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.16 $X2=1.175 $Y2=1.16
r47 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.985
r49 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.995 $X2=0.95
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%B 1 3 6 10 14 15 17 20 22 23 25 26 28 29 30
+ 32 33 35 41 42
c158 42 0 1.03248e-19 $X=4.37 $Y=0.85
c159 32 0 1.85123e-19 $X=4.225 $Y=0.85
c160 25 0 5.53651e-20 $X=4.27 $Y=1.16
c161 6 0 1.08163e-19 $X=2.095 $Y=1.905
r162 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.325
+ $Y=1.16 $X2=4.325 $Y2=1.16
r163 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.16 $X2=1.655 $Y2=1.16
r164 42 50 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=4.365 $Y=0.85
+ $X2=4.365 $Y2=1.16
r165 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0.85
+ $X2=4.37 $Y2=0.85
r166 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=0.85
+ $X2=1.61 $Y2=0.85
r167 32 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=0.85
+ $X2=4.37 $Y2=0.85
r168 32 33 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=4.225 $Y=0.85
+ $X2=1.755 $Y2=0.85
r169 30 46 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.625 $Y=0.85
+ $X2=1.625 $Y2=1.16
r170 30 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0.85
+ $X2=1.61 $Y2=0.85
r171 28 49 126.774 $w=3.3e-07 $l=7.25e-07 $layer=POLY_cond $X=5.05 $Y=1.16
+ $X2=4.325 $Y2=1.16
r172 28 29 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.05 $Y=1.16
+ $X2=5.125 $Y2=1.16
r173 25 49 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.27 $Y=1.16
+ $X2=4.325 $Y2=1.16
r174 25 27 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.127 $Y=1.16
+ $X2=4.127 $Y2=1.325
r175 25 26 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.127 $Y=1.16
+ $X2=4.127 $Y2=0.995
r176 22 45 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=1.655 $Y2=1.16
r177 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=2.095 $Y2=1.16
r178 18 29 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.325
+ $X2=5.125 $Y2=1.16
r179 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.125 $Y=1.325
+ $X2=5.125 $Y2=1.985
r180 15 29 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=0.995
+ $X2=5.125 $Y2=1.16
r181 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.125 $Y=0.995
+ $X2=5.125 $Y2=0.56
r182 14 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.195 $Y=0.565
+ $X2=4.195 $Y2=0.995
r183 10 27 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=4.07 $Y=2.03
+ $X2=4.07 $Y2=1.325
r184 4 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.325
+ $X2=2.095 $Y2=1.16
r185 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.095 $Y=1.325
+ $X2=2.095 $Y2=1.905
r186 1 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.095 $Y2=1.16
r187 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.095 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_489_21# 1 2 7 9 12 14 16 19 23 26 29 30
+ 31 34 38 39 42 46 47 50 53 54 58
c158 31 0 1.03248e-19 $X=3.557 $Y=1.16
c159 14 0 4.5918e-20 $X=3.53 $Y=0.995
c160 12 0 1.08972e-19 $X=2.52 $Y=1.905
c161 7 0 1.21052e-19 $X=2.52 $Y=0.995
r162 54 62 11.1457 $w=4.05e-07 $l=3.7e-07 $layer=LI1_cond $X=4.93 $Y=1.53
+ $X2=4.93 $Y2=1.16
r163 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.845 $Y=1.53
+ $X2=4.845 $Y2=1.53
r164 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.035 $Y=1.53
+ $X2=3.035 $Y2=1.53
r165 47 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.18 $Y=1.53
+ $X2=3.035 $Y2=1.53
r166 46 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.7 $Y=1.53
+ $X2=4.845 $Y2=1.53
r167 46 47 1.88118 $w=1.4e-07 $l=1.52e-06 $layer=MET1_cond $X=4.7 $Y=1.53
+ $X2=3.18 $Y2=1.53
r168 45 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.035 $Y=1.265
+ $X2=3.035 $Y2=1.53
r169 44 45 0.961343 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.035 $Y=1.17
+ $X2=3.035 $Y2=1.265
r170 42 44 15.8531 $w=1.77e-07 $l=2.3e-07 $layer=LI1_cond $X=2.805 $Y=1.17
+ $X2=3.035 $Y2=1.17
r171 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.16 $X2=2.805 $Y2=1.16
r172 39 59 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.16
+ $X2=5.56 $Y2=1.325
r173 39 58 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.16
+ $X2=5.56 $Y2=0.995
r174 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.545
+ $Y=1.16 $X2=5.545 $Y2=1.16
r175 36 62 1.93884 $w=3.3e-07 $l=2.4e-07 $layer=LI1_cond $X=5.17 $Y=1.16
+ $X2=4.93 $Y2=1.16
r176 36 38 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.17 $Y=1.16
+ $X2=5.545 $Y2=1.16
r177 32 62 9.17697 $w=4.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.915 $Y=0.995
+ $X2=4.93 $Y2=1.16
r178 32 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.915 $Y=0.995
+ $X2=4.915 $Y2=0.74
r179 30 43 113.66 $w=3.3e-07 $l=6.5e-07 $layer=POLY_cond $X=3.455 $Y=1.16
+ $X2=2.805 $Y2=1.16
r180 30 31 5.03009 $w=3.3e-07 $l=1.02e-07 $layer=POLY_cond $X=3.455 $Y=1.16
+ $X2=3.557 $Y2=1.16
r181 28 43 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.805 $Y2=1.16
r182 28 29 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.52 $Y2=1.16
r183 26 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.635 $Y=1.985
+ $X2=5.635 $Y2=1.325
r184 23 58 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.635 $Y=0.565
+ $X2=5.635 $Y2=0.995
r185 17 31 37.0704 $w=1.5e-07 $l=1.78452e-07 $layer=POLY_cond $X=3.585 $Y=1.325
+ $X2=3.557 $Y2=1.16
r186 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.585 $Y=1.325
+ $X2=3.585 $Y2=1.905
r187 14 31 37.0704 $w=1.5e-07 $l=1.77989e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.557 $Y2=1.16
r188 14 16 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=0.555
r189 10 29 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=1.325
+ $X2=2.52 $Y2=1.16
r190 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.52 $Y=1.325
+ $X2=2.52 $Y2=1.905
r191 7 29 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=1.16
r192 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=0.565
r193 2 54 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=4.79
+ $Y=1.485 $X2=4.915 $Y2=1.64
r194 1 34 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.605 $X2=4.915 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_434_49# 1 2 9 11 13 14 16 19 21 22 25 29
+ 30 31 32 35 39 41 49 53 54
c192 54 0 1.75206e-19 $X=8.935 $Y=1.16
c193 53 0 9.22668e-20 $X=8.935 $Y=1.16
c194 49 0 2.59669e-19 $X=6.63 $Y=1.16
c195 41 0 9.13617e-20 $X=8.985 $Y=1.19
c196 11 0 1.78045e-19 $X=6.63 $Y=0.995
r197 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.935
+ $Y=1.16 $X2=8.935 $Y2=1.16
r198 48 49 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.575 $Y=1.16
+ $X2=6.63 $Y2=1.16
r199 45 48 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=6.34 $Y=1.16
+ $X2=6.575 $Y2=1.16
r200 41 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.985 $Y=1.19
+ $X2=8.985 $Y2=1.19
r201 39 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.34
+ $Y=1.16 $X2=6.34 $Y2=1.16
r202 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.225 $Y=1.19
+ $X2=6.225 $Y2=1.19
r203 35 62 8.52653 $w=4.03e-07 $l=1.6e-07 $layer=LI1_cond $X=2.187 $Y=1.19
+ $X2=2.187 $Y2=1.35
r204 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.19
r205 32 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.37 $Y=1.19
+ $X2=6.225 $Y2=1.19
r206 31 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.84 $Y=1.19
+ $X2=8.985 $Y2=1.19
r207 31 32 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=8.84 $Y=1.19
+ $X2=6.37 $Y2=1.19
r208 30 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=1.19
+ $X2=2.07 $Y2=1.19
r209 29 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=1.19
+ $X2=6.225 $Y2=1.19
r210 29 30 4.78341 $w=1.4e-07 $l=3.865e-06 $layer=MET1_cond $X=6.08 $Y=1.19
+ $X2=2.215 $Y2=1.19
r211 25 62 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.305 $Y=1.62
+ $X2=2.305 $Y2=1.35
r212 22 35 1.19513 $w=4.03e-07 $l=4.2e-08 $layer=LI1_cond $X=2.187 $Y=1.148
+ $X2=2.187 $Y2=1.19
r213 21 28 3.89425 $w=4.05e-07 $l=1.17e-07 $layer=LI1_cond $X=2.187 $Y=0.877
+ $X2=2.187 $Y2=0.76
r214 21 22 7.71141 $w=4.03e-07 $l=2.71e-07 $layer=LI1_cond $X=2.187 $Y=0.877
+ $X2=2.187 $Y2=1.148
r215 19 53 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.935 $Y=1.995
+ $X2=8.935 $Y2=1.325
r216 14 53 63.3216 $w=2.55e-07 $l=4.45331e-07 $layer=POLY_cond $X=8.6 $Y=0.96
+ $X2=8.935 $Y2=1.217
r217 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.6 $Y=0.96
+ $X2=8.6 $Y2=0.565
r218 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.16
r219 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.565
r220 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.575 $Y=1.325
+ $X2=6.575 $Y2=1.16
r221 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.575 $Y=1.325
+ $X2=6.575 $Y2=1.905
r222 2 25 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.17
+ $Y=1.485 $X2=2.305 $Y2=1.62
r223 1 28 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.245 $X2=2.305 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_721_47# 1 2 9 11 13 16 17 19 21 23 25 26
+ 32 33 34 37 40 41 42 44 45 46 48 51 56 59
c190 51 0 9.22668e-20 $X=7.95 $Y=1.16
c191 32 0 5.53651e-20 $X=3.795 $Y=1.99
c192 17 0 2.15715e-19 $X=8.44 $Y=1.425
c193 9 0 1.73441e-19 $X=6.995 $Y=1.905
r194 58 59 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=7.907 $Y=1.55
+ $X2=7.907 $Y2=1.72
r195 54 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.795 $Y=1.235
+ $X2=3.985 $Y2=1.235
r196 51 58 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.95 $Y=1.16
+ $X2=7.95 $Y2=1.55
r197 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.95
+ $Y=1.16 $X2=7.95 $Y2=1.16
r198 48 59 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.865 $Y=2.295
+ $X2=7.865 $Y2=1.72
r199 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.78 $Y=2.38
+ $X2=7.865 $Y2=2.295
r200 45 46 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=7.78 $Y=2.38
+ $X2=5.995 $Y2=2.38
r201 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.91 $Y=2.295
+ $X2=5.995 $Y2=2.38
r202 43 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.91 $Y=2.065
+ $X2=5.91 $Y2=2.295
r203 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.825 $Y=1.98
+ $X2=5.91 $Y2=2.065
r204 41 42 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.825 $Y=1.98
+ $X2=5.065 $Y2=1.98
r205 39 42 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.94 $Y=2.065
+ $X2=5.065 $Y2=1.98
r206 39 40 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=4.94 $Y=2.065
+ $X2=4.94 $Y2=2.29
r207 35 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=1.15
+ $X2=3.985 $Y2=1.235
r208 35 37 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.985 $Y=1.15
+ $X2=3.985 $Y2=0.76
r209 33 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.815 $Y=2.375
+ $X2=4.94 $Y2=2.29
r210 33 34 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=4.815 $Y=2.375 $X2=3.88
+ $Y2=2.375
r211 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.795 $Y=2.29
+ $X2=3.88 $Y2=2.375
r212 30 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.795 $Y=2.29
+ $X2=3.795 $Y2=1.99
r213 29 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=1.32
+ $X2=3.795 $Y2=1.235
r214 29 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.795 $Y=1.32
+ $X2=3.795 $Y2=1.99
r215 25 52 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=7.995 $Y=1.16
+ $X2=7.95 $Y2=1.16
r216 25 27 68.5835 $w=2.4e-07 $l=2.65e-07 $layer=POLY_cond $X=8.115 $Y=1.16
+ $X2=8.115 $Y2=1.425
r217 25 26 51.39 $w=2.4e-07 $l=1.65e-07 $layer=POLY_cond $X=8.115 $Y=1.16
+ $X2=8.115 $Y2=0.995
r218 22 52 143.386 $w=3.3e-07 $l=8.2e-07 $layer=POLY_cond $X=7.13 $Y=1.16
+ $X2=7.95 $Y2=1.16
r219 22 23 5.03009 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=7.13 $Y=1.16
+ $X2=7.025 $Y2=1.16
r220 19 21 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.515 $Y=1.5
+ $X2=8.515 $Y2=1.995
r221 18 27 13.7767 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=8.235 $Y=1.425
+ $X2=8.115 $Y2=1.425
r222 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.44 $Y=1.425
+ $X2=8.515 $Y2=1.5
r223 17 18 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=8.44 $Y=1.425
+ $X2=8.235 $Y2=1.425
r224 16 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.16 $Y=0.565
+ $X2=8.16 $Y2=0.995
r225 11 23 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=7.055 $Y=0.995
+ $X2=7.025 $Y2=1.16
r226 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.055 $Y=0.995
+ $X2=7.055 $Y2=0.565
r227 7 23 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=6.995 $Y=1.325
+ $X2=7.025 $Y2=1.16
r228 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.995 $Y=1.325
+ $X2=6.995 $Y2=1.905
r229 2 32 600 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.485 $X2=3.795 $Y2=1.99
r230 1 37 182 $w=1.7e-07 $l=6.89293e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.235 $X2=3.985 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_1636_315# 1 2 3 4 15 18 22 24 25 26 31 33
+ 34 36 40 42 44 46 50 55
c124 50 0 2.4093e-19 $X=10.065 $Y=1.16
c125 22 0 1.01924e-19 $X=8.305 $Y=2.12
r126 52 53 8.54777 $w=4.71e-07 $l=3.3e-07 $layer=LI1_cond $X=10.617 $Y=1.63
+ $X2=10.617 $Y2=1.96
r127 50 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.065 $Y=1.16
+ $X2=10.065 $Y2=0.995
r128 49 52 12.1741 $w=4.71e-07 $l=7.51095e-07 $layer=LI1_cond $X=10.065 $Y=1.16
+ $X2=10.617 $Y2=1.63
r129 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.065
+ $Y=1.16 $X2=10.065 $Y2=1.16
r130 42 53 2.5146 $w=4.71e-07 $l=1.21219e-07 $layer=LI1_cond $X=10.71 $Y=2.025
+ $X2=10.617 $Y2=1.96
r131 42 44 9.38418 $w=3.48e-07 $l=2.85e-07 $layer=LI1_cond $X=10.71 $Y=2.025
+ $X2=10.71 $Y2=2.31
r132 38 40 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.72 $Y=0.735
+ $X2=10.72 $Y2=0.4
r133 37 49 8.80679 $w=4.71e-07 $l=4.60977e-07 $layer=LI1_cond $X=10.35 $Y=0.82
+ $X2=10.065 $Y2=1.16
r134 36 38 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=10.53 $Y=0.82
+ $X2=10.72 $Y2=0.735
r135 36 37 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.53 $Y=0.82
+ $X2=10.35 $Y2=0.82
r136 35 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.41 $Y=1.96
+ $X2=9.325 $Y2=1.96
r137 34 53 6.78321 $w=1.7e-07 $l=5.62e-07 $layer=LI1_cond $X=10.055 $Y=1.96
+ $X2=10.617 $Y2=1.96
r138 34 35 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=10.055 $Y=1.96
+ $X2=9.41 $Y2=1.96
r139 32 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=2.045
+ $X2=9.325 $Y2=1.96
r140 32 33 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=9.325 $Y=2.045
+ $X2=9.325 $Y2=2.295
r141 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=1.875
+ $X2=9.325 $Y2=1.96
r142 30 31 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=9.325 $Y=0.765
+ $X2=9.325 $Y2=1.875
r143 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.24 $Y=0.68
+ $X2=9.325 $Y2=0.765
r144 26 28 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=9.24 $Y=0.68
+ $X2=9.23 $Y2=0.68
r145 24 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.24 $Y=2.38
+ $X2=9.325 $Y2=2.295
r146 24 25 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=9.24 $Y=2.38
+ $X2=8.39 $Y2=2.38
r147 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.305 $Y=2.295
+ $X2=8.39 $Y2=2.38
r148 20 22 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.305 $Y=2.295
+ $X2=8.305 $Y2=2.12
r149 16 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.065 $Y=1.325
+ $X2=10.065 $Y2=1.16
r150 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.065 $Y=1.325
+ $X2=10.065 $Y2=1.985
r151 15 55 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.035 $Y=0.565
+ $X2=10.035 $Y2=0.995
r152 4 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.56
+ $Y=1.485 $X2=10.7 $Y2=1.63
r153 4 44 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=10.56
+ $Y=1.485 $X2=10.7 $Y2=2.31
r154 3 22 600 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_PDIFF $count=1 $X=8.18
+ $Y=1.575 $X2=8.305 $Y2=2.12
r155 2 40 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=10.585
+ $Y=0.235 $X2=10.72 $Y2=0.4
r156 1 28 91 $w=1.7e-07 $l=7.41249e-07 $layer=licon1_NDIFF $count=2 $X=8.675
+ $Y=0.245 $X2=9.23 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%CIN 3 5 7 8 10 13 16 17 18 19
c66 19 0 1.5713e-19 $X=10.825 $Y=1.19
c67 5 0 8.32754e-20 $X=10.51 $Y=0.995
c68 3 0 1.46815e-19 $X=10.485 $Y=1.985
r69 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.765
+ $Y=1.16 $X2=10.765 $Y2=1.16
r70 17 22 106.665 $w=3.3e-07 $l=6.1e-07 $layer=POLY_cond $X=11.375 $Y=1.16
+ $X2=10.765 $Y2=1.16
r71 17 18 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.375 $Y=1.16
+ $X2=11.45 $Y2=1.16
r72 15 22 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=10.585 $Y=1.16
+ $X2=10.765 $Y2=1.16
r73 15 16 5.03009 $w=3.3e-07 $l=8.8e-08 $layer=POLY_cond $X=10.585 $Y=1.16
+ $X2=10.497 $Y2=1.16
r74 11 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.45 $Y=1.325
+ $X2=11.45 $Y2=1.16
r75 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.45 $Y=1.325
+ $X2=11.45 $Y2=1.985
r76 8 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.45 $Y=0.995
+ $X2=11.45 $Y2=1.16
r77 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.45 $Y=0.995
+ $X2=11.45 $Y2=0.565
r78 5 16 37.0704 $w=1.5e-07 $l=1.71377e-07 $layer=POLY_cond $X=10.51 $Y=0.995
+ $X2=10.497 $Y2=1.16
r79 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.51 $Y=0.995
+ $X2=10.51 $Y2=0.56
r80 1 16 37.0704 $w=1.5e-07 $l=1.70895e-07 $layer=POLY_cond $X=10.485 $Y=1.325
+ $X2=10.497 $Y2=1.16
r81 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.485 $Y=1.325
+ $X2=10.485 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_1647_49# 1 2 9 13 15 19 22 23 29 33 34 35
+ 42
c106 42 0 9.13617e-20 $X=8.725 $Y=1.7
c107 33 0 1.52424e-19 $X=11.87 $Y=1.16
c108 23 0 2.20632e-19 $X=8.67 $Y=1.53
r109 33 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.87 $Y=1.16
+ $X2=11.87 $Y2=0.995
r110 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.87
+ $Y=1.16 $X2=11.87 $Y2=1.16
r111 30 34 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=11.8 $Y=1.53
+ $X2=11.8 $Y2=1.16
r112 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.765 $Y=1.53
+ $X2=11.765 $Y2=1.53
r113 26 42 10.4686 $w=3.03e-07 $l=2.6e-07 $layer=LI1_cond $X=8.465 $Y=1.615
+ $X2=8.725 $Y2=1.615
r114 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.525 $Y=1.53
+ $X2=8.525 $Y2=1.53
r115 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.67 $Y=1.53
+ $X2=8.525 $Y2=1.53
r116 22 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.62 $Y=1.53
+ $X2=11.765 $Y2=1.53
r117 22 23 3.65098 $w=1.4e-07 $l=2.95e-06 $layer=MET1_cond $X=11.62 $Y=1.53
+ $X2=8.67 $Y2=1.53
r118 19 21 8.52828 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.43 $Y=0.76
+ $X2=8.43 $Y2=0.925
r119 15 26 3.784 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=8.465 $Y=1.445
+ $X2=8.465 $Y2=1.615
r120 15 21 32.0404 $w=1.78e-07 $l=5.2e-07 $layer=LI1_cond $X=8.465 $Y=1.445
+ $X2=8.465 $Y2=0.925
r121 13 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.925 $Y=0.56
+ $X2=11.925 $Y2=0.995
r122 7 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.87 $Y=1.325
+ $X2=11.87 $Y2=1.16
r123 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.87 $Y=1.325
+ $X2=11.87 $Y2=1.985
r124 2 42 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=8.59
+ $Y=1.575 $X2=8.725 $Y2=1.7
r125 1 19 182 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_NDIFF $count=1 $X=8.235
+ $Y=0.245 $X2=8.39 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_27_47# 1 2 3 4 5 6 23 27 29 32 34 35 37
+ 44 46 48 50 52 53 58 59 60 63 65 66
c167 65 0 4.5918e-20 $X=4.405 $Y=0.39
c168 52 0 1.3431e-19 $X=0.265 $Y=1.63
c169 50 0 5.07203e-20 $X=0.257 $Y=0.805
c170 2 0 1.85123e-19 $X=2.595 $Y=0.245
r171 65 66 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=0.365
+ $X2=4.24 $Y2=0.365
r172 57 59 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=2.34
+ $X2=1.97 $Y2=2.34
r173 57 58 5.33595 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.805 $Y=2.34
+ $X2=1.715 $Y2=2.34
r174 54 55 2.75937 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=0.262 $Y=1.925
+ $X2=0.262 $Y2=2.01
r175 52 54 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=1.63
+ $X2=0.262 $Y2=1.925
r176 52 53 7.36284 $w=3.53e-07 $l=1.3e-07 $layer=LI1_cond $X=0.262 $Y=1.63
+ $X2=0.262 $Y2=1.5
r177 50 53 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.17 $Y=0.805
+ $X2=0.17 $Y2=1.5
r178 49 50 5.14454 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.805
r179 48 66 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.73 $Y=0.34
+ $X2=4.24 $Y2=0.34
r180 46 60 18 $w=1.83e-07 $l=2.7e-07 $layer=LI1_cond $X=3.645 $Y=0.79 $X2=3.375
+ $Y2=0.79
r181 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.645 $Y=0.425
+ $X2=3.73 $Y2=0.34
r182 45 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.645 $Y=0.425
+ $X2=3.645 $Y2=0.755
r183 42 63 14.7424 $w=2.41e-07 $l=2.72489e-07 $layer=LI1_cond $X=3.375 $Y=2.11
+ $X2=3.38 $Y2=2.38
r184 42 44 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.375 $Y=2.11
+ $X2=3.375 $Y2=1.62
r185 41 60 1.16186 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.375 $Y=0.925
+ $X2=3.375 $Y2=0.79
r186 41 44 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.375 $Y=0.925
+ $X2=3.375 $Y2=1.62
r187 37 60 24.0793 $w=2.5e-07 $l=4.79974e-07 $layer=LI1_cond $X=2.9 $Y=0.78
+ $X2=3.375 $Y2=0.79
r188 37 39 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.9 $Y=0.78
+ $X2=2.785 $Y2=0.78
r189 35 63 2.78154 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=3.38 $Y2=2.38
r190 35 59 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=1.97 $Y2=2.38
r191 34 58 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.11 $Y=2.3
+ $X2=1.715 $Y2=2.3
r192 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.025 $Y=2.215
+ $X2=1.11 $Y2=2.3
r193 31 32 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.025 $Y=2.01
+ $X2=1.025 $Y2=2.215
r194 30 54 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.44 $Y=1.925
+ $X2=0.262 $Y2=1.925
r195 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.94 $Y=1.925
+ $X2=1.025 $Y2=2.01
r196 29 30 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.94 $Y=1.925
+ $X2=0.44 $Y2=1.925
r197 27 49 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.265 $Y=0.38
+ $X2=0.265 $Y2=0.735
r198 23 55 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=0.257 $Y=2.31
+ $X2=0.257 $Y2=2.01
r199 6 63 600 $w=1.7e-07 $l=9.55458e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.29 $Y2=2.38
r200 6 44 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.375 $Y2=1.62
r201 5 57 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=2.155 $X2=1.805 $Y2=2.3
r202 4 52 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=1.63
r203 4 23 400 $w=1.7e-07 $l=8.87623e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=2.31
r204 3 65 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.245 $X2=4.405 $Y2=0.39
r205 2 39 182 $w=1.7e-07 $l=5.82301e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.245 $X2=2.785 $Y2=0.74
r206 1 27 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%VPWR 1 2 3 4 15 17 21 25 29 31 33 38 46 53
+ 54 57 60 63 66
c128 33 0 1.3431e-19 $X=0.6 $Y=2.72
c129 29 0 1.52424e-19 $X=11.66 $Y=1.95
r130 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r131 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r132 60 61 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 58 61 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 57 58 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 54 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r136 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r137 51 66 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=11.83 $Y=2.72
+ $X2=11.702 $Y2=2.72
r138 51 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.83 $Y=2.72
+ $X2=12.19 $Y2=2.72
r139 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r140 50 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=10.35 $Y2=2.72
r141 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r142 47 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=2.72
+ $X2=10.275 $Y2=2.72
r143 47 49 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=10.36 $Y=2.72
+ $X2=11.27 $Y2=2.72
r144 46 66 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.575 $Y=2.72
+ $X2=11.702 $Y2=2.72
r145 46 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.575 $Y=2.72
+ $X2=11.27 $Y2=2.72
r146 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r147 44 45 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r148 42 45 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=9.89 $Y2=2.72
r149 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r150 41 44 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=9.89 $Y2=2.72
r151 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r152 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=2.72
+ $X2=5.425 $Y2=2.72
r153 39 41 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.59 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 38 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.19 $Y=2.72
+ $X2=10.275 $Y2=2.72
r155 38 44 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.19 $Y=2.72
+ $X2=9.89 $Y2=2.72
r156 33 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.685 $Y2=2.72
r157 33 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r158 31 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r159 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r160 27 66 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.702 $Y=2.635
+ $X2=11.702 $Y2=2.72
r161 27 29 30.9578 $w=2.53e-07 $l=6.85e-07 $layer=LI1_cond $X=11.702 $Y=2.635
+ $X2=11.702 $Y2=1.95
r162 23 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=2.635
+ $X2=10.275 $Y2=2.72
r163 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.275 $Y=2.635
+ $X2=10.275 $Y2=2.36
r164 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=2.635
+ $X2=5.425 $Y2=2.72
r165 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.425 $Y=2.635
+ $X2=5.425 $Y2=2.32
r166 18 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=2.72
+ $X2=0.685 $Y2=2.72
r167 17 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=2.72
+ $X2=5.425 $Y2=2.72
r168 17 18 292.93 $w=1.68e-07 $l=4.49e-06 $layer=LI1_cond $X=5.26 $Y=2.72
+ $X2=0.77 $Y2=2.72
r169 13 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.72
r170 13 15 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.345
r171 4 29 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=11.525
+ $Y=1.485 $X2=11.66 $Y2=1.95
r172 3 25 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.485 $X2=10.275 $Y2=2.36
r173 2 21 600 $w=1.7e-07 $l=9.40798e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.485 $X2=5.425 $Y2=2.32
r174 1 15 600 $w=1.7e-07 $l=9.25041e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.685 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_1142_49# 1 2 3 11 12 15 16 18 19 23 29
c72 29 0 1.73441e-19 $X=6.53 $Y=2.01
c73 19 0 8.41027e-20 $X=7.125 $Y=1.955
c74 18 0 3.53612e-19 $X=7.125 $Y=1.23
r75 28 29 13.0837 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.285 $Y=2.01
+ $X2=6.53 $Y2=2.01
r76 23 25 11.2956 $w=2.88e-07 $l=2.35e-07 $layer=LI1_cond $X=5.825 $Y=0.58
+ $X2=5.825 $Y2=0.815
r77 18 31 26.0563 $w=2.27e-07 $l=5.03786e-07 $layer=LI1_cond $X=7.125 $Y=1.23
+ $X2=7.195 $Y2=0.76
r78 18 19 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.125 $Y=1.23
+ $X2=7.125 $Y2=1.955
r79 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=2.04
+ $X2=7.125 $Y2=1.955
r80 16 29 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.04 $Y=2.04
+ $X2=6.53 $Y2=2.04
r81 15 28 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.285 $Y=1.895
+ $X2=6.285 $Y2=2.01
r82 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.285 $Y=1.725
+ $X2=6.285 $Y2=1.895
r83 13 21 3.40825 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.97 $Y=1.64
+ $X2=5.802 $Y2=1.64
r84 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.2 $Y=1.64
+ $X2=6.285 $Y2=1.725
r85 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.2 $Y=1.64 $X2=5.97
+ $Y2=1.64
r86 11 21 3.40825 $w=1.7e-07 $l=1.19499e-07 $layer=LI1_cond $X=5.885 $Y=1.555
+ $X2=5.802 $Y2=1.64
r87 11 25 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.885 $Y=1.555
+ $X2=5.885 $Y2=0.815
r88 3 28 600 $w=1.7e-07 $l=8.679e-07 $layer=licon1_PDIFF $count=1 $X=5.71
+ $Y=1.485 $X2=6.365 $Y2=1.98
r89 3 21 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.71
+ $Y=1.485 $X2=5.845 $Y2=1.64
r90 2 31 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.245 $X2=7.265 $Y2=0.76
r91 1 23 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=5.71
+ $Y=0.245 $X2=5.845 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%COUT 1 2 7 8 13 18
r28 14 18 0.426831 $w=2.68e-07 $l=1e-08 $layer=LI1_cond $X=6.735 $Y=1.54
+ $X2=6.735 $Y2=1.53
r29 8 24 2.33156 $w=2.25e-07 $l=4.3e-08 $layer=LI1_cond $X=6.735 $Y=1.577
+ $X2=6.735 $Y2=1.62
r30 8 14 2.0467 $w=2.7e-07 $l=3.7e-08 $layer=LI1_cond $X=6.735 $Y=1.577
+ $X2=6.735 $Y2=1.54
r31 8 18 1.62196 $w=2.68e-07 $l=3.8e-08 $layer=LI1_cond $X=6.735 $Y=1.492
+ $X2=6.735 $Y2=1.53
r32 7 13 3.70924 $w=2.7e-07 $l=9.25203e-08 $layer=LI1_cond $X=6.762 $Y=0.845
+ $X2=6.735 $Y2=0.925
r33 7 20 4.16466 $w=2.49e-07 $l=8.5e-08 $layer=LI1_cond $X=6.762 $Y=0.845
+ $X2=6.762 $Y2=0.76
r34 7 8 23.9879 $w=2.68e-07 $l=5.62e-07 $layer=LI1_cond $X=6.735 $Y=0.93
+ $X2=6.735 $Y2=1.492
r35 7 13 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=6.735 $Y=0.93
+ $X2=6.735 $Y2=0.925
r36 2 24 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.65
+ $Y=1.485 $X2=6.785 $Y2=1.62
r37 1 20 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=6.705
+ $Y=0.245 $X2=6.84 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_1251_49# 1 2 3 4 13 17 19 21 27 29 34 38
+ 40 41 44 47 48
c134 41 0 1.52145e-19 $X=7.75 $Y=0.85
r135 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.305 $Y=0.85
+ $X2=11.305 $Y2=0.85
r136 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.605 $Y=0.85
+ $X2=7.605 $Y2=0.85
r137 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.75 $Y=0.85
+ $X2=7.605 $Y2=0.85
r138 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.16 $Y=0.85
+ $X2=11.305 $Y2=0.85
r139 40 41 4.22029 $w=1.4e-07 $l=3.41e-06 $layer=MET1_cond $X=11.16 $Y=0.85
+ $X2=7.75 $Y2=0.85
r140 38 48 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=11.28 $Y=0.805
+ $X2=11.28 $Y2=0.85
r141 38 39 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.28 $Y=0.805
+ $X2=11.28 $Y2=0.68
r142 37 48 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=11.28 $Y=1.455
+ $X2=11.28 $Y2=0.85
r143 35 44 26.9351 $w=1.73e-07 $l=4.25e-07 $layer=LI1_cond $X=7.607 $Y=0.425
+ $X2=7.607 $Y2=0.85
r144 34 44 16.161 $w=1.73e-07 $l=2.55e-07 $layer=LI1_cond $X=7.607 $Y=1.105
+ $X2=7.607 $Y2=0.85
r145 29 32 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.42 $Y=0.34
+ $X2=6.42 $Y2=0.485
r146 27 39 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=11.24 $Y=0.55
+ $X2=11.24 $Y2=0.68
r147 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.24 $Y=1.635
+ $X2=11.24 $Y2=2.315
r148 19 37 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.24 $Y=1.62
+ $X2=11.24 $Y2=1.455
r149 19 21 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.24 $Y=1.62
+ $X2=11.24 $Y2=1.635
r150 15 34 22.5435 $w=2.3e-07 $l=4.90892e-07 $layer=LI1_cond $X=7.465 $Y=1.53
+ $X2=7.607 $Y2=1.105
r151 15 17 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.465 $Y=1.53
+ $X2=7.465 $Y2=1.62
r152 14 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=0.34
+ $X2=6.42 $Y2=0.34
r153 13 35 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=7.52 $Y=0.34
+ $X2=7.607 $Y2=0.425
r154 13 14 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=7.52 $Y=0.34 $X2=6.585
+ $Y2=0.34
r155 4 23 400 $w=1.7e-07 $l=8.90309e-07 $layer=licon1_PDIFF $count=1 $X=11.115
+ $Y=1.485 $X2=11.24 $Y2=2.315
r156 4 21 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=11.115
+ $Y=1.485 $X2=11.24 $Y2=1.635
r157 3 17 300 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=2 $X=7.07
+ $Y=1.485 $X2=7.465 $Y2=1.62
r158 2 27 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=11.115
+ $Y=0.245 $X2=11.24 $Y2=0.55
r159 1 32 182 $w=1.7e-07 $l=3.11769e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.245 $X2=6.42 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%A_1565_49# 1 2 3 12 14 15 16 17 19 22 26
c58 26 0 1.46815e-19 $X=9.845 $Y=1.62
c59 22 0 8.32754e-20 $X=9.81 $Y=0.825
c60 12 0 1.52145e-19 $X=7.95 $Y=0.525
r61 23 26 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=9.725 $Y=1.62
+ $X2=9.845 $Y2=1.62
r62 19 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.725 $Y=1.535
+ $X2=9.725 $Y2=1.62
r63 19 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=9.725 $Y=1.535
+ $X2=9.725 $Y2=0.825
r64 17 22 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=9.81 $Y=0.655
+ $X2=9.81 $Y2=0.825
r65 16 21 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=0.425
+ $X2=9.81 $Y2=0.34
r66 16 17 7.79594 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=9.81 $Y=0.425
+ $X2=9.81 $Y2=0.655
r67 14 21 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.64 $Y=0.34 $X2=9.81
+ $Y2=0.34
r68 14 15 104.711 $w=1.68e-07 $l=1.605e-06 $layer=LI1_cond $X=9.64 $Y=0.34
+ $X2=8.035 $Y2=0.34
r69 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.95 $Y=0.425
+ $X2=8.035 $Y2=0.34
r70 10 12 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=7.95 $Y=0.425 $X2=7.95
+ $Y2=0.525
r71 3 26 600 $w=1.7e-07 $l=8.57205e-07 $layer=licon1_PDIFF $count=1 $X=9.01
+ $Y=1.575 $X2=9.845 $Y2=1.62
r72 2 21 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=9.69
+ $Y=0.245 $X2=9.815 $Y2=0.4
r73 1 12 182 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_NDIFF $count=1 $X=7.825
+ $Y=0.245 $X2=7.95 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%SUM 1 2 7 8 9 10 11 12 24
r19 12 37 8.60032 $w=3.33e-07 $l=2.5e-07 $layer=LI1_cond $X=12.167 $Y=2.21
+ $X2=12.167 $Y2=1.96
r20 11 34 2.88971 $w=3.33e-07 $l=8.4e-08 $layer=LI1_cond $X=12.167 $Y=1.868
+ $X2=12.167 $Y2=1.952
r21 11 37 0.240809 $w=3.33e-07 $l=7e-09 $layer=LI1_cond $X=12.167 $Y=1.953
+ $X2=12.167 $Y2=1.96
r22 11 34 0.0344013 $w=3.33e-07 $l=1e-09 $layer=LI1_cond $X=12.167 $Y=1.953
+ $X2=12.167 $Y2=1.952
r23 10 11 10.0225 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=12.23 $Y=1.53
+ $X2=12.23 $Y2=1.785
r24 9 10 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=12.23 $Y=1.19
+ $X2=12.23 $Y2=1.53
r25 8 41 2.69103 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=12.165 $Y=0.795
+ $X2=12.165 $Y2=0.825
r26 8 22 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=12.165 $Y=0.795
+ $X2=12.165 $Y2=0.655
r27 8 9 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=12.23 $Y=0.88
+ $X2=12.23 $Y2=1.19
r28 8 41 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=12.23 $Y=0.88
+ $X2=12.23 $Y2=0.825
r29 7 22 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=12.165 $Y=0.51
+ $X2=12.165 $Y2=0.655
r30 7 24 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=12.165 $Y=0.51
+ $X2=12.165 $Y2=0.39
r31 2 37 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=11.945
+ $Y=1.485 $X2=12.085 $Y2=1.96
r32 1 24 91 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=2 $X=12
+ $Y=0.235 $X2=12.16 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCIN_1%VGND 1 2 3 4 17 21 25 29 32 33 34 36 51 60
+ 61 64 67 70
c134 25 0 8.37993e-20 $X=10.265 $Y=0.4
c135 17 0 1.50726e-19 $X=0.715 $Y=0.38
r136 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r137 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r138 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r139 61 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r140 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r141 58 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=11.66 $Y2=0
r142 58 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=12.19 $Y2=0
r143 57 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r144 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r145 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r146 53 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r147 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r148 51 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.495 $Y=0
+ $X2=11.66 $Y2=0
r149 51 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.495 $Y=0
+ $X2=11.27 $Y2=0
r150 50 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r151 49 50 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r152 47 50 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=9.89
+ $Y2=0
r153 47 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r154 46 49 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=9.89
+ $Y2=0
r155 46 47 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r156 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=0 $X2=5.345
+ $Y2=0
r157 44 46 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.51 $Y=0 $X2=5.75
+ $Y2=0
r158 43 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r159 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r160 40 43 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r161 40 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r162 39 42 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r163 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r164 37 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.715
+ $Y2=0
r165 37 39 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=1.15
+ $Y2=0
r166 36 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.18 $Y=0 $X2=5.345
+ $Y2=0
r167 36 42 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.18 $Y=0 $X2=4.83
+ $Y2=0
r168 34 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r169 33 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=0
+ $X2=10.35 $Y2=0
r170 32 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.18 $Y=0 $X2=9.89
+ $Y2=0
r171 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.18 $Y=0
+ $X2=10.265 $Y2=0
r172 27 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.66 $Y=0.085
+ $X2=11.66 $Y2=0
r173 27 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=11.66 $Y=0.085
+ $X2=11.66 $Y2=0.39
r174 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=0.085
+ $X2=10.265 $Y2=0
r175 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.265 $Y=0.085
+ $X2=10.265 $Y2=0.4
r176 19 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=0.085
+ $X2=5.345 $Y2=0
r177 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.345 $Y=0.085
+ $X2=5.345 $Y2=0.38
r178 15 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r179 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.38
r180 4 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=11.525
+ $Y=0.245 $X2=11.66 $Y2=0.39
r181 3 25 182 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_NDIFF $count=1 $X=10.11
+ $Y=0.245 $X2=10.265 $Y2=0.4
r182 2 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.2
+ $Y=0.235 $X2=5.345 $Y2=0.38
r183 1 17 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.715 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__nand3_1.pxi.spice
* Created: Thu Aug 27 14:29:25 2020
* 
x_PM_SKY130_FD_SC_HD__NAND3_1%C N_C_c_36_n N_C_M1004_g N_C_M1002_g C C
+ N_C_c_38_n PM_SKY130_FD_SC_HD__NAND3_1%C
x_PM_SKY130_FD_SC_HD__NAND3_1%B N_B_M1001_g N_B_M1000_g B B N_B_c_66_n
+ N_B_c_67_n PM_SKY130_FD_SC_HD__NAND3_1%B
x_PM_SKY130_FD_SC_HD__NAND3_1%A N_A_c_99_n N_A_M1003_g N_A_M1005_g A N_A_c_101_n
+ PM_SKY130_FD_SC_HD__NAND3_1%A
x_PM_SKY130_FD_SC_HD__NAND3_1%VPWR N_VPWR_M1002_s N_VPWR_M1000_d N_VPWR_c_127_n
+ N_VPWR_c_128_n N_VPWR_c_129_n VPWR N_VPWR_c_130_n N_VPWR_c_131_n
+ N_VPWR_c_126_n N_VPWR_c_133_n PM_SKY130_FD_SC_HD__NAND3_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND3_1%Y N_Y_M1003_d N_Y_M1002_d N_Y_M1005_d N_Y_c_158_n
+ N_Y_c_166_n N_Y_c_155_n N_Y_c_156_n N_Y_c_153_n N_Y_c_163_n N_Y_c_154_n
+ N_Y_c_174_n Y PM_SKY130_FD_SC_HD__NAND3_1%Y
x_PM_SKY130_FD_SC_HD__NAND3_1%VGND N_VGND_M1004_s N_VGND_c_206_n N_VGND_c_207_n
+ VGND N_VGND_c_208_n N_VGND_c_209_n PM_SKY130_FD_SC_HD__NAND3_1%VGND
cc_1 VNB N_C_c_36_n 0.0187646f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB C 0.00979336f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_C_c_38_n 0.0438544f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB B 0.0030191f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB N_B_c_66_n 0.0212911f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_B_c_67_n 0.0163546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_c_99_n 0.0227168f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB A 0.0123479f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_9 VNB N_A_c_101_n 0.0328917f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_10 VNB N_VPWR_c_126_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_153_n 0.00247565f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.16
cc_12 VNB N_Y_c_154_n 0.0227006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_206_n 0.00994635f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_14 VNB N_VGND_c_207_n 0.0188538f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_VGND_c_208_n 0.0377585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_209_n 0.123172f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_17 VPB N_C_M1002_g 0.02537f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_18 VPB C 0.00203753f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_19 VPB N_C_c_38_n 0.0114289f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_20 VPB N_B_M1000_g 0.0197775f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_21 VPB B 0.00268241f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_22 VPB N_B_c_66_n 0.00457342f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_23 VPB N_A_M1005_g 0.0269648f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_24 VPB A 0.00158602f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_25 VPB N_A_c_101_n 0.00763104f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_26 VPB N_VPWR_c_127_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_128_n 0.0428281f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_28 VPB N_VPWR_c_129_n 0.00444361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_130_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_131_n 0.0178658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_126_n 0.0431957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_133_n 0.00439144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_Y_c_155_n 0.00752809f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_34 VPB N_Y_c_156_n 0.0312141f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=0.85
cc_35 VPB N_Y_c_153_n 0.00161876f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_36 N_C_M1002_g N_B_M1000_g 0.0229352f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_37 N_C_c_36_n B 5.08642e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_38 N_C_c_38_n N_B_c_66_n 0.0229352f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_39 N_C_c_36_n N_B_c_67_n 0.0229352f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_40 N_C_M1002_g N_VPWR_c_128_n 0.00321527f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_41 C N_VPWR_c_128_n 0.0188755f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_42 N_C_c_38_n N_VPWR_c_128_n 0.00224688f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_43 N_C_M1002_g N_VPWR_c_130_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_44 N_C_M1002_g N_VPWR_c_126_n 0.0104829f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_45 N_C_M1002_g N_Y_c_158_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_46 N_C_c_36_n N_Y_c_153_n 0.0118209f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_47 N_C_M1002_g N_Y_c_153_n 0.00802306f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_48 C N_Y_c_153_n 0.0383894f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_49 N_C_c_38_n N_Y_c_153_n 0.00799491f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_50 N_C_M1002_g N_Y_c_163_n 0.00187637f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_51 N_C_c_36_n Y 0.00861576f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_52 C N_VGND_M1004_s 0.00402836f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_53 N_C_c_36_n N_VGND_c_207_n 0.00450113f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_54 C N_VGND_c_207_n 0.0188142f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_55 N_C_c_38_n N_VGND_c_207_n 0.00137795f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_56 N_C_c_36_n N_VGND_c_208_n 0.00539841f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_57 N_C_c_36_n N_VGND_c_209_n 0.0104859f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_58 C N_VGND_c_209_n 8.97811e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_59 B N_A_c_99_n 0.00635825f $X=1.07 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_60 N_B_c_67_n N_A_c_99_n 0.0318469f $X=0.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_61 N_B_M1000_g N_A_M1005_g 0.0230065f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_62 B A 0.022784f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_63 N_B_c_66_n A 2.52925e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B_c_66_n N_A_c_101_n 0.0206167f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_65 N_B_M1000_g N_VPWR_c_129_n 0.00159126f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_66 N_B_M1000_g N_VPWR_c_130_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_67 N_B_M1000_g N_VPWR_c_126_n 0.00969654f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_68 N_B_M1000_g N_Y_c_158_n 0.0100323f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_69 N_B_M1000_g N_Y_c_166_n 0.0116193f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_70 B N_Y_c_166_n 0.0271843f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_71 N_B_c_66_n N_Y_c_166_n 7.21566e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B_M1000_g N_Y_c_156_n 6.08373e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 B N_Y_c_153_n 0.0424861f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_74 N_B_c_67_n N_Y_c_153_n 0.0109855f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_75 N_B_M1000_g N_Y_c_163_n 0.00196977f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_76 N_B_c_67_n N_Y_c_154_n 0.00102554f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_77 B N_Y_c_174_n 0.0250978f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_78 N_B_c_66_n N_Y_c_174_n 4.33488e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B_c_67_n N_Y_c_174_n 0.0182272f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B_c_67_n N_VGND_c_208_n 0.00357877f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_67_n N_VGND_c_209_n 0.00546655f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_82 B A_193_47# 0.00254132f $X=1.07 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_83 N_A_M1005_g N_VPWR_c_129_n 0.00286079f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_VPWR_c_131_n 0.00541359f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_VPWR_c_126_n 0.0106235f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1005_g N_Y_c_158_n 6.08373e-19 $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1005_g N_Y_c_166_n 0.014647f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1005_g N_Y_c_155_n 0.00125894f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_89 A N_Y_c_155_n 0.0225129f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_101_n N_Y_c_155_n 0.00553375f $X=1.555 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_Y_c_156_n 0.0100323f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_c_99_n N_Y_c_154_n 0.00690727f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_93 A N_Y_c_154_n 0.0221415f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A_c_101_n N_Y_c_154_n 0.00550402f $X=1.555 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_c_99_n N_Y_c_174_n 0.0161709f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_c_99_n N_VGND_c_208_n 0.00359354f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_c_99_n N_VGND_c_209_n 0.00634452f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_98 N_VPWR_c_126_n N_Y_M1002_d 0.00215201f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_99 N_VPWR_c_126_n N_Y_M1005_d 0.00209319f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_100 N_VPWR_c_130_n N_Y_c_158_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_101 N_VPWR_c_126_n N_Y_c_158_n 0.0122217f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_102 N_VPWR_M1000_d N_Y_c_166_n 0.00444864f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_103 N_VPWR_c_129_n N_Y_c_166_n 0.0175734f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_104 N_VPWR_c_131_n N_Y_c_156_n 0.0210382f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_105 N_VPWR_c_126_n N_Y_c_156_n 0.0124268f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_106 N_Y_c_154_n N_VGND_c_208_n 0.0207942f $X=1.58 $Y=0.38 $X2=0 $Y2=0
cc_107 N_Y_c_174_n N_VGND_c_208_n 0.0419481f $X=1.415 $Y=0.425 $X2=0 $Y2=0
cc_108 Y N_VGND_c_208_n 0.0106076f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_109 N_Y_M1003_d N_VGND_c_209_n 0.00209319f $X=1.445 $Y=0.235 $X2=0 $Y2=0
cc_110 N_Y_c_154_n N_VGND_c_209_n 0.0123694f $X=1.58 $Y=0.38 $X2=0 $Y2=0
cc_111 N_Y_c_174_n N_VGND_c_209_n 0.0259983f $X=1.415 $Y=0.425 $X2=0 $Y2=0
cc_112 Y N_VGND_c_209_n 0.00679492f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_113 N_Y_c_153_n A_109_47# 0.00290753f $X=0.605 $Y=1.495 $X2=-0.19 $Y2=-0.24
cc_114 N_Y_c_174_n A_109_47# 0.0031671f $X=1.415 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_115 Y A_109_47# 9.09492e-19 $X=0.61 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_116 N_Y_c_174_n A_193_47# 0.00432137f $X=1.415 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_117 N_VGND_c_209_n A_109_47# 0.00216819f $X=1.61 $Y=0 $X2=-0.19 $Y2=-0.24
cc_118 N_VGND_c_209_n A_193_47# 0.00265018f $X=1.61 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a32o_2.spice.SKY130_FD_SC_HD__A32O_2.pxi
* Created: Thu Aug 27 14:05:24 2020
* 
x_PM_SKY130_FD_SC_HD__A32O_2%A_21_199# N_A_21_199#_M1002_d N_A_21_199#_M1012_d
+ N_A_21_199#_c_69_n N_A_21_199#_M1006_g N_A_21_199#_M1004_g N_A_21_199#_c_70_n
+ N_A_21_199#_M1013_g N_A_21_199#_M1010_g N_A_21_199#_c_71_n N_A_21_199#_c_77_n
+ N_A_21_199#_c_124_p N_A_21_199#_c_72_n N_A_21_199#_c_79_n N_A_21_199#_c_83_p
+ N_A_21_199#_c_89_p N_A_21_199#_c_93_p N_A_21_199#_c_94_p N_A_21_199#_c_84_p
+ N_A_21_199#_c_73_n PM_SKY130_FD_SC_HD__A32O_2%A_21_199#
x_PM_SKY130_FD_SC_HD__A32O_2%B2 N_B2_M1008_g N_B2_M1012_g N_B2_c_165_n
+ N_B2_c_166_n B2 B2 PM_SKY130_FD_SC_HD__A32O_2%B2
x_PM_SKY130_FD_SC_HD__A32O_2%B1 N_B1_M1002_g N_B1_M1011_g N_B1_c_205_n
+ N_B1_c_206_n B1 N_B1_c_208_n PM_SKY130_FD_SC_HD__A32O_2%B1
x_PM_SKY130_FD_SC_HD__A32O_2%A1 N_A1_M1007_g N_A1_M1009_g N_A1_c_250_n
+ N_A1_c_251_n N_A1_c_252_n A1 N_A1_c_253_n PM_SKY130_FD_SC_HD__A32O_2%A1
x_PM_SKY130_FD_SC_HD__A32O_2%A2 N_A2_c_290_n N_A2_M1003_g N_A2_M1001_g A2 A2 A2
+ A2 N_A2_c_293_n PM_SKY130_FD_SC_HD__A32O_2%A2
x_PM_SKY130_FD_SC_HD__A32O_2%A3 N_A3_c_334_n N_A3_M1005_g N_A3_M1000_g A3 A3
+ N_A3_c_336_n PM_SKY130_FD_SC_HD__A32O_2%A3
x_PM_SKY130_FD_SC_HD__A32O_2%X N_X_M1006_s N_X_M1004_d N_X_M1010_d N_X_c_365_n
+ N_X_c_370_n N_X_c_375_n X X X X X N_X_c_360_n X PM_SKY130_FD_SC_HD__A32O_2%X
x_PM_SKY130_FD_SC_HD__A32O_2%VPWR N_VPWR_M1004_s N_VPWR_M1009_d N_VPWR_M1000_d
+ N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n
+ N_VPWR_c_407_n VPWR N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n
+ N_VPWR_c_401_n PM_SKY130_FD_SC_HD__A32O_2%VPWR
x_PM_SKY130_FD_SC_HD__A32O_2%A_299_297# N_A_299_297#_M1012_s
+ N_A_299_297#_M1011_d N_A_299_297#_M1001_d N_A_299_297#_c_463_n
+ N_A_299_297#_c_464_n N_A_299_297#_c_480_n N_A_299_297#_c_469_n
+ N_A_299_297#_c_470_n N_A_299_297#_c_478_n
+ PM_SKY130_FD_SC_HD__A32O_2%A_299_297#
x_PM_SKY130_FD_SC_HD__A32O_2%VGND N_VGND_M1006_d N_VGND_M1013_d N_VGND_M1005_d
+ N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n N_VGND_c_498_n VGND
+ N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ PM_SKY130_FD_SC_HD__A32O_2%VGND
cc_1 VNB N_A_21_199#_c_69_n 0.0182689f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_21_199#_c_70_n 0.0183745f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_21_199#_c_71_n 6.46921e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_4 VNB N_A_21_199#_c_72_n 0.00111496f $X=-0.19 $Y=-0.24 $X2=1.795 $Y2=1.445
cc_5 VNB N_A_21_199#_c_73_n 0.0619839f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_6 VNB N_B2_c_165_n 0.0467187f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_B2_c_166_n 0.0187071f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_8 VNB B2 0.00519049f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_9 VNB N_B1_c_205_n 0.019694f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_10 VNB N_B1_c_206_n 0.00452257f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_11 VNB B1 7.17437e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_12 VNB N_B1_c_208_n 0.0177433f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_13 VNB N_A1_c_250_n 0.00255485f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_14 VNB N_A1_c_251_n 0.0230048f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_A1_c_252_n 0.00115789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_253_n 0.0180843f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_17 VNB N_A2_c_290_n 0.0171124f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=0.235
cc_18 VNB A2 0.0014855f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB A2 0.00256018f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_20 VNB N_A2_c_293_n 0.021893f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_21 VNB N_A3_c_334_n 0.0212957f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=0.235
cc_22 VNB A3 0.0135798f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_23 VNB N_A3_c_336_n 0.0364758f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_24 VNB N_X_c_360_n 0.00687827f $X=-0.19 $Y=-0.24 $X2=2.04 $Y2=1.63
cc_25 VNB X 0.00489318f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.615
cc_26 VNB N_VPWR_c_401_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_495_n 0.0102396f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_28 VNB N_VGND_c_496_n 0.0126038f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_29 VNB N_VGND_c_497_n 0.0102727f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_30 VNB N_VGND_c_498_n 0.0252622f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_31 VNB N_VGND_c_499_n 0.0543071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_500_n 0.0122771f $X=-0.19 $Y=-0.24 $X2=2.42 $Y2=0.615
cc_33 VNB N_VGND_c_501_n 0.0130294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_502_n 0.217717f $X=-0.19 $Y=-0.24 $X2=2.04 $Y2=1.945
cc_35 VPB N_A_21_199#_M1004_g 0.0209564f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB N_A_21_199#_M1010_g 0.024768f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_37 VPB N_A_21_199#_c_71_n 0.00110294f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_38 VPB N_A_21_199#_c_77_n 0.0221865f $X=-0.19 $Y=1.305 $X2=1.7 $Y2=1.53
cc_39 VPB N_A_21_199#_c_72_n 0.00433344f $X=-0.19 $Y=1.305 $X2=1.795 $Y2=1.445
cc_40 VPB N_A_21_199#_c_79_n 0.003468f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.615
cc_41 VPB N_A_21_199#_c_73_n 0.0147792f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_42 VPB N_B2_M1012_g 0.0230609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B2_c_165_n 0.014952f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_44 VPB N_B1_M1011_g 0.0190656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B1_c_205_n 0.0053162f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_46 VPB B1 0.00333547f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_47 VPB N_A1_M1009_g 0.0204128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A1_c_250_n 0.00355917f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_49 VPB N_A1_c_251_n 0.00575562f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_50 VPB N_A2_M1001_g 0.0198325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB A2 5.83477e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_52 VPB A2 0.00153004f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_53 VPB N_A2_c_293_n 0.00460852f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_54 VPB N_A3_M1000_g 0.0212772f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB A3 0.0136664f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_56 VPB N_A3_c_336_n 0.0103896f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_57 VPB X 0.00692367f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_58 VPB X 0.00658948f $X=-0.19 $Y=1.305 $X2=2.42 $Y2=0.615
cc_59 VPB N_VPWR_c_402_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_60 VPB N_VPWR_c_403_n 0.00228535f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_61 VPB N_VPWR_c_404_n 0.0101444f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_VPWR_c_405_n 0.0252999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_406_n 0.0454145f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_64 VPB N_VPWR_c_407_n 0.00507808f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_65 VPB N_VPWR_c_408_n 0.015528f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.53
cc_66 VPB N_VPWR_c_409_n 0.0174538f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_410_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.04 $Y2=2.03
cc_68 VPB N_VPWR_c_401_n 0.0562101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 N_A_21_199#_c_72_n N_B2_M1012_g 0.00500684f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_70 N_A_21_199#_c_79_n N_B2_M1012_g 0.0129811f $X=2 $Y=1.615 $X2=0 $Y2=0
cc_71 N_A_21_199#_c_83_p N_B2_M1012_g 0.00918223f $X=2.04 $Y=1.63 $X2=0 $Y2=0
cc_72 N_A_21_199#_c_84_p N_B2_M1012_g 0.00227571f $X=2.04 $Y=2.03 $X2=0 $Y2=0
cc_73 N_A_21_199#_c_71_n N_B2_c_165_n 4.47682e-19 $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_21_199#_c_77_n N_B2_c_165_n 0.00713356f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_75 N_A_21_199#_c_72_n N_B2_c_165_n 0.0181726f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_76 N_A_21_199#_c_79_n N_B2_c_165_n 0.00744757f $X=2 $Y=1.615 $X2=0 $Y2=0
cc_77 N_A_21_199#_c_89_p N_B2_c_165_n 4.38855e-19 $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_78 N_A_21_199#_c_73_n N_B2_c_165_n 0.016861f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_21_199#_c_70_n N_B2_c_166_n 0.00835312f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_21_199#_c_72_n N_B2_c_166_n 0.0044975f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_81 N_A_21_199#_c_93_p N_B2_c_166_n 0.0107495f $X=1.89 $Y=0.7 $X2=0 $Y2=0
cc_82 N_A_21_199#_c_94_p N_B2_c_166_n 0.00129054f $X=2.42 $Y=0.36 $X2=0 $Y2=0
cc_83 N_A_21_199#_c_70_n B2 0.00883089f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_21_199#_c_71_n B2 0.0112037f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_21_199#_c_77_n B2 0.0328575f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_86 N_A_21_199#_c_72_n B2 0.036593f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_87 N_A_21_199#_c_93_p B2 0.00335214f $X=1.89 $Y=0.7 $X2=0 $Y2=0
cc_88 N_A_21_199#_c_72_n N_B1_M1011_g 4.26124e-19 $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_89 N_A_21_199#_c_79_n N_B1_M1011_g 3.4843e-19 $X=2 $Y=1.615 $X2=0 $Y2=0
cc_90 N_A_21_199#_c_84_p N_B1_M1011_g 0.0033929f $X=2.04 $Y=2.03 $X2=0 $Y2=0
cc_91 N_A_21_199#_c_72_n N_B1_c_205_n 0.00106164f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_92 N_A_21_199#_c_79_n N_B1_c_205_n 2.83298e-19 $X=2 $Y=1.615 $X2=0 $Y2=0
cc_93 N_A_21_199#_c_89_p N_B1_c_205_n 0.00282103f $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_94 N_A_21_199#_c_72_n N_B1_c_206_n 0.0118465f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_95 N_A_21_199#_c_79_n N_B1_c_206_n 0.00264867f $X=2 $Y=1.615 $X2=0 $Y2=0
cc_96 N_A_21_199#_c_89_p N_B1_c_206_n 0.0190498f $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_97 N_A_21_199#_c_72_n B1 0.00655709f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_98 N_A_21_199#_c_79_n B1 0.00270821f $X=2 $Y=1.615 $X2=0 $Y2=0
cc_99 N_A_21_199#_c_89_p B1 8.54474e-19 $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_100 N_A_21_199#_c_72_n N_B1_c_208_n 0.00427939f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_101 N_A_21_199#_c_89_p N_B1_c_208_n 0.0104968f $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_102 N_A_21_199#_c_94_p N_B1_c_208_n 0.00625011f $X=2.42 $Y=0.36 $X2=0 $Y2=0
cc_103 N_A_21_199#_c_77_n N_X_M1010_d 0.00383016f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_104 N_A_21_199#_c_69_n N_X_c_365_n 0.0151812f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_21_199#_c_70_n N_X_c_365_n 0.00680881f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_21_199#_c_71_n N_X_c_365_n 0.010971f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_21_199#_c_77_n N_X_c_365_n 0.00307454f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_108 N_A_21_199#_c_73_n N_X_c_365_n 0.00106268f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_21_199#_M1004_g N_X_c_370_n 0.0135515f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_21_199#_M1010_g N_X_c_370_n 0.00932032f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_21_199#_c_77_n N_X_c_370_n 0.0139464f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_112 N_A_21_199#_c_124_p N_X_c_370_n 0.00903197f $X=0.705 $Y=1.53 $X2=0 $Y2=0
cc_113 N_A_21_199#_c_73_n N_X_c_370_n 2.98348e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_21_199#_c_77_n N_X_c_375_n 0.0132614f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_115 N_A_21_199#_c_69_n X 0.00551704f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_21_199#_M1004_g X 0.00878106f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_21_199#_c_71_n X 0.0287673f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_21_199#_c_124_p X 0.00795336f $X=0.705 $Y=1.53 $X2=0 $Y2=0
cc_119 N_A_21_199#_c_73_n X 0.0331912f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_21_199#_c_77_n N_VPWR_M1004_s 5.54118e-19 $X=1.7 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_21_199#_c_124_p N_VPWR_M1004_s 0.00112835f $X=0.705 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_21_199#_M1004_g N_VPWR_c_402_n 0.0107109f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_21_199#_M1010_g N_VPWR_c_402_n 0.0107254f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_21_199#_M1010_g N_VPWR_c_406_n 0.0046653f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_21_199#_M1004_g N_VPWR_c_408_n 0.0046653f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_21_199#_M1012_d N_VPWR_c_401_n 0.00216833f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_127 N_A_21_199#_M1004_g N_VPWR_c_401_n 0.00515525f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_21_199#_M1010_g N_VPWR_c_401_n 0.00552712f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_21_199#_c_77_n N_A_299_297#_M1012_s 0.00379791f $X=1.7 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_130 N_A_21_199#_c_77_n N_A_299_297#_c_463_n 0.0131801f $X=1.7 $Y=1.53 $X2=0
+ $Y2=0
cc_131 N_A_21_199#_M1012_d N_A_299_297#_c_464_n 0.00316374f $X=1.905 $Y=1.485
+ $X2=0 $Y2=0
cc_132 N_A_21_199#_c_84_p N_A_299_297#_c_464_n 0.0146785f $X=2.04 $Y=2.03 $X2=0
+ $Y2=0
cc_133 N_A_21_199#_c_69_n N_VGND_c_496_n 0.00926215f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_21_199#_c_70_n N_VGND_c_496_n 0.00114456f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_135 N_A_21_199#_c_73_n N_VGND_c_496_n 0.00168205f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_21_199#_c_89_p N_VGND_c_499_n 0.00604929f $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_137 N_A_21_199#_c_93_p N_VGND_c_499_n 0.00319227f $X=1.89 $Y=0.7 $X2=0 $Y2=0
cc_138 N_A_21_199#_c_94_p N_VGND_c_499_n 0.0169571f $X=2.42 $Y=0.36 $X2=0 $Y2=0
cc_139 N_A_21_199#_c_69_n N_VGND_c_500_n 0.00341689f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_140 N_A_21_199#_c_70_n N_VGND_c_500_n 0.00435058f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_21_199#_c_69_n N_VGND_c_501_n 0.00105764f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_A_21_199#_c_70_n N_VGND_c_501_n 0.00992118f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_21_199#_c_94_p N_VGND_c_501_n 0.0046429f $X=2.42 $Y=0.36 $X2=0 $Y2=0
cc_144 N_A_21_199#_M1002_d N_VGND_c_502_n 0.00299085f $X=2.265 $Y=0.235 $X2=0
+ $Y2=0
cc_145 N_A_21_199#_c_69_n N_VGND_c_502_n 0.0040262f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_21_199#_c_70_n N_VGND_c_502_n 0.00694191f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_21_199#_c_89_p N_VGND_c_502_n 0.0097927f $X=2.255 $Y=0.7 $X2=0 $Y2=0
cc_148 N_A_21_199#_c_93_p N_VGND_c_502_n 0.00549371f $X=1.89 $Y=0.7 $X2=0 $Y2=0
cc_149 N_A_21_199#_c_94_p N_VGND_c_502_n 0.0122988f $X=2.42 $Y=0.36 $X2=0 $Y2=0
cc_150 N_A_21_199#_c_72_n A_352_47# 0.00121143f $X=1.795 $Y=1.445 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_21_199#_c_89_p A_352_47# 0.00608077f $X=2.255 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_21_199#_c_93_p A_352_47# 0.00130299f $X=1.89 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_153 N_B2_M1012_g N_B1_M1011_g 0.0259824f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B2_c_165_n N_B1_c_205_n 0.0222403f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B2_c_165_n N_B1_c_206_n 0.00110488f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B2_c_165_n B1 2.26692e-19 $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B2_c_166_n N_B1_c_208_n 0.0295547f $X=1.757 $Y=0.995 $X2=0 $Y2=0
cc_158 B2 N_X_c_365_n 0.00464844f $X=1.125 $Y=0.765 $X2=0 $Y2=0
cc_159 N_B2_M1012_g N_VPWR_c_406_n 0.00357877f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B2_M1012_g N_VPWR_c_401_n 0.00657948f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B2_M1012_g N_A_299_297#_c_464_n 0.0112555f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_162 B2 N_VGND_M1013_d 0.0100518f $X=1.125 $Y=0.765 $X2=0 $Y2=0
cc_163 N_B2_c_166_n N_VGND_c_499_n 0.00401161f $X=1.757 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_165_n N_VGND_c_501_n 0.00279563f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B2_c_166_n N_VGND_c_501_n 0.0116145f $X=1.757 $Y=0.995 $X2=0 $Y2=0
cc_166 B2 N_VGND_c_501_n 0.0209142f $X=1.125 $Y=0.765 $X2=0 $Y2=0
cc_167 N_B2_c_166_n N_VGND_c_502_n 0.00615567f $X=1.757 $Y=0.995 $X2=0 $Y2=0
cc_168 B2 N_VGND_c_502_n 0.0022721f $X=1.125 $Y=0.765 $X2=0 $Y2=0
cc_169 N_B1_M1011_g N_A1_M1009_g 0.0246424f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_170 B1 N_A1_M1009_g 0.00151672f $X=2.355 $Y=1.445 $X2=0 $Y2=0
cc_171 N_B1_c_205_n N_A1_c_250_n 6.71537e-19 $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_172 N_B1_c_206_n N_A1_c_250_n 0.0135529f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_173 B1 N_A1_c_250_n 0.00596835f $X=2.355 $Y=1.445 $X2=0 $Y2=0
cc_174 N_B1_c_205_n N_A1_c_251_n 0.0207793f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B1_c_206_n N_A1_c_251_n 0.00116021f $X=2.43 $Y=1.16 $X2=0 $Y2=0
cc_176 B1 N_A1_c_251_n 0.00323874f $X=2.355 $Y=1.445 $X2=0 $Y2=0
cc_177 N_B1_c_208_n N_A1_c_253_n 0.00965926f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B1_M1011_g N_VPWR_c_403_n 0.00110007f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_179 N_B1_M1011_g N_VPWR_c_406_n 0.00357877f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1011_g N_VPWR_c_401_n 0.00528062f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_181 B1 N_A_299_297#_M1011_d 0.00266867f $X=2.355 $Y=1.445 $X2=0 $Y2=0
cc_182 N_B1_M1011_g N_A_299_297#_c_464_n 0.0112555f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_183 B1 N_A_299_297#_c_469_n 0.0127817f $X=2.355 $Y=1.445 $X2=0 $Y2=0
cc_184 N_B1_c_208_n N_VGND_c_499_n 0.00419584f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B1_c_208_n N_VGND_c_501_n 0.00169718f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_208_n N_VGND_c_502_n 0.00614197f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_252_n N_A2_c_290_n 0.00333931f $X=2.835 $Y=0.955 $X2=-0.19
+ $Y2=-0.24
cc_188 A1 N_A2_c_290_n 0.00190147f $X=2.905 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_189 N_A1_c_253_n N_A2_c_290_n 0.0204014f $X=2.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_190 N_A1_M1009_g N_A2_M1001_g 0.0282973f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A1_c_252_n A2 0.0176409f $X=2.835 $Y=0.955 $X2=0 $Y2=0
cc_192 A1 A2 0.0124253f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_193 N_A1_c_250_n A2 0.0250481f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A1_c_251_n A2 3.24056e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A1_M1009_g A2 0.0013511f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A1_c_250_n N_A2_c_293_n 0.00202486f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A1_c_251_n N_A2_c_293_n 0.0202158f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A1_M1009_g N_VPWR_c_403_n 0.0101679f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A1_M1009_g N_VPWR_c_406_n 0.0035268f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A1_M1009_g N_VPWR_c_401_n 0.00420827f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A1_M1009_g N_A_299_297#_c_470_n 0.0139487f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A1_c_250_n N_A_299_297#_c_470_n 0.00976902f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A1_c_251_n N_A_299_297#_c_470_n 7.09071e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_204 A1 N_VGND_c_498_n 2.56535e-19 $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_205 A1 N_VGND_c_499_n 0.0103948f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_206 N_A1_c_253_n N_VGND_c_499_n 0.00585385f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_207 A1 N_VGND_c_502_n 0.0117623f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_208 N_A1_c_253_n N_VGND_c_502_n 0.0112884f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_252_n A_549_47# 0.0053498f $X=2.835 $Y=0.955 $X2=-0.19 $Y2=-0.24
cc_210 A1 A_549_47# 0.0140793f $X=2.905 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_211 N_A2_c_290_n N_A3_c_334_n 0.0396565f $X=3.25 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_212 A2 N_A3_c_334_n 0.00467581f $X=3.365 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_213 N_A2_M1001_g N_A3_M1000_g 0.0266827f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_214 A2 N_A3_M1000_g 0.0019636f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_215 A2 A3 0.0182501f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_216 A2 A3 0.0129638f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_217 N_A2_c_293_n A3 2.3903e-19 $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_218 A2 N_A3_c_336_n 0.00305966f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_219 N_A2_c_293_n N_A3_c_336_n 0.0207914f $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A2_M1001_g N_VPWR_c_403_n 0.00503117f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A2_M1001_g N_VPWR_c_405_n 6.59159e-19 $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A2_M1001_g N_VPWR_c_409_n 0.00441875f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A2_M1001_g N_VPWR_c_401_n 0.00654032f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_224 A2 N_A_299_297#_M1001_d 0.00190479f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_225 N_A2_M1001_g N_A_299_297#_c_470_n 0.0123221f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_226 A2 N_A_299_297#_c_470_n 0.00426009f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_227 A2 N_A_299_297#_c_470_n 0.00131957f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_228 N_A2_c_293_n N_A_299_297#_c_470_n 9.23185e-19 $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_229 A2 N_A_299_297#_c_478_n 0.013246f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_230 N_A2_c_290_n N_VGND_c_498_n 0.00224948f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A2_c_290_n N_VGND_c_499_n 0.00560723f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_232 A2 N_VGND_c_499_n 0.00682938f $X=3.365 $Y=0.425 $X2=0 $Y2=0
cc_233 N_A2_c_290_n N_VGND_c_502_n 0.0105429f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_234 A2 N_VGND_c_502_n 0.00815638f $X=3.365 $Y=0.425 $X2=0 $Y2=0
cc_235 A2 A_665_47# 0.00277617f $X=3.365 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_236 A3 N_VPWR_M1000_d 0.00540294f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_237 N_A3_M1000_g N_VPWR_c_405_n 0.012699f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_238 A3 N_VPWR_c_405_n 0.0144066f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A3_c_336_n N_VPWR_c_405_n 0.00208124f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A3_M1000_g N_VPWR_c_409_n 0.0046653f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A3_M1000_g N_VPWR_c_401_n 0.007919f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A3_c_334_n N_VGND_c_498_n 0.0149399f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_243 A3 N_VGND_c_498_n 0.018723f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_244 N_A3_c_336_n N_VGND_c_498_n 0.0034472f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A3_c_334_n N_VGND_c_499_n 0.0046653f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A3_c_334_n N_VGND_c_502_n 0.00799591f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_247 N_X_c_370_n N_VPWR_M1004_s 0.00315845f $X=1.015 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_248 N_X_c_370_n N_VPWR_c_402_n 0.0165384f $X=1.015 $Y=1.87 $X2=0 $Y2=0
cc_249 N_X_c_375_n N_VPWR_c_406_n 0.0116048f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_250 X N_VPWR_c_408_n 0.0144177f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_251 N_X_M1004_d N_VPWR_c_401_n 0.00235001f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_252 N_X_M1010_d N_VPWR_c_401_n 0.00378138f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_253 N_X_c_370_n N_VPWR_c_401_n 0.0117708f $X=1.015 $Y=1.87 $X2=0 $Y2=0
cc_254 N_X_c_375_n N_VPWR_c_401_n 0.00646998f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_255 X N_VPWR_c_401_n 0.00801045f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_256 N_X_c_375_n N_A_299_297#_c_463_n 0.0225975f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_257 N_X_c_375_n N_A_299_297#_c_480_n 0.00811593f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_258 N_X_c_360_n N_VGND_M1006_d 0.0105966f $X=0.24 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_259 X N_VGND_M1006_d 0.0023095f $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_260 N_X_c_365_n N_VGND_c_496_n 0.00183815f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_261 N_X_c_360_n N_VGND_c_496_n 0.015569f $X=0.24 $Y=0.825 $X2=0 $Y2=0
cc_262 N_X_c_365_n N_VGND_c_500_n 0.00599455f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_263 N_X_M1006_s N_VGND_c_502_n 0.00323135f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_264 N_X_c_365_n N_VGND_c_502_n 0.011321f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_265 N_X_c_360_n N_VGND_c_502_n 0.00107851f $X=0.24 $Y=0.825 $X2=0 $Y2=0
cc_266 N_VPWR_c_401_n N_A_299_297#_M1012_s 0.00348186f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_267 N_VPWR_c_401_n N_A_299_297#_M1011_d 0.00241761f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_401_n N_A_299_297#_M1001_d 0.00414531f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_406_n N_A_299_297#_c_464_n 0.0472939f $X=2.715 $Y=2.72 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_401_n N_A_299_297#_c_464_n 0.0299868f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_406_n N_A_299_297#_c_480_n 0.0117106f $X=2.715 $Y=2.72 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_401_n N_A_299_297#_c_480_n 0.006547f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_273 N_VPWR_M1009_d N_A_299_297#_c_470_n 0.0125255f $X=2.745 $Y=1.485 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_403_n N_A_299_297#_c_470_n 0.0206595f $X=2.88 $Y=2.225 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_406_n N_A_299_297#_c_470_n 0.0018545f $X=2.715 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_409_n N_A_299_297#_c_470_n 0.00363691f $X=3.715 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_401_n N_A_299_297#_c_470_n 0.0127237f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_409_n N_A_299_297#_c_478_n 0.0113839f $X=3.715 $Y=2.72 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_401_n N_A_299_297#_c_478_n 0.00646745f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VGND_c_502_n A_352_47# 0.00404223f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_281 N_VGND_c_502_n A_549_47# 0.00654476f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_282 N_VGND_c_502_n A_665_47# 0.00415276f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

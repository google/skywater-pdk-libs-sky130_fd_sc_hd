* File: sky130_fd_sc_hd__a32o_1.pxi.spice
* Created: Tue Sep  1 18:55:36 2020
* 
x_PM_SKY130_FD_SC_HD__A32O_1%A_93_21# N_A_93_21#_M1000_d N_A_93_21#_M1006_d
+ N_A_93_21#_M1005_g N_A_93_21#_M1004_g N_A_93_21#_c_65_n N_A_93_21#_c_71_p
+ N_A_93_21#_c_109_p N_A_93_21#_c_70_p N_A_93_21#_c_110_p N_A_93_21#_c_81_p
+ N_A_93_21#_c_82_p N_A_93_21#_c_73_p N_A_93_21#_c_133_p N_A_93_21#_c_60_n
+ N_A_93_21#_c_61_n N_A_93_21#_c_62_n N_A_93_21#_c_63_n
+ PM_SKY130_FD_SC_HD__A32O_1%A_93_21#
x_PM_SKY130_FD_SC_HD__A32O_1%A3 N_A3_M1011_g N_A3_M1008_g A3 N_A3_c_156_n
+ N_A3_c_157_n PM_SKY130_FD_SC_HD__A32O_1%A3
x_PM_SKY130_FD_SC_HD__A32O_1%A2 N_A2_M1009_g N_A2_M1007_g A2 A2 N_A2_c_193_n
+ N_A2_c_194_n PM_SKY130_FD_SC_HD__A32O_1%A2
x_PM_SKY130_FD_SC_HD__A32O_1%A1 N_A1_M1000_g N_A1_M1010_g A1 A1 N_A1_c_230_n
+ N_A1_c_231_n PM_SKY130_FD_SC_HD__A32O_1%A1
x_PM_SKY130_FD_SC_HD__A32O_1%B1 N_B1_M1006_g N_B1_M1002_g B1 B1 N_B1_c_264_n
+ N_B1_c_265_n PM_SKY130_FD_SC_HD__A32O_1%B1
x_PM_SKY130_FD_SC_HD__A32O_1%B2 N_B2_M1003_g N_B2_M1001_g B2 B2 N_B2_c_299_n
+ N_B2_c_300_n PM_SKY130_FD_SC_HD__A32O_1%B2
x_PM_SKY130_FD_SC_HD__A32O_1%X N_X_M1005_s N_X_M1004_s X X X X X X X N_X_c_323_n
+ X PM_SKY130_FD_SC_HD__A32O_1%X
x_PM_SKY130_FD_SC_HD__A32O_1%VPWR N_VPWR_M1004_d N_VPWR_M1007_d N_VPWR_c_341_n
+ N_VPWR_c_342_n VPWR N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_340_n
+ N_VPWR_c_346_n N_VPWR_c_347_n PM_SKY130_FD_SC_HD__A32O_1%VPWR
x_PM_SKY130_FD_SC_HD__A32O_1%A_250_297# N_A_250_297#_M1011_d
+ N_A_250_297#_M1010_d N_A_250_297#_M1001_d N_A_250_297#_c_395_n
+ N_A_250_297#_c_412_n N_A_250_297#_c_396_n N_A_250_297#_c_397_n
+ N_A_250_297#_c_398_n N_A_250_297#_c_422_n N_A_250_297#_c_406_n
+ PM_SKY130_FD_SC_HD__A32O_1%A_250_297#
x_PM_SKY130_FD_SC_HD__A32O_1%VGND N_VGND_M1005_d N_VGND_M1003_d N_VGND_c_424_n
+ N_VGND_c_425_n N_VGND_c_426_n VGND N_VGND_c_427_n N_VGND_c_428_n
+ N_VGND_c_429_n N_VGND_c_430_n PM_SKY130_FD_SC_HD__A32O_1%VGND
cc_1 VNB N_A_93_21#_c_60_n 0.00334019f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_2 VNB N_A_93_21#_c_61_n 0.0274451f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_3 VNB N_A_93_21#_c_62_n 0.00194437f $X=-0.19 $Y=-0.24 $X2=0.722 $Y2=0.995
cc_4 VNB N_A_93_21#_c_63_n 0.020992f $X=-0.19 $Y=-0.24 $X2=0.627 $Y2=0.995
cc_5 VNB A3 0.00233795f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_6 VNB N_A3_c_156_n 0.0220372f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.985
cc_7 VNB N_A3_c_157_n 0.0185846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB A2 0.00388985f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_9 VNB N_A2_c_193_n 0.020678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A2_c_194_n 0.0169206f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.995
cc_11 VNB A1 0.00263615f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_12 VNB N_A1_c_230_n 0.0218583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A1_c_231_n 0.0186152f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.995
cc_14 VNB B1 0.00268297f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_15 VNB N_B1_c_264_n 0.0220377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_c_265_n 0.016623f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.995
cc_17 VNB B2 0.0128601f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_18 VNB N_B2_c_299_n 0.0257796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B2_c_300_n 0.0207477f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.995
cc_20 VNB X 0.0341759f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_21 VNB N_X_c_323_n 0.0104776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_340_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_424_n 0.00287347f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_24 VNB N_VGND_c_425_n 0.0103657f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.985
cc_25 VNB N_VGND_c_426_n 0.0263776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_427_n 0.0171616f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.495
cc_27 VNB N_VGND_c_428_n 0.0581519f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.485
cc_28 VNB N_VGND_c_429_n 0.00513206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_430_n 0.199703f $X=-0.19 $Y=-0.24 $X2=0.722 $Y2=0.995
cc_30 VPB N_A_93_21#_M1004_g 0.0242103f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.985
cc_31 VPB N_A_93_21#_c_65_n 0.00278936f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.495
cc_32 VPB N_A_93_21#_c_60_n 0.00282827f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_33 VPB N_A_93_21#_c_61_n 0.00641059f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_34 VPB N_A3_M1011_g 0.0217949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB A3 4.05393e-19 $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_36 VPB N_A3_c_156_n 0.00413877f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.985
cc_37 VPB N_A2_M1007_g 0.0216147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB A2 0.00119214f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_39 VPB N_A2_c_193_n 0.004301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A1_M1010_g 0.0220179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB A1 0.00189157f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_42 VPB N_A1_c_230_n 0.00461953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B1_M1006_g 0.0203318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB B1 0.00263532f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_45 VPB N_B1_c_264_n 0.00449145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_B2_M1001_g 0.0223177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB B2 0.00108204f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_48 VPB B2 0.0074672f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_49 VPB N_B2_c_299_n 0.0059105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB X 0.0257314f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_51 VPB X 0.0065071f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.985
cc_52 VPB X 0.0136697f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.985
cc_53 VPB N_VPWR_c_341_n 0.00564356f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.985
cc_54 VPB N_VPWR_c_342_n 0.00564356f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=0.995
cc_55 VPB N_VPWR_c_343_n 0.0211763f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=0.74
cc_56 VPB N_VPWR_c_344_n 0.0396882f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=0.4
cc_57 VPB N_VPWR_c_340_n 0.0454843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_346_n 0.0270476f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.96
cc_59 VPB N_VPWR_c_347_n 0.00631679f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_60 N_A_93_21#_M1004_g N_A3_M1011_g 0.0242549f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_93_21#_c_65_n N_A3_M1011_g 0.0017871f $X=0.79 $Y=1.495 $X2=0 $Y2=0
cc_62 N_A_93_21#_c_70_p N_A3_M1011_g 0.0159262f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_63 N_A_93_21#_c_71_p A3 0.0130226f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A_93_21#_c_70_p A3 0.0150596f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_93_21#_c_73_p A3 0.00103508f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_66 N_A_93_21#_c_60_n A3 0.0242383f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_93_21#_c_61_n A3 9.52067e-19 $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_93_21#_c_70_p N_A3_c_156_n 0.0034409f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_69 N_A_93_21#_c_73_p N_A3_c_156_n 0.0016757f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_70 N_A_93_21#_c_60_n N_A3_c_156_n 0.00290133f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_93_21#_c_61_n N_A3_c_156_n 0.0131273f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_93_21#_c_71_p N_A3_c_157_n 0.00814851f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A_93_21#_c_81_p N_A3_c_157_n 0.00575845f $X=1.18 $Y=0.655 $X2=0 $Y2=0
cc_74 N_A_93_21#_c_82_p N_A3_c_157_n 0.00511741f $X=1.265 $Y=0.4 $X2=0 $Y2=0
cc_75 N_A_93_21#_c_73_p N_A3_c_157_n 0.00280533f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_76 N_A_93_21#_c_62_n N_A3_c_157_n 0.00182225f $X=0.722 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_93_21#_c_63_n N_A3_c_157_n 0.0121679f $X=0.627 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_93_21#_c_70_p N_A2_M1007_g 0.0117253f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_79 N_A_93_21#_c_70_p A2 0.0170045f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A_93_21#_c_73_p A2 0.0111382f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_81 N_A_93_21#_c_62_n A2 0.00411674f $X=0.722 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_93_21#_c_70_p N_A2_c_193_n 0.00227792f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_93_21#_c_73_p N_A2_c_193_n 0.00151111f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_84 N_A_93_21#_c_71_p N_A2_c_194_n 2.46613e-19 $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A_93_21#_c_81_p N_A2_c_194_n 0.00101956f $X=1.18 $Y=0.655 $X2=0 $Y2=0
cc_86 N_A_93_21#_c_73_p N_A2_c_194_n 0.0110222f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_87 N_A_93_21#_c_70_p N_A1_M1010_g 0.0134825f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_93_21#_c_70_p A1 0.0205739f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_93_21#_c_73_p A1 0.0164469f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_90 N_A_93_21#_c_70_p N_A1_c_230_n 7.21566e-19 $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_93_21#_c_73_p N_A1_c_230_n 3.46281e-19 $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_92 N_A_93_21#_c_73_p N_A1_c_231_n 0.0129625f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_93 N_A_93_21#_c_70_p N_B1_M1006_g 0.0125783f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_93_21#_M1000_d B1 0.00588959f $X=2.33 $Y=0.235 $X2=0 $Y2=0
cc_95 N_A_93_21#_c_70_p B1 0.0305579f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_93_21#_c_73_p B1 0.0194562f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_97 N_A_93_21#_c_70_p N_B1_c_264_n 6.67961e-19 $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_93_21#_c_73_p N_B1_c_264_n 2.05846e-19 $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_99 N_A_93_21#_c_73_p N_B1_c_265_n 0.00278225f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_100 N_A_93_21#_c_65_n X 0.00775901f $X=0.79 $Y=1.495 $X2=0 $Y2=0
cc_101 N_A_93_21#_c_109_p X 0.00803736f $X=0.875 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_93_21#_c_110_p X 0.00816166f $X=0.875 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A_93_21#_c_60_n X 0.0206287f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_93_21#_c_62_n X 0.00761031f $X=0.722 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_93_21#_c_63_n X 0.0356252f $X=0.627 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_93_21#_c_65_n N_VPWR_M1004_d 2.08871e-19 $X=0.79 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_93_21#_c_70_p N_VPWR_M1004_d 0.00658232f $X=2.905 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_93_21#_c_110_p N_VPWR_M1004_d 0.00534275f $X=0.875 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_93_21#_c_70_p N_VPWR_M1007_d 0.0119524f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_93_21#_M1004_g N_VPWR_c_341_n 0.0114951f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_93_21#_c_70_p N_VPWR_c_341_n 0.0104588f $X=2.905 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A_93_21#_c_110_p N_VPWR_c_341_n 0.0152373f $X=0.875 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A_93_21#_c_60_n N_VPWR_c_341_n 0.00102128f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_93_21#_c_61_n N_VPWR_c_341_n 5.21175e-19 $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_93_21#_M1006_d N_VPWR_c_340_n 0.00224864f $X=2.85 $Y=1.485 $X2=0
+ $Y2=0
cc_116 N_A_93_21#_M1004_g N_VPWR_c_340_n 0.012253f $X=0.54 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_93_21#_M1004_g N_VPWR_c_346_n 0.00585385f $X=0.54 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_93_21#_c_70_p N_A_250_297#_M1011_d 0.0090427f $X=2.905 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_119 N_A_93_21#_c_70_p N_A_250_297#_M1010_d 0.00755311f $X=2.905 $Y=1.58 $X2=0
+ $Y2=0
cc_120 N_A_93_21#_c_70_p N_A_250_297#_c_395_n 0.0148437f $X=2.905 $Y=1.58 $X2=0
+ $Y2=0
cc_121 N_A_93_21#_c_70_p N_A_250_297#_c_396_n 0.0379866f $X=2.905 $Y=1.58 $X2=0
+ $Y2=0
cc_122 N_A_93_21#_c_70_p N_A_250_297#_c_397_n 0.0175925f $X=2.905 $Y=1.58 $X2=0
+ $Y2=0
cc_123 N_A_93_21#_M1006_d N_A_250_297#_c_398_n 0.0033237f $X=2.85 $Y=1.485 $X2=0
+ $Y2=0
cc_124 N_A_93_21#_c_70_p N_A_250_297#_c_398_n 0.00341278f $X=2.905 $Y=1.58 $X2=0
+ $Y2=0
cc_125 N_A_93_21#_c_133_p N_A_250_297#_c_398_n 0.0125742f $X=2.99 $Y=1.96 $X2=0
+ $Y2=0
cc_126 N_A_93_21#_c_71_p N_VGND_M1005_d 0.0076719f $X=1.095 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_93_21#_c_109_p N_VGND_M1005_d 0.0052382f $X=0.875 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_128 N_A_93_21#_c_62_n N_VGND_M1005_d 0.00155546f $X=0.722 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A_93_21#_c_71_p N_VGND_c_424_n 0.00372856f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_93_21#_c_109_p N_VGND_c_424_n 0.014416f $X=0.875 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_93_21#_c_60_n N_VGND_c_424_n 0.00261389f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_93_21#_c_61_n N_VGND_c_424_n 6.60966e-19 $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_93_21#_c_63_n N_VGND_c_424_n 0.0100805f $X=0.627 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_93_21#_c_73_p N_VGND_c_426_n 0.00556752f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_135 N_A_93_21#_c_63_n N_VGND_c_427_n 0.00505556f $X=0.627 $Y=0.995 $X2=0
+ $Y2=0
cc_136 N_A_93_21#_c_71_p N_VGND_c_428_n 0.00267478f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_93_21#_c_82_p N_VGND_c_428_n 0.00737272f $X=1.265 $Y=0.4 $X2=0 $Y2=0
cc_138 N_A_93_21#_c_73_p N_VGND_c_428_n 0.0601675f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_139 N_A_93_21#_M1000_d N_VGND_c_430_n 0.00385123f $X=2.33 $Y=0.235 $X2=0
+ $Y2=0
cc_140 N_A_93_21#_c_71_p N_VGND_c_430_n 0.00498507f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_93_21#_c_109_p N_VGND_c_430_n 8.26975e-19 $X=0.875 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_93_21#_c_82_p N_VGND_c_430_n 0.00565326f $X=1.265 $Y=0.4 $X2=0 $Y2=0
cc_143 N_A_93_21#_c_73_p N_VGND_c_430_n 0.0503517f $X=2.545 $Y=0.4 $X2=0 $Y2=0
cc_144 N_A_93_21#_c_63_n N_VGND_c_430_n 0.00963589f $X=0.627 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_93_21#_c_73_p A_256_47# 0.00833151f $X=2.545 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_93_21#_c_73_p A_346_47# 0.0120661f $X=2.545 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A3_M1011_g N_A2_M1007_g 0.0234228f $X=1.175 $Y=1.985 $X2=0 $Y2=0
cc_148 A3 A2 0.0214645f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A3_c_156_n A2 0.00199283f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A3_c_157_n A2 0.0017374f $X=1.235 $Y=0.995 $X2=0 $Y2=0
cc_151 A3 N_A2_c_193_n 3.4957e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A3_c_156_n N_A2_c_193_n 0.0202813f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A3_c_157_n N_A2_c_194_n 0.0364835f $X=1.235 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A3_M1011_g N_VPWR_c_341_n 0.0106196f $X=1.175 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A3_M1011_g N_VPWR_c_343_n 0.00585385f $X=1.175 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A3_M1011_g N_VPWR_c_340_n 0.0113788f $X=1.175 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A3_c_157_n N_VGND_c_424_n 0.0049358f $X=1.235 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A3_c_157_n N_VGND_c_428_n 0.00369937f $X=1.235 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A3_c_157_n N_VGND_c_430_n 0.00593126f $X=1.235 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_M1007_g N_A1_M1010_g 0.0328384f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_161 A2 A1 0.0475482f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_162 N_A2_c_193_n A1 0.00199358f $X=1.715 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A2_c_194_n A1 0.00110992f $X=1.715 $Y=0.995 $X2=0 $Y2=0
cc_164 A2 N_A1_c_230_n 3.35477e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_165 N_A2_c_193_n N_A1_c_230_n 0.0202262f $X=1.715 $Y=1.16 $X2=0 $Y2=0
cc_166 A2 N_A1_c_231_n 8.43574e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_167 N_A2_c_194_n N_A1_c_231_n 0.0238171f $X=1.715 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_M1007_g N_VPWR_c_342_n 0.00629737f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A2_M1007_g N_VPWR_c_343_n 0.00430895f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A2_M1007_g N_VPWR_c_340_n 0.00642336f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A2_M1007_g N_A_250_297#_c_396_n 0.0109884f $X=1.655 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A2_c_194_n N_VGND_c_428_n 0.00370116f $X=1.715 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_194_n N_VGND_c_430_n 0.00581846f $X=1.715 $Y=0.995 $X2=0 $Y2=0
cc_174 A2 A_346_47# 0.00224772f $X=1.53 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_175 N_A1_M1010_g N_B1_M1006_g 0.0216249f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_176 A1 B1 0.0523772f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_177 N_A1_c_231_n B1 0.00546688f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_178 A1 N_B1_c_264_n 2.86553e-19 $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_179 N_A1_c_230_n N_B1_c_264_n 0.0115654f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_180 A1 N_B1_c_265_n 2.55321e-19 $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_181 N_A1_c_231_n N_B1_c_265_n 0.0229868f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_M1010_g N_VPWR_c_342_n 0.00617297f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A1_M1010_g N_VPWR_c_344_n 0.00430895f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A1_M1010_g N_VPWR_c_340_n 0.00650893f $X=2.255 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A1_M1010_g N_A_250_297#_c_396_n 0.0109884f $X=2.255 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A1_c_231_n N_VGND_c_428_n 0.00370116f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_231_n N_VGND_c_430_n 0.0061191f $X=2.195 $Y=0.995 $X2=0 $Y2=0
cc_188 A1 A_346_47# 0.00354329f $X=1.99 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_189 N_B1_M1006_g N_B2_M1001_g 0.0391628f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_190 B1 B2 0.0156226f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_191 N_B1_c_264_n B2 0.00105949f $X=2.785 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B1_c_264_n N_B2_c_299_n 0.0369225f $X=2.785 $Y=1.16 $X2=0 $Y2=0
cc_193 B1 N_B2_c_300_n 0.00262439f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_194 N_B1_c_265_n N_B2_c_300_n 0.0369225f $X=2.785 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B1_M1006_g N_VPWR_c_344_n 0.00357877f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_M1006_g N_VPWR_c_340_n 0.00553224f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_M1006_g N_A_250_297#_c_398_n 0.00977092f $X=2.775 $Y=1.985 $X2=0
+ $Y2=0
cc_198 B1 N_VGND_c_426_n 0.0057423f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_199 N_B1_c_265_n N_VGND_c_426_n 0.00325933f $X=2.785 $Y=0.995 $X2=0 $Y2=0
cc_200 B1 N_VGND_c_428_n 0.00225695f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_201 N_B1_c_265_n N_VGND_c_428_n 0.00481907f $X=2.785 $Y=0.995 $X2=0 $Y2=0
cc_202 B1 N_VGND_c_430_n 0.0048308f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_203 N_B1_c_265_n N_VGND_c_430_n 0.00786256f $X=2.785 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B2_M1001_g N_VPWR_c_344_n 0.00357877f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B2_M1001_g N_VPWR_c_340_n 0.00623785f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_206 B2 N_A_250_297#_M1001_d 0.00911651f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_207 N_B2_M1001_g N_A_250_297#_c_398_n 0.0121906f $X=3.205 $Y=1.985 $X2=0
+ $Y2=0
cc_208 B2 N_A_250_297#_c_406_n 0.013551f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_209 N_B2_c_299_n N_A_250_297#_c_406_n 2.67591e-19 $X=3.265 $Y=1.16 $X2=0
+ $Y2=0
cc_210 B2 N_VGND_c_426_n 0.0188449f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_211 N_B2_c_299_n N_VGND_c_426_n 0.00258249f $X=3.265 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B2_c_300_n N_VGND_c_426_n 0.0156752f $X=3.265 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B2_c_300_n N_VGND_c_428_n 0.00486043f $X=3.265 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B2_c_300_n N_VGND_c_430_n 0.00814024f $X=3.265 $Y=0.995 $X2=0 $Y2=0
cc_215 X N_VPWR_c_341_n 0.00383937f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_216 N_X_M1004_s N_VPWR_c_340_n 0.00412347f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_217 X N_VPWR_c_340_n 0.0125459f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_218 X N_VPWR_c_346_n 0.0181662f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_219 N_X_c_323_n N_VGND_c_427_n 0.0175601f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_220 N_X_M1005_s N_VGND_c_430_n 0.00412857f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_221 N_X_c_323_n N_VGND_c_430_n 0.012458f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_222 N_VPWR_c_340_n N_A_250_297#_M1011_d 0.00281193f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_223 N_VPWR_c_340_n N_A_250_297#_M1010_d 0.00301425f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_340_n N_A_250_297#_M1001_d 0.00352286f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_341_n N_A_250_297#_c_395_n 0.0113606f $X=0.84 $Y=2 $X2=0 $Y2=0
cc_226 N_VPWR_c_341_n N_A_250_297#_c_412_n 0.0260639f $X=0.84 $Y=2 $X2=0 $Y2=0
cc_227 N_VPWR_c_343_n N_A_250_297#_c_412_n 0.0174097f $X=1.79 $Y=2.72 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_340_n N_A_250_297#_c_412_n 0.0108585f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_M1007_d N_A_250_297#_c_396_n 0.00798574f $X=1.73 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_342_n N_A_250_297#_c_396_n 0.025328f $X=1.955 $Y=2.34 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_343_n N_A_250_297#_c_396_n 0.00317309f $X=1.79 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_344_n N_A_250_297#_c_396_n 0.00290861f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_340_n N_A_250_297#_c_396_n 0.0130124f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_344_n N_A_250_297#_c_398_n 0.0476397f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_340_n N_A_250_297#_c_398_n 0.0296039f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_344_n N_A_250_297#_c_422_n 0.0204419f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_340_n N_A_250_297#_c_422_n 0.0126619f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VGND_c_430_n A_256_47# 0.00246016f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_239 N_VGND_c_430_n A_346_47# 0.00370537f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_240 N_VGND_c_430_n A_584_47# 0.00897657f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

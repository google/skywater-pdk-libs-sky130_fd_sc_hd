* File: sky130_fd_sc_hd__o2111ai_2.spice
* Created: Tue Sep  1 19:20:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2111ai_2.pex.spice"
.subckt sky130_fd_sc_hd__o2111ai_2  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1006 N_A_27_47#_M1006_d N_D1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.22425 AS=0.091 PD=1.99 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.3
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1007_d N_D1_M1007_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1007_d N_C1_M1004_g N_A_298_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75001.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_27_47#_M1016_d N_C1_M1016_g N_A_298_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.19175 AS=0.091 PD=1.89 PS=0.93 NRD=5.532 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_A_497_47#_M1013_d N_B1_M1013_g N_A_298_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1755 AS=0.091 PD=1.84 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1019 N_A_497_47#_M1019_d N_B1_M1019_g N_A_298_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1009 N_A_497_47#_M1019_d N_A2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1018 N_A_497_47#_M1018_d N_A2_M1018_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A1_M1010_g N_A_497_47#_M1018_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1010_d N_A1_M1015_g N_A_497_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.2145 PD=0.93 PS=1.96 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75002.3
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_D1_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.3 A=0.15
+ P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_D1_M1017_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001.9 A=0.15
+ P=2.3 MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001.5 A=0.15
+ P=2.3 MULT=1
MM1012 N_Y_M1000_d N_C1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1014 N_Y_M1002_d N_B1_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75000.2
+ A=0.15 P=2.3 MULT=1
MM1003 N_A_664_297#_M1003_d N_A2_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.14 PD=2.59 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1011 N_A_664_297#_M1011_d N_A2_M1011_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1001 N_A_664_297#_M1011_d N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1008 N_A_664_297#_M1008_d N_A1_M1008_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.33 AS=0.14 PD=2.66 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__o2111ai_2.pxi.spice"
*
.ends
*
*

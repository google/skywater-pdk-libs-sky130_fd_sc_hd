* File: sky130_fd_sc_hd__o21a_1.spice.pex
* Created: Thu Aug 27 14:35:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21A_1%A_79_21# 1 2 7 9 12 17 18 19 20 21 23 27
c57 21 0 1.03558e-19 $X=1.58 $Y=1.69
c58 20 0 5.84632e-20 $X=0.88 $Y=1.582
r59 31 33 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.49
+ $Y2=1.16
r60 21 30 2.8558 $w=3.3e-07 $l=1.08e-07 $layer=LI1_cond $X=1.58 $Y=1.69 $X2=1.58
+ $Y2=1.582
r61 21 23 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=1.58 $Y=1.69
+ $X2=1.58 $Y2=2.34
r62 19 30 4.36303 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=1.582
+ $X2=1.58 $Y2=1.582
r63 19 20 28.6771 $w=2.13e-07 $l=5.35e-07 $layer=LI1_cond $X=1.415 $Y=1.582
+ $X2=0.88 $Y2=1.582
r64 18 33 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.68 $Y=1.16
+ $X2=0.49 $Y2=1.16
r65 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.16 $X2=0.68 $Y2=1.16
r66 15 20 6.99171 $w=2.15e-07 $l=1.89077e-07 $layer=LI1_cond $X=0.737 $Y=1.475
+ $X2=0.88 $Y2=1.582
r67 15 17 12.7375 $w=2.83e-07 $l=3.15e-07 $layer=LI1_cond $X=0.737 $Y=1.475
+ $X2=0.737 $Y2=1.16
r68 14 27 14.983 $w=3.77e-07 $l=6.39397e-07 $layer=LI1_cond $X=0.737 $Y=0.905
+ $X2=1.2 $Y2=0.485
r69 14 17 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.737 $Y=0.905
+ $X2=0.737 $Y2=1.16
r70 10 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r71 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r72 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r73 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r74 2 30 400 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=1.485 $X2=1.58 $Y2=1.66
r75 2 23 400 $w=1.7e-07 $l=9.54241e-07 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=1.485 $X2=1.58 $Y2=2.34
r76 1 27 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.74
r77 1 27 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%B1 3 7 8 11 12 13
c33 13 0 1.80509e-19 $X=1.362 $Y=0.995
c34 11 0 1.22088e-19 $X=1.37 $Y=1.16
r35 11 14 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.362 $Y=1.16
+ $X2=1.362 $Y2=1.325
r36 11 13 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.362 $Y=1.16
+ $X2=1.362 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r38 8 12 11.0234 $w=2.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.15 $Y=1.19 $X2=1.37
+ $Y2=1.19
r39 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.56 $X2=1.41
+ $Y2=0.995
r40 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.295 $Y=1.985
+ $X2=1.295 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%A2 3 5 7 8 12
c39 12 0 1.97717e-19 $X=1.87 $Y=1.16
c40 8 0 1.22088e-19 $X=2.07 $Y=1.19
c41 3 0 1.03558e-19 $X=1.835 $Y=1.985
r42 16 21 0.111026 $w=2.15e-07 $l=1e-07 $layer=LI1_cond $X=2.047 $Y=1.275
+ $X2=2.047 $Y2=1.175
r43 13 21 11.1309 $w=1.94e-07 $l=1.77e-07 $layer=LI1_cond $X=1.87 $Y=1.175
+ $X2=2.047 $Y2=1.175
r44 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.16
+ $X2=1.87 $Y2=1.325
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.87
+ $Y=1.16 $X2=1.87 $Y2=1.16
r46 8 21 1.44639 $w=1.94e-07 $l=2.3e-08 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=2.047 $Y2=1.175
r47 8 16 0.251659 $w=1.113e-06 $l=2.3e-08 $layer=LI1_cond $X=2.07 $Y=1.832
+ $X2=2.047 $Y2=1.832
r48 5 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=0.995
+ $X2=1.87 $Y2=1.16
r49 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.87 $Y=0.995 $X2=1.87
+ $Y2=0.56
r50 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.835 $Y=1.985
+ $X2=1.835 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%A1 1 3 6 10 11 14
c28 14 0 3.61265e-20 $X=2.53 $Y=1.53
c29 10 0 1.61591e-19 $X=2.51 $Y=1.16
r30 13 14 12.7771 $w=2.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.56 $Y=1.275
+ $X2=2.56 $Y2=1.53
r31 11 16 36.2712 $w=3.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.51 $Y=1.17
+ $X2=2.29 $Y2=1.17
r32 10 13 5.08648 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.51 $Y=1.16
+ $X2=2.51 $Y2=1.275
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.16 $X2=2.51 $Y2=1.16
r34 4 16 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.29 $Y=1.345
+ $X2=2.29 $Y2=1.17
r35 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.29 $Y=1.345 $X2=2.29
+ $Y2=1.985
r36 1 16 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.29 $Y=0.995
+ $X2=2.29 $Y2=1.17
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.29 $Y=0.995 $X2=2.29
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%X 1 2 9 12 13 16
r19 13 20 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=2.3
r20 13 16 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.62
r21 12 16 24.2836 $w=2.78e-07 $l=5.9e-07 $layer=LI1_cond $X=0.225 $Y=1.03
+ $X2=0.225 $Y2=1.62
r22 7 12 6.15521 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.86
+ $X2=0.255 $Y2=1.03
r23 7 9 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=0.255 $Y=0.86
+ $X2=0.255 $Y2=0.395
r24 2 20 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r25 2 16 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r26 1 9 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%VPWR 1 2 9 11 13 15 17 22 28 32
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 23 28 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=0.89 $Y2=2.72
r46 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 22 31 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.547 $Y2=2.72
r48 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r49 17 28 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.89 $Y2=2.72
r50 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 15 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 11 31 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.5 $Y=2.635
+ $X2=2.547 $Y2=2.72
r54 11 13 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.5 $Y=2.635
+ $X2=2.5 $Y2=2
r55 7 28 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=2.635 $X2=0.89
+ $Y2=2.72
r56 7 9 10.6973 $w=7.08e-07 $l=6.35e-07 $layer=LI1_cond $X=0.89 $Y=2.635
+ $X2=0.89 $Y2=2
r57 2 13 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.485 $X2=2.5 $Y2=2
r58 1 9 150 $w=1.7e-07 $l=7.2832e-07 $layer=licon1_PDIFF $count=4 $X=0.565
+ $Y=1.485 $X2=1.08 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%VGND 1 2 9 11 15 17 19 26 27 30 33
r40 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r41 31 34 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r42 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r43 27 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r44 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r45 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.08
+ $Y2=0
r46 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.53
+ $Y2=0
r47 19 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r48 19 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r49 17 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r50 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r52 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.38
r53 12 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r54 11 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.08
+ $Y2=0
r55 11 12 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=1.995 $Y=0 $X2=0.765
+ $Y2=0
r56 7 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r57 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0.38
r58 2 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.235 $X2=2.08 $Y2=0.38
r59 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_1%A_297_47# 1 2 7 11 16
c30 16 0 1.80509e-19 $X=1.825 $Y=0.77
r31 14 16 8.06855 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=0.77
+ $X2=1.825 $Y2=0.77
r32 9 11 10.677 $w=3.38e-07 $l=3.15e-07 $layer=LI1_cond $X=2.505 $Y=0.715
+ $X2=2.505 $Y2=0.4
r33 7 9 7.55181 $w=1.9e-07 $l=2.1225e-07 $layer=LI1_cond $X=2.335 $Y=0.81
+ $X2=2.505 $Y2=0.715
r34 7 16 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=2.335 $Y=0.81
+ $X2=1.825 $Y2=0.81
r35 2 11 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.235 $X2=2.5 $Y2=0.4
r36 1 14 182 $w=1.7e-07 $l=5.65774e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.66 $Y2=0.72
.ends


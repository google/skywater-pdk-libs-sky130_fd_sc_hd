* File: sky130_fd_sc_hd__dlxbp_1.spice.pex
* Created: Thu Aug 27 14:18:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLXBP_1%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%A_27_47# 1 2 9 13 17 19 21 23 26 30 31 32 37
+ 40 42 45 46 49 52 53 57 62
c146 62 0 1.79706e-19 $X=2.735 $Y=1.43
c147 53 0 7.75336e-20 $X=2.64 $Y=1.53
c148 13 0 2.6965e-20 $X=0.89 $Y=2.135
c149 9 0 2.6965e-20 $X=0.89 $Y=0.445
r150 60 62 9.60507 $w=2.76e-07 $l=5.5e-08 $layer=POLY_cond $X=2.68 $Y=1.43
+ $X2=2.735 $Y2=1.43
r151 53 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.52 $X2=2.68 $Y2=1.52
r152 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.53
+ $X2=2.64 $Y2=1.53
r153 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r154 46 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r155 45 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=1.53
+ $X2=2.64 $Y2=1.53
r156 45 46 2.04826 $w=1.4e-07 $l=1.655e-06 $layer=MET1_cond $X=2.495 $Y=1.53
+ $X2=0.84 $Y2=1.53
r157 44 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r158 43 49 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r159 41 57 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r160 40 43 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r161 40 42 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r162 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r163 34 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r164 33 37 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r165 32 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r166 32 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r167 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r168 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r169 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r170 24 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r171 23 62 83.8261 $w=2.76e-07 $l=5.9397e-07 $layer=POLY_cond $X=3.215 $Y=1.175
+ $X2=2.735 $Y2=1.43
r172 22 23 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.215 $Y=0.785
+ $X2=3.215 $Y2=1.175
r173 19 22 28.5207 $w=1.69e-07 $l=1.16189e-07 $layer=POLY_cond $X=3.18 $Y=0.685
+ $X2=3.215 $Y2=0.785
r174 19 21 86.76 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.18 $Y=0.685
+ $X2=3.18 $Y2=0.415
r175 15 62 17.0164 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.735 $Y=1.685
+ $X2=2.735 $Y2=1.43
r176 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.735 $Y=1.685
+ $X2=2.735 $Y2=2.275
r177 11 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r178 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r179 7 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r180 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r181 2 37 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r182 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%D 2 3 5 8 11 14 17 19 22 23
c49 17 0 8.04072e-20 $X=1.84 $Y=1.615
r50 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.04 $X2=1.52 $Y2=1.04
r51 19 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.52 $Y=1.19
+ $X2=1.52 $Y2=1.04
r52 15 17 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.58 $Y=1.615
+ $X2=1.84 $Y2=1.615
r53 13 22 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=1.52 $Y=1.07 $X2=1.52
+ $Y2=1.04
r54 13 14 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.52 $Y=1.07
+ $X2=1.52 $Y2=1.205
r55 11 22 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.52 $Y=0.88
+ $X2=1.52 $Y2=1.04
r56 6 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.69 $X2=1.84
+ $Y2=1.615
r57 6 8 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.84 $Y=1.69 $X2=1.84
+ $Y2=2.165
r58 3 11 132.23 $w=1.13e-07 $l=3.1e-07 $layer=POLY_cond $X=1.83 $Y=0.805
+ $X2=1.52 $Y2=0.805
r59 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.73 $X2=1.83
+ $Y2=0.445
r60 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.58 $Y=1.54 $X2=1.58
+ $Y2=1.615
r61 2 14 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.58 $Y=1.54
+ $X2=1.58 $Y2=1.205
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%A_299_47# 1 2 9 13 17 19 20 29
c75 19 0 1.93267e-20 $X=1.985 $Y=1.235
r76 29 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.07
+ $X2=2.22 $Y2=1.235
r77 29 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.07
+ $X2=2.22 $Y2=0.905
r78 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.07 $X2=2.22 $Y2=1.07
r79 26 28 17.0374 $w=4.01e-07 $l=6.94781e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.922 $Y2=1.07
r80 19 28 6.52573 $w=4.01e-07 $l=1.93959e-07 $layer=LI1_cond $X=1.985 $Y=1.235
+ $X2=1.922 $Y2=1.07
r81 19 20 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=1.985 $Y=1.235
+ $X2=1.985 $Y2=1.495
r82 15 20 24.3348 $w=1.68e-07 $l=3.73e-07 $layer=LI1_cond $X=1.612 $Y=1.58
+ $X2=1.985 $Y2=1.58
r83 15 17 10.2615 $w=3.63e-07 $l=3.25e-07 $layer=LI1_cond $X=1.612 $Y=1.665
+ $X2=1.612 $Y2=1.99
r84 13 32 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.26 $Y=2.165
+ $X2=2.26 $Y2=1.235
r85 9 31 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.905
r86 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.505
+ $Y=1.845 $X2=1.63 $Y2=1.99
r87 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%A_193_47# 1 2 7 9 11 13 17 19 25 26 28 29 32
+ 35 41
c126 26 0 1.66933e-20 $X=1.127 $Y=1.797
c127 17 0 6.37139e-20 $X=1.1 $Y=0.51
c128 11 0 7.75336e-20 $X=3.165 $Y=1.88
r129 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.745 $X2=3.205 $Y2=1.745
r130 35 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.05 $Y=1.87
+ $X2=3.05 $Y2=1.87
r131 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r132 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r133 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.905 $Y=1.87
+ $X2=3.05 $Y2=1.87
r134 28 29 1.98638 $w=1.4e-07 $l=1.605e-06 $layer=MET1_cond $X=2.905 $Y=1.87
+ $X2=1.3 $Y2=1.87
r135 26 32 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r136 26 27 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r137 25 41 9.17136 $w=3.05e-07 $l=2.04915e-07 $layer=LI1_cond $X=3.05 $Y=1.575
+ $X2=3.127 $Y2=1.745
r138 24 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.05 $Y=1.065
+ $X2=3.05 $Y2=1.575
r139 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=0.91 $X2=2.75 $Y2=0.91
r140 19 24 8.02311 $w=3.6e-07 $l=2.18403e-07 $layer=LI1_cond $X=2.965 $Y=0.885
+ $X2=3.05 $Y2=1.065
r141 19 21 6.88265 $w=3.58e-07 $l=2.15e-07 $layer=LI1_cond $X=2.965 $Y=0.885
+ $X2=2.75 $Y2=0.885
r142 17 27 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r143 11 40 34.1986 $w=3.29e-07 $l=1.53704e-07 $layer=POLY_cond $X=3.165 $Y=1.88
+ $X2=3.205 $Y2=1.745
r144 11 13 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.165 $Y=1.88
+ $X2=3.165 $Y2=2.275
r145 7 22 40.7934 $w=3.34e-07 $l=1.8735e-07 $layer=POLY_cond $X=2.725 $Y=0.73
+ $X2=2.74 $Y2=0.91
r146 7 9 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.725 $Y=0.73
+ $X2=2.725 $Y2=0.415
r147 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r148 1 17 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%A_716_21# 1 2 9 13 15 17 20 22 24 26 28 31
+ 33 34 35 38 42 45 47 50 51 54 58 59
c116 24 0 6.83847e-20 $X=5.925 $Y=1.325
r117 54 56 7.79652 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.417 $Y=0.58
+ $X2=4.417 $Y2=0.745
r118 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.065
+ $Y=1.16 $X2=5.065 $Y2=1.16
r119 48 59 0.588983 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=4.55 $Y=1.16
+ $X2=4.447 $Y2=1.16
r120 48 50 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=4.55 $Y=1.16
+ $X2=5.065 $Y2=1.16
r121 47 58 7.66117 $w=2e-07 $l=1.79374e-07 $layer=LI1_cond $X=4.43 $Y=1.535
+ $X2=4.4 $Y2=1.7
r122 46 59 8.03064 $w=1.87e-07 $l=1.73292e-07 $layer=LI1_cond $X=4.43 $Y=1.325
+ $X2=4.447 $Y2=1.16
r123 46 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.43 $Y=1.325
+ $X2=4.43 $Y2=1.535
r124 45 59 8.03064 $w=1.87e-07 $l=1.65e-07 $layer=LI1_cond $X=4.447 $Y=0.995
+ $X2=4.447 $Y2=1.16
r125 45 56 13.5255 $w=2.03e-07 $l=2.5e-07 $layer=LI1_cond $X=4.447 $Y=0.995
+ $X2=4.447 $Y2=0.745
r126 40 58 7.66117 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=1.865 $X2=4.4
+ $Y2=1.7
r127 40 42 20.293 $w=2.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.4 $Y=1.865
+ $X2=4.4 $Y2=2.27
r128 38 60 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.905 $Y=1.7
+ $X2=3.655 $Y2=1.7
r129 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.905
+ $Y=1.7 $X2=3.905 $Y2=1.7
r130 35 58 0.381419 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=4.285 $Y=1.7
+ $X2=4.4 $Y2=1.7
r131 35 37 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=4.285 $Y=1.7
+ $X2=3.905 $Y2=1.7
r132 33 34 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.94 $Y=1.62
+ $X2=5.94 $Y2=1.77
r133 31 34 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.955 $Y=2.165
+ $X2=5.955 $Y2=1.77
r134 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.955 $Y=0.73
+ $X2=5.955 $Y2=0.445
r135 24 33 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.925 $Y=1.325
+ $X2=5.925 $Y2=1.62
r136 23 51 5.03009 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.09 $Y=1.16 $X2=5.01
+ $Y2=1.16
r137 22 24 50.6561 $w=1.57e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.94 $Y=1.16
+ $X2=5.925 $Y2=1.325
r138 22 26 132.013 $w=1.57e-07 $l=4.37436e-07 $layer=POLY_cond $X=5.94 $Y=1.16
+ $X2=5.955 $Y2=0.73
r139 22 23 132.895 $w=3.3e-07 $l=7.6e-07 $layer=POLY_cond $X=5.85 $Y=1.16
+ $X2=5.09 $Y2=1.16
r140 18 51 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=5.015 $Y=1.325
+ $X2=5.01 $Y2=1.16
r141 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.015 $Y=1.325
+ $X2=5.015 $Y2=1.985
r142 15 51 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=5.015 $Y=0.995
+ $X2=5.01 $Y2=1.16
r143 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.015 $Y=0.995
+ $X2=5.015 $Y2=0.56
r144 11 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.865
+ $X2=3.655 $Y2=1.7
r145 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.655 $Y=1.865
+ $X2=3.655 $Y2=2.275
r146 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.535
+ $X2=3.655 $Y2=1.7
r147 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.655 $Y=1.535
+ $X2=3.655 $Y2=0.445
r148 2 58 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.26
+ $Y=1.485 $X2=4.385 $Y2=1.755
r149 2 42 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.26
+ $Y=1.485 $X2=4.385 $Y2=2.27
r150 1 54 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.235 $X2=4.385 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%A_560_47# 1 2 7 9 12 14 15 16 20 25 27 29 30
+ 32
c91 30 0 1.45945e-19 $X=3.65 $Y=1.16
c92 20 0 1.60379e-19 $X=3.305 $Y=0.45
c93 15 0 1.26483e-19 $X=4.595 $Y=1.16
r94 35 36 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=1.16
+ $X2=3.555 $Y2=1.16
r95 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.16 $X2=4.09 $Y2=1.16
r96 30 36 4.12602 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.65 $Y=1.16
+ $X2=3.555 $Y2=1.16
r97 30 32 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.65 $Y=1.16
+ $X2=4.09 $Y2=1.16
r98 28 36 2.53051 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=1.325
+ $X2=3.555 $Y2=1.16
r99 28 29 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=3.555 $Y=1.325
+ $X2=3.555 $Y2=1.995
r100 26 29 5.3907 $w=2.15e-07 $l=1.12406e-07 $layer=LI1_cond $X=3.517 $Y=2.09
+ $X2=3.555 $Y2=1.995
r101 26 27 9.89189 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.517 $Y=2.09
+ $X2=3.517 $Y2=2.255
r102 25 35 3.17874 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=0.995
+ $X2=3.39 $Y2=1.16
r103 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.39 $Y=0.535
+ $X2=3.39 $Y2=0.995
r104 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.305 $Y=0.45
+ $X2=3.39 $Y2=0.535
r105 20 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.305 $Y=0.45
+ $X2=2.97 $Y2=0.45
r106 16 27 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.425 $Y=2.34
+ $X2=3.517 $Y2=2.255
r107 16 18 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.425 $Y=2.34
+ $X2=2.95 $Y2=2.34
r108 14 33 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.52 $Y=1.16
+ $X2=4.09 $Y2=1.16
r109 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.52 $Y=1.16
+ $X2=4.595 $Y2=1.16
r110 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=1.325
+ $X2=4.595 $Y2=1.16
r111 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.595 $Y=1.325
+ $X2=4.595 $Y2=1.985
r112 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=0.995
+ $X2=4.595 $Y2=1.16
r113 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.595 $Y=0.995
+ $X2=4.595 $Y2=0.56
r114 2 18 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.065 $X2=2.95 $Y2=2.34
r115 1 22 182 $w=1.7e-07 $l=2.87706e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.97 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%A_1124_47# 1 2 9 12 16 20 24 25 27 29
r48 25 30 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=6.357 $Y=1.16
+ $X2=6.357 $Y2=1.325
r49 25 29 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=6.357 $Y=1.16
+ $X2=6.357 $Y2=0.995
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.345
+ $Y=1.16 $X2=6.345 $Y2=1.16
r51 22 27 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.91 $Y=1.16
+ $X2=5.785 $Y2=1.16
r52 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.91 $Y=1.16
+ $X2=6.345 $Y2=1.16
r53 18 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=1.325
+ $X2=5.785 $Y2=1.16
r54 18 20 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=5.785 $Y=1.325
+ $X2=5.785 $Y2=2.165
r55 14 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0.995
+ $X2=5.785 $Y2=1.16
r56 14 16 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=5.785 $Y=0.995
+ $X2=5.785 $Y2=0.51
r57 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.985
+ $X2=6.43 $Y2=1.325
r58 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.56 $X2=6.43
+ $Y2=0.995
r59 2 20 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=1.845 $X2=5.745 $Y2=2.165
r60 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=5.62
+ $Y=0.235 $X2=5.745 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 39 41 46
+ 58 62 69 70 73 76 79 82
r105 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r106 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r107 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r108 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r109 70 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r110 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r111 67 82 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.237 $Y2=2.72
r112 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.67 $Y2=2.72
r113 66 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 66 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r115 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r116 63 79 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.97 $Y=2.72
+ $X2=4.827 $Y2=2.72
r117 63 65 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.97 $Y=2.72
+ $X2=5.75 $Y2=2.72
r118 62 82 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=6.237 $Y2=2.72
r119 62 65 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 61 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r122 58 79 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.685 $Y=2.72
+ $X2=4.827 $Y2=2.72
r123 58 60 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.685 $Y=2.72
+ $X2=4.37 $Y2=2.72
r124 57 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r127 54 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r128 53 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r130 51 76 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.245 $Y=2.72
+ $X2=2.105 $Y2=2.72
r131 51 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=2.72
+ $X2=2.53 $Y2=2.72
r132 50 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r133 50 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 47 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r136 47 49 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 46 76 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.965 $Y=2.72
+ $X2=2.105 $Y2=2.72
r138 46 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.965 $Y=2.72
+ $X2=1.61 $Y2=2.72
r139 41 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r140 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r141 39 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r142 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r143 37 56 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.45 $Y2=2.72
r144 37 38 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.78 $Y=2.72 $X2=3.88
+ $Y2=2.72
r145 36 60 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.98 $Y=2.72
+ $X2=4.37 $Y2=2.72
r146 36 38 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.98 $Y=2.72 $X2=3.88
+ $Y2=2.72
r147 32 82 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.237 $Y=2.635
+ $X2=6.237 $Y2=2.72
r148 32 34 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=6.237 $Y=2.635
+ $X2=6.237 $Y2=2
r149 28 79 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.827 $Y=2.635
+ $X2=4.827 $Y2=2.72
r150 28 30 36.3929 $w=2.83e-07 $l=9e-07 $layer=LI1_cond $X=4.827 $Y=2.635
+ $X2=4.827 $Y2=1.735
r151 24 38 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.72
r152 24 26 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.34
r153 20 76 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2.72
r154 20 22 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2
r155 16 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r156 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r157 5 34 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=6.03
+ $Y=1.845 $X2=6.22 $Y2=2
r158 4 30 300 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=2 $X=4.67
+ $Y=1.485 $X2=4.805 $Y2=1.735
r159 3 26 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=2.065 $X2=3.865 $Y2=2.34
r160 2 22 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.915
+ $Y=1.845 $X2=2.05 $Y2=2
r161 1 18 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%Q 1 2 10 11 12 13 19 25 31
c28 31 0 1.26483e-19 $X=5.315 $Y=1.67
r29 23 25 0.823174 $w=3.48e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=1.845
+ $X2=5.315 $Y2=1.87
r30 12 23 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=5.315 $Y=1.815
+ $X2=5.315 $Y2=1.845
r31 12 31 7.82994 $w=3.48e-07 $l=1.45e-07 $layer=LI1_cond $X=5.315 $Y=1.815
+ $X2=5.315 $Y2=1.67
r32 12 13 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=5.315 $Y=1.9
+ $X2=5.315 $Y2=2.21
r33 12 25 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=5.315 $Y=1.9
+ $X2=5.315 $Y2=1.87
r34 11 19 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=5.315 $Y=0.51
+ $X2=5.315 $Y2=0.42
r35 10 31 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.405 $Y=0.82
+ $X2=5.405 $Y2=1.67
r36 9 11 4.44514 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.315 $Y=0.645
+ $X2=5.315 $Y2=0.51
r37 9 10 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=5.315 $Y=0.645
+ $X2=5.315 $Y2=0.82
r38 2 12 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.09
+ $Y=1.485 $X2=5.225 $Y2=1.835
r39 1 19 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.235 $X2=5.225 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%Q_N 1 2 10 11 12 13 14 15
r16 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=6.685 $Y=1.82
+ $X2=6.685 $Y2=2.21
r17 11 14 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=6.685 $Y=1.575
+ $X2=6.685 $Y2=1.82
r18 11 12 6.14153 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=6.685 $Y=1.575
+ $X2=6.685 $Y2=1.445
r19 10 12 33.2332 $w=2.13e-07 $l=6.2e-07 $layer=LI1_cond $X=6.707 $Y=0.825
+ $X2=6.707 $Y2=1.445
r20 9 13 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=6.685 $Y=0.695
+ $X2=6.685 $Y2=0.51
r21 9 10 6.14153 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=6.685 $Y=0.695
+ $X2=6.685 $Y2=0.825
r22 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=6.505
+ $Y=1.485 $X2=6.64 $Y2=1.82
r23 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.64 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBP_1%VGND 1 2 3 4 5 18 22 26 30 34 36 38 43 48 56
+ 61 68 69 72 75 78 81 84
c102 69 0 2.71124e-20 $X=6.67 $Y=0
c103 61 0 6.83847e-20 $X=6.09 $Y=0
r104 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r105 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r106 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r107 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r108 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r109 69 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r110 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r111 66 84 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.237 $Y2=0
r112 66 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.67 $Y2=0
r113 65 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r114 65 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=4.83
+ $Y2=0
r115 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r116 62 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.97 $Y=0 $X2=4.845
+ $Y2=0
r117 62 64 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.97 $Y=0 $X2=5.75
+ $Y2=0
r118 61 84 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=6.237
+ $Y2=0
r119 61 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=5.75
+ $Y2=0
r120 60 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r121 60 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r122 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r123 57 78 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.045 $Y=0
+ $X2=3.872 $Y2=0
r124 57 59 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.045 $Y=0
+ $X2=4.37 $Y2=0
r125 56 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=4.845
+ $Y2=0
r126 56 59 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=4.37
+ $Y2=0
r127 55 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r128 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r129 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r130 52 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r131 51 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r132 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r133 49 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r134 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r135 48 78 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.872
+ $Y2=0
r136 48 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.45
+ $Y2=0
r137 47 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r138 47 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r139 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r140 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r141 44 46 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r142 43 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r143 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r144 38 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r145 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r146 36 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r147 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r148 32 84 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.237 $Y=0.085
+ $X2=6.237 $Y2=0
r149 32 34 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=6.237 $Y=0.085
+ $X2=6.237 $Y2=0.38
r150 28 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.845 $Y=0.085
+ $X2=4.845 $Y2=0
r151 28 30 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.845 $Y=0.085
+ $X2=4.845 $Y2=0.55
r152 24 78 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.872 $Y=0.085
+ $X2=3.872 $Y2=0
r153 24 26 12.0255 $w=3.43e-07 $l=3.6e-07 $layer=LI1_cond $X=3.872 $Y=0.085
+ $X2=3.872 $Y2=0.445
r154 20 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r155 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r156 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r157 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r158 5 34 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=6.03
+ $Y=0.235 $X2=6.22 $Y2=0.38
r159 4 30 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.235 $X2=4.805 $Y2=0.55
r160 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.865 $Y2=0.445
r161 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r162 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


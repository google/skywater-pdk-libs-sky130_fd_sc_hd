* File: sky130_fd_sc_hd__nor3b_2.pxi.spice
* Created: Thu Aug 27 14:32:27 2020
* 
x_PM_SKY130_FD_SC_HD__NOR3B_2%A N_A_c_71_n N_A_M1004_g N_A_M1001_g N_A_c_72_n
+ N_A_M1006_g N_A_M1012_g A A N_A_c_74_n PM_SKY130_FD_SC_HD__NOR3B_2%A
x_PM_SKY130_FD_SC_HD__NOR3B_2%B N_B_c_111_n N_B_M1002_g N_B_M1008_g N_B_c_112_n
+ N_B_M1005_g N_B_M1009_g B B B N_B_c_114_n PM_SKY130_FD_SC_HD__NOR3B_2%B
x_PM_SKY130_FD_SC_HD__NOR3B_2%A_531_21# N_A_531_21#_M1011_s N_A_531_21#_M1013_s
+ N_A_531_21#_c_156_n N_A_531_21#_M1007_g N_A_531_21#_M1000_g
+ N_A_531_21#_c_157_n N_A_531_21#_M1010_g N_A_531_21#_M1003_g
+ N_A_531_21#_c_158_n N_A_531_21#_c_159_n N_A_531_21#_c_160_n
+ N_A_531_21#_c_161_n N_A_531_21#_c_162_n N_A_531_21#_c_167_n
+ N_A_531_21#_c_163_n PM_SKY130_FD_SC_HD__NOR3B_2%A_531_21#
x_PM_SKY130_FD_SC_HD__NOR3B_2%C_N N_C_N_M1011_g N_C_N_M1013_g C_N N_C_N_c_219_n
+ N_C_N_c_220_n PM_SKY130_FD_SC_HD__NOR3B_2%C_N
x_PM_SKY130_FD_SC_HD__NOR3B_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1012_s
+ N_A_27_297#_M1009_d N_A_27_297#_c_245_n N_A_27_297#_c_246_n
+ N_A_27_297#_c_247_n N_A_27_297#_c_265_p N_A_27_297#_c_248_n
+ N_A_27_297#_c_249_n N_A_27_297#_c_250_n PM_SKY130_FD_SC_HD__NOR3B_2%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR3B_2%VPWR N_VPWR_M1001_d N_VPWR_M1013_d N_VPWR_c_281_n
+ N_VPWR_c_282_n N_VPWR_c_283_n VPWR N_VPWR_c_284_n N_VPWR_c_285_n
+ N_VPWR_c_286_n N_VPWR_c_280_n PM_SKY130_FD_SC_HD__NOR3B_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR3B_2%A_281_297# N_A_281_297#_M1008_s
+ N_A_281_297#_M1000_d N_A_281_297#_M1003_d N_A_281_297#_c_346_n
+ N_A_281_297#_c_331_n N_A_281_297#_c_356_n N_A_281_297#_c_332_n
+ N_A_281_297#_c_338_n N_A_281_297#_c_360_n N_A_281_297#_c_333_n
+ N_A_281_297#_c_362_n PM_SKY130_FD_SC_HD__NOR3B_2%A_281_297#
x_PM_SKY130_FD_SC_HD__NOR3B_2%Y N_Y_M1004_s N_Y_M1002_d N_Y_M1007_d N_Y_M1000_s
+ N_Y_c_375_n N_Y_c_368_n N_Y_c_369_n N_Y_c_383_n N_Y_c_370_n N_Y_c_371_n
+ N_Y_c_372_n N_Y_c_373_n Y N_Y_c_408_n PM_SKY130_FD_SC_HD__NOR3B_2%Y
x_PM_SKY130_FD_SC_HD__NOR3B_2%VGND N_VGND_M1004_d N_VGND_M1006_d N_VGND_M1005_s
+ N_VGND_M1007_s N_VGND_M1010_s N_VGND_M1011_d N_VGND_c_439_n N_VGND_c_440_n
+ N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n VGND N_VGND_c_449_n
+ N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n PM_SKY130_FD_SC_HD__NOR3B_2%VGND
cc_1 VNB N_A_c_71_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_72_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB A 0.0163753f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_A_c_74_n 0.0382849f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_5 VNB N_B_c_111_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_112_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_7 VNB B 0.0321129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_c_114_n 0.0369647f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_9 VNB N_A_531_21#_c_156_n 0.0214626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_531_21#_c_157_n 0.0196608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_531_21#_c_158_n 0.0108596f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_12 VNB N_A_531_21#_c_159_n 0.0595483f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_13 VNB N_A_531_21#_c_160_n 0.00431685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_531_21#_c_161_n 0.0132286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_531_21#_c_162_n 0.00241416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_531_21#_c_163_n 4.68721e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB C_N 0.0161743f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_18 VNB N_C_N_c_219_n 0.0303785f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.325
cc_19 VNB N_C_N_c_220_n 0.0213916f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_20 VNB N_VPWR_c_280_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_368_n 0.00338427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_369_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_370_n 0.0126676f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_24 VNB N_Y_c_371_n 0.00166887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_372_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_373_n 8.10088e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_439_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_28 VNB N_VGND_c_440_n 0.0330578f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_29 VNB N_VGND_c_441_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_442_n 0.00579864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_443_n 0.0108094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_444_n 0.0348044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_445_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_446_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_447_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_448_n 0.0039398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_449_n 0.0207255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_450_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_451_n 0.0272921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_452_n 0.250926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VPB N_A_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_42 VPB N_A_M1012_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_43 VPB N_A_c_74_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_44 VPB N_B_M1008_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_45 VPB N_B_M1009_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_46 VPB N_B_c_114_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_47 VPB N_A_531_21#_M1000_g 0.0251579f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_48 VPB N_A_531_21#_M1003_g 0.0226362f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_49 VPB N_A_531_21#_c_159_n 0.015261f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_50 VPB N_A_531_21#_c_167_n 0.00981377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_531_21#_c_163_n 0.0039256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_C_N_M1013_g 0.0275674f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_53 VPB N_C_N_c_219_n 0.00551023f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.325
cc_54 VPB N_A_27_297#_c_245_n 0.0103851f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_55 VPB N_A_27_297#_c_246_n 0.0327764f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_56 VPB N_A_27_297#_c_247_n 0.00240493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_297#_c_248_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_297#_c_249_n 0.00322557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_297#_c_250_n 0.00269081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_281_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_61 VPB N_VPWR_c_282_n 0.0112901f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.325
cc_62 VPB N_VPWR_c_283_n 0.048603f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_63 VPB N_VPWR_c_284_n 0.0174963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_285_n 0.0856517f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_65 VPB N_VPWR_c_286_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_280_n 0.0643375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_281_297#_c_331_n 0.0128284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_281_297#_c_332_n 0.00319238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_281_297#_c_333_n 0.00205686f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_70 VPB N_Y_c_371_n 0.00277404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_A_c_72_n N_B_c_111_n 0.0194931f $X=0.91 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_72 N_A_M1012_g N_B_M1008_g 0.0194931f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_73 A B 0.0185436f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_74_n B 0.00160637f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_75 A N_B_c_114_n 2.03927e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_74_n N_B_c_114_n 0.0194931f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_77 A N_A_27_297#_c_245_n 0.0252798f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_A_27_297#_c_247_n 0.0135215f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1012_g N_A_27_297#_c_247_n 0.0135117f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_80 A N_A_27_297#_c_247_n 0.0396361f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_c_74_n N_A_27_297#_c_247_n 0.00211509f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_M1001_g N_VPWR_c_281_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_M1012_g N_VPWR_c_281_n 0.00302074f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1001_g N_VPWR_c_284_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1012_g N_VPWR_c_285_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_VPWR_c_280_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1012_g N_VPWR_c_280_n 0.010464f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_c_71_n N_Y_c_375_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_c_72_n N_Y_c_375_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_c_72_n N_Y_c_368_n 0.00890517f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_91 A N_Y_c_368_n 0.00688575f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A_c_71_n N_Y_c_369_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_72_n N_Y_c_369_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_94 A N_Y_c_369_n 0.0266272f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_c_74_n N_Y_c_369_n 0.00230339f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_c_72_n N_Y_c_383_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_c_71_n N_VGND_c_440_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_98 A N_VGND_c_440_n 0.0217663f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_99 N_A_c_72_n N_VGND_c_441_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_c_71_n N_VGND_c_445_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_c_72_n N_VGND_c_445_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_c_71_n N_VGND_c_452_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_c_72_n N_VGND_c_452_n 0.0057435f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_104 B N_A_531_21#_c_159_n 0.00686059f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_105 N_B_M1008_g N_A_27_297#_c_248_n 0.0132199f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B_M1009_g N_A_27_297#_c_248_n 0.0112055f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_107 B N_A_27_297#_c_248_n 0.0417417f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B_c_114_n N_A_27_297#_c_248_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_109 B N_A_27_297#_c_249_n 0.00942636f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_110 B N_A_27_297#_c_250_n 0.0213978f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B_M1008_g N_VPWR_c_285_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B_M1009_g N_VPWR_c_285_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B_M1008_g N_VPWR_c_280_n 0.0106871f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B_M1009_g N_VPWR_c_280_n 0.00660224f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B_M1009_g N_A_281_297#_c_331_n 0.0119904f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B_M1009_g N_A_281_297#_c_332_n 0.00518348f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_117 B N_A_281_297#_c_332_n 0.0226233f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B_c_111_n N_Y_c_375_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B_c_111_n N_Y_c_368_n 0.00865686f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_120 B N_Y_c_368_n 0.0174927f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_121 N_B_c_111_n N_Y_c_383_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_112_n N_Y_c_383_n 0.0109565f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_112_n N_Y_c_370_n 0.0109318f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_124 B N_Y_c_370_n 0.0709093f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_125 B N_Y_c_371_n 0.0168399f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B_c_111_n N_Y_c_372_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_112_n N_Y_c_372_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_128 B N_Y_c_372_n 0.0266272f $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B_c_114_n N_Y_c_372_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_c_111_n N_VGND_c_441_n 0.00146339f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B_c_111_n N_VGND_c_450_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B_c_112_n N_VGND_c_450_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B_c_112_n N_VGND_c_451_n 0.00336547f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B_c_111_n N_VGND_c_452_n 0.0057435f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B_c_112_n N_VGND_c_452_n 0.0070399f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_531_21#_c_167_n N_C_N_M1013_g 0.00181686f $X=3.92 $Y=1.705 $X2=0
+ $Y2=0
cc_137 N_A_531_21#_c_159_n C_N 4.4116e-19 $X=3.4 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_531_21#_c_161_n C_N 0.0011748f $X=3.92 $Y=0.66 $X2=0 $Y2=0
cc_139 N_A_531_21#_c_162_n C_N 0.01888f $X=3.775 $Y=1.18 $X2=0 $Y2=0
cc_140 N_A_531_21#_c_167_n C_N 0.00115298f $X=3.92 $Y=1.705 $X2=0 $Y2=0
cc_141 N_A_531_21#_c_159_n N_C_N_c_219_n 0.00583755f $X=3.4 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_531_21#_c_162_n N_C_N_c_219_n 8.90581e-19 $X=3.775 $Y=1.18 $X2=0
+ $Y2=0
cc_143 N_A_531_21#_c_163_n N_C_N_c_219_n 0.00520599f $X=3.867 $Y=1.455 $X2=0
+ $Y2=0
cc_144 N_A_531_21#_c_160_n N_C_N_c_220_n 0.00479675f $X=3.775 $Y=1.075 $X2=0
+ $Y2=0
cc_145 N_A_531_21#_c_161_n N_C_N_c_220_n 0.00348716f $X=3.92 $Y=0.66 $X2=0 $Y2=0
cc_146 N_A_531_21#_M1000_g N_VPWR_c_285_n 0.00357877f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_531_21#_M1003_g N_VPWR_c_285_n 0.00357877f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_531_21#_M1000_g N_VPWR_c_280_n 0.00655123f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_531_21#_M1003_g N_VPWR_c_280_n 0.00655123f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_531_21#_c_167_n N_VPWR_c_280_n 0.0133729f $X=3.92 $Y=1.705 $X2=0
+ $Y2=0
cc_151 N_A_531_21#_M1000_g N_A_281_297#_c_332_n 7.02661e-19 $X=2.73 $Y=1.985
+ $X2=0 $Y2=0
cc_152 N_A_531_21#_M1000_g N_A_281_297#_c_338_n 0.0121306f $X=2.73 $Y=1.985
+ $X2=0 $Y2=0
cc_153 N_A_531_21#_M1003_g N_A_281_297#_c_338_n 0.0121747f $X=3.15 $Y=1.985
+ $X2=0 $Y2=0
cc_154 N_A_531_21#_M1003_g N_A_281_297#_c_333_n 7.0048e-19 $X=3.15 $Y=1.985
+ $X2=0 $Y2=0
cc_155 N_A_531_21#_c_158_n N_A_281_297#_c_333_n 0.0198783f $X=3.69 $Y=1.18 $X2=0
+ $Y2=0
cc_156 N_A_531_21#_c_159_n N_A_281_297#_c_333_n 0.0059411f $X=3.4 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A_531_21#_c_167_n N_A_281_297#_c_333_n 0.0287257f $X=3.92 $Y=1.705
+ $X2=0 $Y2=0
cc_158 N_A_531_21#_c_156_n N_Y_c_370_n 0.0145972f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_531_21#_c_156_n N_Y_c_371_n 0.00240809f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_531_21#_M1000_g N_Y_c_371_n 0.00374435f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_531_21#_c_157_n N_Y_c_371_n 0.0012881f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_531_21#_M1003_g N_Y_c_371_n 0.0021084f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_531_21#_c_158_n N_Y_c_371_n 0.0161652f $X=3.69 $Y=1.18 $X2=0 $Y2=0
cc_164 N_A_531_21#_c_159_n N_Y_c_371_n 0.0248813f $X=3.4 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_531_21#_c_160_n N_Y_c_371_n 0.00491768f $X=3.775 $Y=1.075 $X2=0 $Y2=0
cc_166 N_A_531_21#_c_163_n N_Y_c_371_n 0.00508546f $X=3.867 $Y=1.455 $X2=0 $Y2=0
cc_167 N_A_531_21#_c_156_n N_Y_c_373_n 0.00221107f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_531_21#_c_157_n N_Y_c_373_n 0.00380639f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_531_21#_c_161_n N_Y_c_373_n 3.29695e-19 $X=3.92 $Y=0.66 $X2=0 $Y2=0
cc_170 N_A_531_21#_c_156_n N_Y_c_408_n 0.0109565f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_531_21#_c_157_n N_Y_c_408_n 0.00539651f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_531_21#_c_157_n N_VGND_c_442_n 0.00340487f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_531_21#_c_158_n N_VGND_c_442_n 0.0159069f $X=3.69 $Y=1.18 $X2=0 $Y2=0
cc_174 N_A_531_21#_c_159_n N_VGND_c_442_n 0.00518707f $X=3.4 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_531_21#_c_161_n N_VGND_c_442_n 0.0351611f $X=3.92 $Y=0.66 $X2=0 $Y2=0
cc_176 N_A_531_21#_c_161_n N_VGND_c_444_n 0.00696062f $X=3.92 $Y=0.66 $X2=0
+ $Y2=0
cc_177 N_A_531_21#_c_156_n N_VGND_c_447_n 0.00423334f $X=2.73 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_531_21#_c_157_n N_VGND_c_447_n 0.00541359f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_A_531_21#_c_161_n N_VGND_c_449_n 0.0139405f $X=3.92 $Y=0.66 $X2=0 $Y2=0
cc_180 N_A_531_21#_c_156_n N_VGND_c_451_n 0.00336547f $X=2.73 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_531_21#_c_156_n N_VGND_c_452_n 0.0070399f $X=2.73 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_531_21#_c_157_n N_VGND_c_452_n 0.0108276f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_531_21#_c_161_n N_VGND_c_452_n 0.0126218f $X=3.92 $Y=0.66 $X2=0 $Y2=0
cc_184 N_C_N_M1013_g N_VPWR_c_283_n 0.00563018f $X=4.13 $Y=1.695 $X2=0 $Y2=0
cc_185 C_N N_VPWR_c_283_n 0.0135493f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_186 N_C_N_c_219_n N_VPWR_c_283_n 0.00247431f $X=4.195 $Y=1.16 $X2=0 $Y2=0
cc_187 N_C_N_M1013_g N_VPWR_c_285_n 0.00327927f $X=4.13 $Y=1.695 $X2=0 $Y2=0
cc_188 N_C_N_M1013_g N_VPWR_c_280_n 0.00417489f $X=4.13 $Y=1.695 $X2=0 $Y2=0
cc_189 N_C_N_M1013_g N_A_281_297#_c_333_n 0.00411678f $X=4.13 $Y=1.695 $X2=0
+ $Y2=0
cc_190 N_C_N_c_220_n N_VGND_c_442_n 0.00172213f $X=4.192 $Y=0.995 $X2=0 $Y2=0
cc_191 C_N N_VGND_c_444_n 0.0163628f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_192 N_C_N_c_219_n N_VGND_c_444_n 0.0026033f $X=4.195 $Y=1.16 $X2=0 $Y2=0
cc_193 N_C_N_c_220_n N_VGND_c_444_n 0.00395899f $X=4.192 $Y=0.995 $X2=0 $Y2=0
cc_194 N_C_N_c_220_n N_VGND_c_449_n 0.00510437f $X=4.192 $Y=0.995 $X2=0 $Y2=0
cc_195 N_C_N_c_220_n N_VGND_c_452_n 0.00512902f $X=4.192 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_247_n N_VPWR_M1001_d 0.00165831f $X=0.995 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_197 N_A_27_297#_c_247_n N_VPWR_c_281_n 0.0126919f $X=0.995 $Y=1.54 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_246_n N_VPWR_c_284_n 0.0204682f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_199 N_A_27_297#_c_265_p N_VPWR_c_285_n 0.0142343f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_200 N_A_27_297#_M1001_s N_VPWR_c_280_n 0.00260431f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_M1012_s N_VPWR_c_280_n 0.00284632f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_202 N_A_27_297#_M1009_d N_VPWR_c_280_n 0.00226545f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_246_n N_VPWR_c_280_n 0.0120542f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_204 N_A_27_297#_c_265_p N_VPWR_c_280_n 0.00955092f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_205 N_A_27_297#_c_248_n N_A_281_297#_M1008_s 0.00165831f $X=1.835 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_206 N_A_27_297#_c_248_n N_A_281_297#_c_346_n 0.0126766f $X=1.835 $Y=1.54
+ $X2=0 $Y2=0
cc_207 N_A_27_297#_M1009_d N_A_281_297#_c_331_n 0.00593473f $X=1.825 $Y=1.485
+ $X2=0 $Y2=0
cc_208 N_A_27_297#_c_248_n N_A_281_297#_c_331_n 0.00320918f $X=1.835 $Y=1.54
+ $X2=0 $Y2=0
cc_209 N_A_27_297#_c_250_n N_A_281_297#_c_331_n 0.0153739f $X=1.96 $Y=1.62 $X2=0
+ $Y2=0
cc_210 N_A_27_297#_c_250_n N_A_281_297#_c_332_n 0.035828f $X=1.96 $Y=1.62 $X2=0
+ $Y2=0
cc_211 N_A_27_297#_c_247_n N_Y_c_368_n 8.37688e-19 $X=0.995 $Y=1.54 $X2=0 $Y2=0
cc_212 N_A_27_297#_c_249_n N_Y_c_368_n 0.00524452f $X=1.12 $Y=1.62 $X2=0 $Y2=0
cc_213 N_A_27_297#_c_245_n N_VGND_c_440_n 7.84254e-19 $X=0.247 $Y=1.625 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_280_n N_A_281_297#_M1008_s 0.00246446f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_215 N_VPWR_c_280_n N_A_281_297#_M1000_d 0.00225716f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_280_n N_A_281_297#_M1003_d 0.00312505f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_285_n N_A_281_297#_c_331_n 0.0430664f $X=4.215 $Y=2.72 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_280_n N_A_281_297#_c_331_n 0.0256842f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_285_n N_A_281_297#_c_356_n 0.0142933f $X=4.215 $Y=2.72 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_280_n N_A_281_297#_c_356_n 0.00962421f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_285_n N_A_281_297#_c_338_n 0.0330174f $X=4.215 $Y=2.72 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_280_n N_A_281_297#_c_338_n 0.0204627f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_285_n N_A_281_297#_c_360_n 0.0155563f $X=4.215 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_280_n N_A_281_297#_c_360_n 0.00942493f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_285_n N_A_281_297#_c_362_n 0.0173143f $X=4.215 $Y=2.72 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_280_n N_A_281_297#_c_362_n 0.0103877f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_280_n N_Y_M1000_s 0.00216833f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_228 N_A_281_297#_c_338_n N_Y_M1000_s 0.00312348f $X=3.235 $Y=2.38 $X2=0 $Y2=0
cc_229 N_A_281_297#_c_332_n N_Y_c_371_n 0.00232727f $X=2.52 $Y=1.62 $X2=0 $Y2=0
cc_230 N_A_281_297#_c_338_n N_Y_c_371_n 0.0118865f $X=3.235 $Y=2.38 $X2=0 $Y2=0
cc_231 N_A_281_297#_c_333_n N_Y_c_371_n 0.00231016f $X=3.36 $Y=1.62 $X2=0 $Y2=0
cc_232 N_Y_c_368_n N_VGND_M1006_d 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_233 N_Y_c_370_n N_VGND_M1005_s 0.00281828f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_234 N_Y_c_370_n N_VGND_M1007_s 0.00281828f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_235 N_Y_c_369_n N_VGND_c_440_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_236 N_Y_c_368_n N_VGND_c_441_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_237 N_Y_c_373_n N_VGND_c_442_n 0.00751095f $X=2.94 $Y=0.815 $X2=0 $Y2=0
cc_238 N_Y_c_375_n N_VGND_c_445_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_239 N_Y_c_368_n N_VGND_c_445_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_240 N_Y_c_370_n N_VGND_c_447_n 0.00198695f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_241 N_Y_c_408_n N_VGND_c_447_n 0.0188914f $X=2.94 $Y=0.39 $X2=0 $Y2=0
cc_242 N_Y_c_368_n N_VGND_c_450_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_243 N_Y_c_383_n N_VGND_c_450_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_244 N_Y_c_370_n N_VGND_c_450_n 0.00198695f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_245 N_Y_c_370_n N_VGND_c_451_n 0.0568906f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_246 N_Y_M1004_s N_VGND_c_452_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_247 N_Y_M1002_d N_VGND_c_452_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_248 N_Y_M1007_d N_VGND_c_452_n 0.00215201f $X=2.805 $Y=0.235 $X2=0 $Y2=0
cc_249 N_Y_c_375_n N_VGND_c_452_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_250 N_Y_c_368_n N_VGND_c_452_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_251 N_Y_c_383_n N_VGND_c_452_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_252 N_Y_c_370_n N_VGND_c_452_n 0.0104789f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_253 N_Y_c_408_n N_VGND_c_452_n 0.0122184f $X=2.94 $Y=0.39 $X2=0 $Y2=0

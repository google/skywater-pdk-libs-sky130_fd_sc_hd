* File: sky130_fd_sc_hd__o41a_4.pxi.spice
* Created: Tue Sep  1 19:26:33 2020
* 
x_PM_SKY130_FD_SC_HD__O41A_4%A_79_21# N_A_79_21#_M1014_s N_A_79_21#_M1004_s
+ N_A_79_21#_M1006_s N_A_79_21#_M1013_g N_A_79_21#_M1001_g N_A_79_21#_M1018_g
+ N_A_79_21#_M1005_g N_A_79_21#_M1019_g N_A_79_21#_M1020_g N_A_79_21#_M1025_g
+ N_A_79_21#_M1023_g N_A_79_21#_c_136_n N_A_79_21#_c_137_n N_A_79_21#_c_148_p
+ N_A_79_21#_c_144_n N_A_79_21#_c_138_n N_A_79_21#_c_145_n N_A_79_21#_c_139_n
+ PM_SKY130_FD_SC_HD__O41A_4%A_79_21#
x_PM_SKY130_FD_SC_HD__O41A_4%B1 N_B1_M1004_g N_B1_c_255_n N_B1_c_256_n
+ N_B1_M1021_g N_B1_M1014_g N_B1_M1015_g B1 N_B1_c_260_n
+ PM_SKY130_FD_SC_HD__O41A_4%B1
x_PM_SKY130_FD_SC_HD__O41A_4%A4 N_A4_M1002_g N_A4_M1006_g N_A4_M1026_g
+ N_A4_M1010_g A4 A4 N_A4_c_310_n PM_SKY130_FD_SC_HD__O41A_4%A4
x_PM_SKY130_FD_SC_HD__O41A_4%A3 N_A3_M1007_g N_A3_M1003_g N_A3_M1009_g
+ N_A3_M1024_g A3 A3 N_A3_c_361_n PM_SKY130_FD_SC_HD__O41A_4%A3
x_PM_SKY130_FD_SC_HD__O41A_4%A2 N_A2_M1022_g N_A2_M1011_g N_A2_M1027_g
+ N_A2_M1016_g N_A2_c_408_n A2 A2 A2 N_A2_c_410_n N_A2_c_411_n
+ PM_SKY130_FD_SC_HD__O41A_4%A2
x_PM_SKY130_FD_SC_HD__O41A_4%A1 N_A1_M1000_g N_A1_M1008_g N_A1_M1012_g
+ N_A1_M1017_g N_A1_c_462_n A1 A1 A1 N_A1_c_464_n A1
+ PM_SKY130_FD_SC_HD__O41A_4%A1
x_PM_SKY130_FD_SC_HD__O41A_4%VPWR N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_M1023_s
+ N_VPWR_M1021_d N_VPWR_M1008_d N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n
+ N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n VPWR
+ N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_500_n N_VPWR_c_516_n
+ PM_SKY130_FD_SC_HD__O41A_4%VPWR
x_PM_SKY130_FD_SC_HD__O41A_4%X N_X_M1013_s N_X_M1019_s N_X_M1001_d N_X_M1020_d
+ N_X_c_607_n N_X_c_610_n N_X_c_600_n N_X_c_601_n N_X_c_603_n N_X_c_604_n
+ N_X_c_630_n N_X_c_605_n N_X_c_637_n X X X PM_SKY130_FD_SC_HD__O41A_4%X
x_PM_SKY130_FD_SC_HD__O41A_4%A_639_297# N_A_639_297#_M1006_d
+ N_A_639_297#_M1010_d N_A_639_297#_M1024_s N_A_639_297#_c_667_n
+ N_A_639_297#_c_674_n N_A_639_297#_c_668_n N_A_639_297#_c_669_n
+ N_A_639_297#_c_681_n N_A_639_297#_c_670_n N_A_639_297#_c_671_n
+ PM_SKY130_FD_SC_HD__O41A_4%A_639_297#
x_PM_SKY130_FD_SC_HD__O41A_4%A_889_297# N_A_889_297#_M1003_d
+ N_A_889_297#_M1011_s N_A_889_297#_c_730_n N_A_889_297#_c_716_n
+ N_A_889_297#_c_727_n N_A_889_297#_c_720_n
+ PM_SKY130_FD_SC_HD__O41A_4%A_889_297#
x_PM_SKY130_FD_SC_HD__O41A_4%A_1083_297# N_A_1083_297#_M1011_d
+ N_A_1083_297#_M1016_d N_A_1083_297#_M1017_s N_A_1083_297#_c_737_n
+ N_A_1083_297#_c_762_n N_A_1083_297#_c_738_n N_A_1083_297#_c_739_n
+ N_A_1083_297#_c_758_n N_A_1083_297#_c_740_n N_A_1083_297#_c_741_n
+ PM_SKY130_FD_SC_HD__O41A_4%A_1083_297#
x_PM_SKY130_FD_SC_HD__O41A_4%VGND N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1025_d
+ N_VGND_M1002_s N_VGND_M1007_s N_VGND_M1022_d N_VGND_M1000_s N_VGND_c_777_n
+ N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n
+ N_VGND_c_783_n N_VGND_c_784_n N_VGND_c_785_n N_VGND_c_786_n N_VGND_c_787_n
+ N_VGND_c_788_n N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n VGND
+ N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n N_VGND_c_795_n N_VGND_c_796_n
+ N_VGND_c_797_n PM_SKY130_FD_SC_HD__O41A_4%VGND
x_PM_SKY130_FD_SC_HD__O41A_4%A_467_47# N_A_467_47#_M1014_d N_A_467_47#_M1015_d
+ N_A_467_47#_M1026_d N_A_467_47#_M1009_d N_A_467_47#_M1027_s
+ N_A_467_47#_M1012_d N_A_467_47#_c_902_n N_A_467_47#_c_923_n
+ N_A_467_47#_c_915_n N_A_467_47#_c_903_n N_A_467_47#_c_904_n
+ N_A_467_47#_c_976_n N_A_467_47#_c_905_n N_A_467_47#_c_983_n
+ N_A_467_47#_c_906_n N_A_467_47#_c_942_n N_A_467_47#_c_907_n
+ N_A_467_47#_c_951_n N_A_467_47#_c_908_n N_A_467_47#_c_909_n
+ N_A_467_47#_c_910_n PM_SKY130_FD_SC_HD__O41A_4%A_467_47#
cc_1 VNB N_A_79_21#_M1013_g 0.0207742f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_79_21#_M1001_g 4.88014e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_A_79_21#_M1018_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_A_79_21#_M1005_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB N_A_79_21#_M1019_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_6 VNB N_A_79_21#_M1020_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_7 VNB N_A_79_21#_M1025_g 0.0216324f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_A_79_21#_M1023_g 4.65062e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB N_A_79_21#_c_136_n 0.00906818f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=1.185
cc_10 VNB N_A_79_21#_c_137_n 0.00445141f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=1.615
cc_11 VNB N_A_79_21#_c_138_n 0.0025508f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=0.72
cc_12 VNB N_A_79_21#_c_139_n 0.0635513f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_13 VNB N_B1_M1004_g 4.3564e-19 $X=-0.19 $Y=-0.24 $X2=3.605 $Y2=1.485
cc_14 VNB N_B1_c_255_n 0.0214694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_256_n 0.0155438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_M1021_g 6.90363e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_M1014_g 0.0216819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_M1015_g 0.0178808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B1_c_260_n 0.0411861f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_20 VNB N_A4_M1002_g 0.0177606f $X=-0.19 $Y=-0.24 $X2=3.605 $Y2=1.485
cc_21 VNB N_A4_M1006_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A4_M1026_g 0.0175566f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_23 VNB N_A4_M1010_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_24 VNB A4 0.00404201f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_25 VNB N_A4_c_310_n 0.028654f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_26 VNB N_A3_M1007_g 0.0175566f $X=-0.19 $Y=-0.24 $X2=3.605 $Y2=1.485
cc_27 VNB N_A3_M1003_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A3_M1009_g 0.017767f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_29 VNB N_A3_M1024_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_30 VNB A3 0.00301381f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_31 VNB N_A3_c_361_n 0.0298762f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_32 VNB N_A2_M1022_g 0.0205305f $X=-0.19 $Y=-0.24 $X2=3.605 $Y2=1.485
cc_33 VNB N_A2_M1011_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_M1027_g 0.022133f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_35 VNB N_A2_M1016_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_36 VNB N_A2_c_408_n 0.016803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB A2 0.00370972f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_38 VNB N_A2_c_410_n 0.0299385f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_39 VNB N_A2_c_411_n 0.0338971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A1_M1000_g 0.0193695f $X=-0.19 $Y=-0.24 $X2=3.605 $Y2=1.485
cc_41 VNB N_A1_M1008_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A1_M1012_g 0.0238824f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_43 VNB N_A1_M1017_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_44 VNB N_A1_c_462_n 0.0252779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB A1 0.0205413f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_46 VNB N_A1_c_464_n 0.0377344f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_47 VNB N_VPWR_c_500_n 0.326667f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.53
cc_48 VNB N_X_c_600_n 0.004418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_601_n 0.0120919f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_50 VNB X 0.0210175f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_51 VNB N_VGND_c_777_n 0.00988215f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_52 VNB N_VGND_c_778_n 0.0167929f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_53 VNB N_VGND_c_779_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_54 VNB N_VGND_c_780_n 0.0137659f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_55 VNB N_VGND_c_781_n 0.00430662f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_56 VNB N_VGND_c_782_n 0.00401293f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_57 VNB N_VGND_c_783_n 0.00527691f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_58 VNB N_VGND_c_784_n 0.0166611f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.185
cc_59 VNB N_VGND_c_785_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.16
cc_60 VNB N_VGND_c_786_n 0.0370872f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=1.615
cc_61 VNB N_VGND_c_787_n 0.00420034f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=1.66
cc_62 VNB N_VGND_c_788_n 0.0150203f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=2.34
cc_63 VNB N_VGND_c_789_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=2.38 $Y2=2.34
cc_64 VNB N_VGND_c_790_n 0.0206568f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=1.53
cc_65 VNB N_VGND_c_791_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=2.545 $Y2=1.53
cc_66 VNB N_VGND_c_792_n 0.017296f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=0.77
cc_67 VNB N_VGND_c_793_n 0.0254462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_794_n 0.38421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_795_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_796_n 0.0155839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_797_n 0.0155177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_467_47#_c_902_n 0.00245893f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_73 VNB N_A_467_47#_c_903_n 0.00283291f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_74 VNB N_A_467_47#_c_904_n 0.00326596f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_75 VNB N_A_467_47#_c_905_n 0.00337094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_467_47#_c_906_n 0.00630437f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_77 VNB N_A_467_47#_c_907_n 0.0143927f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_78 VNB N_A_467_47#_c_908_n 0.0026015f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=2.34
cc_79 VNB N_A_467_47#_c_909_n 0.00233301f $X=-0.19 $Y=-0.24 $X2=2.38 $Y2=2.34
cc_80 VNB N_A_467_47#_c_910_n 0.00168765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VPB N_A_79_21#_M1001_g 0.0229974f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_82 VPB N_A_79_21#_M1005_g 0.0193321f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_83 VPB N_A_79_21#_M1020_g 0.0193519f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_84 VPB N_A_79_21#_M1023_g 0.0198045f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_85 VPB N_A_79_21#_c_144_n 0.017418f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.53
cc_86 VPB N_A_79_21#_c_145_n 0.0020238f $X=-0.19 $Y=1.305 $X2=3.74 $Y2=1.61
cc_87 VPB N_B1_M1004_g 0.0194056f $X=-0.19 $Y=1.305 $X2=3.605 $Y2=1.485
cc_88 VPB N_B1_M1021_g 0.0263929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A4_M1006_g 0.026721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A4_M1010_g 0.0196623f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_91 VPB N_A3_M1003_g 0.0194853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A3_M1024_g 0.0267067f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_93 VPB N_A2_M1011_g 0.0267252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A2_M1016_g 0.0194911f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_95 VPB N_A1_M1008_g 0.0192639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A1_M1017_g 0.026498f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_97 VPB N_VPWR_c_501_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_98 VPB N_VPWR_c_502_n 0.0297161f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.025
cc_99 VPB N_VPWR_c_503_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_100 VPB N_VPWR_c_504_n 0.00596637f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_101 VPB N_VPWR_c_505_n 0.0111617f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_102 VPB N_VPWR_c_506_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_103 VPB N_VPWR_c_507_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_104 VPB N_VPWR_c_508_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_105 VPB N_VPWR_c_509_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=1.185
cc_106 VPB N_VPWR_c_510_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.185
cc_107 VPB N_VPWR_c_511_n 0.0183907f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_108 VPB N_VPWR_c_512_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_513_n 0.087272f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.77
cc_110 VPB N_VPWR_c_514_n 0.0245821f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.185
cc_111 VPB N_VPWR_c_500_n 0.0592901f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.53
cc_112 VPB N_VPWR_c_516_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_113 VPB N_X_c_603_n 0.00220047f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_114 VPB N_X_c_604_n 0.0125653f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_115 VPB N_X_c_605_n 0.00224287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB X 0.0088204f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_117 VPB N_A_639_297#_c_667_n 0.00480364f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_118 VPB N_A_639_297#_c_668_n 0.00203255f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_119 VPB N_A_639_297#_c_669_n 0.00409472f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_120 VPB N_A_639_297#_c_670_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_121 VPB N_A_639_297#_c_671_n 0.0101002f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_122 VPB N_A_889_297#_c_716_n 0.0119259f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_123 VPB N_A_1083_297#_c_737_n 0.00274954f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_124 VPB N_A_1083_297#_c_738_n 0.00387462f $X=-0.19 $Y=1.305 $X2=0.89
+ $Y2=1.025
cc_125 VPB N_A_1083_297#_c_739_n 0.0096678f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_126 VPB N_A_1083_297#_c_740_n 0.00768346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_1083_297#_c_741_n 0.00236123f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_128 N_A_79_21#_M1023_g N_B1_M1004_g 0.014584f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_137_n N_B1_M1004_g 0.0071507f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_148_p N_B1_M1004_g 0.00909434f $X=2.38 $Y=1.66 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_137_n N_B1_c_255_n 0.0182912f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_136_n N_B1_c_256_n 0.014037f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_137_n N_B1_c_256_n 0.00193329f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_139_n N_B1_c_256_n 0.014584f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_137_n N_B1_M1021_g 0.00734321f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_148_p N_B1_M1021_g 0.0168093f $X=2.38 $Y=1.66 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_144_n N_B1_M1021_g 0.0127536f $X=3.575 $Y=1.53 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_137_n N_B1_M1014_g 0.0131921f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_138_n N_B1_M1014_g 0.00501393f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_137_n N_B1_M1015_g 6.35905e-19 $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_138_n N_B1_M1015_g 0.00396431f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_137_n B1 0.0135702f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_144_n B1 0.0238641f $X=3.575 $Y=1.53 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_138_n B1 0.0156627f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_137_n N_B1_c_260_n 0.0112756f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_144_n N_B1_c_260_n 0.0137331f $X=3.575 $Y=1.53 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_138_n N_B1_c_260_n 0.00208222f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_144_n N_A4_M1006_g 0.0128219f $X=3.575 $Y=1.53 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_145_n N_A4_M1006_g 0.0141102f $X=3.74 $Y=1.61 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_145_n N_A4_M1010_g 3.16391e-19 $X=3.74 $Y=1.61 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_144_n A4 0.0116336f $X=3.575 $Y=1.53 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_145_n A4 0.0202536f $X=3.74 $Y=1.61 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_145_n N_A4_c_310_n 0.00206069f $X=3.74 $Y=1.61 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_144_n N_VPWR_M1021_d 0.00298653f $X=3.575 $Y=1.53 $X2=0
+ $Y2=0
cc_155 N_A_79_21#_M1001_g N_VPWR_c_502_n 0.00321781f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A_79_21#_M1005_g N_VPWR_c_503_n 0.00146448f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_79_21#_M1020_g N_VPWR_c_503_n 0.00146448f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_79_21#_M1023_g N_VPWR_c_504_n 0.00159991f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_79_21#_c_136_n N_VPWR_c_504_n 0.0144431f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_160 N_A_79_21#_c_137_n N_VPWR_c_504_n 0.00703647f $X=2.37 $Y=1.615 $X2=0
+ $Y2=0
cc_161 N_A_79_21#_c_144_n N_VPWR_c_505_n 0.0163834f $X=3.575 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A_79_21#_M1001_g N_VPWR_c_507_n 0.00541359f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_79_21#_M1005_g N_VPWR_c_507_n 0.00541359f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_79_21#_M1020_g N_VPWR_c_509_n 0.00541359f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_79_21#_M1023_g N_VPWR_c_509_n 0.00541359f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_79_21#_c_148_p N_VPWR_c_511_n 0.0203103f $X=2.38 $Y=1.66 $X2=0 $Y2=0
cc_167 N_A_79_21#_M1004_s N_VPWR_c_500_n 0.00231261f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_168 N_A_79_21#_M1006_s N_VPWR_c_500_n 0.00216833f $X=3.605 $Y=1.485 $X2=0
+ $Y2=0
cc_169 N_A_79_21#_M1001_g N_VPWR_c_500_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_79_21#_M1005_g N_VPWR_c_500_n 0.00950154f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_79_21#_M1020_g N_VPWR_c_500_n 0.00950154f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_M1023_g N_VPWR_c_500_n 0.00952874f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_79_21#_c_148_p N_VPWR_c_500_n 0.012992f $X=2.38 $Y=1.66 $X2=0 $Y2=0
cc_174 N_A_79_21#_M1013_g N_X_c_607_n 0.0109535f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_79_21#_M1018_g N_X_c_607_n 0.00631111f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_79_21#_M1019_g N_X_c_607_n 5.2007e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_79_21#_M1001_g N_X_c_610_n 0.0146918f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_79_21#_M1005_g N_X_c_610_n 0.00985707f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_79_21#_M1020_g N_X_c_610_n 6.20279e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_79_21#_M1018_g N_X_c_600_n 0.00890471f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_79_21#_M1019_g N_X_c_600_n 0.0100649f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_79_21#_M1025_g N_X_c_600_n 0.00294852f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_79_21#_c_136_n N_X_c_600_n 0.0267108f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_184 N_A_79_21#_c_137_n N_X_c_600_n 6.73998e-19 $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_185 N_A_79_21#_c_139_n N_X_c_600_n 0.00419427f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_79_21#_M1013_g N_X_c_601_n 0.01335f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A_79_21#_M1018_g N_X_c_601_n 0.0012996f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A_79_21#_c_136_n N_X_c_601_n 0.0605668f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_189 N_A_79_21#_c_139_n N_X_c_601_n 0.00205999f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_79_21#_M1005_g N_X_c_603_n 0.0115138f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_79_21#_M1020_g N_X_c_603_n 0.0115138f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_139_n N_X_c_603_n 0.00194394f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_79_21#_M1001_g N_X_c_604_n 0.0160365f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_79_21#_M1005_g N_X_c_604_n 0.00125262f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_136_n N_X_c_604_n 0.0608108f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_139_n N_X_c_604_n 0.00194394f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_79_21#_M1018_g N_X_c_630_n 5.19281e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_79_21#_M1019_g N_X_c_630_n 0.00620543f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_79_21#_M1025_g N_X_c_630_n 0.0052782f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_79_21#_M1020_g N_X_c_605_n 0.00120279f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_79_21#_M1023_g N_X_c_605_n 0.00275158f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_79_21#_c_136_n N_X_c_605_n 0.0268132f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_139_n N_X_c_605_n 0.00201507f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_79_21#_M1005_g N_X_c_637_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_79_21#_M1020_g N_X_c_637_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_79_21#_M1023_g N_X_c_637_n 0.00857288f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_79_21#_M1013_g X 0.021111f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_136_n X 0.0179682f $X=2.195 $Y=1.185 $X2=0 $Y2=0
cc_209 N_A_79_21#_c_144_n N_A_639_297#_M1006_d 0.00298653f $X=3.575 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_210 N_A_79_21#_c_144_n N_A_639_297#_c_667_n 0.0176815f $X=3.575 $Y=1.53 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_M1006_s N_A_639_297#_c_674_n 0.00312348f $X=3.605 $Y=1.485
+ $X2=0 $Y2=0
cc_212 N_A_79_21#_c_145_n N_A_639_297#_c_674_n 0.0139178f $X=3.74 $Y=1.61 $X2=0
+ $Y2=0
cc_213 N_A_79_21#_c_145_n N_A_639_297#_c_669_n 0.00902116f $X=3.74 $Y=1.61 $X2=0
+ $Y2=0
cc_214 N_A_79_21#_M1013_g N_VGND_c_778_n 0.00321781f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A_79_21#_M1018_g N_VGND_c_779_n 0.00146448f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A_79_21#_M1019_g N_VGND_c_779_n 0.00146448f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A_79_21#_M1025_g N_VGND_c_780_n 0.00321269f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_218 N_A_79_21#_c_136_n N_VGND_c_780_n 0.0189643f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_219 N_A_79_21#_c_137_n N_VGND_c_780_n 0.0200434f $X=2.37 $Y=1.615 $X2=0 $Y2=0
cc_220 N_A_79_21#_M1013_g N_VGND_c_784_n 0.00421248f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A_79_21#_M1018_g N_VGND_c_784_n 0.00421248f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_79_21#_M1019_g N_VGND_c_792_n 0.00422241f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A_79_21#_M1025_g N_VGND_c_792_n 0.00541359f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_79_21#_M1014_s N_VGND_c_794_n 0.00216833f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_M1013_g N_VGND_c_794_n 0.00666524f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A_79_21#_M1018_g N_VGND_c_794_n 0.00571103f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A_79_21#_M1019_g N_VGND_c_794_n 0.00569656f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A_79_21#_M1025_g N_VGND_c_794_n 0.0108276f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A_79_21#_c_137_n N_A_467_47#_M1014_d 0.003096f $X=2.37 $Y=1.615
+ $X2=-0.19 $Y2=-0.24
cc_230 N_A_79_21#_M1014_s N_A_467_47#_c_902_n 0.00304629f $X=2.745 $Y=0.235
+ $X2=0 $Y2=0
cc_231 N_A_79_21#_c_137_n N_A_467_47#_c_902_n 0.024108f $X=2.37 $Y=1.615 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_c_138_n N_A_467_47#_c_902_n 0.0186474f $X=2.88 $Y=0.72 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_c_138_n N_A_467_47#_c_915_n 0.0072979f $X=2.88 $Y=0.72 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_144_n N_A_467_47#_c_904_n 0.00659169f $X=3.575 $Y=1.53 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_c_138_n N_A_467_47#_c_904_n 0.0135776f $X=2.88 $Y=0.72 $X2=0
+ $Y2=0
cc_236 N_B1_M1015_g N_A4_M1002_g 0.0130574f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_237 B1 A4 0.0126301f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_238 N_B1_c_260_n A4 0.00155448f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_239 B1 N_A4_c_310_n 2.34654e-19 $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_240 N_B1_c_260_n N_A4_c_310_n 0.0130574f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B1_M1004_g N_VPWR_c_504_n 0.00282267f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_242 N_B1_M1021_g N_VPWR_c_505_n 0.0044954f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_243 N_B1_M1004_g N_VPWR_c_511_n 0.00541359f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_244 N_B1_M1021_g N_VPWR_c_511_n 0.00541359f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_245 N_B1_M1004_g N_VPWR_c_500_n 0.009581f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_246 N_B1_M1021_g N_VPWR_c_500_n 0.0108799f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_247 N_B1_c_256_n N_VGND_c_780_n 8.28776e-19 $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B1_M1014_g N_VGND_c_780_n 0.00630986f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_249 N_B1_M1014_g N_VGND_c_786_n 0.00357877f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_250 N_B1_M1015_g N_VGND_c_786_n 0.00357877f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_251 N_B1_M1014_g N_VGND_c_794_n 0.00655123f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_252 N_B1_M1015_g N_VGND_c_794_n 0.00530095f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_253 N_B1_c_255_n N_A_467_47#_c_902_n 8.82258e-19 $X=2.515 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_M1014_g N_A_467_47#_c_902_n 0.00866418f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_255 N_B1_M1015_g N_A_467_47#_c_902_n 0.0103285f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_256 B1 N_A_467_47#_c_902_n 0.00288754f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_257 N_B1_M1015_g N_A_467_47#_c_904_n 8.07877e-19 $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A4_M1026_g N_A3_M1007_g 0.0148856f $X=3.95 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A4_M1010_g N_A3_M1003_g 0.0148856f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_260 A4 A3 0.0116851f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_261 N_A4_c_310_n A3 2.32004e-19 $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_262 A4 N_A3_c_361_n 0.00154478f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_263 N_A4_c_310_n N_A3_c_361_n 0.0148856f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A4_M1006_g N_VPWR_c_505_n 0.00229942f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A4_M1006_g N_VPWR_c_513_n 0.00357877f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A4_M1010_g N_VPWR_c_513_n 0.00357835f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A4_M1006_g N_VPWR_c_500_n 0.00655123f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A4_M1010_g N_VPWR_c_500_n 0.00525234f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A4_M1006_g N_A_639_297#_c_674_n 0.0112878f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A4_M1010_g N_A_639_297#_c_674_n 0.0108275f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A4_M1010_g N_A_639_297#_c_669_n 0.00265654f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_272 A4 N_A_639_297#_c_669_n 0.00359221f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_273 N_A4_M1006_g N_A_639_297#_c_681_n 4.72397e-19 $X=3.53 $Y=1.985 $X2=0
+ $Y2=0
cc_274 N_A4_M1010_g N_A_639_297#_c_681_n 0.00846527f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_275 N_A4_M1002_g N_VGND_c_781_n 0.00275964f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A4_M1026_g N_VGND_c_781_n 0.00156096f $X=3.95 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A4_M1002_g N_VGND_c_786_n 0.00422898f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A4_M1026_g N_VGND_c_788_n 0.00438403f $X=3.95 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A4_M1002_g N_VGND_c_794_n 0.00582093f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A4_M1026_g N_VGND_c_794_n 0.00580713f $X=3.95 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A4_M1002_g N_A_467_47#_c_923_n 0.00244813f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A4_M1002_g N_A_467_47#_c_915_n 0.00435425f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A4_M1026_g N_A_467_47#_c_915_n 5.36297e-19 $X=3.95 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A4_M1002_g N_A_467_47#_c_903_n 0.00850187f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A4_M1026_g N_A_467_47#_c_903_n 0.01033f $X=3.95 $Y=0.56 $X2=0 $Y2=0
cc_286 A4 N_A_467_47#_c_903_n 0.0391879f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_287 N_A4_c_310_n N_A_467_47#_c_903_n 0.00205431f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A4_M1002_g N_A_467_47#_c_904_n 0.00106589f $X=3.53 $Y=0.56 $X2=0 $Y2=0
cc_289 A4 N_A_467_47#_c_904_n 0.00613155f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_290 N_A3_M1009_g N_A2_M1022_g 0.0130174f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_291 A3 N_A2_c_408_n 7.95839e-19 $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_292 N_A3_c_361_n N_A2_c_408_n 0.0133308f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_293 A3 A2 0.016126f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_294 N_A3_c_361_n A2 2.11787e-19 $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A3_M1003_g N_VPWR_c_513_n 0.00539841f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A3_M1024_g N_VPWR_c_513_n 0.00357877f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A3_M1003_g N_VPWR_c_500_n 0.00961452f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A3_M1024_g N_VPWR_c_500_n 0.00660224f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A3_M1003_g N_A_639_297#_c_674_n 0.00200982f $X=4.37 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A3_M1003_g N_A_639_297#_c_669_n 0.00173367f $X=4.37 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A3_M1003_g N_A_639_297#_c_681_n 0.00824958f $X=4.37 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A3_M1024_g N_A_639_297#_c_681_n 5.83827e-19 $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A3_M1003_g N_A_639_297#_c_670_n 0.0106641f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A3_M1024_g N_A_639_297#_c_670_n 0.0107189f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_305 A3 N_A_639_297#_c_670_n 0.0356421f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_306 N_A3_c_361_n N_A_639_297#_c_670_n 0.00198252f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A3_M1003_g N_A_639_297#_c_671_n 5.3107e-19 $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A3_M1024_g N_A_639_297#_c_671_n 0.00846753f $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_309 A3 N_A_639_297#_c_671_n 0.0104121f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_310 N_A3_M1024_g N_A_889_297#_c_716_n 0.0134027f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A3_M1024_g N_A_1083_297#_c_740_n 4.42201e-19 $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A3_M1007_g N_VGND_c_782_n 0.00158744f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A3_M1009_g N_VGND_c_782_n 0.00161369f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_314 N_A3_M1007_g N_VGND_c_788_n 0.00438403f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A3_M1007_g N_VGND_c_794_n 0.00580713f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A3_M1009_g N_VGND_c_794_n 0.00585571f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A3_M1009_g N_VGND_c_796_n 0.00438403f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_318 N_A3_M1009_g N_VGND_c_797_n 4.29292e-19 $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_319 N_A3_M1007_g N_A_467_47#_c_905_n 0.0107978f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_320 N_A3_M1009_g N_A_467_47#_c_905_n 0.0103868f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_321 A3 N_A_467_47#_c_905_n 0.0415094f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_322 N_A3_c_361_n N_A_467_47#_c_905_n 0.00205431f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_323 A3 N_A_467_47#_c_909_n 0.00382939f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_324 N_A2_M1027_g N_A1_M1000_g 0.0193433f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A2_M1016_g N_A1_M1008_g 0.0165218f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_326 A2 N_A1_c_462_n 0.00173822f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_327 N_A2_c_411_n N_A1_c_462_n 0.0177243f $X=6.19 $Y=1.16 $X2=0 $Y2=0
cc_328 A2 A1 0.0118168f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_329 N_A2_M1016_g N_VPWR_c_506_n 0.00130512f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A2_M1011_g N_VPWR_c_513_n 0.00357835f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A2_M1016_g N_VPWR_c_513_n 0.00539841f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A2_M1011_g N_VPWR_c_500_n 0.0066022f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A2_M1016_g N_VPWR_c_500_n 0.00961452f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A2_M1011_g N_A_639_297#_c_671_n 4.35828e-19 $X=5.77 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A2_c_408_n N_A_639_297#_c_671_n 3.92905e-19 $X=5.305 $Y=1.16 $X2=0
+ $Y2=0
cc_336 A2 N_A_639_297#_c_671_n 0.0012217f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_337 N_A2_M1011_g N_A_889_297#_c_716_n 0.012922f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A2_M1016_g N_A_889_297#_c_716_n 0.00209036f $X=6.19 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A2_M1011_g N_A_889_297#_c_720_n 0.0118647f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A2_M1016_g N_A_889_297#_c_720_n 0.0057144f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A2_M1011_g N_A_1083_297#_c_737_n 0.0128263f $X=5.77 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A2_M1016_g N_A_1083_297#_c_737_n 0.0124912f $X=6.19 $Y=1.985 $X2=0
+ $Y2=0
cc_343 A2 N_A_1083_297#_c_737_n 0.0472848f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A2_c_410_n N_A_1083_297#_c_737_n 0.00107937f $X=5.695 $Y=1.16 $X2=0
+ $Y2=0
cc_345 N_A2_c_411_n N_A_1083_297#_c_737_n 0.00341937f $X=6.19 $Y=1.16 $X2=0
+ $Y2=0
cc_346 A2 N_A_1083_297#_c_740_n 0.0203601f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_347 N_A2_c_410_n N_A_1083_297#_c_740_n 0.0057216f $X=5.695 $Y=1.16 $X2=0
+ $Y2=0
cc_348 A2 N_A_1083_297#_c_741_n 0.00384327f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_349 N_A2_M1027_g N_VGND_c_790_n 0.00438403f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A2_M1022_g N_VGND_c_794_n 0.00508999f $X=5.23 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A2_M1027_g N_VGND_c_794_n 0.00551776f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_352 N_A2_M1022_g N_VGND_c_796_n 0.00438403f $X=5.23 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A2_M1022_g N_VGND_c_797_n 0.00236143f $X=5.23 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A2_M1027_g N_VGND_c_797_n 0.0039692f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A2_M1022_g N_A_467_47#_c_906_n 0.0117981f $X=5.23 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A2_M1027_g N_A_467_47#_c_906_n 0.0144691f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_357 A2 N_A_467_47#_c_906_n 0.0776664f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_358 N_A2_c_410_n N_A_467_47#_c_906_n 0.0104596f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A2_c_411_n N_A_467_47#_c_906_n 0.0048872f $X=6.19 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A2_M1027_g N_A_467_47#_c_942_n 0.006882f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_361 A2 N_A_467_47#_c_910_n 0.00994057f $X=6.19 $Y=1.105 $X2=0 $Y2=0
cc_362 N_A2_c_411_n N_A_467_47#_c_910_n 0.00178809f $X=6.19 $Y=1.16 $X2=0 $Y2=0
cc_363 N_A1_M1008_g N_VPWR_c_506_n 0.012825f $X=6.61 $Y=1.985 $X2=0 $Y2=0
cc_364 N_A1_M1017_g N_VPWR_c_506_n 0.015466f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A1_M1008_g N_VPWR_c_513_n 0.0046653f $X=6.61 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A1_M1017_g N_VPWR_c_514_n 0.0046653f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A1_M1008_g N_VPWR_c_500_n 0.007919f $X=6.61 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A1_M1017_g N_VPWR_c_500_n 0.00916306f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A1_M1008_g N_A_1083_297#_c_738_n 0.0138858f $X=6.61 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A1_M1017_g N_A_1083_297#_c_738_n 0.0158864f $X=7.03 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_A1_c_462_n N_A_1083_297#_c_738_n 0.00198252f $X=7.105 $Y=1.16 $X2=0
+ $Y2=0
cc_372 A1 N_A_1083_297#_c_738_n 0.0437526f $X=7.55 $Y=1.105 $X2=0 $Y2=0
cc_373 N_A1_c_464_n N_A_1083_297#_c_738_n 0.00350245f $X=7.315 $Y=1.16 $X2=0
+ $Y2=0
cc_374 A1 N_A_1083_297#_c_739_n 0.0273535f $X=7.55 $Y=1.105 $X2=0 $Y2=0
cc_375 N_A1_c_464_n N_A_1083_297#_c_739_n 0.00493159f $X=7.315 $Y=1.16 $X2=0
+ $Y2=0
cc_376 N_A1_M1017_g N_A_1083_297#_c_758_n 0.0207555f $X=7.03 $Y=1.985 $X2=0
+ $Y2=0
cc_377 N_A1_M1000_g N_VGND_c_783_n 0.00306527f $X=6.61 $Y=0.56 $X2=0 $Y2=0
cc_378 N_A1_M1012_g N_VGND_c_783_n 0.00306527f $X=7.03 $Y=0.56 $X2=0 $Y2=0
cc_379 N_A1_M1000_g N_VGND_c_790_n 0.00438403f $X=6.61 $Y=0.56 $X2=0 $Y2=0
cc_380 N_A1_M1012_g N_VGND_c_793_n 0.00438403f $X=7.03 $Y=0.56 $X2=0 $Y2=0
cc_381 N_A1_M1000_g N_VGND_c_794_n 0.00628347f $X=6.61 $Y=0.56 $X2=0 $Y2=0
cc_382 N_A1_M1012_g N_VGND_c_794_n 0.00701993f $X=7.03 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A1_M1000_g N_VGND_c_797_n 8.13483e-19 $X=6.61 $Y=0.56 $X2=0 $Y2=0
cc_384 N_A1_M1000_g N_A_467_47#_c_942_n 0.00724793f $X=6.61 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A1_M1000_g N_A_467_47#_c_907_n 0.0144523f $X=6.61 $Y=0.56 $X2=0 $Y2=0
cc_386 N_A1_M1012_g N_A_467_47#_c_907_n 0.0139787f $X=7.03 $Y=0.56 $X2=0 $Y2=0
cc_387 N_A1_c_462_n N_A_467_47#_c_907_n 0.00205431f $X=7.105 $Y=1.16 $X2=0 $Y2=0
cc_388 A1 N_A_467_47#_c_907_n 0.0710012f $X=7.55 $Y=1.105 $X2=0 $Y2=0
cc_389 N_A1_c_464_n N_A_467_47#_c_907_n 0.00872793f $X=7.315 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A1_M1012_g N_A_467_47#_c_951_n 0.0133575f $X=7.03 $Y=0.56 $X2=0 $Y2=0
cc_391 N_VPWR_c_500_n N_X_M1001_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_500_n N_X_M1020_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_507_n N_X_c_610_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_c_500_n N_X_c_610_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_395 N_VPWR_M1005_s N_X_c_603_n 0.00166664f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_396 N_VPWR_c_503_n N_X_c_603_n 0.0128323f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_397 N_VPWR_M1001_s N_X_c_604_n 0.00296139f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_398 N_VPWR_c_502_n N_X_c_604_n 0.0208833f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_399 N_VPWR_c_504_n N_X_c_605_n 0.00914268f $X=1.94 $Y=1.66 $X2=0 $Y2=0
cc_400 N_VPWR_c_509_n N_X_c_637_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_500_n N_X_c_637_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_500_n N_A_639_297#_M1006_d 0.00209324f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_403 N_VPWR_c_500_n N_A_639_297#_M1010_d 0.00215201f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_500_n N_A_639_297#_M1024_s 0.00226545f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_505_n N_A_639_297#_c_667_n 0.0369016f $X=2.8 $Y=2 $X2=0 $Y2=0
cc_406 N_VPWR_c_513_n N_A_639_297#_c_674_n 0.0512704f $X=6.655 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_500_n N_A_639_297#_c_674_n 0.0329592f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_505_n N_A_639_297#_c_668_n 0.0147456f $X=2.8 $Y=2 $X2=0 $Y2=0
cc_409 N_VPWR_c_513_n N_A_639_297#_c_668_n 0.0187211f $X=6.655 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_500_n N_A_639_297#_c_668_n 0.0103775f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_500_n N_A_889_297#_M1003_d 0.00385313f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_412 N_VPWR_c_500_n N_A_889_297#_M1011_s 0.00215201f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_506_n N_A_889_297#_c_716_n 3.24428e-19 $X=6.82 $Y=1.95 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_513_n N_A_889_297#_c_716_n 0.0870493f $X=6.655 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_500_n N_A_889_297#_c_716_n 0.0538167f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_513_n N_A_889_297#_c_727_n 0.0114668f $X=6.655 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_500_n N_A_889_297#_c_727_n 0.006547f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_500_n N_A_1083_297#_M1011_d 0.00226545f $X=7.59 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_419 N_VPWR_c_500_n N_A_1083_297#_M1016_d 0.00562567f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_500_n N_A_1083_297#_M1017_s 0.00956796f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_513_n N_A_1083_297#_c_762_n 0.0107103f $X=6.655 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_500_n N_A_1083_297#_c_762_n 0.00643939f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_M1008_d N_A_1083_297#_c_738_n 0.00165831f $X=6.685 $Y=1.485 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_506_n N_A_1083_297#_c_738_n 0.0170258f $X=6.82 $Y=1.95 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_506_n N_A_1083_297#_c_758_n 0.0360097f $X=6.82 $Y=1.95 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_514_n N_A_1083_297#_c_758_n 0.0230652f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_500_n N_A_1083_297#_c_758_n 0.0126319f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_X_c_601_n N_VGND_M1013_d 0.00285834f $X=0.845 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_429 N_X_c_600_n N_VGND_M1018_d 0.00162148f $X=1.355 $Y=0.81 $X2=0 $Y2=0
cc_430 N_X_c_601_n N_VGND_c_778_n 0.0199638f $X=0.845 $Y=0.81 $X2=0 $Y2=0
cc_431 N_X_c_600_n N_VGND_c_779_n 0.0122675f $X=1.355 $Y=0.81 $X2=0 $Y2=0
cc_432 N_X_c_607_n N_VGND_c_784_n 0.0184921f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_433 N_X_c_601_n N_VGND_c_784_n 0.0041083f $X=0.845 $Y=0.81 $X2=0 $Y2=0
cc_434 N_X_c_600_n N_VGND_c_792_n 0.00203746f $X=1.355 $Y=0.81 $X2=0 $Y2=0
cc_435 N_X_c_630_n N_VGND_c_792_n 0.0188551f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_436 N_X_M1013_s N_VGND_c_794_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_437 N_X_M1019_s N_VGND_c_794_n 0.00215201f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_438 N_X_c_607_n N_VGND_c_794_n 0.012098f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_439 N_X_c_600_n N_VGND_c_794_n 0.00455756f $X=1.355 $Y=0.81 $X2=0 $Y2=0
cc_440 N_X_c_601_n N_VGND_c_794_n 0.00886193f $X=0.845 $Y=0.81 $X2=0 $Y2=0
cc_441 N_X_c_630_n N_VGND_c_794_n 0.0122069f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_442 N_A_639_297#_c_670_n N_A_889_297#_M1003_d 0.00165831f $X=4.835 $Y=1.53
+ $X2=-0.19 $Y2=1.305
cc_443 N_A_639_297#_c_670_n N_A_889_297#_c_730_n 0.0126919f $X=4.835 $Y=1.53
+ $X2=0 $Y2=0
cc_444 N_A_639_297#_M1024_s N_A_889_297#_c_716_n 0.00545241f $X=4.865 $Y=1.485
+ $X2=0 $Y2=0
cc_445 N_A_639_297#_c_671_n N_A_889_297#_c_716_n 0.0195167f $X=5 $Y=1.61 $X2=0
+ $Y2=0
cc_446 N_A_639_297#_c_671_n N_A_1083_297#_c_740_n 0.0458157f $X=5 $Y=1.61 $X2=0
+ $Y2=0
cc_447 N_A_639_297#_c_669_n N_A_467_47#_c_903_n 0.00130635f $X=4.16 $Y=1.615
+ $X2=0 $Y2=0
cc_448 N_A_639_297#_c_669_n N_A_467_47#_c_905_n 0.0027567f $X=4.16 $Y=1.615
+ $X2=0 $Y2=0
cc_449 N_A_639_297#_c_671_n N_A_467_47#_c_906_n 0.00243757f $X=5 $Y=1.61 $X2=0
+ $Y2=0
cc_450 N_A_639_297#_c_669_n N_A_467_47#_c_908_n 0.0070861f $X=4.16 $Y=1.615
+ $X2=0 $Y2=0
cc_451 N_A_639_297#_c_671_n N_A_467_47#_c_909_n 0.00520448f $X=5 $Y=1.61 $X2=0
+ $Y2=0
cc_452 N_A_889_297#_c_716_n N_A_1083_297#_M1011_d 0.00545241f $X=5.815 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_453 N_A_889_297#_M1011_s N_A_1083_297#_c_737_n 0.00165831f $X=5.845 $Y=1.485
+ $X2=0 $Y2=0
cc_454 N_A_889_297#_c_720_n N_A_1083_297#_c_737_n 0.0170258f $X=5.98 $Y=1.95
+ $X2=0 $Y2=0
cc_455 N_A_889_297#_c_716_n N_A_1083_297#_c_740_n 0.0175913f $X=5.815 $Y=2.38
+ $X2=0 $Y2=0
cc_456 N_A_1083_297#_c_738_n N_A_467_47#_c_907_n 0.00469518f $X=7.265 $Y=1.53
+ $X2=0 $Y2=0
cc_457 N_A_1083_297#_c_741_n N_A_467_47#_c_907_n 0.00281867f $X=6.4 $Y=1.61
+ $X2=0 $Y2=0
cc_458 N_A_1083_297#_c_741_n N_A_467_47#_c_910_n 0.0020842f $X=6.4 $Y=1.61 $X2=0
+ $Y2=0
cc_459 N_VGND_c_794_n N_A_467_47#_M1014_d 0.00209344f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_460 N_VGND_c_794_n N_A_467_47#_M1015_d 0.00231267f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_794_n N_A_467_47#_M1026_d 0.00263776f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_794_n N_A_467_47#_M1009_d 0.00290077f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_794_n N_A_467_47#_M1027_s 0.00531264f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_794_n N_A_467_47#_M1012_d 0.00478998f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_465 N_VGND_c_780_n N_A_467_47#_c_902_n 0.0166761f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_466 N_VGND_c_786_n N_A_467_47#_c_902_n 0.0532068f $X=3.655 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_794_n N_A_467_47#_c_902_n 0.0336592f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_c_786_n N_A_467_47#_c_923_n 0.015453f $X=3.655 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_794_n N_A_467_47#_c_923_n 0.00940698f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_M1002_s N_A_467_47#_c_903_n 0.00169589f $X=3.605 $Y=0.235 $X2=0
+ $Y2=0
cc_471 N_VGND_c_781_n N_A_467_47#_c_903_n 0.0111177f $X=3.74 $Y=0.38 $X2=0 $Y2=0
cc_472 N_VGND_c_786_n N_A_467_47#_c_903_n 0.00193763f $X=3.655 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_788_n N_A_467_47#_c_903_n 0.00233081f $X=4.445 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_794_n N_A_467_47#_c_903_n 0.0091145f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_788_n N_A_467_47#_c_976_n 0.0113595f $X=4.445 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_794_n N_A_467_47#_c_976_n 0.0064623f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_M1007_s N_A_467_47#_c_905_n 0.00169589f $X=4.445 $Y=0.235 $X2=0
+ $Y2=0
cc_478 N_VGND_c_782_n N_A_467_47#_c_905_n 0.0111177f $X=4.58 $Y=0.38 $X2=0 $Y2=0
cc_479 N_VGND_c_788_n N_A_467_47#_c_905_n 0.00233081f $X=4.445 $Y=0 $X2=0 $Y2=0
cc_480 N_VGND_c_794_n N_A_467_47#_c_905_n 0.00994094f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_481 N_VGND_c_796_n N_A_467_47#_c_905_n 0.00233081f $X=5.305 $Y=0.23 $X2=0
+ $Y2=0
cc_482 N_VGND_c_794_n N_A_467_47#_c_983_n 0.0064623f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_796_n N_A_467_47#_c_983_n 0.0115672f $X=5.305 $Y=0.23 $X2=0
+ $Y2=0
cc_484 N_VGND_c_797_n N_A_467_47#_c_983_n 0.0197649f $X=5.915 $Y=0.23 $X2=0
+ $Y2=0
cc_485 N_VGND_M1022_d N_A_467_47#_c_906_n 0.00746577f $X=5.305 $Y=0.235 $X2=0
+ $Y2=0
cc_486 N_VGND_c_790_n N_A_467_47#_c_906_n 0.00405733f $X=6.685 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_794_n N_A_467_47#_c_906_n 0.015104f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_796_n N_A_467_47#_c_906_n 0.0025616f $X=5.305 $Y=0.23 $X2=0
+ $Y2=0
cc_489 N_VGND_c_797_n N_A_467_47#_c_906_n 0.0351821f $X=5.915 $Y=0.23 $X2=0
+ $Y2=0
cc_490 N_VGND_c_783_n N_A_467_47#_c_942_n 0.0157558f $X=6.82 $Y=0.38 $X2=0 $Y2=0
cc_491 N_VGND_c_790_n N_A_467_47#_c_942_n 0.0117748f $X=6.685 $Y=0 $X2=0 $Y2=0
cc_492 N_VGND_c_794_n N_A_467_47#_c_942_n 0.0064623f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_493 N_VGND_c_797_n N_A_467_47#_c_942_n 0.0149815f $X=5.915 $Y=0.23 $X2=0
+ $Y2=0
cc_494 N_VGND_M1000_s N_A_467_47#_c_907_n 0.00169589f $X=6.685 $Y=0.235 $X2=0
+ $Y2=0
cc_495 N_VGND_c_783_n N_A_467_47#_c_907_n 0.0111177f $X=6.82 $Y=0.38 $X2=0 $Y2=0
cc_496 N_VGND_c_790_n N_A_467_47#_c_907_n 0.00334772f $X=6.685 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_793_n N_A_467_47#_c_907_n 0.00384444f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_498 N_VGND_c_794_n N_A_467_47#_c_907_n 0.0148867f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_499 N_VGND_c_783_n N_A_467_47#_c_951_n 0.0151751f $X=6.82 $Y=0.38 $X2=0 $Y2=0
cc_500 N_VGND_c_793_n N_A_467_47#_c_951_n 0.022989f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_501 N_VGND_c_794_n N_A_467_47#_c_951_n 0.0126169f $X=7.59 $Y=0 $X2=0 $Y2=0

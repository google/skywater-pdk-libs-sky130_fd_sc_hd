* File: sky130_fd_sc_hd__mux2_2.spice
* Created: Tue Sep  1 19:14:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2_2.pex.spice"
.subckt sky130_fd_sc_hd__mux2_2  VNB VPB A0 A1 S VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_79_21#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_79_21#_M1011_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.08775 PD=1.18458 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1004 A_288_47# N_A_257_199#_M1004_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.0761495 PD=0.745 PS=0.765421 NRD=30.708 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1008 N_A_79_21#_M1008_d N_A0_M1008_g A_288_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.17325 AS=0.06825 PD=1.245 PS=0.745 NRD=0 NRS=30.708 M=1 R=2.8 SA=75001.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_578_47# N_A1_M1002_g N_A_79_21#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.17325 PD=0.695 PS=1.245 NRD=23.568 NRS=9.996 M=1 R=2.8
+ SA=75002.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_S_M1010_g A_578_47# VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.05775 PD=0.69 PS=0.695 NRD=0 NRS=23.568 M=1 R=2.8 SA=75003 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_257_199#_M1013_d N_S_M1013_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0567 PD=1.38 PS=0.69 NRD=1.428 NRS=0 M=1 R=2.8 SA=75003.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_79_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_79_21#_M1009_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.216829 AS=0.135 PD=1.72561 PS=1.27 NRD=8.8453 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1012 A_306_369# N_A_257_199#_M1012_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2288 AS=0.138771 PD=1.355 PS=1.10439 NRD=93.1022 NRS=27.6982 M=1
+ R=4.26667 SA=75001.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1005 N_A_79_21#_M1005_d N_A1_M1005_g A_306_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1312 AS=0.2288 PD=1.05 PS=1.355 NRD=29.2348 NRS=93.1022 M=1 R=4.26667
+ SA=75002 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1001 A_591_369# N_A0_M1001_g N_A_79_21#_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1312 PD=0.85 PS=1.05 NRD=15.3857 NRS=10.7562 M=1 R=4.26667
+ SA=75002.6 SB=75001 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_S_M1003_g A_591_369# VPB PHIGHVT L=0.15 W=0.64 AD=0.0864
+ AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75003 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1000 N_A_257_199#_M1000_d N_S_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1728 AS=0.0864 PD=1.82 PS=0.91 NRD=1.5366 NRS=0 M=1 R=4.26667 SA=75003.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_73 VPB 0 1.28281e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__mux2_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdlclkp_4.pex.spice
* Created: Thu Aug 27 14:47:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%SCE 3 7 9 10 17
r27 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r28 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.16
+ $X2=0.215 $Y2=1.53
r29 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r30 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r31 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.165
r32 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r33 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%GATE 3 7 9 10 15 16
c42 16 0 2.81318e-20 $X=0.94 $Y=1.16
c43 15 0 9.56754e-20 $X=0.94 $Y=1.16
r44 15 18 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.915 $Y2=1.325
r45 15 17 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.915 $Y2=0.995
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r47 9 10 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.047 $Y=1.53
+ $X2=1.047 $Y2=1.87
r48 9 16 8.21746 $w=4.63e-07 $l=2.85e-07 $layer=LI1_cond $X=1.025 $Y=1.445
+ $X2=1.025 $Y2=1.16
r49 7 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.995
r50 3 18 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.83 $Y=2.165
+ $X2=0.83 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%A_257_147# 1 2 9 13 17 21 24 25 28 30 33
+ 35 37 41 44 53 54 57 60 68 74
c173 68 0 1.23968e-19 $X=1.78 $Y=1.74
c174 57 0 3.38573e-20 $X=1.615 $Y=1.53
c175 44 0 9.25246e-21 $X=4.1 $Y=1.19
c176 41 0 2.00517e-19 $X=1.615 $Y=1.325
c177 24 0 3.18278e-20 $X=1.45 $Y=0.87
c178 9 0 2.35132e-20 $X=1.375 $Y=0.415
r179 68 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.74
+ $X2=1.78 $Y2=1.905
r180 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=1.74 $X2=1.78 $Y2=1.74
r181 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.395 $Y=1.53
+ $X2=4.395 $Y2=1.53
r182 57 69 5.52036 $w=4.53e-07 $l=2.1e-07 $layer=LI1_cond $X=1.637 $Y=1.53
+ $X2=1.637 $Y2=1.74
r183 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.53
r184 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=1.53
+ $X2=1.615 $Y2=1.53
r185 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.25 $Y=1.53
+ $X2=4.395 $Y2=1.53
r186 53 54 3.08168 $w=1.4e-07 $l=2.49e-06 $layer=MET1_cond $X=4.25 $Y=1.53
+ $X2=1.76 $Y2=1.53
r187 44 74 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.1 $Y=1.19
+ $X2=4.1 $Y2=1.325
r188 44 73 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.1 $Y=1.19
+ $X2=4.1 $Y2=1.055
r189 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=1.19 $X2=4.1 $Y2=1.19
r190 41 57 5.38892 $w=4.53e-07 $l=2.05e-07 $layer=LI1_cond $X=1.637 $Y=1.325
+ $X2=1.637 $Y2=1.53
r191 40 41 3.94479 $w=4.53e-07 $l=1.2e-07 $layer=LI1_cond $X=1.615 $Y=1.205
+ $X2=1.615 $Y2=1.325
r192 35 37 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=4.72 $Y=0.615
+ $X2=4.72 $Y2=0.465
r193 31 61 3.79964 $w=2.5e-07 $l=1.53e-07 $layer=LI1_cond $X=4.48 $Y=1.62
+ $X2=4.327 $Y2=1.62
r194 31 33 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=4.48 $Y=1.62
+ $X2=4.81 $Y2=1.62
r195 29 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.335 $Y=0.7
+ $X2=4.72 $Y2=0.7
r196 29 30 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=4.335 $Y=0.785
+ $X2=4.335 $Y2=1.105
r197 28 61 3.10428 $w=3.05e-07 $l=1.25e-07 $layer=LI1_cond $X=4.327 $Y=1.495
+ $X2=4.327 $Y2=1.62
r198 27 30 0.521925 $w=1.68e-07 $l=8e-09 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.335 $Y2=1.19
r199 27 43 14.8096 $w=1.68e-07 $l=2.27e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.1 $Y2=1.19
r200 27 28 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=4.327 $Y=1.275
+ $X2=4.327 $Y2=1.495
r201 25 63 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=0.87
+ $X2=1.375 $Y2=0.87
r202 24 40 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0.87
+ $X2=1.535 $Y2=1.205
r203 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=0.87 $X2=1.45 $Y2=0.87
r204 21 74 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.05 $Y=1.835
+ $X2=4.05 $Y2=1.325
r205 17 73 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.05 $Y=0.445
+ $X2=4.05 $Y2=1.055
r206 13 71 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.84 $Y=2.275
+ $X2=1.84 $Y2=1.905
r207 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.375 $Y=0.735
+ $X2=1.375 $Y2=0.87
r208 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.375 $Y=0.735
+ $X2=1.375 $Y2=0.415
r209 2 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.675
+ $Y=1.515 $X2=4.81 $Y2=1.66
r210 1 37 182 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.68 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%A_257_243# 1 2 9 11 12 15 17 20 23 27 29
+ 30 36 37 40 41 42
c115 41 0 1.47482e-19 $X=1.96 $Y=0.87
c116 37 0 1.34642e-19 $X=3.935 $Y=0.85
c117 36 0 5.98268e-21 $X=3.935 $Y=0.85
c118 27 0 1.20845e-19 $X=3.84 $Y=1.66
c119 17 0 2.81318e-20 $X=1.9 $Y=1.215
c120 12 0 2.67301e-20 $X=1.435 $Y=1.29
c121 9 0 3.17216e-20 $X=1.36 $Y=2.275
r122 40 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=0.87
+ $X2=1.96 $Y2=1.035
r123 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=0.87
+ $X2=1.96 $Y2=0.705
r124 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=0.87 $X2=1.96 $Y2=0.87
r125 37 49 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.807 $Y=0.85
+ $X2=3.807 $Y2=0.935
r126 37 48 2.91128 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.807 $Y=0.85
+ $X2=3.807 $Y2=0.765
r127 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=0.85
+ $X2=3.935 $Y2=0.85
r128 32 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.075 $Y=0.85
+ $X2=2.075 $Y2=0.85
r129 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.22 $Y=0.85
+ $X2=2.075 $Y2=0.85
r130 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.79 $Y=0.85
+ $X2=3.935 $Y2=0.85
r131 29 30 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=3.79 $Y=0.85
+ $X2=2.22 $Y2=0.85
r132 24 27 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.68 $Y=1.66
+ $X2=3.84 $Y2=1.66
r133 23 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.575
+ $X2=3.68 $Y2=1.66
r134 23 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.68 $Y=1.575
+ $X2=3.68 $Y2=0.935
r135 20 48 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.76 $Y=0.465
+ $X2=3.76 $Y2=0.765
r136 17 43 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.9 $Y=1.215
+ $X2=1.9 $Y2=1.035
r137 15 42 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.9 $Y=0.415
+ $X2=1.9 $Y2=0.705
r138 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.9 $Y2=1.215
r139 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.435 $Y2=1.29
r140 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.36 $Y=1.365
+ $X2=1.435 $Y2=1.29
r141 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.36 $Y=1.365
+ $X2=1.36 $Y2=2.275
r142 2 27 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=1.515 $X2=3.84 $Y2=1.66
r143 1 20 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=3.715
+ $Y=0.235 $X2=3.84 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%A_465_315# 1 2 9 13 17 20 22 26 30 32 36
+ 37 41 43 44 49
c129 41 0 1.77265e-19 $X=2.46 $Y=1.74
c130 32 0 5.5315e-20 $X=5.165 $Y=2
c131 13 0 1.38699e-19 $X=2.51 $Y=0.445
r132 41 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.74
+ $X2=2.46 $Y2=1.905
r133 41 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.74
+ $X2=2.46 $Y2=1.575
r134 40 43 3.38343 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.74
+ $X2=2.545 $Y2=1.74
r135 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.74 $X2=2.46 $Y2=1.74
r136 37 50 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.445 $Y=1.16
+ $X2=5.445 $Y2=1.325
r137 37 49 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.445 $Y=1.16
+ $X2=5.445 $Y2=0.995
r138 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.39
+ $Y=1.16 $X2=5.39 $Y2=1.16
r139 34 36 24.8598 $w=3.48e-07 $l=7.55e-07 $layer=LI1_cond $X=5.34 $Y=1.915
+ $X2=5.34 $Y2=1.16
r140 33 44 3.05 $w=1.7e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.405 $Y=2
+ $X2=3.295 $Y2=1.86
r141 32 34 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.165 $Y=2
+ $X2=5.34 $Y2=1.915
r142 32 33 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=5.165 $Y=2
+ $X2=3.405 $Y2=2
r143 28 44 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.295 $Y=2.085
+ $X2=3.295 $Y2=1.86
r144 28 30 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=3.295 $Y=2.085
+ $X2=3.295 $Y2=2.205
r145 24 44 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.295 $Y=1.635
+ $X2=3.295 $Y2=1.86
r146 24 26 63.6463 $w=2.18e-07 $l=1.215e-06 $layer=LI1_cond $X=3.295 $Y=1.635
+ $X2=3.295 $Y2=0.42
r147 22 44 3.05 $w=2.7e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.185 $Y=1.77
+ $X2=3.295 $Y2=1.86
r148 22 43 27.3172 $w=2.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.185 $Y=1.77
+ $X2=2.545 $Y2=1.77
r149 20 50 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.56 $Y=1.985
+ $X2=5.56 $Y2=1.325
r150 17 49 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.56 $Y=0.56
+ $X2=5.56 $Y2=0.995
r151 13 46 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.51 $Y=0.445
+ $X2=2.51 $Y2=1.575
r152 9 47 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.43 $Y=2.275
+ $X2=2.43 $Y2=1.905
r153 2 30 600 $w=1.7e-07 $l=7.84602e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=2.205
r154 1 26 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.235 $X2=3.32 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%A_287_413# 1 2 7 9 12 14 18 23 25 26 28 35
c99 28 0 1.77265e-19 $X=2.93 $Y=1.16
c100 26 0 3.17216e-20 $X=2.5 $Y=1.185
c101 25 0 3.18278e-20 $X=2.415 $Y=0.995
c102 14 0 2.67301e-20 $X=2.33 $Y=0.395
r103 31 32 14.6301 $w=2.46e-07 $l=2.95e-07 $layer=LI1_cond $X=2.12 $Y=1.205
+ $X2=2.415 $Y2=1.205
r104 29 35 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.93 $Y=1.16
+ $X2=3.11 $Y2=1.16
r105 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.16 $X2=2.93 $Y2=1.16
r106 26 32 4.2431 $w=3.8e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.5 $Y=1.185
+ $X2=2.415 $Y2=1.205
r107 26 28 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.5 $Y=1.185
+ $X2=2.93 $Y2=1.185
r108 25 32 2.90119 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.415 $Y=0.995
+ $X2=2.415 $Y2=1.205
r109 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.415 $Y=0.535
+ $X2=2.415 $Y2=0.995
r110 22 31 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.12 $Y=1.375
+ $X2=2.12 $Y2=1.205
r111 22 23 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.12 $Y=1.375
+ $X2=2.12 $Y2=2.125
r112 18 23 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.035 $Y=2.295
+ $X2=2.12 $Y2=2.125
r113 18 20 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=2.035 $Y=2.295
+ $X2=1.6 $Y2=2.295
r114 14 24 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.33 $Y=0.395
+ $X2=2.415 $Y2=0.535
r115 14 16 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=2.33 $Y=0.395
+ $X2=1.635 $Y2=0.395
r116 10 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r117 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.985
r118 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=1.16
r119 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=0.56
r120 2 20 600 $w=1.7e-07 $l=3.22102e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=2.065 $X2=1.6 $Y2=2.315
r121 1 16 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.635 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%CLK 3 5 8 11 14 16 17 18 20 21 27 31 33 35
+ 36 37
c97 35 0 7.75798e-20 $X=5.98 $Y=1.16
c98 33 0 1.20845e-19 $X=4.735 $Y=1.325
c99 21 0 9.25246e-21 $X=5 $Y=1.19
c100 18 0 1.33709e-19 $X=4.855 $Y=1.19
c101 17 0 1.40624e-19 $X=4.67 $Y=0.88
c102 14 0 5.5315e-20 $X=5.98 $Y=1.985
r103 35 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.98 $Y=1.16
+ $X2=5.98 $Y2=0.995
r104 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.98
+ $Y=1.16 $X2=5.98 $Y2=1.16
r105 31 33 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.16
+ $X2=4.735 $Y2=1.325
r106 28 36 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=5.795 $Y=1.16
+ $X2=5.98 $Y2=1.16
r107 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.795 $Y=1.19
+ $X2=5.795 $Y2=1.19
r108 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5 $Y=1.19
+ $X2=4.855 $Y2=1.19
r109 20 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.65 $Y=1.19
+ $X2=5.795 $Y2=1.19
r110 20 21 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=5.65 $Y=1.19 $X2=5
+ $Y2=1.19
r111 18 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.81
+ $Y=1.16 $X2=4.81 $Y2=1.16
r112 18 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.855 $Y=1.19
+ $X2=4.855 $Y2=1.19
r113 16 17 44.1654 $w=4.2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.67 $Y=0.73
+ $X2=4.67 $Y2=0.88
r114 12 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.98 $Y=1.325
+ $X2=5.98 $Y2=1.16
r115 12 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.98 $Y=1.325
+ $X2=5.98 $Y2=1.985
r116 11 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.92 $Y=0.56
+ $X2=5.92 $Y2=0.995
r117 8 33 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.6 $Y=1.835 $X2=4.6
+ $Y2=1.325
r118 5 31 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=4.735 $Y=1.115
+ $X2=4.735 $Y2=1.16
r119 5 17 31.1181 $w=4.2e-07 $l=2.35e-07 $layer=POLY_cond $X=4.735 $Y=1.115
+ $X2=4.735 $Y2=0.88
r120 3 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.47 $Y=0.445
+ $X2=4.47 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%A_1045_47# 1 2 9 13 17 21 25 29 33 37 39
+ 41 45 47 48 53 59 61 67
c136 67 0 1.27353e-19 $X=7.715 $Y=1.16
c137 61 0 5.45858e-20 $X=6.325 $Y=1.185
c138 47 0 7.75798e-20 $X=6.325 $Y=1.495
c139 37 0 1.09886e-19 $X=7.715 $Y=1.985
c140 33 0 1.24697e-19 $X=7.715 $Y=0.56
c141 21 0 1.33408e-19 $X=6.875 $Y=1.985
r142 66 67 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.295 $Y=1.16
+ $X2=7.715 $Y2=1.16
r143 65 66 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.875 $Y=1.16
+ $X2=7.295 $Y2=1.16
r144 57 59 11.2512 $w=5.88e-07 $l=5.55e-07 $layer=LI1_cond $X=5.77 $Y=1.79
+ $X2=6.325 $Y2=1.79
r145 53 55 6.58539 $w=4.18e-07 $l=2.4e-07 $layer=LI1_cond $X=5.225 $Y=0.46
+ $X2=5.225 $Y2=0.7
r146 51 65 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=6.545 $Y=1.16
+ $X2=6.875 $Y2=1.16
r147 51 62 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.545 $Y=1.16
+ $X2=6.455 $Y2=1.16
r148 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.545
+ $Y=1.16 $X2=6.545 $Y2=1.16
r149 48 61 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=1.185
+ $X2=6.325 $Y2=1.185
r150 48 50 6.33462 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=6.41 $Y=1.185
+ $X2=6.545 $Y2=1.185
r151 47 59 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.325 $Y=1.495
+ $X2=6.325 $Y2=1.79
r152 46 61 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.325 $Y=1.315
+ $X2=6.325 $Y2=1.185
r153 46 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.325 $Y=1.315
+ $X2=6.325 $Y2=1.495
r154 45 61 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.325 $Y=1.055
+ $X2=6.325 $Y2=1.185
r155 44 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.325 $Y=0.785
+ $X2=6.325 $Y2=1.055
r156 41 57 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=5.77 $Y=2.085
+ $X2=5.77 $Y2=1.79
r157 41 43 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=5.77 $Y=2.085 $X2=5.77
+ $Y2=2.125
r158 40 55 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.435 $Y=0.7
+ $X2=5.225 $Y2=0.7
r159 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.24 $Y=0.7
+ $X2=6.325 $Y2=0.785
r160 39 40 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=6.24 $Y=0.7
+ $X2=5.435 $Y2=0.7
r161 35 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.715 $Y=1.295
+ $X2=7.715 $Y2=1.16
r162 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.715 $Y=1.295
+ $X2=7.715 $Y2=1.985
r163 31 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.715 $Y=1.025
+ $X2=7.715 $Y2=1.16
r164 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.715 $Y=1.025
+ $X2=7.715 $Y2=0.56
r165 27 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.295 $Y=1.295
+ $X2=7.295 $Y2=1.16
r166 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.295 $Y=1.295
+ $X2=7.295 $Y2=1.985
r167 23 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.295 $Y=1.025
+ $X2=7.295 $Y2=1.16
r168 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.295 $Y=1.025
+ $X2=7.295 $Y2=0.56
r169 19 65 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.875 $Y=1.295
+ $X2=6.875 $Y2=1.16
r170 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.875 $Y=1.295
+ $X2=6.875 $Y2=1.985
r171 15 65 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.875 $Y=1.025
+ $X2=6.875 $Y2=1.16
r172 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.875 $Y=1.025
+ $X2=6.875 $Y2=0.56
r173 11 62 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.455 $Y=1.295
+ $X2=6.455 $Y2=1.16
r174 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.455 $Y=1.295
+ $X2=6.455 $Y2=1.985
r175 7 62 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.455 $Y=1.025
+ $X2=6.455 $Y2=1.16
r176 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.455 $Y=1.025
+ $X2=6.455 $Y2=0.56
r177 2 43 600 $w=1.7e-07 $l=7.04273e-07 $layer=licon1_PDIFF $count=1 $X=5.635
+ $Y=1.485 $X2=5.77 $Y2=2.125
r178 1 53 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.225
+ $Y=0.235 $X2=5.35 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 34 36 40 42
+ 43 57 63 68 73 84 87 93 95 98 102
c116 32 0 1.27353e-19 $X=7.085 $Y=2
r117 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r118 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 92 93 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=2.53
+ $X2=5.515 $Y2=2.53
r121 89 92 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=5.29 $Y=2.53 $X2=5.35
+ $Y2=2.53
r122 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r123 86 87 11.8978 $w=7.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.795 $Y=2.44
+ $X2=3.015 $Y2=2.44
r124 82 86 4.34193 $w=7.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.795 $Y2=2.44
r125 82 84 10.8328 $w=7.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.375 $Y2=2.44
r126 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r127 77 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r128 77 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r129 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r130 74 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.25 $Y=2.72
+ $X2=7.125 $Y2=2.72
r131 74 76 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.25 $Y=2.72
+ $X2=7.59 $Y2=2.72
r132 73 101 4.56302 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=7.89 $Y=2.72
+ $X2=8.085 $Y2=2.72
r133 73 76 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.89 $Y=2.72 $X2=7.59
+ $Y2=2.72
r134 72 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r135 72 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r136 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r137 69 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.22 $Y2=2.72
r138 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.67 $Y2=2.72
r139 68 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7 $Y=2.72 $X2=7.125
+ $Y2=2.72
r140 68 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7 $Y=2.72 $X2=6.67
+ $Y2=2.72
r141 67 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r142 67 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r143 66 93 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=5.515 $Y2=2.72
r144 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r145 63 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=6.22 $Y2=2.72
r146 63 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=5.75 $Y2=2.72
r147 60 90 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r148 59 62 9.02495 $w=5.48e-07 $l=4.15e-07 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=4.325 $Y2=2.53
r149 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r150 57 89 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=5.24 $Y=2.53 $X2=5.29
+ $Y2=2.53
r151 57 62 19.8984 $w=5.48e-07 $l=9.15e-07 $layer=LI1_cond $X=5.24 $Y=2.53
+ $X2=4.325 $Y2=2.53
r152 56 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r153 56 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r154 55 87 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.015 $Y2=2.72
r155 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r156 52 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r157 51 84 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.375 $Y2=2.72
r158 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 49 52 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r160 48 51 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r161 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r162 46 79 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r163 46 48 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r164 43 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r165 43 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r166 42 55 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.45 $Y2=2.72
r167 40 59 0.869875 $w=5.48e-07 $l=4e-08 $layer=LI1_cond $X=3.87 $Y=2.53
+ $X2=3.91 $Y2=2.53
r168 40 42 12.2241 $w=5.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.87 $Y=2.53
+ $X2=3.595 $Y2=2.53
r169 36 39 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=8.042 $Y=1.66
+ $X2=8.042 $Y2=2.34
r170 34 101 2.99522 $w=3.05e-07 $l=1.04307e-07 $layer=LI1_cond $X=8.042 $Y=2.635
+ $X2=8.085 $Y2=2.72
r171 34 39 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=8.042 $Y=2.635
+ $X2=8.042 $Y2=2.34
r172 30 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=2.635
+ $X2=7.125 $Y2=2.72
r173 30 32 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.125 $Y=2.635
+ $X2=7.125 $Y2=2
r174 26 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2.72
r175 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2.36
r176 22 79 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r177 22 24 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r178 7 39 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=7.79
+ $Y=1.485 $X2=7.975 $Y2=2.34
r179 7 36 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=7.79
+ $Y=1.485 $X2=7.975 $Y2=1.66
r180 6 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.95
+ $Y=1.485 $X2=7.085 $Y2=2
r181 5 28 600 $w=1.7e-07 $l=9.53939e-07 $layer=licon1_PDIFF $count=1 $X=6.055
+ $Y=1.485 $X2=6.22 $Y2=2.36
r182 4 92 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=5.205
+ $Y=1.485 $X2=5.35 $Y2=2.36
r183 3 62 600 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=1.515 $X2=4.325 $Y2=2.34
r184 2 86 600 $w=1.7e-07 $l=4.15421e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=2.065 $X2=2.795 $Y2=2.36
r185 1 24 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%A_27_47# 1 2 3 12 15 16 17 18 20 24
r49 22 24 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.105 $Y=0.615
+ $X2=1.105 $Y2=0.42
r50 18 20 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=0.685 $Y=2.295
+ $X2=1.095 $Y2=2.295
r51 17 28 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.7 $X2=0.6
+ $Y2=0.7
r52 16 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.015 $Y=0.7
+ $X2=1.105 $Y2=0.615
r53 16 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.015 $Y=0.7
+ $X2=0.685 $Y2=0.7
r54 15 18 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.6 $Y=2.125
+ $X2=0.685 $Y2=2.295
r55 14 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=0.785 $X2=0.6
+ $Y2=0.7
r56 14 15 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=0.6 $Y=0.785
+ $X2=0.6 $Y2=2.125
r57 10 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.6 $Y2=0.7
r58 10 12 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.43
r59 3 20 600 $w=1.7e-07 $l=5.31578e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.845 $X2=1.095 $Y2=2.29
r60 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%GCLK 1 2 3 4 13 14 15 16 18 20 23 24 25 26
+ 27 28 29 30 31 32 47 57 73
c74 28 0 1.93102e-19 $X=7.635 $Y=1.19
c75 15 0 1.09886e-19 $X=7.05 $Y=1.57
c76 13 0 1.24697e-19 $X=7.05 $Y=0.8
r77 47 80 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=6.705 $Y=0.51
+ $X2=6.705 $Y2=0.445
r78 32 73 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=8.095 $Y=1.185
+ $X2=8.05 $Y2=1.185
r79 30 31 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=7.57 $Y=1.87 $X2=7.57
+ $Y2=2.21
r80 30 65 2.11281 $w=2.98e-07 $l=5.5e-08 $layer=LI1_cond $X=7.57 $Y=1.87
+ $X2=7.57 $Y2=1.815
r81 29 65 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=7.57 $Y=1.53
+ $X2=7.57 $Y2=1.815
r82 29 55 8.25918 $w=2.98e-07 $l=2.15e-07 $layer=LI1_cond $X=7.57 $Y=1.53
+ $X2=7.57 $Y2=1.315
r83 28 55 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=7.635 $Y=1.185
+ $X2=7.57 $Y2=1.185
r84 28 73 10.6322 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=7.72 $Y=1.185
+ $X2=8.05 $Y2=1.185
r85 27 55 7.87503 $w=2.98e-07 $l=2.05e-07 $layer=LI1_cond $X=7.57 $Y=0.85
+ $X2=7.57 $Y2=1.055
r86 27 57 16.5184 $w=2.98e-07 $l=4.3e-07 $layer=LI1_cond $X=7.57 $Y=0.85
+ $X2=7.57 $Y2=0.42
r87 26 55 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=7.175 $Y=1.185
+ $X2=7.57 $Y2=1.185
r88 26 81 1.77299 $w=2.58e-07 $l=4e-08 $layer=LI1_cond $X=7.175 $Y=1.185
+ $X2=7.135 $Y2=1.185
r89 24 25 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.705 $Y=1.815
+ $X2=6.705 $Y2=2.21
r90 23 80 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.665 $Y=0.36
+ $X2=6.665 $Y2=0.445
r91 23 47 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.705 $Y=0.52
+ $X2=6.705 $Y2=0.51
r92 22 24 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=6.705 $Y=1.655
+ $X2=6.705 $Y2=1.815
r93 21 23 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=6.705 $Y=0.715
+ $X2=6.705 $Y2=0.52
r94 19 81 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.135 $Y=1.315
+ $X2=7.135 $Y2=1.185
r95 19 20 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.135 $Y=1.315
+ $X2=7.135 $Y2=1.485
r96 18 81 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.135 $Y=1.055
+ $X2=7.135 $Y2=1.185
r97 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.135 $Y=0.885
+ $X2=7.135 $Y2=1.055
r98 16 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.83 $Y=1.57
+ $X2=6.705 $Y2=1.655
r99 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=1.57
+ $X2=7.135 $Y2=1.485
r100 15 16 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.05 $Y=1.57
+ $X2=6.83 $Y2=1.57
r101 14 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.83 $Y=0.8
+ $X2=6.705 $Y2=0.715
r102 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=0.8
+ $X2=7.135 $Y2=0.885
r103 13 14 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.05 $Y=0.8
+ $X2=6.83 $Y2=0.8
r104 4 65 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=7.37
+ $Y=1.485 $X2=7.505 $Y2=1.815
r105 3 24 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=6.53
+ $Y=1.485 $X2=6.665 $Y2=1.815
r106 2 57 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.37
+ $Y=0.235 $X2=7.505 $Y2=0.42
r107 1 23 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.53
+ $Y=0.235 $X2=6.665 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_4%VGND 1 2 3 4 5 6 21 25 29 33 35 37 39 41
+ 46 54 64 69 75 78 81 86 92 94 98
r129 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r130 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r131 90 92 8.68883 $w=5.28e-07 $l=1.2e-07 $layer=LI1_cond $X=6.21 $Y=0.18
+ $X2=6.33 $Y2=0.18
r132 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r133 88 90 1.01554 $w=5.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.165 $Y=0.18
+ $X2=6.21 $Y2=0.18
r134 85 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r135 84 88 9.36552 $w=5.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.75 $Y=0.18
+ $X2=6.165 $Y2=0.18
r136 84 86 9.25302 $w=5.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.75 $Y=0.18
+ $X2=5.605 $Y2=0.18
r137 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r138 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r139 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r140 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r141 73 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r142 73 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r143 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r144 70 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.25 $Y=0 $X2=7.125
+ $Y2=0
r145 70 72 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.25 $Y=0 $X2=7.59
+ $Y2=0
r146 69 97 4.56302 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=7.89 $Y=0 $X2=8.085
+ $Y2=0
r147 69 72 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.89 $Y=0 $X2=7.59
+ $Y2=0
r148 68 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r149 68 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r150 67 92 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.33
+ $Y2=0
r151 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r152 64 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7 $Y=0 $X2=7.125
+ $Y2=0
r153 64 67 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7 $Y=0 $X2=6.67
+ $Y2=0
r154 63 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r155 63 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r156 62 86 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.605 $Y2=0
r157 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r158 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.26
+ $Y2=0
r159 60 62 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.425 $Y=0
+ $X2=5.29 $Y2=0
r160 58 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r161 58 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r162 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r163 55 78 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.015 $Y=0
+ $X2=2.842 $Y2=0
r164 55 57 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.015 $Y=0
+ $X2=3.91 $Y2=0
r165 54 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0 $X2=4.26
+ $Y2=0
r166 54 57 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=3.91 $Y2=0
r167 53 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r168 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r169 50 53 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.53 $Y2=0
r170 50 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r171 49 52 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r172 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r173 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r174 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r175 46 78 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.842
+ $Y2=0
r176 46 52 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.53
+ $Y2=0
r177 41 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r178 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r179 39 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r180 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r181 35 97 2.99522 $w=3.05e-07 $l=1.04307e-07 $layer=LI1_cond $X=8.042 $Y=0.085
+ $X2=8.085 $Y2=0
r182 35 37 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=8.042 $Y=0.085
+ $X2=8.042 $Y2=0.38
r183 31 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.085
+ $X2=7.125 $Y2=0
r184 31 33 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.125 $Y=0.085
+ $X2=7.125 $Y2=0.38
r185 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0
r186 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0.36
r187 23 78 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.842 $Y=0.085
+ $X2=2.842 $Y2=0
r188 23 25 14.1968 $w=3.43e-07 $l=4.25e-07 $layer=LI1_cond $X=2.842 $Y=0.085
+ $X2=2.842 $Y2=0.51
r189 19 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r190 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r191 6 37 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.235 $X2=7.975 $Y2=0.38
r192 5 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.235 $X2=7.085 $Y2=0.38
r193 4 88 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=5.995
+ $Y=0.235 $X2=6.165 $Y2=0.36
r194 3 29 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.125
+ $Y=0.235 $X2=4.26 $Y2=0.36
r195 2 25 182 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.815 $Y2=0.51
r196 1 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__sdfsbp_1.spice
* Created: Thu Aug 27 14:46:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfsbp_1.spice.pex"
.subckt sky130_fd_sc_hd__sdfsbp_1  VNB VPB SCD SCE D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1039 A_109_47# N_SCD_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1012 N_A_181_47#_M1012_d N_SCE_M1012_g A_109_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1022 A_265_47# N_D_M1022_g N_A_181_47#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_319_21#_M1031_g A_265_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1218 AS=0.0567 PD=1.42 PS=0.69 NRD=7.14 NRS=22.848 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_SCE_M1013_g N_A_319_21#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_CLK_M1000_g N_A_643_369#_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1036 N_A_809_369#_M1036_d N_A_643_369#_M1036_g N_VGND_M1000_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_997_413#_M1023_d N_A_643_369#_M1023_g N_A_181_47#_M1023_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1024 A_1087_47# N_A_809_369#_M1024_g N_A_997_413#_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_1129_21#_M1025_g A_1087_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_1347_47# N_A_997_413#_M1009_g N_A_1129_21#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1041 N_VGND_M1041_d N_SET_B_M1041_g A_1347_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0758774 AS=0.0441 PD=0.764717 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1014 A_1514_47# N_A_997_413#_M1014_g N_VGND_M1041_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2224 AS=0.115623 PD=1.335 PS=1.16528 NRD=54.84 NRS=9.372 M=1 R=4.26667
+ SA=75000.7 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1006 N_A_1587_329#_M1006_d N_A_809_369#_M1006_g A_1514_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.152392 AS=0.2224 PD=1.34038 PS=1.335 NRD=3.744 NRS=54.84 M=1
+ R=4.26667 SA=75001.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1015 A_1807_47# N_A_643_369#_M1015_g N_A_1587_329#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.100008 PD=0.63 PS=0.879623 NRD=14.28 NRS=48.564 M=1
+ R=2.8 SA=75002.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1018 A_1879_47# N_A_1770_295#_M1018_g A_1807_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1029 AS=0.0441 PD=0.91 PS=0.63 NRD=54.276 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_SET_B_M1010_g A_1879_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.08505 AS=0.1029 PD=0.825 PS=0.91 NRD=37.14 NRS=54.276 M=1 R=2.8
+ SA=75003.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1020 N_A_1770_295#_M1020_d N_A_1587_329#_M1020_g N_VGND_M1010_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.08505 PD=1.36 PS=0.825 NRD=0 NRS=0 M=1 R=2.8
+ SA=75004 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_Q_N_M1005_d N_A_1587_329#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1033 N_VGND_M1033_d N_A_1587_329#_M1033_g N_A_2412_47#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_Q_M1019_d N_A_2412_47#_M1019_g N_VGND_M1033_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1021 N_VPWR_M1021_d N_SCD_M1021_g N_A_27_369#_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 A_193_369# N_SCE_M1002_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1004 N_A_181_47#_M1004_d N_D_M1004_g A_193_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_27_369#_M1001_d N_A_319_21#_M1001_g N_A_181_47#_M1004_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_VPWR_M1026_d N_SCE_M1026_g N_A_319_21#_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.1664 PD=1.8 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_CLK_M1034_g N_A_643_369#_M1034_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1030 N_A_809_369#_M1030_d N_A_643_369#_M1030_g N_VPWR_M1034_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_997_413#_M1007_d N_A_809_369#_M1007_g N_A_181_47#_M1007_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1035 A_1081_413# N_A_643_369#_M1035_g N_A_997_413#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0756 AS=0.0567 PD=0.78 PS=0.69 NRD=58.6272 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1037 N_VPWR_M1037_d N_A_1129_21#_M1037_g A_1081_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0924 AS=0.0756 PD=0.86 PS=0.78 NRD=25.7873 NRS=58.6272 M=1 R=2.8
+ SA=75001.1 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_1129_21#_M1008_d N_A_997_413#_M1008_g N_VPWR_M1037_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.07035 AS=0.0924 PD=0.755 PS=0.86 NRD=7.0329 NRS=49.25 M=1
+ R=2.8 SA=75001.7 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_SET_B_M1032_g N_A_1129_21#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0952 AS=0.07035 PD=0.846667 PS=0.755 NRD=18.7544 NRS=18.7544 M=1
+ R=2.8 SA=75002.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1016 A_1514_329# N_A_997_413#_M1016_g N_VPWR_M1032_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.0903 AS=0.1904 PD=1.055 PS=1.69333 NRD=12.2928 NRS=25.7873 M=1 R=5.6
+ SA=75001.5 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1017 N_A_1587_329#_M1017_d N_A_643_369#_M1017_g A_1514_329# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.203 AS=0.0903 PD=1.75333 PS=1.055 NRD=32.8202 NRS=12.2928 M=1
+ R=5.6 SA=75001.8 SB=75001 A=0.126 P=1.98 MULT=1
MM1040 A_1712_413# N_A_809_369#_M1040_g N_A_1587_329#_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0609 AS=0.1015 PD=0.71 PS=0.876667 NRD=42.1974 NRS=25.7873 M=1
+ R=2.8 SA=75003.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_1770_295#_M1011_g A_1712_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.10395 AS=0.0609 PD=0.915 PS=0.71 NRD=103.189 NRS=42.1974 M=1 R=2.8
+ SA=75004.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1028 N_A_1587_329#_M1028_d N_SET_B_M1028_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.10395 PD=1.36 PS=0.915 NRD=0 NRS=0 M=1 R=2.8 SA=75004.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 N_A_1770_295#_M1038_d N_A_1587_329#_M1038_g N_VPWR_M1038_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_Q_N_M1029_d N_A_1587_329#_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1027 N_VPWR_M1027_d N_A_1587_329#_M1027_g N_A_2412_47#_M1027_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_Q_M1003_d N_A_2412_47#_M1003_g N_VPWR_M1027_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX42_noxref VNB VPB NWDIODE A=22.0206 P=30.65
c_131 VNB 0 1.07953e-19 $X=0.15 $Y=-0.085
c_282 VPB 0 1.93782e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__sdfsbp_1.spice.SKY130_FD_SC_HD__SDFSBP_1.pxi"
*
.ends
*
*

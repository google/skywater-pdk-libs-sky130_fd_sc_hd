* File: sky130_fd_sc_hd__o31ai_2.spice
* Created: Tue Sep  1 19:25:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o31ai_2.pex.spice"
.subckt sky130_fd_sc_hd__o31ai_2  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_47#_M1003_d N_A1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_A1_M1005_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_27_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.08775 PD=1.26 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1002_d N_A2_M1009_g N_A_27_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.12675 PD=1.26 PS=1.04 NRD=0 NRS=6.456 M=1 R=4.33333 SA=75001.8
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1009_s N_A3_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.11375 PD=1.04 PS=1 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1015 N_A_27_47#_M1015_d N_A3_M1015_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75002.8
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1015_d N_B1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75003.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_27_47#_M1010_d N_B1_M1010_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12675 PD=1.82 PS=1.04 NRD=0 NRS=6.456 M=1 R=4.33333 SA=75003.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1001_d N_A1_M1013_g N_A_27_297#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1006 N_A_27_297#_M1013_s N_A2_M1006_g N_A_281_297#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_297#_M1008_d N_A2_M1008_g N_A_281_297#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_A3_M1007_g N_A_281_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1011 N_Y_M1011_d N_A3_M1011_g N_A_281_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1011_d VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.135 PD=1.39 PS=1.27 NRD=14.7553 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1000_d N_B1_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.26 PD=1.39 PS=2.52 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75001.6 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__o31ai_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__and4bb_1.pxi.spice
* Created: Thu Aug 27 14:09:01 2020
* 
x_PM_SKY130_FD_SC_HD__AND4BB_1%A_N N_A_N_M1007_g N_A_N_M1006_g A_N N_A_N_c_101_n
+ N_A_N_c_102_n PM_SKY130_FD_SC_HD__AND4BB_1%A_N
x_PM_SKY130_FD_SC_HD__AND4BB_1%B_N N_B_N_M1009_g N_B_N_M1012_g N_B_N_c_135_n
+ N_B_N_c_136_n B_N PM_SKY130_FD_SC_HD__AND4BB_1%B_N
x_PM_SKY130_FD_SC_HD__AND4BB_1%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1006_s
+ N_A_27_47#_c_181_n N_A_27_47#_c_182_n N_A_27_47#_M1011_g N_A_27_47#_M1008_g
+ N_A_27_47#_c_183_n N_A_27_47#_c_191_n N_A_27_47#_c_192_n N_A_27_47#_c_184_n
+ N_A_27_47#_c_193_n N_A_27_47#_c_185_n N_A_27_47#_c_195_n N_A_27_47#_c_186_n
+ N_A_27_47#_c_187_n N_A_27_47#_c_197_n N_A_27_47#_c_188_n
+ PM_SKY130_FD_SC_HD__AND4BB_1%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4BB_1%A_223_47# N_A_223_47#_M1009_d N_A_223_47#_M1012_d
+ N_A_223_47#_M1001_g N_A_223_47#_M1002_g N_A_223_47#_c_290_n
+ N_A_223_47#_c_273_n N_A_223_47#_c_282_n N_A_223_47#_c_283_n
+ N_A_223_47#_c_274_n N_A_223_47#_c_275_n N_A_223_47#_c_276_n
+ N_A_223_47#_c_286_n N_A_223_47#_c_277_n N_A_223_47#_c_278_n
+ N_A_223_47#_c_279_n N_A_223_47#_c_280_n PM_SKY130_FD_SC_HD__AND4BB_1%A_223_47#
x_PM_SKY130_FD_SC_HD__AND4BB_1%C N_C_M1000_g N_C_M1004_g C C C C N_C_c_374_n
+ N_C_c_375_n PM_SKY130_FD_SC_HD__AND4BB_1%C
x_PM_SKY130_FD_SC_HD__AND4BB_1%D N_D_c_417_n N_D_M1010_g N_D_M1003_g D D D D
+ N_D_c_420_n PM_SKY130_FD_SC_HD__AND4BB_1%D
x_PM_SKY130_FD_SC_HD__AND4BB_1%A_343_93# N_A_343_93#_M1011_s N_A_343_93#_M1008_d
+ N_A_343_93#_M1004_d N_A_343_93#_M1005_g N_A_343_93#_M1013_g
+ N_A_343_93#_c_462_n N_A_343_93#_c_463_n N_A_343_93#_c_482_n
+ N_A_343_93#_c_469_n N_A_343_93#_c_503_n N_A_343_93#_c_470_n
+ N_A_343_93#_c_464_n N_A_343_93#_c_465_n N_A_343_93#_c_473_n
+ N_A_343_93#_c_474_n N_A_343_93#_c_466_n PM_SKY130_FD_SC_HD__AND4BB_1%A_343_93#
x_PM_SKY130_FD_SC_HD__AND4BB_1%VPWR N_VPWR_M1006_d N_VPWR_M1008_s N_VPWR_M1002_d
+ N_VPWR_M1003_d N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n VPWR
+ N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_553_n N_VPWR_c_565_n N_VPWR_c_566_n
+ PM_SKY130_FD_SC_HD__AND4BB_1%VPWR
x_PM_SKY130_FD_SC_HD__AND4BB_1%X N_X_M1005_d N_X_M1013_d X X X X X N_X_c_630_n
+ PM_SKY130_FD_SC_HD__AND4BB_1%X
x_PM_SKY130_FD_SC_HD__AND4BB_1%VGND N_VGND_M1007_d N_VGND_M1010_d N_VGND_c_642_n
+ N_VGND_c_643_n VGND N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n
+ N_VGND_c_647_n N_VGND_c_648_n PM_SKY130_FD_SC_HD__AND4BB_1%VGND
cc_1 VNB N_A_N_M1007_g 0.0485608f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.445
cc_2 VNB N_B_N_M1009_g 0.0269569f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.445
cc_3 VNB N_B_N_M1012_g 0.00876222f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=2.275
cc_4 VNB N_B_N_c_135_n 0.0034985f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.74
cc_5 VNB N_B_N_c_136_n 0.0294168f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.74
cc_6 VNB B_N 0.00441802f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.605
cc_7 VNB N_A_27_47#_c_181_n 0.0195365f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=2.275
cc_8 VNB N_A_27_47#_c_182_n 0.0116556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_183_n 0.0322341f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.74
cc_10 VNB N_A_27_47#_c_184_n 0.0339472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_185_n 0.0119841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_186_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_187_n 9.40304e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_188_n 7.42329e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_223_47#_c_273_n 0.0111109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_223_47#_c_274_n 0.0234873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_223_47#_c_275_n 0.00693987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_223_47#_c_276_n 0.00115074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_223_47#_c_277_n 0.00107416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_223_47#_c_278_n 0.0245205f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_223_47#_c_279_n 0.0159573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_223_47#_c_280_n 0.0274056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB C 0.00267896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB C 0.00379285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_C_c_374_n 0.0217254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_C_c_375_n 0.0298708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_D_c_417_n 0.0323823f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.605
cc_28 VNB D 0.00204978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB D 0.00238997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_D_c_420_n 0.0217406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_343_93#_c_462_n 0.00248341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_343_93#_c_463_n 0.00223177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_343_93#_c_464_n 0.00213406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_343_93#_c_465_n 0.0495199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_343_93#_c_466_n 0.0206453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_553_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_630_n 0.0405911f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.87
cc_38 VNB N_VGND_c_642_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.74
cc_39 VNB N_VGND_c_643_n 0.00536564f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.875
cc_40 VNB N_VGND_c_644_n 0.0702445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_645_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_646_n 0.273097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_647_n 0.0238568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_648_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VPB N_A_N_M1007_g 0.0174512f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.445
cc_46 VPB N_A_N_M1006_g 0.0241623f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=2.275
cc_47 VPB N_A_N_c_101_n 0.0281827f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.74
cc_48 VPB N_A_N_c_102_n 0.00678501f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.74
cc_49 VPB N_B_N_M1012_g 0.0525232f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=2.275
cc_50 VPB N_A_27_47#_c_182_n 0.0148747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_M1008_g 0.0253614f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.605
cc_52 VPB N_A_27_47#_c_191_n 0.0438528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_192_n 0.022989f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.87
cc_54 VPB N_A_27_47#_c_193_n 0.032102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_185_n 0.0141184f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_195_n 0.00511147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_187_n 0.00704895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_197_n 0.0129899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_188_n 0.00671189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_223_47#_M1002_g 0.0508144f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.74
cc_61 VPB N_A_223_47#_c_282_n 0.00862973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_223_47#_c_283_n 0.00399188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_223_47#_c_275_n 0.00168007f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_223_47#_c_276_n 0.00224508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_223_47#_c_286_n 0.00184235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_223_47#_c_277_n 0.00112043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_223_47#_c_278_n 0.00491745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_C_M1004_g 0.050576f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=2.275
cc_69 VPB C 8.41709e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB C 0.005924f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.74
cc_71 VPB N_C_c_374_n 0.00459387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_D_M1003_g 0.0551466f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=2.275
cc_73 VPB D 2.76307e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB D 0.00335703f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.74
cc_75 VPB N_D_c_420_n 0.0047381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_343_93#_M1013_g 0.0228013f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.875
cc_77 VPB N_A_343_93#_c_463_n 0.00557738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_343_93#_c_469_n 0.011417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_343_93#_c_470_n 0.0073307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_343_93#_c_464_n 0.00136695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_343_93#_c_465_n 0.0171282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_343_93#_c_473_n 0.00273854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_343_93#_c_474_n 0.00639189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_554_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_555_n 0.00765163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_556_n 0.00285986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_557_n 0.00281836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_558_n 0.0176408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_559_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_560_n 0.0144076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_561_n 0.00518085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_562_n 0.0225035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_563_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_553_n 0.0465904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_565_n 0.0238568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_566_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_X_c_630_n 0.0450095f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.87
cc_98 N_A_N_M1007_g N_B_N_M1009_g 0.0199063f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_N_M1007_g N_B_N_M1012_g 0.0204873f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_N_M1006_g N_B_N_M1012_g 0.0179558f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_101 N_A_N_c_101_n N_B_N_M1012_g 0.0161134f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_102 N_A_N_c_102_n N_B_N_M1012_g 0.00497199f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_103 N_A_N_M1007_g N_B_N_c_136_n 0.0174541f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_N_M1007_g B_N 0.0115479f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_N_M1007_g N_A_27_47#_c_184_n 0.0170868f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_N_M1007_g N_A_27_47#_c_193_n 0.00453467f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_N_M1006_g N_A_27_47#_c_193_n 0.00590661f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_108 N_A_N_c_101_n N_A_27_47#_c_193_n 0.00635646f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_109 N_A_N_c_102_n N_A_27_47#_c_193_n 0.0252461f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_110 N_A_N_M1007_g N_A_27_47#_c_185_n 0.014302f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_N_c_101_n N_A_27_47#_c_185_n 0.00397826f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_112 N_A_N_c_102_n N_A_27_47#_c_185_n 0.0258004f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_113 N_A_N_M1007_g N_A_27_47#_c_186_n 0.00850046f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_N_M1006_g N_A_27_47#_c_197_n 0.00850046f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_115 N_A_N_M1007_g N_A_27_47#_c_188_n 8.94388e-19 $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_N_c_101_n N_A_27_47#_c_188_n 2.50711e-19 $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_117 N_A_N_c_102_n N_A_27_47#_c_188_n 0.00646019f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_118 N_A_N_c_102_n N_A_223_47#_c_283_n 0.00179773f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_119 N_A_N_M1006_g N_VPWR_c_554_n 0.00929121f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_120 N_A_N_c_101_n N_VPWR_c_554_n 2.43281e-19 $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_121 N_A_N_c_102_n N_VPWR_c_554_n 0.00418254f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_122 N_A_N_M1006_g N_VPWR_c_553_n 0.00534909f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_123 N_A_N_c_102_n N_VPWR_c_553_n 0.00864222f $X=0.59 $Y=1.74 $X2=0 $Y2=0
cc_124 N_A_N_M1006_g N_VPWR_c_565_n 0.0046653f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_125 N_A_N_M1007_g N_VGND_c_642_n 0.00929121f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_N_M1007_g N_VGND_c_646_n 0.00753396f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_127 N_A_N_M1007_g N_VGND_c_647_n 0.0046653f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_128 N_B_N_c_136_n N_A_27_47#_c_181_n 0.00283603f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_129 N_B_N_M1012_g N_A_27_47#_c_182_n 0.00364862f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_130 N_B_N_M1012_g N_A_27_47#_c_191_n 0.0218357f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_131 B_N N_A_27_47#_c_184_n 0.0148521f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_132 N_B_N_M1012_g N_A_27_47#_c_185_n 0.00838864f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_133 N_B_N_c_135_n N_A_27_47#_c_185_n 0.0164529f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_134 N_B_N_c_136_n N_A_27_47#_c_185_n 0.0015978f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_135 B_N N_A_27_47#_c_185_n 0.0160213f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_136 N_B_N_c_135_n N_A_27_47#_c_195_n 3.40116e-19 $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_137 N_B_N_M1012_g N_A_27_47#_c_188_n 0.0150352f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_138 N_B_N_c_135_n N_A_27_47#_c_188_n 0.0128119f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_139 N_B_N_c_136_n N_A_27_47#_c_188_n 0.00232299f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_140 N_B_N_M1012_g N_A_223_47#_c_290_n 0.00429957f $X=1.04 $Y=2.275 $X2=0
+ $Y2=0
cc_141 N_B_N_M1009_g N_A_223_47#_c_273_n 0.0029049f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_142 N_B_N_M1012_g N_A_223_47#_c_273_n 0.00145594f $X=1.04 $Y=2.275 $X2=0
+ $Y2=0
cc_143 N_B_N_c_135_n N_A_223_47#_c_273_n 0.0129015f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_144 N_B_N_c_136_n N_A_223_47#_c_273_n 0.00334594f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_145 B_N N_A_223_47#_c_273_n 0.00587766f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_146 N_B_N_M1012_g N_A_223_47#_c_283_n 0.00675059f $X=1.04 $Y=2.275 $X2=0
+ $Y2=0
cc_147 N_B_N_M1012_g N_A_223_47#_c_276_n 0.00176506f $X=1.04 $Y=2.275 $X2=0
+ $Y2=0
cc_148 N_B_N_M1012_g N_A_223_47#_c_286_n 0.00219804f $X=1.04 $Y=2.275 $X2=0
+ $Y2=0
cc_149 N_B_N_M1009_g N_A_223_47#_c_279_n 0.0120126f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_150 N_B_N_c_135_n N_A_223_47#_c_279_n 0.00426445f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_151 N_B_N_c_136_n N_A_223_47#_c_279_n 0.00137363f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_152 N_B_N_M1012_g N_VPWR_c_554_n 0.00881093f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_153 N_B_N_M1012_g N_VPWR_c_555_n 0.00250714f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_154 N_B_N_M1012_g N_VPWR_c_558_n 0.00505556f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_155 N_B_N_M1012_g N_VPWR_c_553_n 0.00983214f $X=1.04 $Y=2.275 $X2=0 $Y2=0
cc_156 N_B_N_M1009_g N_VGND_c_642_n 0.00802059f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_157 N_B_N_c_135_n N_VGND_c_642_n 0.00495747f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_158 N_B_N_c_136_n N_VGND_c_642_n 0.0010875f $X=1.06 $Y=1.03 $X2=0 $Y2=0
cc_159 B_N N_VGND_c_642_n 0.00625365f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_160 N_B_N_M1009_g N_VGND_c_644_n 0.00505556f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_161 N_B_N_M1009_g N_VGND_c_646_n 0.00995901f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_162 B_N N_VGND_c_646_n 0.00236747f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_192_n N_A_223_47#_M1002_g 0.0305118f $X=1.965 $Y=1.66 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1008_g N_A_223_47#_c_290_n 0.00294634f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_181_n N_A_223_47#_c_273_n 0.00329188f $X=1.965 $Y=1.155
+ $X2=0 $Y2=0
cc_166 N_A_27_47#_c_183_n N_A_223_47#_c_273_n 8.53847e-19 $X=1.965 $Y=0.975
+ $X2=0 $Y2=0
cc_167 N_A_27_47#_M1008_g N_A_223_47#_c_282_n 0.00395448f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_191_n N_A_223_47#_c_282_n 0.0100768f $X=1.785 $Y=1.66 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_195_n N_A_223_47#_c_282_n 0.0149809f $X=1.46 $Y=1.66 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_191_n N_A_223_47#_c_283_n 0.00229181f $X=1.785 $Y=1.66 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_195_n N_A_223_47#_c_283_n 0.0154314f $X=1.46 $Y=1.66 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_183_n N_A_223_47#_c_274_n 0.0113457f $X=1.965 $Y=0.975 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_182_n N_A_223_47#_c_275_n 0.0110563f $X=1.965 $Y=1.495 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_191_n N_A_223_47#_c_275_n 0.0060558f $X=1.785 $Y=1.66 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_195_n N_A_223_47#_c_275_n 0.00425338f $X=1.46 $Y=1.66 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_191_n N_A_223_47#_c_276_n 0.0043649f $X=1.785 $Y=1.66 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_195_n N_A_223_47#_c_276_n 0.0137147f $X=1.46 $Y=1.66 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_188_n N_A_223_47#_c_276_n 0.00959073f $X=1.13 $Y=1.37 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_182_n N_A_223_47#_c_286_n 0.00379184f $X=1.965 $Y=1.495
+ $X2=0 $Y2=0
cc_180 N_A_27_47#_M1008_g N_A_223_47#_c_286_n 0.0020133f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_192_n N_A_223_47#_c_286_n 0.0184626f $X=1.965 $Y=1.66 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_195_n N_A_223_47#_c_286_n 0.012273f $X=1.46 $Y=1.66 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_188_n N_A_223_47#_c_286_n 0.00483681f $X=1.13 $Y=1.37 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_183_n N_A_223_47#_c_277_n 0.00162973f $X=1.965 $Y=0.975
+ $X2=0 $Y2=0
cc_185 N_A_27_47#_c_181_n N_A_223_47#_c_278_n 0.0305118f $X=1.965 $Y=1.155 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_183_n N_A_223_47#_c_279_n 0.00565593f $X=1.965 $Y=0.975
+ $X2=0 $Y2=0
cc_187 N_A_27_47#_c_183_n N_A_223_47#_c_280_n 0.0305118f $X=1.965 $Y=0.975 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_181_n N_A_343_93#_c_462_n 0.00747878f $X=1.965 $Y=1.155
+ $X2=0 $Y2=0
cc_189 N_A_27_47#_c_183_n N_A_343_93#_c_462_n 0.0165287f $X=1.965 $Y=0.975 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_181_n N_A_343_93#_c_463_n 0.00554823f $X=1.965 $Y=1.155
+ $X2=0 $Y2=0
cc_191 N_A_27_47#_c_182_n N_A_343_93#_c_463_n 0.00814416f $X=1.965 $Y=1.495
+ $X2=0 $Y2=0
cc_192 N_A_27_47#_M1008_g N_A_343_93#_c_463_n 0.00152683f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_183_n N_A_343_93#_c_463_n 0.00129648f $X=1.965 $Y=0.975
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_c_192_n N_A_343_93#_c_463_n 0.00731784f $X=1.965 $Y=1.66 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1008_g N_A_343_93#_c_482_n 0.00408662f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1008_g N_A_343_93#_c_473_n 0.0038429f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_197_n N_VPWR_c_554_n 0.0100793f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_198 N_A_27_47#_M1008_g N_VPWR_c_555_n 0.0034507f $X=2.07 $Y=2.275 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_192_n N_VPWR_c_555_n 9.22729e-19 $X=1.965 $Y=1.66 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_M1008_g N_VPWR_c_556_n 5.04416e-19 $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_M1008_g N_VPWR_c_560_n 0.00572911f $X=2.07 $Y=2.275 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_M1006_s N_VPWR_c_553_n 0.00662376f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1008_g N_VPWR_c_553_n 0.0114771f $X=2.07 $Y=2.275 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_197_n N_VPWR_c_553_n 0.00982816f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_197_n N_VPWR_c_565_n 0.0173041f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_186_n N_VGND_c_642_n 0.0100793f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_183_n N_VGND_c_644_n 0.00357877f $X=1.965 $Y=0.975 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_M1007_s N_VGND_c_646_n 0.00984512f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_183_n N_VGND_c_646_n 0.00669482f $X=1.965 $Y=0.975 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_186_n N_VGND_c_646_n 0.00982816f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_186_n N_VGND_c_647_n 0.0173041f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_212 N_A_223_47#_M1002_g N_C_M1004_g 0.0324496f $X=2.5 $Y=2.275 $X2=0 $Y2=0
cc_213 N_A_223_47#_c_274_n C 6.48139e-19 $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_214 N_A_223_47#_c_277_n C 0.0382002f $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_223_47#_c_280_n C 7.86361e-19 $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_223_47#_c_278_n C 0.00195547f $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_223_47#_M1002_g C 0.00250344f $X=2.5 $Y=2.275 $X2=0 $Y2=0
cc_218 N_A_223_47#_c_277_n N_C_c_374_n 3.83742e-19 $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_223_47#_c_278_n N_C_c_374_n 0.0204055f $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_223_47#_c_274_n N_C_c_375_n 0.00401384f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_221 N_A_223_47#_c_277_n N_C_c_375_n 0.00189153f $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_223_47#_c_280_n N_C_c_375_n 0.0302321f $X=2.56 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_223_47#_c_274_n N_A_343_93#_c_462_n 0.035698f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_224 N_A_223_47#_c_275_n N_A_343_93#_c_462_n 0.0111143f $X=1.795 $Y=1.32 $X2=0
+ $Y2=0
cc_225 N_A_223_47#_c_277_n N_A_343_93#_c_462_n 0.025658f $X=2.56 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_223_47#_c_279_n N_A_343_93#_c_462_n 0.0253926f $X=1.365 $Y=0.34 $X2=0
+ $Y2=0
cc_227 N_A_223_47#_c_280_n N_A_343_93#_c_462_n 0.00226568f $X=2.56 $Y=0.995
+ $X2=0 $Y2=0
cc_228 N_A_223_47#_c_273_n N_A_343_93#_c_463_n 0.00882702f $X=1.48 $Y=1.235
+ $X2=0 $Y2=0
cc_229 N_A_223_47#_c_275_n N_A_343_93#_c_463_n 0.0127601f $X=1.795 $Y=1.32 $X2=0
+ $Y2=0
cc_230 N_A_223_47#_c_286_n N_A_343_93#_c_463_n 0.0346969f $X=1.88 $Y=1.915 $X2=0
+ $Y2=0
cc_231 N_A_223_47#_c_277_n N_A_343_93#_c_463_n 0.0285363f $X=2.56 $Y=1.16 $X2=0
+ $Y2=0
cc_232 N_A_223_47#_c_280_n N_A_343_93#_c_463_n 0.0120897f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_223_47#_M1002_g N_A_343_93#_c_469_n 0.0149218f $X=2.5 $Y=2.275 $X2=0
+ $Y2=0
cc_234 N_A_223_47#_c_277_n N_A_343_93#_c_469_n 0.00482177f $X=2.56 $Y=1.16 $X2=0
+ $Y2=0
cc_235 N_A_223_47#_c_278_n N_A_343_93#_c_469_n 0.00159061f $X=2.56 $Y=1.16 $X2=0
+ $Y2=0
cc_236 N_A_223_47#_c_282_n N_A_343_93#_c_473_n 0.0141708f $X=1.795 $Y=2 $X2=0
+ $Y2=0
cc_237 N_A_223_47#_c_282_n N_VPWR_M1008_s 0.00268439f $X=1.795 $Y=2 $X2=0 $Y2=0
cc_238 N_A_223_47#_c_290_n N_VPWR_c_554_n 0.0119937f $X=1.31 $Y=2.3 $X2=0 $Y2=0
cc_239 N_A_223_47#_c_290_n N_VPWR_c_555_n 0.0125193f $X=1.31 $Y=2.3 $X2=0 $Y2=0
cc_240 N_A_223_47#_c_282_n N_VPWR_c_555_n 0.0219734f $X=1.795 $Y=2 $X2=0 $Y2=0
cc_241 N_A_223_47#_M1002_g N_VPWR_c_556_n 0.00545865f $X=2.5 $Y=2.275 $X2=0
+ $Y2=0
cc_242 N_A_223_47#_c_290_n N_VPWR_c_558_n 0.0130174f $X=1.31 $Y=2.3 $X2=0 $Y2=0
cc_243 N_A_223_47#_c_282_n N_VPWR_c_558_n 0.00453603f $X=1.795 $Y=2 $X2=0 $Y2=0
cc_244 N_A_223_47#_M1002_g N_VPWR_c_560_n 0.00410216f $X=2.5 $Y=2.275 $X2=0
+ $Y2=0
cc_245 N_A_223_47#_M1012_d N_VPWR_c_553_n 0.00646873f $X=1.115 $Y=2.065 $X2=0
+ $Y2=0
cc_246 N_A_223_47#_M1002_g N_VPWR_c_553_n 0.00470902f $X=2.5 $Y=2.275 $X2=0
+ $Y2=0
cc_247 N_A_223_47#_c_290_n N_VPWR_c_553_n 0.00720049f $X=1.31 $Y=2.3 $X2=0 $Y2=0
cc_248 N_A_223_47#_c_282_n N_VPWR_c_553_n 0.00854597f $X=1.795 $Y=2 $X2=0 $Y2=0
cc_249 N_A_223_47#_c_274_n N_VGND_c_644_n 0.0698554f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_250 N_A_223_47#_c_279_n N_VGND_c_644_n 0.0275958f $X=1.365 $Y=0.34 $X2=0
+ $Y2=0
cc_251 N_A_223_47#_c_280_n N_VGND_c_644_n 0.00357738f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_223_47#_M1009_d N_VGND_c_646_n 0.00444558f $X=1.115 $Y=0.235 $X2=0
+ $Y2=0
cc_253 N_A_223_47#_c_274_n N_VGND_c_646_n 0.0390701f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_254 N_A_223_47#_c_279_n N_VGND_c_646_n 0.0152582f $X=1.365 $Y=0.34 $X2=0
+ $Y2=0
cc_255 N_A_223_47#_c_280_n N_VGND_c_646_n 0.00553714f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_A_223_47#_c_277_n A_515_93# 0.00427981f $X=2.56 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_257 C N_D_c_417_n 7.7368e-19 $X=2.9 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_258 N_C_c_375_n N_D_c_417_n 0.0291435f $X=3.04 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_259 N_C_M1004_g N_D_M1003_g 0.0357201f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_260 C N_D_M1003_g 9.31547e-19 $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_261 C D 0.019566f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_262 N_C_c_375_n D 0.00210817f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_263 C D 0.0202173f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_264 N_C_c_374_n D 0.00197826f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_265 N_C_M1004_g D 0.00113488f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_266 C D 0.0171476f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_267 C N_D_c_420_n 3.63217e-19 $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_268 N_C_c_374_n N_D_c_420_n 0.0203259f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_269 C N_A_343_93#_c_463_n 0.00978322f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_270 N_C_M1004_g N_A_343_93#_c_469_n 0.0132612f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_271 C N_A_343_93#_c_469_n 0.00129035f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_272 C N_A_343_93#_c_469_n 0.00962195f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_273 N_C_c_374_n N_A_343_93#_c_469_n 0.00117241f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_274 N_C_M1004_g N_A_343_93#_c_503_n 0.00411901f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_275 N_C_c_374_n N_A_343_93#_c_474_n 4.17784e-19 $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_276 N_C_M1004_g N_VPWR_c_556_n 0.00314432f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_277 N_C_M1004_g N_VPWR_c_562_n 0.00425094f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_278 N_C_M1004_g N_VPWR_c_553_n 0.00607026f $X=3 $Y=2.275 $X2=0 $Y2=0
cc_279 C N_VGND_c_644_n 0.00606925f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_280 N_C_c_375_n N_VGND_c_644_n 0.00388886f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_281 C N_VGND_c_646_n 0.00568835f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_282 N_C_c_375_n N_VGND_c_646_n 0.00589495f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_283 N_D_M1003_g N_A_343_93#_M1013_g 0.0240974f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_284 D N_A_343_93#_M1013_g 3.06136e-19 $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_285 N_D_M1003_g N_A_343_93#_c_503_n 0.00606986f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_286 N_D_M1003_g N_A_343_93#_c_470_n 0.0141729f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_287 D N_A_343_93#_c_470_n 0.00154436f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_288 D N_A_343_93#_c_470_n 0.0106564f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_289 N_D_c_420_n N_A_343_93#_c_470_n 0.00149935f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_290 N_D_M1003_g N_A_343_93#_c_464_n 0.00744911f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_291 D N_A_343_93#_c_464_n 0.0142753f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_292 D N_A_343_93#_c_464_n 0.0123147f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_293 N_D_c_420_n N_A_343_93#_c_464_n 0.0010689f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_294 D N_A_343_93#_c_465_n 0.00123839f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_295 N_D_c_420_n N_A_343_93#_c_465_n 0.0212063f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_296 N_D_c_417_n N_A_343_93#_c_466_n 0.0159661f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_297 D N_A_343_93#_c_466_n 0.00237991f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_298 N_D_M1003_g N_VPWR_c_557_n 0.00531701f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_299 N_D_M1003_g N_VPWR_c_562_n 0.00425094f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_300 N_D_M1003_g N_VPWR_c_553_n 0.006581f $X=3.52 $Y=2.275 $X2=0 $Y2=0
cc_301 N_D_c_417_n N_VGND_c_643_n 0.00753552f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_302 D N_VGND_c_643_n 0.00292986f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_303 N_D_c_417_n N_VGND_c_644_n 0.00456292f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_304 D N_VGND_c_644_n 0.00645623f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_305 N_D_c_417_n N_VGND_c_646_n 0.00795744f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_306 D N_VGND_c_646_n 0.00626842f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_307 D A_615_93# 0.00443277f $X=3.36 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_308 N_A_343_93#_c_469_n N_VPWR_M1002_d 0.00241353f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_309 N_A_343_93#_c_470_n N_VPWR_M1003_d 0.00853586f $X=3.915 $Y=2 $X2=0 $Y2=0
cc_310 N_A_343_93#_c_464_n N_VPWR_M1003_d 0.0054989f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_343_93#_c_482_n N_VPWR_c_555_n 0.0140523f $X=2.29 $Y=2.3 $X2=0 $Y2=0
cc_312 N_A_343_93#_c_469_n N_VPWR_c_556_n 0.0182509f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_313 N_A_343_93#_M1013_g N_VPWR_c_557_n 0.00864708f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_343_93#_c_503_n N_VPWR_c_557_n 0.00815282f $X=3.245 $Y=2.3 $X2=0
+ $Y2=0
cc_315 N_A_343_93#_c_470_n N_VPWR_c_557_n 0.0213052f $X=3.915 $Y=2 $X2=0 $Y2=0
cc_316 N_A_343_93#_c_482_n N_VPWR_c_560_n 0.0115368f $X=2.29 $Y=2.3 $X2=0 $Y2=0
cc_317 N_A_343_93#_c_469_n N_VPWR_c_560_n 0.00285218f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_318 N_A_343_93#_c_473_n N_VPWR_c_560_n 7.88667e-19 $X=2.255 $Y=2 $X2=0 $Y2=0
cc_319 N_A_343_93#_c_469_n N_VPWR_c_562_n 0.00372949f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_320 N_A_343_93#_c_503_n N_VPWR_c_562_n 0.0116326f $X=3.245 $Y=2.3 $X2=0 $Y2=0
cc_321 N_A_343_93#_c_470_n N_VPWR_c_562_n 0.00637056f $X=3.915 $Y=2 $X2=0 $Y2=0
cc_322 N_A_343_93#_M1013_g N_VPWR_c_563_n 0.0046653f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_343_93#_M1008_d N_VPWR_c_553_n 0.00260941f $X=2.145 $Y=2.065 $X2=0
+ $Y2=0
cc_324 N_A_343_93#_M1004_d N_VPWR_c_553_n 0.00367297f $X=3.075 $Y=2.065 $X2=0
+ $Y2=0
cc_325 N_A_343_93#_M1013_g N_VPWR_c_553_n 0.008846f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_343_93#_c_482_n N_VPWR_c_553_n 0.0064554f $X=2.29 $Y=2.3 $X2=0 $Y2=0
cc_327 N_A_343_93#_c_469_n N_VPWR_c_553_n 0.0127664f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_328 N_A_343_93#_c_503_n N_VPWR_c_553_n 0.00643448f $X=3.245 $Y=2.3 $X2=0
+ $Y2=0
cc_329 N_A_343_93#_c_470_n N_VPWR_c_553_n 0.0128685f $X=3.915 $Y=2 $X2=0 $Y2=0
cc_330 N_A_343_93#_c_473_n N_VPWR_c_553_n 0.00200712f $X=2.255 $Y=2 $X2=0 $Y2=0
cc_331 N_A_343_93#_M1013_g N_X_c_630_n 0.0089479f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_343_93#_c_464_n N_X_c_630_n 0.0494302f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_343_93#_c_465_n N_X_c_630_n 0.0279795f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_343_93#_c_466_n N_X_c_630_n 0.00967574f $X=4.177 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_343_93#_c_464_n N_VGND_c_643_n 0.00476568f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_343_93#_c_465_n N_VGND_c_643_n 0.00214632f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_343_93#_c_466_n N_VGND_c_643_n 0.00899988f $X=4.177 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_343_93#_c_466_n N_VGND_c_645_n 0.0046653f $X=4.177 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_A_343_93#_c_466_n N_VGND_c_646_n 0.008846f $X=4.177 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_A_343_93#_c_462_n A_429_93# 0.00355432f $X=2.135 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_341 N_VPWR_c_553_n N_X_M1013_d 0.00382897f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_342 N_VPWR_c_563_n N_X_c_630_n 0.018001f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_343 N_VPWR_c_553_n N_X_c_630_n 0.00993603f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_344 N_X_c_630_n N_VGND_c_645_n 0.0180148f $X=4.34 $Y=0.42 $X2=0 $Y2=0
cc_345 N_X_M1005_d N_VGND_c_646_n 0.00374699f $X=4.205 $Y=0.235 $X2=0 $Y2=0
cc_346 N_X_c_630_n N_VGND_c_646_n 0.00993603f $X=4.34 $Y=0.42 $X2=0 $Y2=0

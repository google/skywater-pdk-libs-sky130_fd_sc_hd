* File: sky130_fd_sc_hd__and4_1.spice
* Created: Tue Sep  1 18:58:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4_1.pex.spice"
.subckt sky130_fd_sc_hd__and4_1  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1008 A_109_47# N_A_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.1092 PD=0.71 PS=1.36 NRD=25.704 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1003 A_197_47# N_B_M1003_g A_109_47# VNB NSHORT L=0.15 W=0.42 AD=0.0798
+ AS=0.0609 PD=0.8 PS=0.71 NRD=38.568 NRS=25.704 M=1 R=2.8 SA=75000.6 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1001 A_303_47# N_C_M1001_g A_197_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0798 PD=0.75 PS=0.8 NRD=31.428 NRS=38.568 M=1 R=2.8 SA=75001.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_D_M1006_g A_303_47# VNB NSHORT L=0.15 W=0.42 AD=0.154085
+ AS=0.0693 PD=1.04411 PS=0.75 NRD=94.992 NRS=31.428 M=1 R=2.8 SA=75001.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_27_47#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.238465 PD=1.82 PS=1.61589 NRD=0 NRS=12.912 M=1 R=4.33333
+ SA=75001.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1092 PD=0.77 PS=1.36 NRD=16.4101 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_27_47#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0777 AS=0.0735 PD=0.79 PS=0.77 NRD=21.0987 NRS=16.4101 M=1 R=2.8
+ SA=75000.7 SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_A_27_47#_M1000_d N_C_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0777 PD=0.7 PS=0.79 NRD=0 NRS=21.0987 M=1 R=2.8 SA=75001.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_D_M1007_g N_A_27_47#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.18483 AS=0.0588 PD=0.993803 PS=0.7 NRD=153.601 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_27_47#_M1009_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.44007 PD=2.52 PS=2.3662 NRD=0 NRS=14.7553 M=1 R=6.66667
+ SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_59 VPB 0 1.22265e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__and4_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__xnor2_4.pxi.spice
* Created: Tue Sep  1 19:32:55 2020
* 
x_PM_SKY130_FD_SC_HD__XNOR2_4%B N_B_c_153_n N_B_M1025_g N_B_M1007_g N_B_c_154_n
+ N_B_M1027_g N_B_M1018_g N_B_c_155_n N_B_M1035_g N_B_M1020_g N_B_c_156_n
+ N_B_M1038_g N_B_M1028_g N_B_c_157_n N_B_M1002_g N_B_M1000_g N_B_c_158_n
+ N_B_M1006_g N_B_M1001_g N_B_c_159_n N_B_M1015_g N_B_M1013_g N_B_c_160_n
+ N_B_M1034_g N_B_M1017_g N_B_c_172_n N_B_c_173_n N_B_c_174_n N_B_c_175_n
+ N_B_c_197_p N_B_c_161_n N_B_c_194_p B N_B_c_162_n N_B_c_163_n
+ PM_SKY130_FD_SC_HD__XNOR2_4%B
x_PM_SKY130_FD_SC_HD__XNOR2_4%A N_A_c_356_n N_A_M1003_g N_A_M1005_g N_A_c_357_n
+ N_A_M1030_g N_A_M1011_g N_A_c_358_n N_A_M1032_g N_A_M1016_g N_A_c_359_n
+ N_A_M1036_g N_A_M1021_g N_A_c_360_n N_A_M1004_g N_A_M1008_g N_A_c_361_n
+ N_A_M1009_g N_A_M1012_g N_A_c_362_n N_A_M1033_g N_A_M1022_g N_A_c_363_n
+ N_A_M1039_g N_A_M1026_g A N_A_c_364_n N_A_c_365_n N_A_c_366_n
+ PM_SKY130_FD_SC_HD__XNOR2_4%A
x_PM_SKY130_FD_SC_HD__XNOR2_4%A_38_297# N_A_38_297#_M1025_d N_A_38_297#_M1035_d
+ N_A_38_297#_M1007_s N_A_38_297#_M1018_s N_A_38_297#_M1028_s
+ N_A_38_297#_M1011_d N_A_38_297#_M1021_d N_A_38_297#_c_508_n
+ N_A_38_297#_M1019_g N_A_38_297#_M1010_g N_A_38_297#_c_509_n
+ N_A_38_297#_M1023_g N_A_38_297#_M1014_g N_A_38_297#_c_510_n
+ N_A_38_297#_M1024_g N_A_38_297#_M1029_g N_A_38_297#_c_511_n
+ N_A_38_297#_M1031_g N_A_38_297#_M1037_g N_A_38_297#_c_512_n
+ N_A_38_297#_c_524_n N_A_38_297#_c_513_n N_A_38_297#_c_514_n
+ N_A_38_297#_c_525_n N_A_38_297#_c_526_n N_A_38_297#_c_554_n
+ N_A_38_297#_c_560_n N_A_38_297#_c_561_n N_A_38_297#_c_515_n
+ N_A_38_297#_c_516_n N_A_38_297#_c_517_n N_A_38_297#_c_528_n
+ N_A_38_297#_c_625_p N_A_38_297#_c_565_n N_A_38_297#_c_566_n
+ N_A_38_297#_c_529_n N_A_38_297#_c_530_n N_A_38_297#_c_531_n
+ N_A_38_297#_c_532_n N_A_38_297#_c_533_n N_A_38_297#_c_518_n
+ PM_SKY130_FD_SC_HD__XNOR2_4%A_38_297#
x_PM_SKY130_FD_SC_HD__XNOR2_4%VPWR N_VPWR_M1007_d N_VPWR_M1020_d N_VPWR_M1005_s
+ N_VPWR_M1016_s N_VPWR_M1008_s N_VPWR_M1022_s N_VPWR_M1010_s N_VPWR_M1029_s
+ N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n
+ N_VPWR_c_726_n N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n
+ N_VPWR_c_731_n N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n
+ N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_738_n VPWR N_VPWR_c_739_n
+ N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_720_n N_VPWR_c_743_n N_VPWR_c_744_n
+ N_VPWR_c_745_n PM_SKY130_FD_SC_HD__XNOR2_4%VPWR
x_PM_SKY130_FD_SC_HD__XNOR2_4%A_820_297# N_A_820_297#_M1008_d
+ N_A_820_297#_M1012_d N_A_820_297#_M1026_d N_A_820_297#_M1001_s
+ N_A_820_297#_M1017_s N_A_820_297#_c_883_n N_A_820_297#_c_884_n
+ N_A_820_297#_c_886_n N_A_820_297#_c_926_n N_A_820_297#_c_879_n
+ N_A_820_297#_c_880_n N_A_820_297#_c_892_n
+ PM_SKY130_FD_SC_HD__XNOR2_4%A_820_297#
x_PM_SKY130_FD_SC_HD__XNOR2_4%Y N_Y_M1019_d N_Y_M1024_d N_Y_M1000_d N_Y_M1013_d
+ N_Y_M1010_d N_Y_M1014_d N_Y_M1037_d N_Y_c_942_n N_Y_c_943_n N_Y_c_944_n
+ N_Y_c_940_n N_Y_c_994_n N_Y_c_945_n N_Y_c_941_n N_Y_c_947_n N_Y_c_948_n
+ N_Y_c_949_n Y PM_SKY130_FD_SC_HD__XNOR2_4%Y
x_PM_SKY130_FD_SC_HD__XNOR2_4%A_38_47# N_A_38_47#_M1025_s N_A_38_47#_M1027_s
+ N_A_38_47#_M1038_s N_A_38_47#_M1030_d N_A_38_47#_M1036_d N_A_38_47#_c_1016_n
+ N_A_38_47#_c_1028_n N_A_38_47#_c_1017_n N_A_38_47#_c_1018_n
+ N_A_38_47#_c_1036_n N_A_38_47#_c_1019_n N_A_38_47#_c_1020_n
+ N_A_38_47#_c_1021_n PM_SKY130_FD_SC_HD__XNOR2_4%A_38_47#
x_PM_SKY130_FD_SC_HD__XNOR2_4%VGND N_VGND_M1003_s N_VGND_M1032_s N_VGND_M1004_d
+ N_VGND_M1009_d N_VGND_M1039_d N_VGND_M1006_d N_VGND_M1034_d N_VGND_c_1084_n
+ N_VGND_c_1085_n N_VGND_c_1086_n N_VGND_c_1087_n N_VGND_c_1088_n
+ N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n N_VGND_c_1092_n
+ N_VGND_c_1093_n N_VGND_c_1094_n N_VGND_c_1095_n N_VGND_c_1096_n
+ N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n N_VGND_c_1100_n
+ N_VGND_c_1101_n VGND N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n
+ N_VGND_c_1105_n N_VGND_c_1106_n PM_SKY130_FD_SC_HD__XNOR2_4%VGND
x_PM_SKY130_FD_SC_HD__XNOR2_4%A_902_47# N_A_902_47#_M1004_s N_A_902_47#_M1033_s
+ N_A_902_47#_M1002_s N_A_902_47#_M1015_s N_A_902_47#_M1019_s
+ N_A_902_47#_M1023_s N_A_902_47#_M1031_s N_A_902_47#_c_1276_n
+ N_A_902_47#_c_1239_n N_A_902_47#_c_1240_n N_A_902_47#_c_1250_n
+ N_A_902_47#_c_1241_n N_A_902_47#_c_1254_n N_A_902_47#_c_1242_n
+ N_A_902_47#_c_1261_n N_A_902_47#_c_1243_n N_A_902_47#_c_1244_n
+ N_A_902_47#_c_1245_n N_A_902_47#_c_1246_n N_A_902_47#_c_1247_n
+ N_A_902_47#_c_1248_n N_A_902_47#_c_1249_n
+ PM_SKY130_FD_SC_HD__XNOR2_4%A_902_47#
cc_1 VNB N_B_c_153_n 0.0192188f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_2 VNB N_B_c_154_n 0.0157855f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.995
cc_3 VNB N_B_c_155_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=0.995
cc_4 VNB N_B_c_156_n 0.0161471f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.995
cc_5 VNB N_B_c_157_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=0.995
cc_6 VNB N_B_c_158_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=0.995
cc_7 VNB N_B_c_159_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=0.995
cc_8 VNB N_B_c_160_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=0.995
cc_9 VNB N_B_c_161_n 0.00499013f $X=-0.19 $Y=-0.24 $X2=7.26 $Y2=1.16
cc_10 VNB N_B_c_162_n 0.0667627f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_11 VNB N_B_c_163_n 0.0677764f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=1.16
cc_12 VNB N_A_c_356_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_13 VNB N_A_c_357_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=0.995
cc_14 VNB N_A_c_358_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=0.995
cc_15 VNB N_A_c_359_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.995
cc_16 VNB N_A_c_360_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=0.995
cc_17 VNB N_A_c_361_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=0.995
cc_18 VNB N_A_c_362_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=0.995
cc_19 VNB N_A_c_363_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=0.995
cc_20 VNB N_A_c_364_n 0.0705732f $X=-0.19 $Y=-0.24 $X2=7.26 $Y2=1.16
cc_21 VNB N_A_c_365_n 0.0224696f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_22 VNB N_A_c_366_n 0.0692681f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=1.16
cc_23 VNB N_A_38_297#_c_508_n 0.0213688f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.995
cc_24 VNB N_A_38_297#_c_509_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=0.995
cc_25 VNB N_A_38_297#_c_510_n 0.0157854f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=0.995
cc_26 VNB N_A_38_297#_c_511_n 0.0192138f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=0.995
cc_27 VNB N_A_38_297#_c_512_n 0.0205747f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=0.56
cc_28 VNB N_A_38_297#_c_513_n 0.0129845f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.445
cc_29 VNB N_A_38_297#_c_514_n 0.00828076f $X=-0.19 $Y=-0.24 $X2=5.645 $Y2=1.445
cc_30 VNB N_A_38_297#_c_515_n 7.92547e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_38_297#_c_516_n 0.00395418f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=1.16
cc_32 VNB N_A_38_297#_c_517_n 0.0126159f $X=-0.19 $Y=-0.24 $X2=7.26 $Y2=1.16
cc_33 VNB N_A_38_297#_c_518_n 0.0717961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_720_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_940_n 0.021012f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=1.985
cc_36 VNB N_Y_c_941_n 0.0201724f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=1.985
cc_37 VNB N_A_38_47#_c_1016_n 0.00936711f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=0.56
cc_38 VNB N_A_38_47#_c_1017_n 0.00320487f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.56
cc_39 VNB N_A_38_47#_c_1018_n 0.00205567f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.56
cc_40 VNB N_A_38_47#_c_1019_n 0.00635542f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=0.56
cc_41 VNB N_A_38_47#_c_1020_n 0.00439026f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=1.985
cc_42 VNB N_A_38_47#_c_1021_n 0.00209731f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=1.985
cc_43 VNB N_VGND_c_1084_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.56
cc_44 VNB N_VGND_c_1085_n 0.0035943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_1086_n 0.0133337f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=1.325
cc_46 VNB N_VGND_c_1087_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=0.995
cc_47 VNB N_VGND_c_1088_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=1.985
cc_48 VNB N_VGND_c_1089_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1090_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=1.325
cc_50 VNB N_VGND_c_1091_n 0.0087688f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=0.995
cc_51 VNB N_VGND_c_1092_n 0.0564265f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=1.325
cc_52 VNB N_VGND_c_1093_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=1.985
cc_53 VNB N_VGND_c_1094_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1095_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.275
cc_55 VNB N_VGND_c_1096_n 0.0175644f $X=-0.19 $Y=-0.24 $X2=5.56 $Y2=1.53
cc_56 VNB N_VGND_c_1097_n 0.00528623f $X=-0.19 $Y=-0.24 $X2=1.855 $Y2=1.53
cc_57 VNB N_VGND_c_1098_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=5.645 $Y2=1.445
cc_58 VNB N_VGND_c_1099_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=5.73 $Y2=1.175
cc_59 VNB N_VGND_c_1100_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=6.24 $Y2=1.175
cc_60 VNB N_VGND_c_1101_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=6.24 $Y2=1.16
cc_61 VNB N_VGND_c_1102_n 0.0166727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1103_n 0.0588343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1104_n 0.477734f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=1.175
cc_64 VNB N_VGND_c_1105_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1106_n 0.00516249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_902_47#_c_1239_n 0.00205567f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.985
cc_67 VNB N_A_902_47#_c_1240_n 0.00209731f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.985
cc_68 VNB N_A_902_47#_c_1241_n 0.00234038f $X=-0.19 $Y=-0.24 $X2=6.115 $Y2=1.325
cc_69 VNB N_A_902_47#_c_1242_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=6.535 $Y2=0.56
cc_70 VNB N_A_902_47#_c_1243_n 0.0131996f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=0.56
cc_71 VNB N_A_902_47#_c_1244_n 0.00186471f $X=-0.19 $Y=-0.24 $X2=6.955 $Y2=1.325
cc_72 VNB N_A_902_47#_c_1245_n 0.00286122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_902_47#_c_1246_n 0.00730526f $X=-0.19 $Y=-0.24 $X2=7.375 $Y2=1.985
cc_74 VNB N_A_902_47#_c_1247_n 0.00274656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_902_47#_c_1248_n 0.00213756f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.275
cc_76 VNB N_A_902_47#_c_1249_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.445
cc_77 VPB N_B_M1007_g 0.022018f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.985
cc_78 VPB N_B_M1018_g 0.0179788f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_79 VPB N_B_M1020_g 0.0182751f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.985
cc_80 VPB N_B_M1028_g 0.0178886f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_81 VPB N_B_M1000_g 0.0182444f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=1.985
cc_82 VPB N_B_M1001_g 0.0181379f $X=-0.19 $Y=1.305 $X2=6.535 $Y2=1.985
cc_83 VPB N_B_M1013_g 0.0181184f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=1.985
cc_84 VPB N_B_M1017_g 0.022018f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=1.985
cc_85 VPB N_B_c_172_n 0.00101843f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.445
cc_86 VPB N_B_c_173_n 0.0356055f $X=-0.19 $Y=1.305 $X2=5.56 $Y2=1.53
cc_87 VPB N_B_c_174_n 2.62327e-19 $X=-0.19 $Y=1.305 $X2=1.855 $Y2=1.53
cc_88 VPB N_B_c_175_n 0.0011758f $X=-0.19 $Y=1.305 $X2=5.645 $Y2=1.445
cc_89 VPB N_B_c_162_n 0.0108204f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.16
cc_90 VPB N_B_c_163_n 0.0102625f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=1.16
cc_91 VPB N_A_M1005_g 0.0183686f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.985
cc_92 VPB N_A_M1011_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_93 VPB N_A_M1016_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.985
cc_94 VPB N_A_M1021_g 0.025044f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_95 VPB N_A_M1008_g 0.025044f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=1.985
cc_96 VPB N_A_M1012_g 0.0181194f $X=-0.19 $Y=1.305 $X2=6.535 $Y2=1.985
cc_97 VPB N_A_M1022_g 0.0180981f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=1.985
cc_98 VPB N_A_M1026_g 0.0179955f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=1.985
cc_99 VPB N_A_c_364_n 0.0108499f $X=-0.19 $Y=1.305 $X2=7.26 $Y2=1.16
cc_100 VPB N_A_c_366_n 0.0108529f $X=-0.19 $Y=1.305 $X2=1.675 $Y2=1.16
cc_101 VPB N_A_38_297#_M1010_g 0.0227299f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_102 VPB N_A_38_297#_M1014_g 0.018138f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=1.985
cc_103 VPB N_A_38_297#_M1029_g 0.0181184f $X=-0.19 $Y=1.305 $X2=6.535 $Y2=1.985
cc_104 VPB N_A_38_297#_M1037_g 0.0220113f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=1.985
cc_105 VPB N_A_38_297#_c_512_n 0.00738835f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=0.56
cc_106 VPB N_A_38_297#_c_524_n 0.0361631f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=1.985
cc_107 VPB N_A_38_297#_c_525_n 0.00233345f $X=-0.19 $Y=1.305 $X2=6.24 $Y2=1.175
cc_108 VPB N_A_38_297#_c_526_n 0.00125163f $X=-0.19 $Y=1.305 $X2=6.24 $Y2=1.16
cc_109 VPB N_A_38_297#_c_515_n 0.00379876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_38_297#_c_528_n 0.00958327f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.175
cc_111 VPB N_A_38_297#_c_529_n 0.00175452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_38_297#_c_530_n 0.0118681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_38_297#_c_531_n 0.00254455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_38_297#_c_532_n 0.00207063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_38_297#_c_533_n 0.0016129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_38_297#_c_518_n 0.0105282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_721_n 0.00454762f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=0.995
cc_118 VPB N_VPWR_c_722_n 0.00393015f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=1.985
cc_119 VPB N_VPWR_c_723_n 0.00393015f $X=-0.19 $Y=1.305 $X2=6.535 $Y2=0.56
cc_120 VPB N_VPWR_c_724_n 0.00454762f $X=-0.19 $Y=1.305 $X2=6.535 $Y2=1.985
cc_121 VPB N_VPWR_c_725_n 0.00454762f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=0.56
cc_122 VPB N_VPWR_c_726_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_727_n 0.00454762f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=1.325
cc_124 VPB N_VPWR_c_728_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.275
cc_125 VPB N_VPWR_c_729_n 0.0150723f $X=-0.19 $Y=1.305 $X2=1.855 $Y2=1.53
cc_126 VPB N_VPWR_c_730_n 0.00478085f $X=-0.19 $Y=1.305 $X2=5.645 $Y2=1.275
cc_127 VPB N_VPWR_c_731_n 0.0150723f $X=-0.19 $Y=1.305 $X2=5.73 $Y2=1.175
cc_128 VPB N_VPWR_c_732_n 0.00478085f $X=-0.19 $Y=1.305 $X2=6.24 $Y2=1.175
cc_129 VPB N_VPWR_c_733_n 0.0289933f $X=-0.19 $Y=1.305 $X2=6.24 $Y2=1.16
cc_130 VPB N_VPWR_c_734_n 0.00478085f $X=-0.19 $Y=1.305 $X2=7.26 $Y2=1.175
cc_131 VPB N_VPWR_c_735_n 0.0150723f $X=-0.19 $Y=1.305 $X2=7.26 $Y2=1.16
cc_132 VPB N_VPWR_c_736_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_737_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_134 VPB N_VPWR_c_738_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_739_n 0.0157253f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_136 VPB N_VPWR_c_740_n 0.0661083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_741_n 0.0182338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_720_n 0.0583141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_743_n 0.0234649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_744_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_745_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_820_297#_c_879_n 0.00297825f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=0.56
cc_143 VPB N_A_820_297#_c_880_n 0.00781334f $X=-0.19 $Y=1.305 $X2=6.115
+ $Y2=1.985
cc_144 VPB N_Y_c_942_n 0.00947509f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=0.995
cc_145 VPB N_Y_c_943_n 0.00470887f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=0.56
cc_146 VPB N_Y_c_944_n 0.00247713f $X=-0.19 $Y=1.305 $X2=6.115 $Y2=1.325
cc_147 VPB N_Y_c_945_n 0.00239552f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=0.56
cc_148 VPB N_Y_c_941_n 0.00723025f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=1.985
cc_149 VPB N_Y_c_947_n 0.00756442f $X=-0.19 $Y=1.305 $X2=6.955 $Y2=1.985
cc_150 VPB N_Y_c_948_n 0.00204415f $X=-0.19 $Y=1.305 $X2=7.375 $Y2=1.985
cc_151 VPB N_Y_c_949_n 0.011585f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.275
cc_152 VPB Y 0.0331391f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.445
cc_153 N_B_c_156_n N_A_c_356_n 0.0196735f $X=1.805 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_154 N_B_M1028_g N_A_M1005_g 0.0196735f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B_c_173_n N_A_M1005_g 0.010626f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B_c_173_n N_A_M1011_g 0.0103677f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B_c_173_n N_A_M1016_g 0.0103677f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_158 N_B_c_173_n N_A_M1021_g 0.0124706f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B_c_173_n N_A_M1008_g 0.0124706f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_160 N_B_c_173_n N_A_M1012_g 0.0103677f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_161 N_B_c_173_n N_A_M1022_g 0.0103677f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_162 N_B_c_175_n N_A_M1022_g 0.0023324f $X=5.645 $Y=1.445 $X2=0 $Y2=0
cc_163 N_B_c_157_n N_A_c_363_n 0.0240355f $X=6.115 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B_M1000_g N_A_M1026_g 0.0240355f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B_c_173_n N_A_M1026_g 0.0056919f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_166 N_B_c_175_n N_A_M1026_g 0.0031027f $X=5.645 $Y=1.445 $X2=0 $Y2=0
cc_167 N_B_c_172_n N_A_c_364_n 0.00106864f $X=1.77 $Y=1.445 $X2=0 $Y2=0
cc_168 N_B_c_173_n N_A_c_364_n 0.00642092f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_169 N_B_c_194_p N_A_c_364_n 8.71509e-19 $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_170 N_B_c_162_n N_A_c_364_n 0.0196735f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B_c_173_n N_A_c_365_n 0.210898f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_172 N_B_c_197_p N_A_c_365_n 0.0167609f $X=5.73 $Y=1.175 $X2=0 $Y2=0
cc_173 N_B_c_194_p N_A_c_365_n 0.0100567f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_174 N_B_c_162_n N_A_c_365_n 8.57456e-19 $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B_c_173_n N_A_c_366_n 0.00679673f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_176 N_B_c_175_n N_A_c_366_n 0.00359368f $X=5.645 $Y=1.445 $X2=0 $Y2=0
cc_177 N_B_c_197_p N_A_c_366_n 0.0084991f $X=5.73 $Y=1.175 $X2=0 $Y2=0
cc_178 N_B_c_161_n N_A_c_366_n 0.00445487f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_c_163_n N_A_c_366_n 0.0240355f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B_c_173_n N_A_38_297#_M1028_s 0.00165831f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_181 N_B_c_173_n N_A_38_297#_M1011_d 0.00165831f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_182 N_B_c_173_n N_A_38_297#_M1021_d 0.00272914f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_183 N_B_c_153_n N_A_38_297#_c_512_n 0.0187167f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_194_p N_A_38_297#_c_512_n 0.0162001f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_185 N_B_c_153_n N_A_38_297#_c_514_n 0.0136978f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B_c_154_n N_A_38_297#_c_514_n 0.01096f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_c_155_n N_A_38_297#_c_514_n 0.0109547f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B_c_156_n N_A_38_297#_c_514_n 0.00372402f $X=1.805 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B_c_194_p N_A_38_297#_c_514_n 0.0918942f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_190 N_B_c_162_n N_A_38_297#_c_514_n 0.00672641f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B_M1007_g N_A_38_297#_c_525_n 0.0139421f $X=0.545 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B_M1018_g N_A_38_297#_c_525_n 0.0124082f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B_c_194_p N_A_38_297#_c_525_n 0.0390663f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_194 N_B_c_162_n N_A_38_297#_c_525_n 0.00214031f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_195 N_B_M1020_g N_A_38_297#_c_526_n 8.33719e-19 $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B_c_174_n N_A_38_297#_c_526_n 0.00330694f $X=1.855 $Y=1.53 $X2=0 $Y2=0
cc_197 N_B_c_194_p N_A_38_297#_c_526_n 0.0163165f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_198 N_B_c_162_n N_A_38_297#_c_526_n 0.00213602f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B_M1020_g N_A_38_297#_c_554_n 0.0127541f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B_M1028_g N_A_38_297#_c_554_n 0.0112323f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B_c_173_n N_A_38_297#_c_554_n 0.00150426f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_202 N_B_c_174_n N_A_38_297#_c_554_n 0.00866684f $X=1.855 $Y=1.53 $X2=0 $Y2=0
cc_203 N_B_c_194_p N_A_38_297#_c_554_n 0.00442469f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_204 N_B_c_162_n N_A_38_297#_c_554_n 0.00167017f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B_c_173_n N_A_38_297#_c_560_n 0.0292185f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_206 N_B_c_173_n N_A_38_297#_c_561_n 0.0292185f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_207 N_B_c_163_n N_A_38_297#_c_515_n 0.00626632f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B_c_161_n N_A_38_297#_c_516_n 0.0176521f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_209 N_B_c_163_n N_A_38_297#_c_516_n 0.00561847f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B_c_173_n N_A_38_297#_c_565_n 0.0114165f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_211 N_B_c_173_n N_A_38_297#_c_566_n 0.0114165f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_212 N_B_c_173_n N_A_38_297#_c_529_n 0.0148561f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_213 N_B_M1000_g N_A_38_297#_c_530_n 0.00951001f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B_M1001_g N_A_38_297#_c_530_n 0.0103235f $X=6.535 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B_M1013_g N_A_38_297#_c_530_n 0.0103677f $X=6.955 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B_M1017_g N_A_38_297#_c_530_n 0.0120981f $X=7.375 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B_c_173_n N_A_38_297#_c_530_n 0.0120296f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_218 N_B_c_161_n N_A_38_297#_c_530_n 0.105384f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B_c_163_n N_A_38_297#_c_530_n 0.00638706f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B_M1020_g N_A_38_297#_c_531_n 0.00406924f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B_c_173_n N_A_38_297#_c_531_n 0.158668f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_222 N_B_c_174_n N_A_38_297#_c_531_n 0.0131089f $X=1.855 $Y=1.53 $X2=0 $Y2=0
cc_223 N_B_c_161_n N_A_38_297#_c_531_n 0.00607479f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B_c_194_p N_A_38_297#_c_531_n 0.0104195f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_225 N_B_c_162_n N_A_38_297#_c_531_n 0.00221769f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_226 N_B_M1007_g N_A_38_297#_c_532_n 2.84901e-19 $X=0.545 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B_M1018_g N_A_38_297#_c_532_n 0.0027915f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B_M1020_g N_A_38_297#_c_532_n 5.09574e-19 $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B_c_172_n N_A_38_297#_c_532_n 0.00116315f $X=1.77 $Y=1.445 $X2=0 $Y2=0
cc_230 N_B_c_174_n N_A_38_297#_c_532_n 2.40981e-19 $X=1.855 $Y=1.53 $X2=0 $Y2=0
cc_231 N_B_c_194_p N_A_38_297#_c_532_n 0.00798985f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_232 N_B_c_162_n N_A_38_297#_c_532_n 0.00244142f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B_M1000_g N_A_38_297#_c_533_n 0.00376143f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_234 N_B_M1001_g N_A_38_297#_c_533_n 9.85556e-19 $X=6.535 $Y=1.985 $X2=0 $Y2=0
cc_235 N_B_c_175_n N_A_38_297#_c_533_n 0.00100671f $X=5.645 $Y=1.445 $X2=0 $Y2=0
cc_236 N_B_c_161_n N_A_38_297#_c_533_n 0.00764793f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B_c_163_n N_A_38_297#_c_533_n 0.00203452f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_238 N_B_c_173_n N_VPWR_M1005_s 0.00166235f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_239 N_B_c_173_n N_VPWR_M1016_s 0.00166235f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_240 N_B_c_173_n N_VPWR_M1008_s 0.00166235f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_241 N_B_c_173_n N_VPWR_M1022_s 0.00161973f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_242 N_B_M1007_g N_VPWR_c_721_n 0.00302074f $X=0.545 $Y=1.985 $X2=0 $Y2=0
cc_243 N_B_M1018_g N_VPWR_c_721_n 0.00157837f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_244 N_B_M1020_g N_VPWR_c_722_n 0.00157837f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_245 N_B_M1028_g N_VPWR_c_722_n 0.00157837f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_246 N_B_M1028_g N_VPWR_c_729_n 0.00436487f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_247 N_B_M1018_g N_VPWR_c_739_n 0.00585385f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_248 N_B_M1020_g N_VPWR_c_739_n 0.00436487f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B_M1000_g N_VPWR_c_740_n 0.00357877f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_250 N_B_M1001_g N_VPWR_c_740_n 0.00357877f $X=6.535 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B_M1013_g N_VPWR_c_740_n 0.00357877f $X=6.955 $Y=1.985 $X2=0 $Y2=0
cc_252 N_B_M1017_g N_VPWR_c_740_n 0.00357877f $X=7.375 $Y=1.985 $X2=0 $Y2=0
cc_253 N_B_M1007_g N_VPWR_c_720_n 0.0114555f $X=0.545 $Y=1.985 $X2=0 $Y2=0
cc_254 N_B_M1018_g N_VPWR_c_720_n 0.0104367f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B_M1020_g N_VPWR_c_720_n 0.00576179f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_256 N_B_M1028_g N_VPWR_c_720_n 0.00578899f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B_M1000_g N_VPWR_c_720_n 0.00525237f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B_M1001_g N_VPWR_c_720_n 0.00522516f $X=6.535 $Y=1.985 $X2=0 $Y2=0
cc_259 N_B_M1013_g N_VPWR_c_720_n 0.00522516f $X=6.955 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B_M1017_g N_VPWR_c_720_n 0.00655123f $X=7.375 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B_M1007_g N_VPWR_c_743_n 0.00585385f $X=0.545 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B_c_173_n N_A_820_297#_M1008_d 0.00272914f $X=5.56 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_263 N_B_c_173_n N_A_820_297#_M1012_d 0.00165831f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_264 N_B_c_173_n N_A_820_297#_c_883_n 0.0292185f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_265 N_B_c_173_n N_A_820_297#_c_884_n 0.0274531f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_266 N_B_c_161_n N_A_820_297#_c_884_n 5.61731e-19 $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B_c_161_n N_A_820_297#_c_886_n 0.00157122f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B_M1000_g N_A_820_297#_c_879_n 0.0112879f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B_M1001_g N_A_820_297#_c_879_n 0.00964167f $X=6.535 $Y=1.985 $X2=0
+ $Y2=0
cc_270 N_B_M1013_g N_A_820_297#_c_879_n 0.00970685f $X=6.955 $Y=1.985 $X2=0
+ $Y2=0
cc_271 N_B_M1017_g N_A_820_297#_c_879_n 0.00970685f $X=7.375 $Y=1.985 $X2=0
+ $Y2=0
cc_272 N_B_c_173_n N_A_820_297#_c_880_n 0.0197936f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_273 N_B_c_173_n N_A_820_297#_c_892_n 0.0114165f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_274 N_B_M1000_g N_Y_c_942_n 0.00347766f $X=6.115 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B_M1001_g N_Y_c_942_n 0.0107426f $X=6.535 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B_M1013_g N_Y_c_942_n 0.0107426f $X=6.955 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B_M1017_g N_Y_c_942_n 0.0135897f $X=7.375 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B_M1017_g N_Y_c_947_n 0.00867664f $X=7.375 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B_c_153_n N_A_38_47#_c_1016_n 0.00892725f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B_c_154_n N_A_38_47#_c_1016_n 0.00892725f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B_c_155_n N_A_38_47#_c_1016_n 0.00892725f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_c_156_n N_A_38_47#_c_1016_n 0.0109954f $X=1.805 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B_c_194_p N_A_38_47#_c_1016_n 0.00253946f $X=1.685 $Y=1.175 $X2=0 $Y2=0
cc_284 N_B_c_173_n N_A_38_47#_c_1017_n 0.00701044f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_285 N_B_c_157_n N_VGND_c_1088_n 0.00146448f $X=6.115 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B_c_157_n N_VGND_c_1089_n 0.00423334f $X=6.115 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B_c_158_n N_VGND_c_1089_n 0.00423334f $X=6.535 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B_c_158_n N_VGND_c_1090_n 0.00146448f $X=6.535 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B_c_159_n N_VGND_c_1090_n 0.00146448f $X=6.955 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B_c_160_n N_VGND_c_1091_n 0.00322276f $X=7.375 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B_c_153_n N_VGND_c_1092_n 0.00357877f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B_c_154_n N_VGND_c_1092_n 0.00357877f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B_c_155_n N_VGND_c_1092_n 0.00357877f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B_c_156_n N_VGND_c_1092_n 0.00357877f $X=1.805 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B_c_159_n N_VGND_c_1102_n 0.00423334f $X=6.955 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B_c_160_n N_VGND_c_1102_n 0.00423423f $X=7.375 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B_c_153_n N_VGND_c_1104_n 0.00624395f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B_c_154_n N_VGND_c_1104_n 0.00522516f $X=0.965 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B_c_155_n N_VGND_c_1104_n 0.00522516f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B_c_156_n N_VGND_c_1104_n 0.00525237f $X=1.805 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B_c_157_n N_VGND_c_1104_n 0.0057435f $X=6.115 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B_c_158_n N_VGND_c_1104_n 0.0057163f $X=6.535 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B_c_159_n N_VGND_c_1104_n 0.0057163f $X=6.955 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B_c_160_n N_VGND_c_1104_n 0.00704386f $X=7.375 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B_c_157_n N_A_902_47#_c_1250_n 5.22228e-19 $X=6.115 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_B_c_157_n N_A_902_47#_c_1241_n 0.00864883f $X=6.115 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_B_c_197_p N_A_902_47#_c_1241_n 0.00581326f $X=5.73 $Y=1.175 $X2=0 $Y2=0
cc_308 N_B_c_161_n N_A_902_47#_c_1241_n 0.0306946f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_309 N_B_c_157_n N_A_902_47#_c_1254_n 0.00630972f $X=6.115 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_B_c_158_n N_A_902_47#_c_1254_n 0.00630972f $X=6.535 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_B_c_159_n N_A_902_47#_c_1254_n 5.22228e-19 $X=6.955 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_B_c_158_n N_A_902_47#_c_1242_n 0.00870364f $X=6.535 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_B_c_159_n N_A_902_47#_c_1242_n 0.00870364f $X=6.955 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_B_c_161_n N_A_902_47#_c_1242_n 0.036111f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_315 N_B_c_163_n N_A_902_47#_c_1242_n 0.00222133f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_316 N_B_c_158_n N_A_902_47#_c_1261_n 5.22228e-19 $X=6.535 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_B_c_159_n N_A_902_47#_c_1261_n 0.00630972f $X=6.955 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_B_c_160_n N_A_902_47#_c_1261_n 0.00724186f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_B_c_160_n N_A_902_47#_c_1243_n 0.00532457f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_B_c_160_n N_A_902_47#_c_1245_n 0.00262222f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_B_c_173_n N_A_902_47#_c_1247_n 0.00493013f $X=5.56 $Y=1.53 $X2=0 $Y2=0
cc_322 N_B_c_197_p N_A_902_47#_c_1247_n 0.00750378f $X=5.73 $Y=1.175 $X2=0 $Y2=0
cc_323 N_B_c_157_n N_A_902_47#_c_1248_n 0.00113067f $X=6.115 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_B_c_158_n N_A_902_47#_c_1248_n 0.00113286f $X=6.535 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_B_c_161_n N_A_902_47#_c_1248_n 0.0259404f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_326 N_B_c_163_n N_A_902_47#_c_1248_n 0.00230339f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_327 N_B_c_159_n N_A_902_47#_c_1249_n 0.00113286f $X=6.955 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_B_c_160_n N_A_902_47#_c_1249_n 0.00687246f $X=7.375 $Y=0.995 $X2=0
+ $Y2=0
cc_329 N_B_c_161_n N_A_902_47#_c_1249_n 0.0334729f $X=7.26 $Y=1.16 $X2=0 $Y2=0
cc_330 N_B_c_163_n N_A_902_47#_c_1249_n 0.00230339f $X=7.375 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_M1005_g N_A_38_297#_c_560_n 0.0113077f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_M1011_g N_A_38_297#_c_560_n 0.0113077f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A_M1016_g N_A_38_297#_c_561_n 0.0112504f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A_M1021_g N_A_38_297#_c_561_n 0.0113077f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A_M1026_g N_A_38_297#_c_530_n 9.11257e-19 $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_M1026_g N_A_38_297#_c_531_n 0.00158448f $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_c_365_n N_A_38_297#_c_531_n 0.0232559f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_M1026_g N_A_38_297#_c_533_n 3.16155e-19 $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_M1005_g N_VPWR_c_723_n 0.00157837f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A_M1011_g N_VPWR_c_723_n 0.00157837f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A_M1016_g N_VPWR_c_724_n 0.00157837f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_M1021_g N_VPWR_c_724_n 0.00302074f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A_M1008_g N_VPWR_c_725_n 0.00302074f $X=4.435 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_M1012_g N_VPWR_c_725_n 0.00157837f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A_M1022_g N_VPWR_c_726_n 0.00157837f $X=5.275 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A_M1026_g N_VPWR_c_726_n 0.00302074f $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A_M1005_g N_VPWR_c_729_n 0.00436487f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A_M1011_g N_VPWR_c_731_n 0.00436487f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A_M1016_g N_VPWR_c_731_n 0.00436487f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A_M1021_g N_VPWR_c_733_n 0.00436487f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_351 N_A_M1008_g N_VPWR_c_733_n 0.00436487f $X=4.435 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A_M1012_g N_VPWR_c_735_n 0.00436487f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A_M1022_g N_VPWR_c_735_n 0.00436487f $X=5.275 $Y=1.985 $X2=0 $Y2=0
cc_354 N_A_M1026_g N_VPWR_c_740_n 0.00436487f $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_355 N_A_M1005_g N_VPWR_c_720_n 0.00578899f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A_M1011_g N_VPWR_c_720_n 0.00576179f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A_M1016_g N_VPWR_c_720_n 0.00576179f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A_M1021_g N_VPWR_c_720_n 0.00708786f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A_M1008_g N_VPWR_c_720_n 0.00708786f $X=4.435 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A_M1012_g N_VPWR_c_720_n 0.00576179f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A_M1022_g N_VPWR_c_720_n 0.00576179f $X=5.275 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A_M1026_g N_VPWR_c_720_n 0.00578899f $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A_M1008_g N_A_820_297#_c_883_n 0.0113077f $X=4.435 $Y=1.985 $X2=0 $Y2=0
cc_364 N_A_M1012_g N_A_820_297#_c_883_n 0.0113077f $X=4.855 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A_M1022_g N_A_820_297#_c_884_n 0.0112504f $X=5.275 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A_M1026_g N_A_820_297#_c_884_n 0.0116687f $X=5.695 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A_c_356_n N_A_38_47#_c_1028_n 0.00255288f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A_c_356_n N_A_38_47#_c_1017_n 0.0051603f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A_c_357_n N_A_38_47#_c_1017_n 4.58193e-19 $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A_c_365_n N_A_38_47#_c_1017_n 3.71806e-19 $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_371 N_A_c_356_n N_A_38_47#_c_1018_n 0.00869748f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A_c_357_n N_A_38_47#_c_1018_n 0.0086507f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A_c_364_n N_A_38_47#_c_1018_n 0.00222133f $X=3.485 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_c_365_n N_A_38_47#_c_1018_n 0.0350477f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_375 N_A_c_356_n N_A_38_47#_c_1036_n 5.22228e-19 $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A_c_357_n N_A_38_47#_c_1036_n 0.00630972f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A_c_358_n N_A_38_47#_c_1036_n 0.00630972f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A_c_359_n N_A_38_47#_c_1036_n 5.22228e-19 $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A_c_358_n N_A_38_47#_c_1019_n 0.00869748f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_c_359_n N_A_38_47#_c_1019_n 0.00999129f $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_c_364_n N_A_38_47#_c_1019_n 0.00222133f $X=3.485 $Y=1.16 $X2=0 $Y2=0
cc_382 N_A_c_365_n N_A_38_47#_c_1019_n 0.0620128f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_c_358_n N_A_38_47#_c_1020_n 5.22228e-19 $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A_c_359_n N_A_38_47#_c_1020_n 0.00630972f $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_385 N_A_c_357_n N_A_38_47#_c_1021_n 0.00113127f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A_c_358_n N_A_38_47#_c_1021_n 0.00113127f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A_c_364_n N_A_38_47#_c_1021_n 0.00230339f $X=3.485 $Y=1.16 $X2=0 $Y2=0
cc_388 N_A_c_365_n N_A_38_47#_c_1021_n 0.0256833f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_c_356_n N_VGND_c_1084_n 0.00268723f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_390 N_A_c_357_n N_VGND_c_1084_n 0.00146448f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_391 N_A_c_358_n N_VGND_c_1085_n 0.00146448f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_392 N_A_c_359_n N_VGND_c_1085_n 0.00146992f $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_393 N_A_c_359_n N_VGND_c_1086_n 0.00245379f $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_394 N_A_c_360_n N_VGND_c_1086_n 0.00366968f $X=4.435 $Y=0.995 $X2=0 $Y2=0
cc_395 N_A_c_365_n N_VGND_c_1086_n 0.0225889f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_396 N_A_c_361_n N_VGND_c_1087_n 0.00146448f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A_c_362_n N_VGND_c_1087_n 0.00146448f $X=5.275 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A_c_363_n N_VGND_c_1088_n 0.00146448f $X=5.695 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A_c_356_n N_VGND_c_1092_n 0.00421816f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A_c_357_n N_VGND_c_1094_n 0.00423334f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_c_358_n N_VGND_c_1094_n 0.00423334f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_c_359_n N_VGND_c_1096_n 0.00423334f $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A_c_360_n N_VGND_c_1098_n 0.00541359f $X=4.435 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A_c_361_n N_VGND_c_1098_n 0.00423334f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A_c_362_n N_VGND_c_1100_n 0.00423334f $X=5.275 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A_c_363_n N_VGND_c_1100_n 0.00423334f $X=5.695 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A_c_356_n N_VGND_c_1104_n 0.00575258f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A_c_357_n N_VGND_c_1104_n 0.0057163f $X=2.645 $Y=0.995 $X2=0 $Y2=0
cc_409 N_A_c_358_n N_VGND_c_1104_n 0.0057163f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A_c_359_n N_VGND_c_1104_n 0.00704237f $X=3.485 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A_c_360_n N_VGND_c_1104_n 0.0108276f $X=4.435 $Y=0.995 $X2=0 $Y2=0
cc_412 N_A_c_361_n N_VGND_c_1104_n 0.0057163f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_413 N_A_c_362_n N_VGND_c_1104_n 0.0057163f $X=5.275 $Y=0.995 $X2=0 $Y2=0
cc_414 N_A_c_363_n N_VGND_c_1104_n 0.0057435f $X=5.695 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A_c_360_n N_A_902_47#_c_1276_n 0.00539651f $X=4.435 $Y=0.995 $X2=0
+ $Y2=0
cc_416 N_A_c_361_n N_A_902_47#_c_1276_n 0.00630972f $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_A_c_362_n N_A_902_47#_c_1276_n 5.22228e-19 $X=5.275 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A_c_361_n N_A_902_47#_c_1239_n 0.00869748f $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_A_c_362_n N_A_902_47#_c_1239_n 0.00869748f $X=5.275 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A_c_365_n N_A_902_47#_c_1239_n 0.0350477f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_421 N_A_c_366_n N_A_902_47#_c_1239_n 0.00222133f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_422 N_A_c_360_n N_A_902_47#_c_1240_n 0.00262649f $X=4.435 $Y=0.995 $X2=0
+ $Y2=0
cc_423 N_A_c_361_n N_A_902_47#_c_1240_n 0.00113127f $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_424 N_A_c_365_n N_A_902_47#_c_1240_n 0.0256833f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_425 N_A_c_366_n N_A_902_47#_c_1240_n 0.00230339f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_426 N_A_c_361_n N_A_902_47#_c_1250_n 5.22228e-19 $X=4.855 $Y=0.995 $X2=0
+ $Y2=0
cc_427 N_A_c_362_n N_A_902_47#_c_1250_n 0.00630972f $X=5.275 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A_c_363_n N_A_902_47#_c_1250_n 0.00630972f $X=5.695 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_A_c_363_n N_A_902_47#_c_1241_n 0.00864748f $X=5.695 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A_c_363_n N_A_902_47#_c_1254_n 5.22228e-19 $X=5.695 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_A_c_362_n N_A_902_47#_c_1247_n 0.00113127f $X=5.275 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_A_c_363_n N_A_902_47#_c_1247_n 0.00113002f $X=5.695 $Y=0.995 $X2=0
+ $Y2=0
cc_433 N_A_c_365_n N_A_902_47#_c_1247_n 0.00537533f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A_c_366_n N_A_902_47#_c_1247_n 0.0028467f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_435 N_A_38_297#_c_525_n N_VPWR_M1007_d 0.00185611f $X=1.05 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_436 N_A_38_297#_c_554_n N_VPWR_M1020_d 0.00383085f $X=1.89 $Y=1.895 $X2=0
+ $Y2=0
cc_437 N_A_38_297#_c_531_n N_VPWR_M1020_d 0.00179738f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_438 N_A_38_297#_c_560_n N_VPWR_M1005_s 0.00304824f $X=2.73 $Y=1.895 $X2=0
+ $Y2=0
cc_439 N_A_38_297#_c_561_n N_VPWR_M1016_s 0.00304824f $X=3.57 $Y=1.895 $X2=0
+ $Y2=0
cc_440 N_A_38_297#_c_525_n N_VPWR_c_721_n 0.0104788f $X=1.05 $Y=1.53 $X2=0 $Y2=0
cc_441 N_A_38_297#_c_554_n N_VPWR_c_722_n 0.0120197f $X=1.89 $Y=1.895 $X2=0
+ $Y2=0
cc_442 N_A_38_297#_c_560_n N_VPWR_c_723_n 0.0120197f $X=2.73 $Y=1.895 $X2=0
+ $Y2=0
cc_443 N_A_38_297#_c_561_n N_VPWR_c_724_n 0.0120197f $X=3.57 $Y=1.895 $X2=0
+ $Y2=0
cc_444 N_A_38_297#_M1010_g N_VPWR_c_727_n 0.00302074f $X=8.335 $Y=1.985 $X2=0
+ $Y2=0
cc_445 N_A_38_297#_M1014_g N_VPWR_c_727_n 0.00157837f $X=8.755 $Y=1.985 $X2=0
+ $Y2=0
cc_446 N_A_38_297#_M1029_g N_VPWR_c_728_n 0.00157837f $X=9.175 $Y=1.985 $X2=0
+ $Y2=0
cc_447 N_A_38_297#_M1037_g N_VPWR_c_728_n 0.00302074f $X=9.595 $Y=1.985 $X2=0
+ $Y2=0
cc_448 N_A_38_297#_c_554_n N_VPWR_c_729_n 0.00223194f $X=1.89 $Y=1.895 $X2=0
+ $Y2=0
cc_449 N_A_38_297#_c_560_n N_VPWR_c_729_n 0.00223194f $X=2.73 $Y=1.895 $X2=0
+ $Y2=0
cc_450 N_A_38_297#_c_565_n N_VPWR_c_729_n 0.0142343f $X=2.015 $Y=1.96 $X2=0
+ $Y2=0
cc_451 N_A_38_297#_c_560_n N_VPWR_c_731_n 0.00223194f $X=2.73 $Y=1.895 $X2=0
+ $Y2=0
cc_452 N_A_38_297#_c_561_n N_VPWR_c_731_n 0.00223194f $X=3.57 $Y=1.895 $X2=0
+ $Y2=0
cc_453 N_A_38_297#_c_566_n N_VPWR_c_731_n 0.0142343f $X=2.855 $Y=1.96 $X2=0
+ $Y2=0
cc_454 N_A_38_297#_c_561_n N_VPWR_c_733_n 0.00223194f $X=3.57 $Y=1.895 $X2=0
+ $Y2=0
cc_455 N_A_38_297#_c_529_n N_VPWR_c_733_n 0.0158369f $X=3.695 $Y=1.96 $X2=0
+ $Y2=0
cc_456 N_A_38_297#_M1014_g N_VPWR_c_737_n 0.00585385f $X=8.755 $Y=1.985 $X2=0
+ $Y2=0
cc_457 N_A_38_297#_M1029_g N_VPWR_c_737_n 0.00585385f $X=9.175 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_A_38_297#_c_554_n N_VPWR_c_739_n 0.00223194f $X=1.89 $Y=1.895 $X2=0
+ $Y2=0
cc_459 N_A_38_297#_c_625_p N_VPWR_c_739_n 0.0142343f $X=1.175 $Y=1.96 $X2=0
+ $Y2=0
cc_460 N_A_38_297#_M1010_g N_VPWR_c_740_n 0.00585385f $X=8.335 $Y=1.985 $X2=0
+ $Y2=0
cc_461 N_A_38_297#_M1037_g N_VPWR_c_741_n 0.00585385f $X=9.595 $Y=1.985 $X2=0
+ $Y2=0
cc_462 N_A_38_297#_M1007_s N_VPWR_c_720_n 0.00260431f $X=0.19 $Y=1.485 $X2=0
+ $Y2=0
cc_463 N_A_38_297#_M1018_s N_VPWR_c_720_n 0.00253454f $X=1.04 $Y=1.485 $X2=0
+ $Y2=0
cc_464 N_A_38_297#_M1028_s N_VPWR_c_720_n 0.00222276f $X=1.88 $Y=1.485 $X2=0
+ $Y2=0
cc_465 N_A_38_297#_M1011_d N_VPWR_c_720_n 0.00222276f $X=2.72 $Y=1.485 $X2=0
+ $Y2=0
cc_466 N_A_38_297#_M1021_d N_VPWR_c_720_n 0.00212053f $X=3.56 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_A_38_297#_M1010_g N_VPWR_c_720_n 0.0117628f $X=8.335 $Y=1.985 $X2=0
+ $Y2=0
cc_468 N_A_38_297#_M1014_g N_VPWR_c_720_n 0.0104367f $X=8.755 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_A_38_297#_M1029_g N_VPWR_c_720_n 0.0104367f $X=9.175 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_A_38_297#_M1037_g N_VPWR_c_720_n 0.0114397f $X=9.595 $Y=1.985 $X2=0
+ $Y2=0
cc_471 N_A_38_297#_c_524_n N_VPWR_c_720_n 0.0143649f $X=0.335 $Y=1.62 $X2=0
+ $Y2=0
cc_472 N_A_38_297#_c_554_n N_VPWR_c_720_n 0.00843576f $X=1.89 $Y=1.895 $X2=0
+ $Y2=0
cc_473 N_A_38_297#_c_560_n N_VPWR_c_720_n 0.00843576f $X=2.73 $Y=1.895 $X2=0
+ $Y2=0
cc_474 N_A_38_297#_c_561_n N_VPWR_c_720_n 0.00843576f $X=3.57 $Y=1.895 $X2=0
+ $Y2=0
cc_475 N_A_38_297#_c_625_p N_VPWR_c_720_n 0.00955092f $X=1.175 $Y=1.96 $X2=0
+ $Y2=0
cc_476 N_A_38_297#_c_565_n N_VPWR_c_720_n 0.00955092f $X=2.015 $Y=1.96 $X2=0
+ $Y2=0
cc_477 N_A_38_297#_c_566_n N_VPWR_c_720_n 0.00955092f $X=2.855 $Y=1.96 $X2=0
+ $Y2=0
cc_478 N_A_38_297#_c_529_n N_VPWR_c_720_n 0.00955092f $X=3.695 $Y=1.96 $X2=0
+ $Y2=0
cc_479 N_A_38_297#_c_524_n N_VPWR_c_743_n 0.0247699f $X=0.335 $Y=1.62 $X2=0
+ $Y2=0
cc_480 N_A_38_297#_c_530_n N_A_820_297#_M1026_d 0.0015431f $X=7.6 $Y=1.53 $X2=0
+ $Y2=0
cc_481 N_A_38_297#_c_531_n N_A_820_297#_M1026_d 0.00104207f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_482 N_A_38_297#_c_530_n N_A_820_297#_M1001_s 0.00166235f $X=7.6 $Y=1.53 $X2=0
+ $Y2=0
cc_483 N_A_38_297#_c_530_n N_A_820_297#_M1017_s 0.00276773f $X=7.6 $Y=1.53 $X2=0
+ $Y2=0
cc_484 N_A_38_297#_c_531_n N_A_820_297#_c_883_n 0.00434997f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_485 N_A_38_297#_c_531_n N_A_820_297#_c_884_n 0.00525976f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_486 N_A_38_297#_c_530_n N_A_820_297#_c_886_n 0.00607416f $X=7.6 $Y=1.53 $X2=0
+ $Y2=0
cc_487 N_A_38_297#_c_531_n N_A_820_297#_c_886_n 0.00456848f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_488 N_A_38_297#_c_530_n N_A_820_297#_c_879_n 0.00166404f $X=7.6 $Y=1.53 $X2=0
+ $Y2=0
cc_489 N_A_38_297#_c_531_n N_A_820_297#_c_879_n 4.50181e-19 $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_490 N_A_38_297#_c_533_n N_A_820_297#_c_879_n 0.0019336f $X=6.21 $Y=1.53 $X2=0
+ $Y2=0
cc_491 N_A_38_297#_c_529_n N_A_820_297#_c_880_n 0.0479914f $X=3.695 $Y=1.96
+ $X2=0 $Y2=0
cc_492 N_A_38_297#_c_531_n N_A_820_297#_c_880_n 0.00264177f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_493 N_A_38_297#_c_531_n N_A_820_297#_c_892_n 0.00209664f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_494 N_A_38_297#_c_530_n N_Y_M1000_d 0.00102351f $X=7.6 $Y=1.53 $X2=0 $Y2=0
cc_495 N_A_38_297#_c_533_n N_Y_M1000_d 0.00184953f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_496 N_A_38_297#_c_530_n N_Y_M1013_d 0.00166235f $X=7.6 $Y=1.53 $X2=0 $Y2=0
cc_497 N_A_38_297#_c_517_n N_Y_c_942_n 0.00697711f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_498 N_A_38_297#_c_530_n N_Y_c_942_n 0.0893769f $X=7.6 $Y=1.53 $X2=0 $Y2=0
cc_499 N_A_38_297#_c_533_n N_Y_c_942_n 0.00545811f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_500 N_A_38_297#_M1010_g N_Y_c_944_n 0.014983f $X=8.335 $Y=1.985 $X2=0 $Y2=0
cc_501 N_A_38_297#_M1014_g N_Y_c_944_n 0.0148339f $X=8.755 $Y=1.985 $X2=0 $Y2=0
cc_502 N_A_38_297#_c_517_n N_Y_c_944_n 0.0424318f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_503 N_A_38_297#_c_518_n N_Y_c_944_n 0.00215368f $X=9.595 $Y=1.16 $X2=0 $Y2=0
cc_504 N_A_38_297#_c_508_n N_Y_c_940_n 0.00387177f $X=8.335 $Y=0.995 $X2=0 $Y2=0
cc_505 N_A_38_297#_c_509_n N_Y_c_940_n 0.0109625f $X=8.755 $Y=0.995 $X2=0 $Y2=0
cc_506 N_A_38_297#_c_510_n N_Y_c_940_n 0.0109625f $X=9.175 $Y=0.995 $X2=0 $Y2=0
cc_507 N_A_38_297#_c_511_n N_Y_c_940_n 0.0136878f $X=9.595 $Y=0.995 $X2=0 $Y2=0
cc_508 N_A_38_297#_c_517_n N_Y_c_940_n 0.0929387f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_509 N_A_38_297#_c_518_n N_Y_c_940_n 0.00672641f $X=9.595 $Y=1.16 $X2=0 $Y2=0
cc_510 N_A_38_297#_M1029_g N_Y_c_945_n 0.0148912f $X=9.175 $Y=1.985 $X2=0 $Y2=0
cc_511 N_A_38_297#_M1037_g N_Y_c_945_n 0.0155329f $X=9.595 $Y=1.985 $X2=0 $Y2=0
cc_512 N_A_38_297#_c_517_n N_Y_c_945_n 0.0399041f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_513 N_A_38_297#_c_518_n N_Y_c_945_n 0.00215368f $X=9.595 $Y=1.16 $X2=0 $Y2=0
cc_514 N_A_38_297#_c_511_n N_Y_c_941_n 0.018715f $X=9.595 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A_38_297#_c_517_n N_Y_c_941_n 0.0161218f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_516 N_A_38_297#_M1010_g N_Y_c_947_n 7.38343e-19 $X=8.335 $Y=1.985 $X2=0 $Y2=0
cc_517 N_A_38_297#_c_517_n N_Y_c_947_n 0.0245969f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_518 N_A_38_297#_c_530_n N_Y_c_947_n 0.0137728f $X=7.6 $Y=1.53 $X2=0 $Y2=0
cc_519 N_A_38_297#_c_517_n N_Y_c_948_n 0.0203891f $X=9.465 $Y=1.16 $X2=0 $Y2=0
cc_520 N_A_38_297#_c_518_n N_Y_c_948_n 0.00222737f $X=9.595 $Y=1.16 $X2=0 $Y2=0
cc_521 N_A_38_297#_c_513_n N_A_38_47#_M1025_s 0.00271814f $X=0.32 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_522 N_A_38_297#_c_514_n N_A_38_47#_M1025_s 9.57256e-19 $X=1.595 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_523 N_A_38_297#_c_514_n N_A_38_47#_M1027_s 0.00162317f $X=1.595 $Y=0.73 $X2=0
+ $Y2=0
cc_524 N_A_38_297#_M1025_d N_A_38_47#_c_1016_n 0.00305026f $X=0.62 $Y=0.235
+ $X2=0 $Y2=0
cc_525 N_A_38_297#_M1035_d N_A_38_47#_c_1016_n 0.00305026f $X=1.46 $Y=0.235
+ $X2=0 $Y2=0
cc_526 N_A_38_297#_c_513_n N_A_38_47#_c_1016_n 0.011822f $X=0.32 $Y=0.775 $X2=0
+ $Y2=0
cc_527 N_A_38_297#_c_514_n N_A_38_47#_c_1016_n 0.0730521f $X=1.595 $Y=0.73 $X2=0
+ $Y2=0
cc_528 N_A_38_297#_c_514_n N_A_38_47#_c_1017_n 0.00841895f $X=1.595 $Y=0.73
+ $X2=0 $Y2=0
cc_529 N_A_38_297#_c_531_n N_A_38_47#_c_1017_n 0.00185567f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_530 N_A_38_297#_c_508_n N_VGND_c_1091_n 0.00300306f $X=8.335 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_38_297#_c_513_n N_VGND_c_1092_n 0.00169073f $X=0.32 $Y=0.775 $X2=0
+ $Y2=0
cc_532 N_A_38_297#_c_508_n N_VGND_c_1103_n 0.00368123f $X=8.335 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_A_38_297#_c_509_n N_VGND_c_1103_n 0.00368123f $X=8.755 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_A_38_297#_c_510_n N_VGND_c_1103_n 0.00368123f $X=9.175 $Y=0.995 $X2=0
+ $Y2=0
cc_535 N_A_38_297#_c_511_n N_VGND_c_1103_n 0.00368123f $X=9.595 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_A_38_297#_M1025_d N_VGND_c_1104_n 0.00216833f $X=0.62 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_A_38_297#_M1035_d N_VGND_c_1104_n 0.00216833f $X=1.46 $Y=0.235 $X2=0
+ $Y2=0
cc_538 N_A_38_297#_c_508_n N_VGND_c_1104_n 0.00657241f $X=8.335 $Y=0.995 $X2=0
+ $Y2=0
cc_539 N_A_38_297#_c_509_n N_VGND_c_1104_n 0.00524634f $X=8.755 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_A_38_297#_c_510_n N_VGND_c_1104_n 0.00524634f $X=9.175 $Y=0.995 $X2=0
+ $Y2=0
cc_541 N_A_38_297#_c_511_n N_VGND_c_1104_n 0.00624931f $X=9.595 $Y=0.995 $X2=0
+ $Y2=0
cc_542 N_A_38_297#_c_513_n N_VGND_c_1104_n 0.00291453f $X=0.32 $Y=0.775 $X2=0
+ $Y2=0
cc_543 N_A_38_297#_c_531_n N_A_902_47#_c_1241_n 2.60979e-19 $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_544 N_A_38_297#_c_508_n N_A_902_47#_c_1243_n 4.83058e-19 $X=8.335 $Y=0.995
+ $X2=0 $Y2=0
cc_545 N_A_38_297#_c_516_n N_A_902_47#_c_1243_n 0.0140881f $X=7.77 $Y=1.175
+ $X2=0 $Y2=0
cc_546 N_A_38_297#_c_517_n N_A_902_47#_c_1243_n 0.0355439f $X=9.465 $Y=1.16
+ $X2=0 $Y2=0
cc_547 N_A_38_297#_c_530_n N_A_902_47#_c_1243_n 0.00556609f $X=7.6 $Y=1.53 $X2=0
+ $Y2=0
cc_548 N_A_38_297#_c_508_n N_A_902_47#_c_1246_n 0.00957565f $X=8.335 $Y=0.995
+ $X2=0 $Y2=0
cc_549 N_A_38_297#_c_509_n N_A_902_47#_c_1246_n 0.00795669f $X=8.755 $Y=0.995
+ $X2=0 $Y2=0
cc_550 N_A_38_297#_c_510_n N_A_902_47#_c_1246_n 0.00795669f $X=9.175 $Y=0.995
+ $X2=0 $Y2=0
cc_551 N_A_38_297#_c_511_n N_A_902_47#_c_1246_n 0.00795669f $X=9.595 $Y=0.995
+ $X2=0 $Y2=0
cc_552 N_A_38_297#_c_517_n N_A_902_47#_c_1246_n 0.00369351f $X=9.465 $Y=1.16
+ $X2=0 $Y2=0
cc_553 N_A_38_297#_c_531_n N_A_902_47#_c_1247_n 0.0017748f $X=6.065 $Y=1.53
+ $X2=0 $Y2=0
cc_554 N_VPWR_c_720_n N_A_820_297#_M1008_d 0.00212856f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_555 N_VPWR_c_720_n N_A_820_297#_M1012_d 0.00222276f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_720_n N_A_820_297#_M1026_d 0.00219546f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_720_n N_A_820_297#_M1001_s 0.00215227f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_720_n N_A_820_297#_M1017_s 0.00209344f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_559 N_VPWR_M1008_s N_A_820_297#_c_883_n 0.00304824f $X=4.51 $Y=1.485 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_725_n N_A_820_297#_c_883_n 0.0120197f $X=4.645 $Y=2.34 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_733_n N_A_820_297#_c_883_n 0.00223194f $X=4.52 $Y=2.72 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_735_n N_A_820_297#_c_883_n 0.00223194f $X=5.36 $Y=2.72 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_720_n N_A_820_297#_c_883_n 0.00843576f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_564 N_VPWR_M1022_s N_A_820_297#_c_884_n 0.00301886f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_726_n N_A_820_297#_c_884_n 0.0120197f $X=5.485 $Y=2.34 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_735_n N_A_820_297#_c_884_n 0.00223194f $X=5.36 $Y=2.72 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_740_n N_A_820_297#_c_884_n 0.00223194f $X=8.42 $Y=2.72 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_720_n N_A_820_297#_c_884_n 0.00843576f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_740_n N_A_820_297#_c_926_n 0.012886f $X=8.42 $Y=2.72 $X2=0 $Y2=0
cc_570 N_VPWR_c_720_n N_A_820_297#_c_926_n 0.00808224f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_740_n N_A_820_297#_c_879_n 0.0999013f $X=8.42 $Y=2.72 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_720_n N_A_820_297#_c_879_n 0.0630837f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_733_n N_A_820_297#_c_880_n 0.0204957f $X=4.52 $Y=2.72 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_720_n N_A_820_297#_c_880_n 0.0120542f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_735_n N_A_820_297#_c_892_n 0.0142343f $X=5.36 $Y=2.72 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_720_n N_A_820_297#_c_892_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_720_n N_Y_M1000_d 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_578 N_VPWR_c_720_n N_Y_M1013_d 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_579 N_VPWR_c_720_n N_Y_M1010_d 0.00260431f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_580 N_VPWR_c_720_n N_Y_M1014_d 0.00284632f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_581 N_VPWR_c_720_n N_Y_M1037_d 0.00260431f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_582 N_VPWR_c_740_n N_Y_c_942_n 0.00364434f $X=8.42 $Y=2.72 $X2=0 $Y2=0
cc_583 N_VPWR_c_720_n N_Y_c_942_n 0.00882371f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_584 N_VPWR_c_740_n N_Y_c_943_n 0.0186759f $X=8.42 $Y=2.72 $X2=0 $Y2=0
cc_585 N_VPWR_c_720_n N_Y_c_943_n 0.0110914f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_586 N_VPWR_M1010_s N_Y_c_944_n 0.00167154f $X=8.41 $Y=1.485 $X2=0 $Y2=0
cc_587 N_VPWR_c_727_n N_Y_c_944_n 0.0129161f $X=8.545 $Y=2 $X2=0 $Y2=0
cc_588 N_VPWR_c_737_n N_Y_c_994_n 0.0142343f $X=9.26 $Y=2.72 $X2=0 $Y2=0
cc_589 N_VPWR_c_720_n N_Y_c_994_n 0.00955092f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_590 N_VPWR_M1029_s N_Y_c_945_n 0.00167154f $X=9.25 $Y=1.485 $X2=0 $Y2=0
cc_591 N_VPWR_c_728_n N_Y_c_945_n 0.0129161f $X=9.385 $Y=2 $X2=0 $Y2=0
cc_592 N_VPWR_c_741_n Y 0.023336f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_593 N_VPWR_c_720_n Y 0.0135946f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_594 N_A_820_297#_c_879_n N_Y_M1000_d 0.00314678f $X=7.585 $Y=2.3 $X2=0 $Y2=0
cc_595 N_A_820_297#_c_879_n N_Y_M1013_d 0.00316492f $X=7.585 $Y=2.3 $X2=0 $Y2=0
cc_596 N_A_820_297#_M1001_s N_Y_c_942_n 0.00319635f $X=6.61 $Y=1.485 $X2=0 $Y2=0
cc_597 N_A_820_297#_M1017_s N_Y_c_942_n 0.00545425f $X=7.45 $Y=1.485 $X2=0 $Y2=0
cc_598 N_A_820_297#_c_879_n N_Y_c_942_n 0.0850862f $X=7.585 $Y=2.3 $X2=0 $Y2=0
cc_599 N_A_820_297#_c_879_n N_Y_c_943_n 0.0187296f $X=7.585 $Y=2.3 $X2=0 $Y2=0
cc_600 N_Y_c_940_n N_VGND_c_1103_n 0.00129291f $X=9.815 $Y=0.775 $X2=0 $Y2=0
cc_601 N_Y_M1019_d N_VGND_c_1104_n 0.00220248f $X=8.41 $Y=0.235 $X2=0 $Y2=0
cc_602 N_Y_M1024_d N_VGND_c_1104_n 0.00220248f $X=9.25 $Y=0.235 $X2=0 $Y2=0
cc_603 N_Y_c_940_n N_VGND_c_1104_n 0.0023297f $X=9.815 $Y=0.775 $X2=0 $Y2=0
cc_604 N_Y_c_940_n N_A_902_47#_M1023_s 0.00162317f $X=9.815 $Y=0.775 $X2=0 $Y2=0
cc_605 N_Y_c_940_n N_A_902_47#_M1031_s 0.00367682f $X=9.815 $Y=0.775 $X2=0 $Y2=0
cc_606 N_Y_c_940_n N_A_902_47#_c_1243_n 0.00799569f $X=9.815 $Y=0.775 $X2=0
+ $Y2=0
cc_607 N_Y_M1019_d N_A_902_47#_c_1246_n 0.00318958f $X=8.41 $Y=0.235 $X2=0 $Y2=0
cc_608 N_Y_M1024_d N_A_902_47#_c_1246_n 0.00318958f $X=9.25 $Y=0.235 $X2=0 $Y2=0
cc_609 N_Y_c_940_n N_A_902_47#_c_1246_n 0.0832295f $X=9.815 $Y=0.775 $X2=0 $Y2=0
cc_610 N_A_38_47#_c_1018_n N_VGND_M1003_s 0.00162089f $X=2.69 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_611 N_A_38_47#_c_1019_n N_VGND_M1032_s 0.00162089f $X=3.53 $Y=0.815 $X2=0
+ $Y2=0
cc_612 N_A_38_47#_c_1018_n N_VGND_c_1084_n 0.0122559f $X=2.69 $Y=0.815 $X2=0
+ $Y2=0
cc_613 N_A_38_47#_c_1019_n N_VGND_c_1085_n 0.0122559f $X=3.53 $Y=0.815 $X2=0
+ $Y2=0
cc_614 N_A_38_47#_c_1019_n N_VGND_c_1086_n 0.0153977f $X=3.53 $Y=0.815 $X2=0
+ $Y2=0
cc_615 N_A_38_47#_c_1020_n N_VGND_c_1086_n 0.0377811f $X=3.695 $Y=0.39 $X2=0
+ $Y2=0
cc_616 N_A_38_47#_c_1016_n N_VGND_c_1092_n 0.0991547f $X=1.93 $Y=0.365 $X2=0
+ $Y2=0
cc_617 N_A_38_47#_c_1028_n N_VGND_c_1092_n 0.0152108f $X=2.055 $Y=0.475 $X2=0
+ $Y2=0
cc_618 N_A_38_47#_c_1018_n N_VGND_c_1092_n 0.00198695f $X=2.69 $Y=0.815 $X2=0
+ $Y2=0
cc_619 N_A_38_47#_c_1018_n N_VGND_c_1094_n 0.00198695f $X=2.69 $Y=0.815 $X2=0
+ $Y2=0
cc_620 N_A_38_47#_c_1036_n N_VGND_c_1094_n 0.0188551f $X=2.855 $Y=0.39 $X2=0
+ $Y2=0
cc_621 N_A_38_47#_c_1019_n N_VGND_c_1094_n 0.00198695f $X=3.53 $Y=0.815 $X2=0
+ $Y2=0
cc_622 N_A_38_47#_c_1019_n N_VGND_c_1096_n 0.00198695f $X=3.53 $Y=0.815 $X2=0
+ $Y2=0
cc_623 N_A_38_47#_c_1020_n N_VGND_c_1096_n 0.0209752f $X=3.695 $Y=0.39 $X2=0
+ $Y2=0
cc_624 N_A_38_47#_M1025_s N_VGND_c_1104_n 0.00225742f $X=0.19 $Y=0.235 $X2=0
+ $Y2=0
cc_625 N_A_38_47#_M1027_s N_VGND_c_1104_n 0.00215227f $X=1.04 $Y=0.235 $X2=0
+ $Y2=0
cc_626 N_A_38_47#_M1038_s N_VGND_c_1104_n 0.00215206f $X=1.88 $Y=0.235 $X2=0
+ $Y2=0
cc_627 N_A_38_47#_M1030_d N_VGND_c_1104_n 0.00215201f $X=2.72 $Y=0.235 $X2=0
+ $Y2=0
cc_628 N_A_38_47#_M1036_d N_VGND_c_1104_n 0.00209319f $X=3.56 $Y=0.235 $X2=0
+ $Y2=0
cc_629 N_A_38_47#_c_1016_n N_VGND_c_1104_n 0.0628989f $X=1.93 $Y=0.365 $X2=0
+ $Y2=0
cc_630 N_A_38_47#_c_1028_n N_VGND_c_1104_n 0.00940698f $X=2.055 $Y=0.475 $X2=0
+ $Y2=0
cc_631 N_A_38_47#_c_1018_n N_VGND_c_1104_n 0.00835832f $X=2.69 $Y=0.815 $X2=0
+ $Y2=0
cc_632 N_A_38_47#_c_1036_n N_VGND_c_1104_n 0.0122069f $X=2.855 $Y=0.39 $X2=0
+ $Y2=0
cc_633 N_A_38_47#_c_1019_n N_VGND_c_1104_n 0.00835832f $X=3.53 $Y=0.815 $X2=0
+ $Y2=0
cc_634 N_A_38_47#_c_1020_n N_VGND_c_1104_n 0.0124119f $X=3.695 $Y=0.39 $X2=0
+ $Y2=0
cc_635 N_VGND_c_1104_n N_A_902_47#_M1004_s 0.00215201f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_636 N_VGND_c_1104_n N_A_902_47#_M1033_s 0.00215201f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_637 N_VGND_c_1104_n N_A_902_47#_M1002_s 0.00215201f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_638 N_VGND_c_1104_n N_A_902_47#_M1015_s 0.00215201f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_639 N_VGND_c_1104_n N_A_902_47#_M1019_s 0.00212536f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_640 N_VGND_c_1104_n N_A_902_47#_M1023_s 0.00218617f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_641 N_VGND_c_1104_n N_A_902_47#_M1031_s 0.00229271f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_642 N_VGND_c_1098_n N_A_902_47#_c_1276_n 0.0188551f $X=4.98 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1104_n N_A_902_47#_c_1276_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_644 N_VGND_M1009_d N_A_902_47#_c_1239_n 0.00162089f $X=4.93 $Y=0.235 $X2=0
+ $Y2=0
cc_645 N_VGND_c_1087_n N_A_902_47#_c_1239_n 0.0122559f $X=5.065 $Y=0.39 $X2=0
+ $Y2=0
cc_646 N_VGND_c_1098_n N_A_902_47#_c_1239_n 0.00198695f $X=4.98 $Y=0 $X2=0 $Y2=0
cc_647 N_VGND_c_1100_n N_A_902_47#_c_1239_n 0.00198695f $X=5.82 $Y=0 $X2=0 $Y2=0
cc_648 N_VGND_c_1104_n N_A_902_47#_c_1239_n 0.00835832f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1086_n N_A_902_47#_c_1240_n 0.00835456f $X=4.225 $Y=0.39 $X2=0
+ $Y2=0
cc_650 N_VGND_c_1100_n N_A_902_47#_c_1250_n 0.0188551f $X=5.82 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1104_n N_A_902_47#_c_1250_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_M1039_d N_A_902_47#_c_1241_n 0.00162089f $X=5.77 $Y=0.235 $X2=0
+ $Y2=0
cc_653 N_VGND_c_1088_n N_A_902_47#_c_1241_n 0.0122559f $X=5.905 $Y=0.39 $X2=0
+ $Y2=0
cc_654 N_VGND_c_1089_n N_A_902_47#_c_1241_n 0.00198695f $X=6.66 $Y=0 $X2=0 $Y2=0
cc_655 N_VGND_c_1100_n N_A_902_47#_c_1241_n 0.00198695f $X=5.82 $Y=0 $X2=0 $Y2=0
cc_656 N_VGND_c_1104_n N_A_902_47#_c_1241_n 0.00835832f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_657 N_VGND_c_1089_n N_A_902_47#_c_1254_n 0.0188551f $X=6.66 $Y=0 $X2=0 $Y2=0
cc_658 N_VGND_c_1104_n N_A_902_47#_c_1254_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_659 N_VGND_M1006_d N_A_902_47#_c_1242_n 0.00162089f $X=6.61 $Y=0.235 $X2=0
+ $Y2=0
cc_660 N_VGND_c_1089_n N_A_902_47#_c_1242_n 0.00198695f $X=6.66 $Y=0 $X2=0 $Y2=0
cc_661 N_VGND_c_1090_n N_A_902_47#_c_1242_n 0.0122559f $X=6.745 $Y=0.39 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1102_n N_A_902_47#_c_1242_n 0.00198695f $X=7.5 $Y=0 $X2=0 $Y2=0
cc_663 N_VGND_c_1104_n N_A_902_47#_c_1242_n 0.00835832f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1102_n N_A_902_47#_c_1261_n 0.0188551f $X=7.5 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1104_n N_A_902_47#_c_1261_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_666 N_VGND_M1034_d N_A_902_47#_c_1243_n 0.00281754f $X=7.45 $Y=0.235 $X2=0
+ $Y2=0
cc_667 N_VGND_c_1091_n N_A_902_47#_c_1243_n 0.0197489f $X=7.585 $Y=0.39 $X2=0
+ $Y2=0
cc_668 N_VGND_c_1102_n N_A_902_47#_c_1243_n 6.27034e-19 $X=7.5 $Y=0 $X2=0 $Y2=0
cc_669 N_VGND_c_1103_n N_A_902_47#_c_1243_n 0.00282598f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_670 N_VGND_c_1104_n N_A_902_47#_c_1243_n 0.00773162f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1091_n N_A_902_47#_c_1244_n 0.0137035f $X=7.585 $Y=0.39 $X2=0
+ $Y2=0
cc_672 N_VGND_c_1103_n N_A_902_47#_c_1244_n 0.0130441f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_673 N_VGND_c_1104_n N_A_902_47#_c_1244_n 0.00935125f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_674 N_VGND_c_1091_n N_A_902_47#_c_1245_n 0.00590433f $X=7.585 $Y=0.39 $X2=0
+ $Y2=0
cc_675 N_VGND_c_1103_n N_A_902_47#_c_1246_n 0.0743048f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_676 N_VGND_c_1104_n N_A_902_47#_c_1246_n 0.0604695f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_677 N_VGND_c_1102_n N_A_902_47#_c_1249_n 0.00134771f $X=7.5 $Y=0 $X2=0 $Y2=0
cc_678 N_VGND_c_1104_n N_A_902_47#_c_1249_n 0.002153f $X=9.89 $Y=0 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
M1000 VGND A a_32_297# VNB nshort w=650000u l=150000u
+  ad=9.4575e+11p pd=9.41e+06u as=4.225e+11p ps=3.9e+06u
M1001 X a_32_297# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=0p ps=0u
M1002 a_114_297# D a_32_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.8e+11p pd=2.76e+06u as=2.6e+11p ps=2.52e+06u
M1003 VGND a_32_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_32_297# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_304_297# VPB phighvt w=1e+06u l=150000u
+  ad=9.2e+11p pd=7.84e+06u as=2.7e+11p ps=2.54e+06u
M1006 VGND a_32_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_32_297# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1008 a_304_297# B a_220_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1009 a_220_297# C a_114_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_32_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_32_297# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C a_32_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_32_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_32_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_32_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__o32a_2.spice.SKY130_FD_SC_HD__O32A_2.pxi
* Created: Thu Aug 27 14:40:56 2020
* 
x_PM_SKY130_FD_SC_HD__O32A_2%A_79_21# N_A_79_21#_M1007_d N_A_79_21#_M1000_d
+ N_A_79_21#_c_60_n N_A_79_21#_M1005_g N_A_79_21#_M1002_g N_A_79_21#_c_61_n
+ N_A_79_21#_M1012_g N_A_79_21#_M1008_g N_A_79_21#_c_62_n N_A_79_21#_c_63_n
+ N_A_79_21#_c_72_p N_A_79_21#_c_107_p N_A_79_21#_c_81_p N_A_79_21#_c_91_p
+ N_A_79_21#_c_64_n N_A_79_21#_c_86_p N_A_79_21#_c_100_p
+ PM_SKY130_FD_SC_HD__O32A_2%A_79_21#
x_PM_SKY130_FD_SC_HD__O32A_2%A1 N_A1_M1013_g N_A1_M1006_g A1 N_A1_c_144_n
+ N_A1_c_145_n PM_SKY130_FD_SC_HD__O32A_2%A1
x_PM_SKY130_FD_SC_HD__O32A_2%A2 N_A2_c_177_n N_A2_M1010_g N_A2_M1001_g A2
+ N_A2_c_179_n PM_SKY130_FD_SC_HD__O32A_2%A2
x_PM_SKY130_FD_SC_HD__O32A_2%A3 N_A3_M1009_g N_A3_M1000_g A3 N_A3_c_217_n
+ N_A3_c_218_n PM_SKY130_FD_SC_HD__O32A_2%A3
x_PM_SKY130_FD_SC_HD__O32A_2%B2 N_B2_c_254_n N_B2_M1007_g N_B2_M1004_g B2
+ N_B2_c_256_n PM_SKY130_FD_SC_HD__O32A_2%B2
x_PM_SKY130_FD_SC_HD__O32A_2%B1 N_B1_M1011_g N_B1_M1003_g B1 N_B1_c_296_n
+ PM_SKY130_FD_SC_HD__O32A_2%B1
x_PM_SKY130_FD_SC_HD__O32A_2%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_M1003_d
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n VPWR
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_319_n
+ PM_SKY130_FD_SC_HD__O32A_2%VPWR
x_PM_SKY130_FD_SC_HD__O32A_2%X N_X_M1005_s N_X_M1002_s X X X X X X N_X_c_367_n
+ PM_SKY130_FD_SC_HD__O32A_2%X
x_PM_SKY130_FD_SC_HD__O32A_2%VGND N_VGND_M1005_d N_VGND_M1012_d N_VGND_M1010_d
+ N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n
+ N_VGND_c_393_n N_VGND_c_394_n VGND N_VGND_c_395_n N_VGND_c_396_n
+ N_VGND_c_397_n PM_SKY130_FD_SC_HD__O32A_2%VGND
x_PM_SKY130_FD_SC_HD__O32A_2%A_345_47# N_A_345_47#_M1013_d N_A_345_47#_M1009_d
+ N_A_345_47#_M1011_d N_A_345_47#_c_447_n N_A_345_47#_c_451_n
+ N_A_345_47#_c_448_n N_A_345_47#_c_462_n N_A_345_47#_c_457_n
+ N_A_345_47#_c_444_n N_A_345_47#_c_443_n PM_SKY130_FD_SC_HD__O32A_2%A_345_47#
cc_1 VNB N_A_79_21#_c_60_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_61_n 0.0182509f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_62_n 0.00723034f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.16
cc_4 VNB N_A_79_21#_c_63_n 0.0593438f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.16
cc_5 VNB N_A_79_21#_c_64_n 0.00872092f $X=-0.19 $Y=-0.24 $X2=3.425 $Y2=1.785
cc_6 VNB N_A1_c_144_n 0.0260847f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_7 VNB N_A1_c_145_n 0.0189678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_177_n 0.0178306f $X=-0.19 $Y=-0.24 $X2=3.145 $Y2=0.235
cc_9 VNB A2 2.15474e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A2_c_179_n 0.0221035f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_11 VNB A3 0.00149073f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_12 VNB N_A3_c_217_n 0.024989f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_13 VNB N_A3_c_218_n 0.0178286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B2_c_254_n 0.0173976f $X=-0.19 $Y=-0.24 $X2=3.145 $Y2=0.235
cc_15 VNB B2 0.00243579f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_B2_c_256_n 0.0217129f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_17 VNB N_B1_M1011_g 0.024216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB B1 0.00882068f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB N_B1_c_296_n 0.0400235f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_20 VNB N_VPWR_c_319_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_388_n 0.00991007f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_22 VNB N_VGND_c_389_n 0.0339415f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_23 VNB N_VGND_c_390_n 0.0204915f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_24 VNB N_VGND_c_391_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_25 VNB N_VGND_c_392_n 0.00552413f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.16
cc_26 VNB N_VGND_c_393_n 0.0203935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_394_n 0.0063086f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=1.87
cc_28 VNB N_VGND_c_395_n 0.03962f $X=-0.19 $Y=-0.24 $X2=3.36 $Y2=0.71
cc_29 VNB N_VGND_c_396_n 0.217941f $X=-0.19 $Y=-0.24 $X2=3.36 $Y2=0.72
cc_30 VNB N_VGND_c_397_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_31 VNB N_A_345_47#_c_443_n 0.0289176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_79_21#_M1002_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB N_A_79_21#_M1008_g 0.0208957f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_34 VPB N_A_79_21#_c_62_n 0.00205725f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_35 VPB N_A_79_21#_c_63_n 0.0145282f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_36 VPB N_A_79_21#_c_64_n 0.00388469f $X=-0.19 $Y=1.305 $X2=3.425 $Y2=1.785
cc_37 VPB N_A1_M1006_g 0.020996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB A1 0.00116592f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_39 VPB N_A1_c_144_n 0.005029f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_40 VPB N_A2_M1001_g 0.0188666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB A2 0.00241175f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_42 VPB N_A2_c_179_n 0.00477593f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_43 VPB N_A3_M1000_g 0.0197804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB A3 0.00116047f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_45 VPB N_A3_c_217_n 0.00586668f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_46 VPB N_B2_M1004_g 0.0184295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB B2 0.00235037f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_48 VPB N_B2_c_256_n 0.00467716f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_49 VPB N_B1_M1003_g 0.0285192f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_50 VPB B1 0.00389979f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_51 VPB N_B1_c_296_n 0.0106223f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_52 VPB N_VPWR_c_320_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_53 VPB N_VPWR_c_321_n 0.0429874f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_54 VPB N_VPWR_c_322_n 0.011811f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_55 VPB N_VPWR_c_323_n 0.0451224f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_56 VPB N_VPWR_c_324_n 0.0179805f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_57 VPB N_VPWR_c_325_n 0.0656944f $X=-0.19 $Y=1.305 $X2=2.86 $Y2=2
cc_58 VPB N_VPWR_c_326_n 0.0158646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_319_n 0.0424765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_A_79_21#_M1008_g N_A1_M1006_g 0.0131246f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_62_n N_A1_M1006_g 0.00507161f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_72_p N_A1_M1006_g 0.0130903f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_62_n A1 0.04826f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_63_n A1 3.15549e-19 $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_72_p A1 0.0123779f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_62_n N_A1_c_144_n 0.00200274f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_63_n N_A1_c_144_n 0.0203372f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_72_p N_A1_c_144_n 0.00160939f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_61_n N_A1_c_145_n 0.0129346f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_72_p N_A2_M1001_g 0.0123027f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_81_p N_A2_M1001_g 0.00233207f $X=2.86 $Y=2 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_72_p A2 0.0113381f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_72_p N_A2_c_179_n 0.00152251f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_72_p N_A3_M1000_g 0.0106448f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_81_p N_A3_M1000_g 0.0108649f $X=2.86 $Y=2 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_86_p N_A3_M1000_g 0.00219785f $X=2.86 $Y=1.87 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_72_p A3 0.0126959f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_72_p N_A3_c_217_n 5.18848e-19 $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_64_n N_B2_c_254_n 0.00375117f $X=3.425 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_79_21#_c_81_p N_B2_M1004_g 0.0106666f $X=2.86 $Y=2 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_91_p N_B2_M1004_g 0.00860088f $X=3.325 $Y=1.87 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_64_n N_B2_M1004_g 0.00475572f $X=3.425 $Y=1.785 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_86_p N_B2_M1004_g 0.00111269f $X=2.86 $Y=1.87 $X2=0 $Y2=0
cc_84 N_A_79_21#_M1000_d B2 0.00164025f $X=2.725 $Y=1.485 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_91_p B2 0.00899128f $X=3.325 $Y=1.87 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_64_n B2 0.0419889f $X=3.425 $Y=1.785 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_86_p B2 0.00500489f $X=2.86 $Y=1.87 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_91_p N_B2_c_256_n 7.83613e-19 $X=3.325 $Y=1.87 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_64_n N_B2_c_256_n 0.00240848f $X=3.425 $Y=1.785 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_100_p N_B2_c_256_n 2.58039e-19 $X=3.425 $Y=0.71 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_64_n N_B1_M1011_g 0.0137685f $X=3.425 $Y=1.785 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_81_p N_B1_M1003_g 0.0016154f $X=2.86 $Y=2 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_91_p N_B1_M1003_g 0.00178326f $X=3.325 $Y=1.87 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_64_n B1 0.0185769f $X=3.425 $Y=1.785 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_62_n N_VPWR_M1008_d 0.00800199f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_72_p N_VPWR_M1008_d 0.0081412f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_107_p N_VPWR_M1008_d 0.00610823f $X=1.325 $Y=1.87 $X2=0 $Y2=0
cc_98 N_A_79_21#_M1002_g N_VPWR_c_321_n 0.00321781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_79_21#_M1002_g N_VPWR_c_324_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_79_21#_M1008_g N_VPWR_c_324_n 0.00541359f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_c_81_p N_VPWR_c_325_n 0.0189039f $X=2.86 $Y=2 $X2=0 $Y2=0
cc_102 N_A_79_21#_M1008_g N_VPWR_c_326_n 0.00205456f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_c_72_p N_VPWR_c_326_n 0.0152204f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_107_p N_VPWR_c_326_n 0.026419f $X=1.325 $Y=1.87 $X2=0 $Y2=0
cc_105 N_A_79_21#_M1000_d N_VPWR_c_319_n 0.00215201f $X=2.725 $Y=1.485 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_M1002_g N_VPWR_c_319_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_79_21#_M1008_g N_VPWR_c_319_n 0.0101559f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_72_p N_VPWR_c_319_n 0.0405197f $X=2.695 $Y=1.87 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_107_p N_VPWR_c_319_n 0.00125007f $X=1.325 $Y=1.87 $X2=0
+ $Y2=0
cc_110 N_A_79_21#_c_81_p N_VPWR_c_319_n 0.0122217f $X=2.86 $Y=2 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_91_p N_VPWR_c_319_n 0.0184337f $X=3.325 $Y=1.87 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_60_n N_X_c_367_n 0.0131951f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_79_21#_M1002_g N_X_c_367_n 0.0201414f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_61_n N_X_c_367_n 0.0163489f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_79_21#_M1008_g N_X_c_367_n 0.0201698f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_62_n N_X_c_367_n 0.0484225f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_63_n N_X_c_367_n 0.0326728f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_72_p A_345_297# 0.00878422f $X=2.695 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_79_21#_c_72_p A_429_297# 0.0156213f $X=2.695 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_79_21#_c_91_p A_629_297# 0.0113582f $X=3.325 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_79_21#_c_64_n A_629_297# 0.005451f $X=3.425 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_79_21#_c_60_n N_VGND_c_389_n 0.00450677f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_60_n N_VGND_c_390_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_61_n N_VGND_c_390_n 0.00541359f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_61_n N_VGND_c_391_n 0.00952644f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_62_n N_VGND_c_391_n 0.020331f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_63_n N_VGND_c_391_n 0.00110015f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_79_21#_M1007_d N_VGND_c_396_n 0.00304369f $X=3.145 $Y=0.235 $X2=0
+ $Y2=0
cc_129 N_A_79_21#_c_60_n N_VGND_c_396_n 0.0104557f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_61_n N_VGND_c_396_n 0.0103797f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_79_21#_M1007_d N_A_345_47#_c_444_n 0.00548683f $X=3.145 $Y=0.235
+ $X2=0 $Y2=0
cc_132 N_A_79_21#_c_100_p N_A_345_47#_c_444_n 0.0185943f $X=3.425 $Y=0.71 $X2=0
+ $Y2=0
cc_133 N_A_79_21#_c_64_n N_A_345_47#_c_443_n 0.00384746f $X=3.425 $Y=1.785 $X2=0
+ $Y2=0
cc_134 N_A1_c_145_n N_A2_c_177_n 0.0125313f $X=1.585 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A1_M1006_g N_A2_M1001_g 0.0620481f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_136 A1 N_A2_M1001_g 3.64771e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A1_M1006_g A2 0.00123459f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_138 A1 A2 0.0272271f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A1_c_144_n A2 0.00104616f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_140 A1 N_A2_c_179_n 0.00113485f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A1_c_144_n N_A2_c_179_n 0.0197752f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_142 A1 N_VPWR_M1008_d 0.00149498f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A1_M1006_g N_VPWR_c_325_n 0.00585385f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A1_M1006_g N_VPWR_c_326_n 0.00345545f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1006_g N_VPWR_c_319_n 0.00671297f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_c_145_n N_VGND_c_391_n 0.00932203f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A1_c_145_n N_VGND_c_393_n 0.00541359f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A1_c_145_n N_VGND_c_396_n 0.0104069f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A1_c_145_n N_A_345_47#_c_447_n 0.0056663f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_150 A1 N_A_345_47#_c_448_n 0.00165159f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A1_c_145_n N_A_345_47#_c_448_n 0.00305045f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A2_M1001_g N_A3_M1000_g 0.0368518f $X=2.07 $Y=1.985 $X2=0 $Y2=0
cc_153 A2 N_A3_M1000_g 5.098e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A2_M1001_g A3 0.00109128f $X=2.07 $Y=1.985 $X2=0 $Y2=0
cc_155 A2 A3 0.0294353f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A2_c_179_n A3 0.00115025f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_157 A2 N_A3_c_217_n 0.00106587f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A2_c_179_n N_A3_c_217_n 0.0198769f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_c_177_n N_A3_c_218_n 0.0227875f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_M1001_g N_VPWR_c_325_n 0.00585385f $X=2.07 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A2_M1001_g N_VPWR_c_319_n 0.00661129f $X=2.07 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A2_c_177_n N_VGND_c_392_n 0.00463199f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_177_n N_VGND_c_393_n 0.00415469f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_177_n N_VGND_c_396_n 0.00603429f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_177_n N_A_345_47#_c_447_n 0.00620061f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A2_c_177_n N_A_345_47#_c_451_n 0.00899381f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_167 A2 N_A_345_47#_c_451_n 0.00961793f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A2_c_179_n N_A_345_47#_c_451_n 9.82446e-19 $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A2_c_177_n N_A_345_47#_c_448_n 8.65818e-19 $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_170 A2 N_A_345_47#_c_448_n 0.00282369f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A2_c_179_n N_A_345_47#_c_448_n 0.00110149f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_c_177_n N_A_345_47#_c_457_n 5.47014e-19 $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A3_c_218_n N_B2_c_254_n 0.0121662f $X=2.57 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_174 N_A3_M1000_g N_B2_M1004_g 0.0284506f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_175 A3 N_B2_M1004_g 2.87966e-19 $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_176 A3 B2 0.0323095f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_177 N_A3_c_217_n B2 0.00409502f $X=2.55 $Y=1.16 $X2=0 $Y2=0
cc_178 A3 N_B2_c_256_n 3.50527e-19 $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A3_c_217_n N_B2_c_256_n 0.0205659f $X=2.55 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A3_M1000_g N_VPWR_c_325_n 0.00541359f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A3_M1000_g N_VPWR_c_319_n 0.00637543f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_182 A3 A_429_297# 0.00246954f $X=2.45 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_183 N_A3_c_218_n N_VGND_c_392_n 0.00463199f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A3_c_218_n N_VGND_c_395_n 0.00413951f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A3_c_218_n N_VGND_c_396_n 0.00604337f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A3_c_218_n N_A_345_47#_c_447_n 5.80627e-19 $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_187 A3 N_A_345_47#_c_451_n 0.0147844f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A3_c_217_n N_A_345_47#_c_451_n 9.96495e-19 $X=2.55 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A3_c_218_n N_A_345_47#_c_451_n 0.0127684f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A3_c_218_n N_A_345_47#_c_462_n 0.00206937f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A3_c_218_n N_A_345_47#_c_457_n 0.00413665f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B2_c_254_n N_B1_M1011_g 0.0200591f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B2_c_256_n N_B1_M1011_g 0.0108193f $X=3.07 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B2_M1004_g N_B1_M1003_g 0.0362781f $X=3.07 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B2_M1004_g N_VPWR_c_325_n 0.00541359f $X=3.07 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B2_M1004_g N_VPWR_c_319_n 0.00627491f $X=3.07 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B2_c_254_n N_VGND_c_395_n 0.00357835f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B2_c_254_n N_VGND_c_396_n 0.00553668f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B2_c_254_n N_A_345_47#_c_451_n 0.00221533f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_200 B2 N_A_345_47#_c_451_n 0.00729955f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_201 N_B2_c_256_n N_A_345_47#_c_451_n 0.00122358f $X=3.07 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B2_c_254_n N_A_345_47#_c_462_n 7.12665e-19 $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B2_c_254_n N_A_345_47#_c_457_n 0.00409601f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B2_c_254_n N_A_345_47#_c_444_n 0.00855061f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_205 B2 N_A_345_47#_c_444_n 0.00347297f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_206 N_B2_c_256_n N_A_345_47#_c_444_n 6.70009e-19 $X=3.07 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B1_M1003_g N_VPWR_c_323_n 0.004853f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_208 B1 N_VPWR_c_323_n 0.0278621f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_209 N_B1_c_296_n N_VPWR_c_323_n 0.00230437f $X=3.86 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B1_M1003_g N_VPWR_c_325_n 0.00585385f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1003_g N_VPWR_c_319_n 0.011837f $X=3.6 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1011_g N_VGND_c_395_n 0.00357877f $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_213 N_B1_M1011_g N_VGND_c_396_n 0.00652442f $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_214 N_B1_M1011_g N_A_345_47#_c_457_n 3.69453e-19 $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_215 N_B1_M1011_g N_A_345_47#_c_444_n 0.0127122f $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_216 N_B1_M1011_g N_A_345_47#_c_443_n 4.65807e-19 $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_217 B1 N_A_345_47#_c_443_n 0.0296768f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_218 N_B1_c_296_n N_A_345_47#_c_443_n 0.00824702f $X=3.86 $Y=1.16 $X2=0 $Y2=0
cc_219 N_VPWR_c_319_n N_X_M1002_s 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_324_n N_X_c_367_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_319_n N_X_c_367_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_319_n A_345_297# 0.0036717f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_223 N_VPWR_c_319_n A_429_297# 0.00585928f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_224 N_VPWR_c_319_n A_629_297# 0.00516458f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_225 N_VPWR_c_321_n N_VGND_c_389_n 0.00886897f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_226 N_X_c_367_n N_VGND_c_390_n 0.0189039f $X=0.68 $Y=0.38 $X2=0.89 $Y2=0.995
cc_227 N_X_c_367_n N_VGND_c_391_n 0.032916f $X=0.68 $Y=0.38 $X2=0.89 $Y2=1.985
cc_228 N_X_M1005_s N_VGND_c_396_n 0.00215201f $X=0.545 $Y=0.235 $X2=3.36
+ $Y2=0.72
cc_229 N_X_c_367_n N_VGND_c_396_n 0.0122217f $X=0.68 $Y=0.38 $X2=3.36 $Y2=0.72
cc_230 N_VGND_c_396_n N_A_345_47#_M1013_d 0.00215201f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_231 N_VGND_c_396_n N_A_345_47#_M1009_d 0.00215201f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_396_n N_A_345_47#_M1011_d 0.00266707f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_391_n N_A_345_47#_c_447_n 0.0217537f $X=1.26 $Y=0.38 $X2=0 $Y2=0
cc_234 N_VGND_c_393_n N_A_345_47#_c_447_n 0.018715f $X=2.195 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_396_n N_A_345_47#_c_447_n 0.0121647f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_M1010_d N_A_345_47#_c_451_n 0.012762f $X=2.145 $Y=0.235 $X2=0
+ $Y2=0
cc_237 N_VGND_c_392_n N_A_345_47#_c_451_n 0.0242585f $X=2.36 $Y=0.38 $X2=0 $Y2=0
cc_238 N_VGND_c_393_n N_A_345_47#_c_451_n 0.00232396f $X=2.195 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_395_n N_A_345_47#_c_451_n 0.00232396f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_396_n N_A_345_47#_c_451_n 0.0096743f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_391_n N_A_345_47#_c_448_n 0.00980138f $X=1.26 $Y=0.38 $X2=0
+ $Y2=0
cc_242 N_VGND_c_395_n N_A_345_47#_c_462_n 0.0188496f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_396_n N_A_345_47#_c_462_n 0.0122322f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_395_n N_A_345_47#_c_444_n 0.0381452f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_245 N_VGND_c_396_n N_A_345_47#_c_444_n 0.0236493f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_246 N_VGND_c_395_n N_A_345_47#_c_443_n 0.0240197f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_396_n N_A_345_47#_c_443_n 0.0138479f $X=3.91 $Y=0 $X2=0 $Y2=0

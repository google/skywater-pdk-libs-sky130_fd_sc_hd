# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__mux2_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.180000 0.645000 6.895000 0.815000 ;
        RECT 5.180000 0.815000 5.350000 1.325000 ;
        RECT 5.305000 0.425000 5.890000 0.645000 ;
        RECT 6.725000 0.815000 6.895000 0.995000 ;
        RECT 6.725000 0.995000 7.195000 1.165000 ;
        RECT 7.025000 1.165000 7.195000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.105000 4.475000 1.275000 ;
        RECT 4.305000 0.995000 4.475000 1.105000 ;
        RECT 4.305000 1.275000 4.475000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.960000 0.995000 8.245000 1.325000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.230000 1.075000 4.520000 1.120000 ;
        RECT 4.230000 1.120000 8.190000 1.260000 ;
        RECT 4.230000 1.260000 4.520000 1.305000 ;
        RECT 7.900000 1.075000 8.190000 1.120000 ;
        RECT 7.900000 1.260000 8.190000 1.305000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.739500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795000 0.995000 3.965000 1.495000 ;
        RECT 3.795000 1.495000 6.035000 1.665000 ;
        RECT 5.670000 0.995000 6.035000 1.495000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.215000 0.995000 9.510000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.610000 1.415000 5.900000 1.460000 ;
        RECT 5.610000 1.460000 9.570000 1.600000 ;
        RECT 5.610000 1.600000 5.900000 1.645000 ;
        RECT 9.280000 1.415000 9.570000 1.460000 ;
        RECT 9.280000 1.600000 9.570000 1.645000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 0.635000 3.285000 0.805000 ;
        RECT 0.595000 0.805000 0.815000 1.575000 ;
        RECT 0.595000 1.575000 3.285000 1.745000 ;
        RECT 0.595000 1.745000 0.765000 2.465000 ;
        RECT 1.435000 0.295000 1.605000 0.635000 ;
        RECT 1.435000 1.745000 1.605000 2.465000 ;
        RECT 2.275000 0.255000 2.445000 0.635000 ;
        RECT 2.275000 1.745000 2.445000 2.465000 ;
        RECT 3.115000 0.295000 3.285000 0.635000 ;
        RECT 3.115000 1.745000 3.285000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.090000  0.085000 0.425000 0.465000 ;
        RECT 0.935000  0.085000 1.265000 0.465000 ;
        RECT 1.775000  0.085000 2.105000 0.465000 ;
        RECT 2.615000  0.085000 2.945000 0.465000 ;
        RECT 3.455000  0.085000 3.785000 0.465000 ;
        RECT 6.060000  0.085000 6.390000 0.465000 ;
        RECT 8.815000  0.085000 9.145000 0.465000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.090000 1.915000 0.425000 2.635000 ;
        RECT 0.935000 1.915000 1.265000 2.635000 ;
        RECT 1.775000 1.915000 2.105000 2.635000 ;
        RECT 2.615000 1.915000 2.945000 2.635000 ;
        RECT 3.455000 2.255000 3.785000 2.635000 ;
        RECT 6.075000 2.175000 6.245000 2.635000 ;
        RECT 8.815000 2.255000 9.145000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.985000 1.075000 3.625000 1.245000 ;
      RECT 3.455000 0.635000 4.920000 0.805000 ;
      RECT 3.455000 0.805000 3.625000 1.075000 ;
      RECT 3.455000 1.245000 3.625000 1.835000 ;
      RECT 3.455000 1.835000 8.225000 2.005000 ;
      RECT 3.955000 0.295000 5.125000 0.465000 ;
      RECT 3.955000 2.255000 5.905000 2.425000 ;
      RECT 4.750000 0.805000 4.920000 0.935000 ;
      RECT 6.345000 0.995000 6.515000 1.495000 ;
      RECT 6.345000 1.495000 8.855000 1.665000 ;
      RECT 6.480000 2.255000 8.645000 2.425000 ;
      RECT 6.575000 0.295000 7.865000 0.465000 ;
      RECT 7.115000 0.635000 7.670000 0.805000 ;
      RECT 7.500000 0.805000 7.670000 0.935000 ;
      RECT 8.685000 0.645000 9.485000 0.815000 ;
      RECT 8.685000 0.815000 8.855000 1.495000 ;
      RECT 8.685000 1.665000 8.855000 1.915000 ;
      RECT 8.685000 1.915000 9.485000 2.085000 ;
      RECT 9.315000 0.295000 9.485000 0.645000 ;
      RECT 9.315000 1.795000 9.485000 1.915000 ;
      RECT 9.315000 2.085000 9.485000 2.465000 ;
    LAYER mcon ;
      RECT 4.750000 0.765000 4.920000 0.935000 ;
      RECT 7.500000 0.765000 7.670000 0.935000 ;
    LAYER met1 ;
      RECT 4.690000 0.735000 4.980000 0.780000 ;
      RECT 4.690000 0.780000 7.730000 0.920000 ;
      RECT 4.690000 0.920000 4.980000 0.965000 ;
      RECT 7.440000 0.735000 7.730000 0.780000 ;
      RECT 7.440000 0.920000 7.730000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2_8

* File: sky130_fd_sc_hd__and4_1.spice.pex
* Created: Thu Aug 27 14:08:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4_1%A 3 7 9 15
r30 12 15 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r31 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r32 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r34 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%B 3 7 9 10 14
r36 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.16
+ $X2=0.97 $Y2=0.995
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.16 $X2=0.97 $Y2=1.16
r38 10 15 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=1.06 $Y=0.85
+ $X2=1.06 $Y2=1.16
r39 9 10 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=0.51 $X2=1.06
+ $Y2=0.85
r40 5 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.325
+ $X2=0.97 $Y2=1.16
r41 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.97 $Y=1.325 $X2=0.97
+ $Y2=2.275
r42 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.91 $Y=0.445
+ $X2=0.91 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%C 3 7 9 10 11 16
c34 9 0 6.08002e-20 $X=1.61 $Y=0.51
r35 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.16 $X2=1.5
+ $Y2=1.325
r36 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.16 $X2=1.5
+ $Y2=0.995
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.16 $X2=1.5 $Y2=1.16
r38 11 17 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=1.565 $Y=1.19
+ $X2=1.565 $Y2=1.16
r39 10 17 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=1.565 $Y=0.85
+ $X2=1.565 $Y2=1.16
r40 9 10 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.565 $Y=0.51
+ $X2=1.565 $Y2=0.85
r41 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.49 $Y=2.275
+ $X2=1.49 $Y2=1.325
r42 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.44 $Y=0.445
+ $X2=1.44 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%D 3 7 9 12
r35 12 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.16
+ $X2=2.005 $Y2=1.325
r36 12 14 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.16
+ $X2=2.005 $Y2=0.995
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.16 $X2=1.98 $Y2=1.16
r38 9 13 1.13196 $w=9.68e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=0.84 $X2=1.98
+ $Y2=0.84
r39 7 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.92 $Y=2.275
+ $X2=1.92 $Y2=1.325
r40 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.92 $Y=0.445
+ $X2=1.92 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%A_27_47# 1 2 3 10 12 15 18 21 23 27 29 32 36
+ 38 39 41 47
c85 41 0 1.54239e-19 $X=2.535 $Y=1.16
c86 32 0 1.33435e-19 $X=2.527 $Y=1.495
r87 42 47 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.535 $Y=1.16
+ $X2=2.75 $Y2=1.16
r88 41 44 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.535 $Y2=1.325
r89 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=1.16 $X2=2.535 $Y2=1.16
r90 34 36 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.26 $Y=0.42
+ $X2=0.58 $Y2=0.42
r91 32 44 6.21953 $w=3.13e-07 $l=1.7e-07 $layer=LI1_cond $X=2.527 $Y=1.495
+ $X2=2.527 $Y2=1.325
r92 30 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=1.58
+ $X2=1.705 $Y2=1.58
r93 29 32 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=2.37 $Y=1.58
+ $X2=2.527 $Y2=1.495
r94 29 30 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.37 $Y=1.58
+ $X2=1.83 $Y2=1.58
r95 25 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.58
r96 25 27 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=2.3
r97 24 38 2.11342 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.67 $Y2=1.58
r98 23 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.58 $Y=1.58
+ $X2=1.705 $Y2=1.58
r99 23 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.58 $Y=1.58
+ $X2=0.845 $Y2=1.58
r100 19 38 4.3182 $w=2.1e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.67 $Y2=1.58
r101 19 21 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=2.3
r102 18 38 4.3182 $w=2.1e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.58 $Y=1.495
+ $X2=0.67 $Y2=1.58
r103 17 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0.585
+ $X2=0.58 $Y2=0.42
r104 17 18 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.58 $Y=0.585
+ $X2=0.58 $Y2=1.495
r105 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.325
+ $X2=2.75 $Y2=1.16
r106 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.325
+ $X2=2.75 $Y2=1.985
r107 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=0.995
+ $X2=2.75 $Y2=1.16
r108 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.995
+ $X2=2.75 $Y2=0.56
r109 3 27 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=2.065 $X2=1.705 $Y2=2.3
r110 2 21 600 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.72 $Y2=2.3
r111 1 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%VPWR 1 2 3 10 12 16 20 22 24 29 36 37 43 46
c46 3 0 1.33435e-19 $X=1.995 $Y=2.065
r47 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=2.72
+ $X2=2.46 $Y2=2.72
r52 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.23 $Y2=2.72
r57 30 32 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.46 $Y2=2.72
r59 29 32 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 25 40 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r63 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.23 $Y2=2.72
r65 24 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 22 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.72
r69 18 20 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2
r70 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.72
r71 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.34
r72 10 40 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r73 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r74 3 20 300 $w=1.7e-07 $l=4.96437e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=2.065 $X2=2.46 $Y2=2
r75 2 16 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=2.065 $X2=1.23 $Y2=2.34
r76 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%X 1 2 7 8 9 10 11 12 24 36 43
r15 43 44 0.8362 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.965 $Y=2.21 $X2=2.965
+ $Y2=2.205
r16 24 41 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.005 $Y=0.85
+ $X2=3.005 $Y2=0.805
r17 12 47 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=2.965 $Y=2.25
+ $X2=2.965 $Y2=2.34
r18 12 43 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=2.965 $Y=2.25
+ $X2=2.965 $Y2=2.21
r19 12 44 1.77299 $w=2.58e-07 $l=4e-08 $layer=LI1_cond $X=3.005 $Y=2.165
+ $X2=3.005 $Y2=2.205
r20 11 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.005 $Y=1.87
+ $X2=3.005 $Y2=2.165
r21 11 31 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=3.005 $Y=1.87
+ $X2=3.005 $Y2=1.66
r22 10 31 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.005 $Y=1.53
+ $X2=3.005 $Y2=1.66
r23 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.005 $Y=1.19
+ $X2=3.005 $Y2=1.53
r24 8 41 1.34463 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=2.965 $Y=0.785
+ $X2=2.965 $Y2=0.805
r25 8 9 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=3.005 $Y=0.87
+ $X2=3.005 $Y2=1.19
r26 8 24 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.005 $Y=0.87
+ $X2=3.005 $Y2=0.85
r27 7 8 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=2.965 $Y=0.51
+ $X2=2.965 $Y2=0.785
r28 7 36 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=2.965 $Y=0.51
+ $X2=2.965 $Y2=0.38
r29 2 47 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=2.34
r30 2 31 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.66
r31 1 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_1%VGND 1 6 8 10 20 21 24
c38 6 0 2.88263e-20 $X=2.465 $Y=0.38
r39 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r40 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r41 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r42 18 24 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.49
+ $Y2=0
r43 18 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.99
+ $Y2=0
r44 17 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r45 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r46 12 16 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r47 10 24 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.49
+ $Y2=0
r48 10 16 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.07
+ $Y2=0
r49 8 17 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r50 8 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 4 24 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0
r52 4 6 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0.38
r53 1 6 91 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_NDIFF $count=2 $X=1.995
+ $Y=0.235 $X2=2.465 $Y2=0.38
.ends


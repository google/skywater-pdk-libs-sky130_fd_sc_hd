* File: sky130_fd_sc_hd__a221oi_1.spice
* Created: Thu Aug 27 14:01:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a221oi_1.spice.pex"
.subckt sky130_fd_sc_hd__a221oi_1  VNB VPB C1 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.169 PD=0.975 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 A_204_47# N_B2_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.069875 AS=0.105625 PD=0.865 PS=0.975 NRD=9.684 NRS=9.228 M=1 R=4.33333
+ SA=75000.7 SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g A_204_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.069875 PD=1.82 PS=0.865 NRD=0 NRS=9.684 M=1 R=4.33333 SA=75001 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1003 A_465_47# N_A1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.099125
+ AS=0.169 PD=0.955 PS=1.82 NRD=18 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.7
+ A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_465_47# VNB NSHORT L=0.15 W=0.65 AD=0.19825
+ AS=0.099125 PD=1.91 PS=0.955 NRD=0 NRS=18 M=1 R=4.33333 SA=75000.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1005 N_A_109_297#_M1005_d N_C1_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1002 N_A_193_297#_M1002_d N_B2_M1002_g N_A_109_297#_M1005_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_109_297#_M1000_d N_B1_M1000_g N_A_193_297#_M1002_d VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_193_297#_M1006_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.26 PD=1.305 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_193_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.305 AS=0.1525 PD=2.61 PS=1.305 NRD=7.8603 NRS=5.8903 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_56 VPB 0 1.48028e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a221oi_1.spice.SKY130_FD_SC_HD__A221OI_1.pxi"
*
.ends
*
*

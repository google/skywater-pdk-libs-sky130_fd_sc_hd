* File: sky130_fd_sc_hd__o32a_4.pxi.spice
* Created: Tue Sep  1 19:25:55 2020
* 
x_PM_SKY130_FD_SC_HD__O32A_4%A1 N_A1_M1012_g N_A1_M1007_g N_A1_M1027_g
+ N_A1_M1019_g A1 A1 N_A1_c_135_n N_A1_c_136_n PM_SKY130_FD_SC_HD__O32A_4%A1
x_PM_SKY130_FD_SC_HD__O32A_4%A2 N_A2_M1016_g N_A2_M1003_g N_A2_M1018_g
+ N_A2_M1026_g A2 A2 N_A2_c_177_n PM_SKY130_FD_SC_HD__O32A_4%A2
x_PM_SKY130_FD_SC_HD__O32A_4%A3 N_A3_M1014_g N_A3_M1017_g N_A3_M1009_g
+ N_A3_M1015_g A3 N_A3_c_217_n N_A3_c_218_n PM_SKY130_FD_SC_HD__O32A_4%A3
x_PM_SKY130_FD_SC_HD__O32A_4%B1 N_B1_M1001_g N_B1_M1011_g N_B1_M1023_g
+ N_B1_M1013_g B1 N_B1_c_262_n N_B1_c_263_n PM_SKY130_FD_SC_HD__O32A_4%B1
x_PM_SKY130_FD_SC_HD__O32A_4%B2 N_B2_M1005_g N_B2_M1008_g N_B2_M1006_g
+ N_B2_M1010_g N_B2_c_319_n N_B2_c_320_n N_B2_c_321_n B2 N_B2_c_322_n
+ PM_SKY130_FD_SC_HD__O32A_4%B2
x_PM_SKY130_FD_SC_HD__O32A_4%A_549_297# N_A_549_297#_M1001_d
+ N_A_549_297#_M1023_d N_A_549_297#_M1006_d N_A_549_297#_M1009_s
+ N_A_549_297#_M1008_d N_A_549_297#_M1000_g N_A_549_297#_M1002_g
+ N_A_549_297#_M1021_g N_A_549_297#_M1004_g N_A_549_297#_M1024_g
+ N_A_549_297#_M1020_g N_A_549_297#_M1025_g N_A_549_297#_M1022_g
+ N_A_549_297#_c_389_n N_A_549_297#_c_374_n N_A_549_297#_c_396_n
+ N_A_549_297#_c_375_n N_A_549_297#_c_376_n N_A_549_297#_c_377_n
+ N_A_549_297#_c_378_n N_A_549_297#_c_420_n N_A_549_297#_c_391_n
+ N_A_549_297#_c_414_n N_A_549_297#_c_428_n N_A_549_297#_c_379_n
+ N_A_549_297#_c_380_n N_A_549_297#_c_381_n N_A_549_297#_c_382_n
+ N_A_549_297#_c_474_p N_A_549_297#_c_416_n N_A_549_297#_c_383_n
+ N_A_549_297#_c_384_n PM_SKY130_FD_SC_HD__O32A_4%A_549_297#
x_PM_SKY130_FD_SC_HD__O32A_4%A_27_297# N_A_27_297#_M1007_d N_A_27_297#_M1019_d
+ N_A_27_297#_M1026_s N_A_27_297#_c_540_n N_A_27_297#_c_541_n
+ N_A_27_297#_c_542_n N_A_27_297#_c_543_n N_A_27_297#_c_556_n
+ N_A_27_297#_c_544_n N_A_27_297#_c_545_n PM_SKY130_FD_SC_HD__O32A_4%A_27_297#
x_PM_SKY130_FD_SC_HD__O32A_4%VPWR N_VPWR_M1007_s N_VPWR_M1011_s N_VPWR_M1002_s
+ N_VPWR_M1004_s N_VPWR_M1022_s N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_591_n
+ N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n
+ N_VPWR_c_597_n N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n
+ VPWR N_VPWR_c_602_n N_VPWR_c_603_n N_VPWR_c_588_n N_VPWR_c_605_n
+ PM_SKY130_FD_SC_HD__O32A_4%VPWR
x_PM_SKY130_FD_SC_HD__O32A_4%A_277_297# N_A_277_297#_M1003_d
+ N_A_277_297#_M1009_d N_A_277_297#_M1015_d N_A_277_297#_c_725_n
+ N_A_277_297#_c_694_n N_A_277_297#_c_695_n N_A_277_297#_c_696_n
+ N_A_277_297#_c_697_n N_A_277_297#_c_713_n N_A_277_297#_c_698_n
+ N_A_277_297#_c_699_n PM_SKY130_FD_SC_HD__O32A_4%A_277_297#
x_PM_SKY130_FD_SC_HD__O32A_4%A_739_297# N_A_739_297#_M1011_d
+ N_A_739_297#_M1013_d N_A_739_297#_M1010_s N_A_739_297#_c_746_n
+ N_A_739_297#_c_747_n N_A_739_297#_c_758_n N_A_739_297#_c_762_n
+ N_A_739_297#_c_769_n N_A_739_297#_c_764_n N_A_739_297#_c_748_n
+ N_A_739_297#_c_749_n N_A_739_297#_c_750_n
+ PM_SKY130_FD_SC_HD__O32A_4%A_739_297#
x_PM_SKY130_FD_SC_HD__O32A_4%X N_X_M1000_d N_X_M1024_d N_X_M1002_d N_X_M1020_d
+ N_X_c_817_n N_X_c_820_n N_X_c_824_n N_X_c_812_n N_X_c_813_n N_X_c_836_n
+ N_X_c_840_n N_X_c_843_n X X X PM_SKY130_FD_SC_HD__O32A_4%X
x_PM_SKY130_FD_SC_HD__O32A_4%A_27_47# N_A_27_47#_M1012_d N_A_27_47#_M1027_d
+ N_A_27_47#_M1018_d N_A_27_47#_M1017_d N_A_27_47#_M1001_s N_A_27_47#_M1005_s
+ N_A_27_47#_c_881_n N_A_27_47#_c_882_n N_A_27_47#_c_883_n N_A_27_47#_c_884_n
+ N_A_27_47#_c_885_n N_A_27_47#_c_886_n PM_SKY130_FD_SC_HD__O32A_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O32A_4%VGND N_VGND_M1012_s N_VGND_M1016_s N_VGND_M1014_s
+ N_VGND_M1000_s N_VGND_M1021_s N_VGND_M1025_s N_VGND_c_945_n N_VGND_c_946_n
+ N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n
+ N_VGND_c_952_n N_VGND_c_953_n VGND N_VGND_c_954_n N_VGND_c_955_n
+ N_VGND_c_956_n N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n
+ PM_SKY130_FD_SC_HD__O32A_4%VGND
cc_1 VNB N_A1_M1012_g 0.0241044f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A1_M1007_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_A1_M1027_g 0.0168056f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_A1_M1019_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB N_A1_c_135_n 0.0367002f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_6 VNB N_A1_c_136_n 0.025781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_7 VNB N_A2_M1016_g 0.0168056f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_8 VNB N_A2_M1003_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_9 VNB N_A2_M1018_g 0.0170173f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_10 VNB N_A2_M1026_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_11 VNB A2 0.00451123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_177_n 0.0299286f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_13 VNB N_A3_M1014_g 0.0170173f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_14 VNB N_A3_M1017_g 0.0241044f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_15 VNB N_A3_M1009_g 7.17862e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_16 VNB N_A3_M1015_g 7.17862e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_17 VNB N_A3_c_217_n 0.00310996f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_18 VNB N_A3_c_218_n 0.0748688f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_19 VNB N_B1_M1001_g 0.0212292f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_20 VNB N_B1_M1011_g 7.19366e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_21 VNB N_B1_M1023_g 0.0169639f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_22 VNB N_B1_M1013_g 4.13233e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_23 VNB N_B1_c_262_n 0.00263632f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_24 VNB N_B1_c_263_n 0.0370846f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_25 VNB N_B2_M1005_g 0.0180967f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_26 VNB N_B2_M1008_g 4.74715e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_27 VNB N_B2_M1006_g 0.0211959f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_28 VNB N_B2_M1010_g 7.31445e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_29 VNB N_B2_c_319_n 0.00824007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_B2_c_320_n 0.0142786f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_31 VNB N_B2_c_321_n 0.011472f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_32 VNB N_B2_c_322_n 0.00136859f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_33 VNB N_A_549_297#_M1000_g 0.021414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_549_297#_M1002_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_549_297#_M1021_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_36 VNB N_A_549_297#_M1004_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_549_297#_M1024_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_549_297#_M1020_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_549_297#_M1025_g 0.0207742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_549_297#_M1022_g 4.88014e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_549_297#_c_374_n 0.0178491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_549_297#_c_375_n 0.0120406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_549_297#_c_376_n 0.00169196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_549_297#_c_377_n 0.00530411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_549_297#_c_378_n 0.00340237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_549_297#_c_379_n 0.00338168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_549_297#_c_380_n 0.00609746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_549_297#_c_381_n 0.0079406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_549_297#_c_382_n 0.00756596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_549_297#_c_383_n 0.0360636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_549_297#_c_384_n 0.0598782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VPWR_c_588_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_X_c_812_n 0.00218776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_X_c_813_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB X 0.0443776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_27_47#_c_881_n 0.0147612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_27_47#_c_882_n 0.00598208f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_58 VNB N_A_27_47#_c_883_n 0.0125434f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_59 VNB N_A_27_47#_c_884_n 0.00629395f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.175
cc_60 VNB N_A_27_47#_c_885_n 6.01562e-19 $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_61 VNB N_A_27_47#_c_886_n 0.0229995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_945_n 0.0051816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_946_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.16
cc_64 VNB N_VGND_c_947_n 0.0166345f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_65 VNB N_VGND_c_948_n 0.0780906f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=1.175
cc_66 VNB N_VGND_c_949_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_67 VNB N_VGND_c_950_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_951_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_952_n 0.0166611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_953_n 0.00487366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_954_n 0.0159491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_955_n 0.00755071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_956_n 0.0133492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_957_n 0.408917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_958_n 0.0142881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_959_n 0.00390482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VPB N_A1_M1007_g 0.0267067f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_78 VPB N_A1_M1019_g 0.0194853f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_79 VPB N_A2_M1003_g 0.0196623f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_80 VPB N_A2_M1026_g 0.0267252f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_81 VPB N_A3_M1009_g 0.0268425f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.025
cc_82 VPB N_A3_M1015_g 0.0268425f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_83 VPB N_B1_M1011_g 0.0268725f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_84 VPB N_B1_M1013_g 0.0188305f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_85 VPB N_B2_M1008_g 0.0198202f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_86 VPB N_B2_M1010_g 0.027261f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_87 VPB N_A_549_297#_M1002_g 0.0269034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_549_297#_M1004_g 0.019557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_549_297#_M1020_g 0.0195491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_549_297#_M1022_g 0.0230153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_549_297#_c_389_n 0.00304637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_549_297#_c_378_n 0.00138178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_549_297#_c_391_n 0.00474864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_297#_c_540_n 0.0116735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_297#_c_541_n 0.0316915f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_96 VPB N_A_27_297#_c_542_n 0.00241638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_297#_c_543_n 0.00320917f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_98 VPB N_A_27_297#_c_544_n 0.00181581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_297#_c_545_n 0.00421657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_589_n 0.00462218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_590_n 0.00462218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_591_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_103 VPB N_VPWR_c_592_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_593_n 0.0294655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_594_n 0.0819029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_595_n 0.00323699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_596_n 0.0404364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_597_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_598_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_599_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_600_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_601_n 0.00487564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_602_n 0.0177718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_603_n 0.0142356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_588_n 0.0832498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_605_n 0.00323699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_277_297#_c_694_n 0.0148708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_277_297#_c_695_n 0.00154215f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_119 VPB N_A_277_297#_c_696_n 0.00226708f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_120 VPB N_A_277_297#_c_697_n 0.00826596f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_121 VPB N_A_277_297#_c_698_n 0.00182586f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_122 VPB N_A_277_297#_c_699_n 0.0104897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_739_297#_c_746_n 0.00736243f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_124 VPB N_A_739_297#_c_747_n 0.0048178f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_125 VPB N_A_739_297#_c_748_n 0.0020947f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_126 VPB N_A_739_297#_c_749_n 0.0135798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_739_297#_c_750_n 0.0015346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB X 0.0126193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB X 0.0178552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 N_A1_M1027_g N_A2_M1016_g 0.0193304f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A1_M1019_g N_A2_M1003_g 0.0193304f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_132 A1 A2 0.0116776f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_133 N_A1_c_136_n A2 0.00212278f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A1_c_136_n N_A2_c_177_n 0.0193304f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A1_M1007_g N_A_27_297#_c_540_n 0.00183031f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_136 A1 N_A_27_297#_c_540_n 0.0222544f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A1_c_135_n N_A_27_297#_c_540_n 0.00689231f $X=0.465 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_M1007_g N_A_27_297#_c_541_n 0.00975139f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_M1019_g N_A_27_297#_c_541_n 6.1925e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_M1007_g N_A_27_297#_c_542_n 0.0120357f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_M1019_g N_A_27_297#_c_542_n 0.013558f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_142 A1 N_A_27_297#_c_542_n 0.0257313f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A1_c_136_n N_A_27_297#_c_542_n 0.0019951f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A1_M1019_g N_A_27_297#_c_543_n 0.00188655f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1007_g N_A_27_297#_c_556_n 5.69091e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1019_g N_A_27_297#_c_556_n 0.00975726f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_M1007_g N_VPWR_c_589_n 0.00268723f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A1_M1019_g N_VPWR_c_589_n 0.00268723f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A1_M1019_g N_VPWR_c_594_n 0.00539841f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A1_M1007_g N_VPWR_c_602_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A1_M1007_g N_VPWR_c_588_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1019_g N_VPWR_c_588_n 0.00949176f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A1_M1012_g N_A_27_47#_c_882_n 0.0154462f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A1_M1027_g N_A_27_47#_c_882_n 0.0123913f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_155 A1 N_A_27_47#_c_882_n 0.0242556f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_136_n N_A_27_47#_c_882_n 0.00205022f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_157 A1 N_A_27_47#_c_883_n 0.0139018f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A1_c_135_n N_A_27_47#_c_883_n 0.00584782f $X=0.465 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_M1012_g N_VGND_c_955_n 0.00844723f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A1_M1027_g N_VGND_c_955_n 0.0154735f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_161 N_A1_M1012_g N_VGND_c_957_n 0.00496232f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A1_M1012_g N_VGND_c_958_n 0.00339367f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A2_M1018_g N_A3_M1014_g 0.0191123f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_164 A2 N_A3_c_217_n 0.0110929f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A2_c_177_n N_A3_c_217_n 0.00180164f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A2_c_177_n N_A3_c_218_n 0.0191123f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A2_M1003_g N_A_27_297#_c_543_n 0.00317142f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_168 A2 N_A_27_297#_c_543_n 0.0164031f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A2_M1003_g N_A_27_297#_c_556_n 0.00899034f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A2_M1026_g N_A_27_297#_c_556_n 8.14766e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A2_M1003_g N_A_27_297#_c_544_n 0.0101149f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A2_M1026_g N_A_27_297#_c_544_n 0.00881754f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_M1003_g N_A_27_297#_c_545_n 7.5534e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A2_M1026_g N_A_27_297#_c_545_n 0.00666655f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A2_M1003_g N_VPWR_c_594_n 0.00357835f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A2_M1026_g N_VPWR_c_594_n 0.00357835f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1003_g N_VPWR_c_588_n 0.00525234f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_M1026_g N_VPWR_c_588_n 0.0065512f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_M1026_g N_A_277_297#_c_694_n 0.0183978f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_180 A2 N_A_277_297#_c_694_n 0.0068644f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A2_M1003_g N_A_277_297#_c_695_n 0.00107984f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_182 A2 N_A_277_297#_c_695_n 0.0137181f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_183 N_A2_c_177_n N_A_277_297#_c_695_n 0.00205276f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A2_M1026_g N_A_277_297#_c_697_n 0.00382857f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A2_M1016_g N_A_27_47#_c_882_n 0.0105972f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A2_M1018_g N_A_27_47#_c_882_n 0.0118499f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_187 A2 N_A_27_47#_c_882_n 0.0364031f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A2_c_177_n N_A_27_47#_c_882_n 0.00205022f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_M1016_g N_VGND_c_954_n 0.0154735f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A2_M1018_g N_VGND_c_954_n 0.0157269f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A3_M1009_g N_A_549_297#_c_389_n 0.00461391f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A3_M1015_g N_A_549_297#_c_389_n 0.0046145f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A3_c_218_n N_A_549_297#_c_389_n 0.0040847f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A3_c_218_n N_A_549_297#_c_374_n 0.0184924f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A3_c_217_n N_A_549_297#_c_396_n 0.0141975f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A3_c_218_n N_A_549_297#_c_396_n 0.00660782f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A3_c_218_n N_A_549_297#_c_375_n 0.00293666f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A3_M1009_g N_VPWR_c_594_n 0.00357835f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A3_M1015_g N_VPWR_c_594_n 0.00357835f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A3_M1009_g N_VPWR_c_588_n 0.0065512f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A3_M1015_g N_VPWR_c_588_n 0.0065512f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A3_c_217_n N_A_277_297#_c_694_n 0.0215291f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A3_c_218_n N_A_277_297#_c_694_n 0.00543343f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A3_M1009_g N_A_277_297#_c_696_n 0.00394447f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A3_c_217_n N_A_277_297#_c_696_n 0.0267742f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A3_c_218_n N_A_277_297#_c_696_n 0.00792212f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A3_M1009_g N_A_277_297#_c_697_n 0.00873792f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A3_M1015_g N_A_277_297#_c_697_n 8.05149e-19 $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A3_M1009_g N_A_277_297#_c_713_n 0.0101149f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A3_M1015_g N_A_277_297#_c_713_n 0.0101149f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A3_M1015_g N_A_277_297#_c_698_n 7.12665e-19 $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A3_M1009_g N_A_277_297#_c_699_n 8.77653e-19 $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A3_M1015_g N_A_277_297#_c_699_n 0.0117993f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A3_M1015_g N_A_739_297#_c_746_n 6.26407e-19 $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A3_M1014_g N_A_27_47#_c_882_n 0.0105972f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A3_M1017_g N_A_27_47#_c_882_n 0.0166781f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A3_c_217_n N_A_27_47#_c_882_n 0.034918f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A3_c_218_n N_A_27_47#_c_882_n 0.0102904f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A3_c_218_n N_A_27_47#_c_886_n 0.00395772f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A3_M1017_g N_VGND_c_948_n 0.00339367f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A3_M1014_g N_VGND_c_954_n 0.0157269f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A3_M1017_g N_VGND_c_957_n 0.00534848f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A3_M1017_g N_VGND_c_959_n 0.00844185f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_224 N_B1_M1023_g N_B2_M1005_g 0.0233529f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_225 N_B1_M1013_g N_B2_M1008_g 0.0233529f $X=4.45 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B1_c_263_n N_B2_c_319_n 0.0233529f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B1_c_263_n N_B2_c_322_n 5.82394e-19 $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_228 N_B1_c_262_n N_A_549_297#_c_374_n 0.0123937f $X=4.065 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B1_c_263_n N_A_549_297#_c_374_n 0.00119472f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B1_M1001_g N_A_549_297#_c_375_n 0.0053779f $X=4.03 $Y=0.56 $X2=0 $Y2=0
cc_231 N_B1_c_262_n N_A_549_297#_c_375_n 0.00189339f $X=4.065 $Y=1.16 $X2=0
+ $Y2=0
cc_232 N_B1_c_263_n N_A_549_297#_c_375_n 0.00209453f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B1_M1001_g N_A_549_297#_c_376_n 0.00893253f $X=4.03 $Y=0.56 $X2=0 $Y2=0
cc_234 N_B1_M1023_g N_A_549_297#_c_376_n 0.00371007f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B1_c_262_n N_A_549_297#_c_376_n 0.0147322f $X=4.065 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B1_c_263_n N_A_549_297#_c_376_n 0.00265771f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B1_M1001_g N_A_549_297#_c_378_n 0.00131437f $X=4.03 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B1_M1011_g N_A_549_297#_c_378_n 8.9314e-19 $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B1_M1023_g N_A_549_297#_c_378_n 0.00625559f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B1_M1013_g N_A_549_297#_c_378_n 0.00456119f $X=4.45 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_B1_c_262_n N_A_549_297#_c_378_n 0.014586f $X=4.065 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B1_c_263_n N_A_549_297#_c_378_n 0.0105179f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B1_M1011_g N_A_549_297#_c_414_n 5.79286e-19 $X=4.03 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_B1_M1013_g N_A_549_297#_c_414_n 0.00746964f $X=4.45 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_B1_M1023_g N_A_549_297#_c_416_n 0.00376185f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_246 N_B1_M1011_g N_VPWR_c_590_n 0.00268723f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_247 N_B1_M1013_g N_VPWR_c_590_n 0.00268723f $X=4.45 $Y=1.985 $X2=0 $Y2=0
cc_248 N_B1_M1011_g N_VPWR_c_594_n 0.00541359f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B1_M1013_g N_VPWR_c_596_n 0.00539841f $X=4.45 $Y=1.985 $X2=0 $Y2=0
cc_250 N_B1_M1011_g N_VPWR_c_588_n 0.00712156f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B1_M1013_g N_VPWR_c_588_n 0.00583177f $X=4.45 $Y=1.985 $X2=0 $Y2=0
cc_252 N_B1_M1011_g N_A_277_297#_c_699_n 0.00142513f $X=4.03 $Y=1.985 $X2=0
+ $Y2=0
cc_253 N_B1_M1011_g N_A_739_297#_c_746_n 0.00700015f $X=4.03 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_B1_M1013_g N_A_739_297#_c_746_n 0.00131467f $X=4.45 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_B1_c_262_n N_A_739_297#_c_746_n 0.00928116f $X=4.065 $Y=1.16 $X2=0
+ $Y2=0
cc_256 N_B1_c_263_n N_A_739_297#_c_746_n 0.00126157f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B1_M1011_g N_A_739_297#_c_747_n 0.0067269f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B1_M1013_g N_A_739_297#_c_747_n 5.34018e-19 $X=4.45 $Y=1.985 $X2=0
+ $Y2=0
cc_259 N_B1_M1011_g N_A_739_297#_c_758_n 0.00941328f $X=4.03 $Y=1.985 $X2=0
+ $Y2=0
cc_260 N_B1_M1013_g N_A_739_297#_c_758_n 0.0099353f $X=4.45 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B1_c_262_n N_A_739_297#_c_758_n 0.00621006f $X=4.065 $Y=1.16 $X2=0
+ $Y2=0
cc_262 N_B1_c_263_n N_A_739_297#_c_758_n 0.00203906f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_M1011_g N_A_739_297#_c_762_n 4.80671e-19 $X=4.03 $Y=1.985 $X2=0
+ $Y2=0
cc_264 N_B1_M1013_g N_A_739_297#_c_762_n 0.00459933f $X=4.45 $Y=1.985 $X2=0
+ $Y2=0
cc_265 N_B1_M1013_g N_A_739_297#_c_764_n 0.00213389f $X=4.45 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_B1_M1011_g N_A_739_297#_c_750_n 4.64231e-19 $X=4.03 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_B1_M1001_g N_A_27_47#_c_886_n 0.0112708f $X=4.03 $Y=0.56 $X2=0 $Y2=0
cc_268 N_B1_M1023_g N_A_27_47#_c_886_n 0.00860718f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_269 N_B1_M1001_g N_VGND_c_948_n 0.00357877f $X=4.03 $Y=0.56 $X2=0 $Y2=0
cc_270 N_B1_M1023_g N_VGND_c_948_n 0.00357877f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_271 N_B1_M1001_g N_VGND_c_957_n 0.00660224f $X=4.03 $Y=0.56 $X2=0 $Y2=0
cc_272 N_B1_M1023_g N_VGND_c_957_n 0.00525341f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_273 N_B2_M1005_g N_A_549_297#_c_378_n 0.00561058f $X=4.87 $Y=0.56 $X2=0 $Y2=0
cc_274 N_B2_c_319_n N_A_549_297#_c_378_n 0.00431235f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_275 N_B2_c_322_n N_A_549_297#_c_378_n 0.0165182f $X=5.095 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B2_M1005_g N_A_549_297#_c_420_n 0.00911499f $X=4.87 $Y=0.56 $X2=0 $Y2=0
cc_277 N_B2_M1006_g N_A_549_297#_c_420_n 0.0122409f $X=5.32 $Y=0.56 $X2=0 $Y2=0
cc_278 N_B2_c_320_n N_A_549_297#_c_420_n 0.00256095f $X=5.245 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_B2_c_322_n N_A_549_297#_c_420_n 0.0199021f $X=5.095 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B2_M1008_g N_A_549_297#_c_391_n 0.0118828f $X=4.87 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B2_M1010_g N_A_549_297#_c_391_n 9.21719e-19 $X=5.32 $Y=1.985 $X2=0
+ $Y2=0
cc_282 N_B2_c_320_n N_A_549_297#_c_391_n 0.00274632f $X=5.245 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_B2_c_322_n N_A_549_297#_c_391_n 0.0302425f $X=5.095 $Y=1.16 $X2=0 $Y2=0
cc_284 N_B2_M1008_g N_A_549_297#_c_428_n 0.00483324f $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_285 N_B2_M1006_g N_A_549_297#_c_380_n 0.00823039f $X=5.32 $Y=0.56 $X2=0 $Y2=0
cc_286 N_B2_c_321_n N_A_549_297#_c_382_n 0.00249748f $X=5.32 $Y=1.16 $X2=0 $Y2=0
cc_287 N_B2_c_322_n N_A_549_297#_c_382_n 0.0119158f $X=5.095 $Y=1.16 $X2=0 $Y2=0
cc_288 N_B2_c_321_n N_A_549_297#_c_383_n 0.00566067f $X=5.32 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B2_M1010_g N_VPWR_c_591_n 0.00194637f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_290 N_B2_M1008_g N_VPWR_c_596_n 0.00357835f $X=4.87 $Y=1.985 $X2=0 $Y2=0
cc_291 N_B2_M1010_g N_VPWR_c_596_n 0.00357835f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_292 N_B2_M1008_g N_VPWR_c_588_n 0.00533296f $X=4.87 $Y=1.985 $X2=0 $Y2=0
cc_293 N_B2_M1010_g N_VPWR_c_588_n 0.00663183f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_294 N_B2_M1008_g N_A_739_297#_c_758_n 0.00257035f $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_B2_M1008_g N_A_739_297#_c_762_n 0.00482758f $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_B2_M1010_g N_A_739_297#_c_762_n 4.93332e-19 $X=5.32 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_B2_M1008_g N_A_739_297#_c_769_n 0.00871845f $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_B2_M1010_g N_A_739_297#_c_769_n 0.0105709f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_299 N_B2_M1008_g N_A_739_297#_c_764_n 7.39973e-19 $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_B2_M1010_g N_A_739_297#_c_748_n 7.39973e-19 $X=5.32 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_B2_M1008_g N_A_739_297#_c_749_n 7.04912e-19 $X=4.87 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_B2_M1010_g N_A_739_297#_c_749_n 0.0117137f $X=5.32 $Y=1.985 $X2=0 $Y2=0
cc_303 N_B2_M1005_g N_A_27_47#_c_886_n 0.00861238f $X=4.87 $Y=0.56 $X2=0 $Y2=0
cc_304 N_B2_M1006_g N_A_27_47#_c_886_n 0.0104463f $X=5.32 $Y=0.56 $X2=0 $Y2=0
cc_305 N_B2_M1006_g N_VGND_c_945_n 0.0055724f $X=5.32 $Y=0.56 $X2=0 $Y2=0
cc_306 N_B2_M1005_g N_VGND_c_948_n 0.00357877f $X=4.87 $Y=0.56 $X2=0 $Y2=0
cc_307 N_B2_M1006_g N_VGND_c_948_n 0.00357877f $X=5.32 $Y=0.56 $X2=0 $Y2=0
cc_308 N_B2_M1005_g N_VGND_c_957_n 0.00533105f $X=4.87 $Y=0.56 $X2=0 $Y2=0
cc_309 N_B2_M1006_g N_VGND_c_957_n 0.00667988f $X=5.32 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A_549_297#_M1002_g N_VPWR_c_591_n 0.00316354f $X=6.26 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_549_297#_c_381_n N_VPWR_c_591_n 0.00507078f $X=6.04 $Y=1.17 $X2=0
+ $Y2=0
cc_312 N_A_549_297#_c_383_n N_VPWR_c_591_n 0.00295642f $X=6.185 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A_549_297#_M1004_g N_VPWR_c_592_n 0.00146448f $X=6.68 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_549_297#_M1020_g N_VPWR_c_592_n 0.00146448f $X=7.1 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_549_297#_M1022_g N_VPWR_c_593_n 0.00321527f $X=7.52 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_549_297#_M1002_g N_VPWR_c_598_n 0.00541359f $X=6.26 $Y=1.985 $X2=0
+ $Y2=0
cc_317 N_A_549_297#_M1004_g N_VPWR_c_598_n 0.00541359f $X=6.68 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_549_297#_M1020_g N_VPWR_c_600_n 0.00541359f $X=7.1 $Y=1.985 $X2=0
+ $Y2=0
cc_319 N_A_549_297#_M1022_g N_VPWR_c_600_n 0.00541359f $X=7.52 $Y=1.985 $X2=0
+ $Y2=0
cc_320 N_A_549_297#_M1009_s N_VPWR_c_588_n 0.00216833f $X=2.745 $Y=1.485 $X2=0
+ $Y2=0
cc_321 N_A_549_297#_M1008_d N_VPWR_c_588_n 0.00240926f $X=4.945 $Y=1.485 $X2=0
+ $Y2=0
cc_322 N_A_549_297#_M1002_g N_VPWR_c_588_n 0.0108276f $X=6.26 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_549_297#_M1004_g N_VPWR_c_588_n 0.00950154f $X=6.68 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_549_297#_M1020_g N_VPWR_c_588_n 0.00950154f $X=7.1 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_549_297#_M1022_g N_VPWR_c_588_n 0.0106413f $X=7.52 $Y=1.985 $X2=0
+ $Y2=0
cc_326 N_A_549_297#_c_389_n N_A_277_297#_c_696_n 0.0117939f $X=2.88 $Y=1.865
+ $X2=0 $Y2=0
cc_327 N_A_549_297#_M1009_s N_A_277_297#_c_713_n 0.0034358f $X=2.745 $Y=1.485
+ $X2=0 $Y2=0
cc_328 N_A_549_297#_c_389_n N_A_277_297#_c_713_n 0.0085321f $X=2.88 $Y=1.865
+ $X2=0 $Y2=0
cc_329 N_A_549_297#_c_389_n N_A_277_297#_c_699_n 0.0239807f $X=2.88 $Y=1.865
+ $X2=0 $Y2=0
cc_330 N_A_549_297#_c_374_n N_A_277_297#_c_699_n 0.0275043f $X=3.455 $Y=1.19
+ $X2=0 $Y2=0
cc_331 N_A_549_297#_c_391_n N_A_739_297#_M1013_d 0.00124373f $X=5.025 $Y=1.53
+ $X2=0 $Y2=0
cc_332 N_A_549_297#_c_414_n N_A_739_297#_M1013_d 4.20517e-19 $X=4.62 $Y=1.53
+ $X2=0 $Y2=0
cc_333 N_A_549_297#_c_376_n N_A_739_297#_c_746_n 0.00688653f $X=4.4 $Y=0.72
+ $X2=0 $Y2=0
cc_334 N_A_549_297#_c_414_n N_A_739_297#_c_746_n 0.00658484f $X=4.62 $Y=1.53
+ $X2=0 $Y2=0
cc_335 N_A_549_297#_c_391_n N_A_739_297#_c_758_n 0.0118491f $X=5.025 $Y=1.53
+ $X2=0 $Y2=0
cc_336 N_A_549_297#_c_414_n N_A_739_297#_c_758_n 0.0131261f $X=4.62 $Y=1.53
+ $X2=0 $Y2=0
cc_337 N_A_549_297#_c_428_n N_A_739_297#_c_758_n 0.0117759f $X=5.11 $Y=1.95
+ $X2=0 $Y2=0
cc_338 N_A_549_297#_c_428_n N_A_739_297#_c_762_n 0.010389f $X=5.11 $Y=1.95 $X2=0
+ $Y2=0
cc_339 N_A_549_297#_M1008_d N_A_739_297#_c_769_n 0.00396155f $X=4.945 $Y=1.485
+ $X2=0 $Y2=0
cc_340 N_A_549_297#_c_391_n N_A_739_297#_c_769_n 0.00316936f $X=5.025 $Y=1.53
+ $X2=0 $Y2=0
cc_341 N_A_549_297#_c_428_n N_A_739_297#_c_769_n 0.0124067f $X=5.11 $Y=1.95
+ $X2=0 $Y2=0
cc_342 N_A_549_297#_M1002_g N_A_739_297#_c_749_n 0.00754979f $X=6.26 $Y=1.985
+ $X2=0 $Y2=0
cc_343 N_A_549_297#_c_420_n N_A_739_297#_c_749_n 0.00392771f $X=5.52 $Y=0.72
+ $X2=0 $Y2=0
cc_344 N_A_549_297#_c_391_n N_A_739_297#_c_749_n 0.00822727f $X=5.025 $Y=1.53
+ $X2=0 $Y2=0
cc_345 N_A_549_297#_c_382_n N_A_739_297#_c_749_n 0.0155624f $X=5.775 $Y=1.17
+ $X2=0 $Y2=0
cc_346 N_A_549_297#_M1000_g N_X_c_817_n 0.0052782f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A_549_297#_M1021_g N_X_c_817_n 0.00620543f $X=6.68 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A_549_297#_M1024_g N_X_c_817_n 5.19281e-19 $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A_549_297#_M1002_g N_X_c_820_n 0.00418271f $X=6.26 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A_549_297#_M1004_g N_X_c_820_n 9.81519e-19 $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_351 N_A_549_297#_c_474_p N_X_c_820_n 0.0152982f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A_549_297#_c_384_n N_X_c_820_n 0.00205364f $X=7.52 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A_549_297#_M1002_g N_X_c_824_n 0.0108021f $X=6.26 $Y=1.985 $X2=0 $Y2=0
cc_354 N_A_549_297#_M1004_g N_X_c_824_n 0.00975139f $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_355 N_A_549_297#_M1020_g N_X_c_824_n 6.1949e-19 $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A_549_297#_M1021_g N_X_c_812_n 0.00890471f $X=6.68 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_549_297#_M1024_g N_X_c_812_n 0.00890471f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_549_297#_c_474_p N_X_c_812_n 0.0594155f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A_549_297#_c_384_n N_X_c_812_n 0.00205999f $X=7.52 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A_549_297#_M1000_g N_X_c_813_n 0.00291527f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_549_297#_M1021_g N_X_c_813_n 0.00116017f $X=6.68 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_549_297#_c_380_n N_X_c_813_n 6.95047e-19 $X=5.647 $Y=1.075 $X2=0
+ $Y2=0
cc_363 N_A_549_297#_c_474_p N_X_c_813_n 0.0262563f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_364 N_A_549_297#_c_384_n N_X_c_813_n 0.00213429f $X=7.52 $Y=1.16 $X2=0 $Y2=0
cc_365 N_A_549_297#_M1004_g N_X_c_836_n 0.0110913f $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A_549_297#_M1020_g N_X_c_836_n 0.0110913f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A_549_297#_c_474_p N_X_c_836_n 0.0368171f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_368 N_A_549_297#_c_384_n N_X_c_836_n 0.00194825f $X=7.52 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A_549_297#_M1021_g N_X_c_840_n 5.2007e-19 $X=6.68 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_549_297#_M1024_g N_X_c_840_n 0.00631111f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_549_297#_M1025_g N_X_c_840_n 0.0109535f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_549_297#_M1004_g N_X_c_843_n 6.20279e-19 $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_373 N_A_549_297#_M1020_g N_X_c_843_n 0.00985707f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A_549_297#_M1022_g N_X_c_843_n 0.0146918f $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A_549_297#_M1024_g X 0.0012996f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A_549_297#_M1025_g X 0.0384512f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A_549_297#_c_474_p X 0.0145279f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A_549_297#_c_384_n X 0.00205999f $X=7.52 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_549_297#_M1020_g X 0.00103475f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A_549_297#_M1022_g X 0.0152974f $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A_549_297#_c_384_n X 0.00194825f $X=7.52 $Y=1.16 $X2=0 $Y2=0
cc_382 N_A_549_297#_c_376_n N_A_27_47#_M1001_s 0.00431257f $X=4.4 $Y=0.72 $X2=0
+ $Y2=0
cc_383 N_A_549_297#_c_420_n N_A_27_47#_M1005_s 0.00400597f $X=5.52 $Y=0.72 $X2=0
+ $Y2=0
cc_384 N_A_549_297#_c_396_n N_A_27_47#_c_882_n 0.0121626f $X=2.965 $Y=1.19 $X2=0
+ $Y2=0
cc_385 N_A_549_297#_c_375_n N_A_27_47#_c_882_n 0.0032466f $X=3.55 $Y=1.105 $X2=0
+ $Y2=0
cc_386 N_A_549_297#_c_377_n N_A_27_47#_c_882_n 0.00761768f $X=3.645 $Y=0.72
+ $X2=0 $Y2=0
cc_387 N_A_549_297#_M1001_d N_A_27_47#_c_886_n 0.00501743f $X=3.695 $Y=0.235
+ $X2=0 $Y2=0
cc_388 N_A_549_297#_M1023_d N_A_27_47#_c_886_n 0.00313628f $X=4.525 $Y=0.235
+ $X2=0 $Y2=0
cc_389 N_A_549_297#_M1006_d N_A_27_47#_c_886_n 0.00500321f $X=5.395 $Y=0.235
+ $X2=0 $Y2=0
cc_390 N_A_549_297#_c_374_n N_A_27_47#_c_886_n 0.0140981f $X=3.455 $Y=1.19 $X2=0
+ $Y2=0
cc_391 N_A_549_297#_c_376_n N_A_27_47#_c_886_n 0.0400874f $X=4.4 $Y=0.72 $X2=0
+ $Y2=0
cc_392 N_A_549_297#_c_377_n N_A_27_47#_c_886_n 0.0153145f $X=3.645 $Y=0.72 $X2=0
+ $Y2=0
cc_393 N_A_549_297#_c_420_n N_A_27_47#_c_886_n 0.0455132f $X=5.52 $Y=0.72 $X2=0
+ $Y2=0
cc_394 N_A_549_297#_c_379_n N_A_27_47#_c_886_n 0.0136888f $X=5.647 $Y=0.805
+ $X2=0 $Y2=0
cc_395 N_A_549_297#_c_416_n N_A_27_47#_c_886_n 0.0120569f $X=4.51 $Y=0.72 $X2=0
+ $Y2=0
cc_396 N_A_549_297#_M1000_g N_VGND_c_945_n 0.00316354f $X=6.26 $Y=0.56 $X2=0
+ $Y2=0
cc_397 N_A_549_297#_c_379_n N_VGND_c_945_n 0.0130371f $X=5.647 $Y=0.805 $X2=0
+ $Y2=0
cc_398 N_A_549_297#_c_380_n N_VGND_c_945_n 0.00560016f $X=5.647 $Y=1.075 $X2=0
+ $Y2=0
cc_399 N_A_549_297#_c_381_n N_VGND_c_945_n 0.0119798f $X=6.04 $Y=1.17 $X2=0
+ $Y2=0
cc_400 N_A_549_297#_c_383_n N_VGND_c_945_n 0.00393791f $X=6.185 $Y=1.16 $X2=0
+ $Y2=0
cc_401 N_A_549_297#_M1021_g N_VGND_c_946_n 0.00146448f $X=6.68 $Y=0.56 $X2=0
+ $Y2=0
cc_402 N_A_549_297#_M1024_g N_VGND_c_946_n 0.00146448f $X=7.1 $Y=0.56 $X2=0
+ $Y2=0
cc_403 N_A_549_297#_M1025_g N_VGND_c_947_n 0.00321527f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_404 N_A_549_297#_c_379_n N_VGND_c_948_n 0.00161476f $X=5.647 $Y=0.805 $X2=0
+ $Y2=0
cc_405 N_A_549_297#_M1000_g N_VGND_c_950_n 0.00541359f $X=6.26 $Y=0.56 $X2=0
+ $Y2=0
cc_406 N_A_549_297#_M1021_g N_VGND_c_950_n 0.00422241f $X=6.68 $Y=0.56 $X2=0
+ $Y2=0
cc_407 N_A_549_297#_M1024_g N_VGND_c_952_n 0.00421248f $X=7.1 $Y=0.56 $X2=0
+ $Y2=0
cc_408 N_A_549_297#_M1025_g N_VGND_c_952_n 0.00421248f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_409 N_A_549_297#_M1001_d N_VGND_c_957_n 0.00210147f $X=3.695 $Y=0.235 $X2=0
+ $Y2=0
cc_410 N_A_549_297#_M1023_d N_VGND_c_957_n 0.00216833f $X=4.525 $Y=0.235 $X2=0
+ $Y2=0
cc_411 N_A_549_297#_M1006_d N_VGND_c_957_n 0.00210147f $X=5.395 $Y=0.235 $X2=0
+ $Y2=0
cc_412 N_A_549_297#_M1000_g N_VGND_c_957_n 0.0108276f $X=6.26 $Y=0.56 $X2=0
+ $Y2=0
cc_413 N_A_549_297#_M1021_g N_VGND_c_957_n 0.00569656f $X=6.68 $Y=0.56 $X2=0
+ $Y2=0
cc_414 N_A_549_297#_M1024_g N_VGND_c_957_n 0.00571103f $X=7.1 $Y=0.56 $X2=0
+ $Y2=0
cc_415 N_A_549_297#_M1025_g N_VGND_c_957_n 0.00685076f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_416 N_A_549_297#_c_379_n N_VGND_c_957_n 0.00283774f $X=5.647 $Y=0.805 $X2=0
+ $Y2=0
cc_417 N_A_27_297#_c_542_n N_VPWR_M1007_s 0.00167154f $X=0.935 $Y=1.555
+ $X2=-0.19 $Y2=1.305
cc_418 N_A_27_297#_c_542_n N_VPWR_c_589_n 0.0129161f $X=0.935 $Y=1.555 $X2=0
+ $Y2=0
cc_419 N_A_27_297#_c_556_n N_VPWR_c_594_n 0.0190403f $X=1.1 $Y=2.295 $X2=0 $Y2=0
cc_420 N_A_27_297#_c_544_n N_VPWR_c_594_n 0.0496369f $X=1.775 $Y=2.38 $X2=0
+ $Y2=0
cc_421 N_A_27_297#_c_541_n N_VPWR_c_602_n 0.0217551f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_422 N_A_27_297#_M1007_d N_VPWR_c_588_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_423 N_A_27_297#_M1019_d N_VPWR_c_588_n 0.00215201f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_424 N_A_27_297#_M1026_s N_VPWR_c_588_n 0.00209319f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_425 N_A_27_297#_c_541_n N_VPWR_c_588_n 0.0128119f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_426 N_A_27_297#_c_556_n N_VPWR_c_588_n 0.0122896f $X=1.1 $Y=2.295 $X2=0 $Y2=0
cc_427 N_A_27_297#_c_544_n N_VPWR_c_588_n 0.0303579f $X=1.775 $Y=2.38 $X2=0
+ $Y2=0
cc_428 N_A_27_297#_c_544_n N_A_277_297#_M1003_d 0.0034358f $X=1.775 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_429 N_A_27_297#_c_544_n N_A_277_297#_c_725_n 0.00845382f $X=1.775 $Y=2.38
+ $X2=0 $Y2=0
cc_430 N_A_27_297#_M1026_s N_A_277_297#_c_694_n 0.00308569f $X=1.805 $Y=1.485
+ $X2=0 $Y2=0
cc_431 N_A_27_297#_c_544_n N_A_277_297#_c_694_n 0.00290214f $X=1.775 $Y=2.38
+ $X2=0 $Y2=0
cc_432 N_A_27_297#_c_545_n N_A_277_297#_c_694_n 0.0223255f $X=1.94 $Y=2 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_c_543_n N_A_277_297#_c_695_n 0.0111374f $X=1.1 $Y=1.665 $X2=0
+ $Y2=0
cc_434 N_A_27_297#_c_544_n N_A_277_297#_c_697_n 0.0147157f $X=1.775 $Y=2.38
+ $X2=0 $Y2=0
cc_435 N_A_27_297#_c_545_n N_A_277_297#_c_697_n 0.033419f $X=1.94 $Y=2 $X2=0
+ $Y2=0
cc_436 N_A_27_297#_c_542_n N_A_27_47#_c_882_n 0.00379316f $X=0.935 $Y=1.555
+ $X2=0 $Y2=0
cc_437 N_A_27_297#_c_543_n N_A_27_47#_c_882_n 0.0037624f $X=1.1 $Y=1.665 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_c_540_n N_A_27_47#_c_883_n 0.00258654f $X=0.255 $Y=1.665
+ $X2=0 $Y2=0
cc_439 N_VPWR_c_588_n N_A_277_297#_M1003_d 0.00216833f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_440 N_VPWR_c_588_n N_A_277_297#_M1009_d 0.00209319f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_588_n N_A_277_297#_M1015_d 0.00209319f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_594_n N_A_277_297#_c_697_n 0.021178f $X=4.155 $Y=2.72 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_588_n N_A_277_297#_c_697_n 0.0124992f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_594_n N_A_277_297#_c_713_n 0.0286211f $X=4.155 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_588_n N_A_277_297#_c_713_n 0.0178969f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_594_n N_A_277_297#_c_698_n 0.021178f $X=4.155 $Y=2.72 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_588_n N_A_277_297#_c_698_n 0.0124992f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_588_n N_A_739_297#_M1011_d 0.00209319f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_449 N_VPWR_c_588_n N_A_739_297#_M1013_d 0.00215201f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_588_n N_A_739_297#_M1010_s 0.00209319f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_594_n N_A_739_297#_c_747_n 0.0210382f $X=4.155 $Y=2.72 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_588_n N_A_739_297#_c_747_n 0.0124268f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_M1011_s N_A_739_297#_c_758_n 0.00486285f $X=4.105 $Y=1.485 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_590_n N_A_739_297#_c_758_n 0.0123301f $X=4.24 $Y=2.29 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_588_n N_A_739_297#_c_758_n 0.0112186f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_596_n N_A_739_297#_c_769_n 0.0306231f $X=5.965 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_588_n N_A_739_297#_c_769_n 0.0190382f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_596_n N_A_739_297#_c_764_n 0.0190403f $X=5.965 $Y=2.72 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_588_n N_A_739_297#_c_764_n 0.0122896f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_591_n N_A_739_297#_c_748_n 0.0107408f $X=6.05 $Y=2 $X2=0 $Y2=0
cc_461 N_VPWR_c_596_n N_A_739_297#_c_748_n 0.021178f $X=5.965 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_588_n N_A_739_297#_c_748_n 0.0124992f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_591_n N_A_739_297#_c_749_n 0.0251781f $X=6.05 $Y=2 $X2=0 $Y2=0
cc_464 N_VPWR_c_588_n N_X_M1002_d 0.00215201f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_c_588_n N_X_M1020_d 0.00215201f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_466 N_VPWR_c_598_n N_X_c_824_n 0.0189039f $X=6.805 $Y=2.72 $X2=0 $Y2=0
cc_467 N_VPWR_c_588_n N_X_c_824_n 0.0122217f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_468 N_VPWR_M1004_s N_X_c_836_n 0.00338137f $X=6.755 $Y=1.485 $X2=0 $Y2=0
cc_469 N_VPWR_c_592_n N_X_c_836_n 0.0126919f $X=6.89 $Y=2 $X2=0 $Y2=0
cc_470 N_VPWR_c_600_n N_X_c_843_n 0.0189039f $X=7.645 $Y=2.72 $X2=0 $Y2=0
cc_471 N_VPWR_c_588_n N_X_c_843_n 0.0122217f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_472 N_VPWR_M1022_s X 6.44532e-19 $X=7.595 $Y=1.485 $X2=0 $Y2=0
cc_473 N_VPWR_M1022_s X 0.00350209f $X=7.595 $Y=1.485 $X2=0 $Y2=0
cc_474 N_VPWR_c_593_n X 0.020232f $X=7.73 $Y=2 $X2=0 $Y2=0
cc_475 N_A_277_297#_c_699_n N_A_739_297#_c_746_n 0.0261423f $X=3.3 $Y=1.66 $X2=0
+ $Y2=0
cc_476 N_A_277_297#_c_698_n N_A_739_297#_c_747_n 0.0139f $X=3.3 $Y=2.295 $X2=0
+ $Y2=0
cc_477 N_A_277_297#_c_699_n N_A_739_297#_c_747_n 0.0261038f $X=3.3 $Y=1.66 $X2=0
+ $Y2=0
cc_478 N_A_277_297#_c_699_n N_A_739_297#_c_750_n 0.0139f $X=3.3 $Y=1.66 $X2=0
+ $Y2=0
cc_479 N_A_277_297#_c_694_n N_A_27_47#_c_882_n 0.00872848f $X=2.295 $Y=1.567
+ $X2=0 $Y2=0
cc_480 N_A_739_297#_c_749_n N_X_c_820_n 0.00538452f $X=5.53 $Y=1.66 $X2=0 $Y2=0
cc_481 N_A_739_297#_c_749_n N_X_c_824_n 0.00510446f $X=5.53 $Y=1.66 $X2=0 $Y2=0
cc_482 N_X_c_812_n N_VGND_M1021_s 0.00162148f $X=7.145 $Y=0.81 $X2=0 $Y2=0
cc_483 X N_VGND_M1025_s 0.00285834f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_484 N_X_c_812_n N_VGND_c_946_n 0.0122675f $X=7.145 $Y=0.81 $X2=0 $Y2=0
cc_485 X N_VGND_c_947_n 0.0195556f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_486 N_X_c_817_n N_VGND_c_950_n 0.0188551f $X=6.47 $Y=0.38 $X2=0 $Y2=0
cc_487 N_X_c_812_n N_VGND_c_950_n 0.00203746f $X=7.145 $Y=0.81 $X2=0 $Y2=0
cc_488 N_X_c_812_n N_VGND_c_952_n 0.0041083f $X=7.145 $Y=0.81 $X2=0 $Y2=0
cc_489 N_X_c_840_n N_VGND_c_952_n 0.0184921f $X=7.31 $Y=0.38 $X2=0 $Y2=0
cc_490 X N_VGND_c_956_n 0.00367389f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_491 N_X_M1000_d N_VGND_c_957_n 0.00215201f $X=6.335 $Y=0.235 $X2=0 $Y2=0
cc_492 N_X_M1024_d N_VGND_c_957_n 0.00215201f $X=7.175 $Y=0.235 $X2=0 $Y2=0
cc_493 N_X_c_817_n N_VGND_c_957_n 0.0122069f $X=6.47 $Y=0.38 $X2=0 $Y2=0
cc_494 N_X_c_812_n N_VGND_c_957_n 0.0124122f $X=7.145 $Y=0.81 $X2=0 $Y2=0
cc_495 N_X_c_840_n N_VGND_c_957_n 0.012098f $X=7.31 $Y=0.38 $X2=0 $Y2=0
cc_496 X N_VGND_c_957_n 0.00731285f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_497 N_A_27_47#_c_882_n N_VGND_M1012_s 0.00315199f $X=2.715 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_498 N_A_27_47#_c_882_n N_VGND_M1016_s 0.00315199f $X=2.715 $Y=0.76 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_882_n N_VGND_M1014_s 0.00315199f $X=2.715 $Y=0.76 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_886_n N_VGND_c_945_n 0.0124116f $X=5.11 $Y=0.38 $X2=0 $Y2=0
cc_501 N_A_27_47#_c_882_n N_VGND_c_948_n 0.00248431f $X=2.715 $Y=0.76 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_c_885_n N_VGND_c_948_n 0.0172951f $X=2.965 $Y=0.36 $X2=0 $Y2=0
cc_503 N_A_27_47#_c_886_n N_VGND_c_948_n 0.161839f $X=5.11 $Y=0.38 $X2=0 $Y2=0
cc_504 N_A_27_47#_M1027_d N_VGND_c_954_n 0.00119315f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_M1018_d N_VGND_c_954_n 0.00194439f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_M1027_d N_VGND_c_955_n 4.7505e-19 $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_882_n N_VGND_c_955_n 0.109936f $X=2.715 $Y=0.76 $X2=0 $Y2=0
cc_508 N_A_27_47#_M1012_d N_VGND_c_957_n 0.0022756f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_M1017_d N_VGND_c_957_n 0.00228363f $X=2.665 $Y=0.235 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_M1001_s N_VGND_c_957_n 0.00215227f $X=4.105 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_M1005_s N_VGND_c_957_n 0.00239319f $X=4.945 $Y=0.235 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_c_881_n N_VGND_c_957_n 0.00991615f $X=0.26 $Y=0.505 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_c_882_n N_VGND_c_957_n 0.0176107f $X=2.715 $Y=0.76 $X2=0 $Y2=0
cc_514 N_A_27_47#_c_885_n N_VGND_c_957_n 0.00960867f $X=2.965 $Y=0.36 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_c_886_n N_VGND_c_957_n 0.0991252f $X=5.11 $Y=0.38 $X2=0 $Y2=0
cc_516 N_A_27_47#_c_881_n N_VGND_c_958_n 0.0179011f $X=0.26 $Y=0.505 $X2=0 $Y2=0
cc_517 N_A_27_47#_c_882_n N_VGND_c_958_n 0.00248431f $X=2.715 $Y=0.76 $X2=0
+ $Y2=0

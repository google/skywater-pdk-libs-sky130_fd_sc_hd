* File: sky130_fd_sc_hd__lpflow_bleeder_1.pxi.spice
* Created: Thu Aug 27 14:23:07 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%SHORT N_SHORT_c_22_n N_SHORT_M1000_g
+ N_SHORT_c_23_n N_SHORT_M1004_g N_SHORT_c_24_n N_SHORT_M1001_g N_SHORT_c_25_n
+ N_SHORT_M1003_g N_SHORT_c_26_n N_SHORT_M1002_g SHORT N_SHORT_c_27_n
+ N_SHORT_c_28_n PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%SHORT
x_PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%VGND N_VGND_M1000_s N_VGND_c_48_n
+ N_VGND_c_49_n N_VGND_c_50_n VGND N_VGND_c_51_n N_VGND_c_52_n
+ PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%VPWR N_VPWR_M1002_d N_VPWR_c_68_n
+ N_VPWR_c_71_n N_VPWR_c_72_n N_VPWR_c_73_n VPWR N_VPWR_c_69_n
+ PM_SKY130_FD_SC_HD__LPFLOW_BLEEDER_1%VPWR
cc_1 VNB N_SHORT_c_22_n 0.0203602f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.995
cc_2 VNB N_SHORT_c_23_n 0.0150145f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=0.995
cc_3 VNB N_SHORT_c_24_n 0.0150214f $X=-0.19 $Y=-0.24 $X2=1.38 $Y2=0.995
cc_4 VNB N_SHORT_c_25_n 0.0150157f $X=-0.19 $Y=-0.24 $X2=1.74 $Y2=0.995
cc_5 VNB N_SHORT_c_26_n 0.0207836f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=0.995
cc_6 VNB N_SHORT_c_27_n 0.0152784f $X=-0.19 $Y=-0.24 $X2=1.74 $Y2=1.16
cc_7 VNB N_SHORT_c_28_n 0.0773592f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=1.16
cc_8 VNB N_VGND_c_48_n 0.0370138f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=0.705
cc_9 VNB N_VGND_c_49_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=1.38 $Y2=0.705
cc_10 VNB N_VGND_c_50_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=1.74 $Y2=0.995
cc_11 VNB N_VGND_c_51_n 0.0686387f $X=-0.19 $Y=-0.24 $X2=0.72 $Y2=1.16
cc_12 VNB N_VGND_c_52_n 0.226699f $X=-0.19 $Y=-0.24 $X2=0.72 $Y2=1.16
cc_13 VNB N_VPWR_c_68_n 0.0313115f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=0.705
cc_14 VNB N_VPWR_c_69_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.72 $Y2=1.16
cc_15 VPB N_SHORT_c_27_n 0.105444f $X=-0.19 $Y=1.305 $X2=1.74 $Y2=1.16
cc_16 VPB N_SHORT_c_28_n 0.0544707f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=1.16
cc_17 VPB N_VPWR_c_68_n 0.0940676f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=0.705
cc_18 VPB N_VPWR_c_71_n 0.0112126f $X=-0.19 $Y=1.305 $X2=1.38 $Y2=0.705
cc_19 VPB N_VPWR_c_72_n 0.0704015f $X=-0.19 $Y=1.305 $X2=1.38 $Y2=0.705
cc_20 VPB N_VPWR_c_73_n 0.00632158f $X=-0.19 $Y=1.305 $X2=1.74 $Y2=0.995
cc_21 VPB N_VPWR_c_69_n 0.135719f $X=-0.19 $Y=1.305 $X2=0.72 $Y2=1.16
cc_22 N_SHORT_c_22_n N_VGND_c_48_n 0.0120533f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_23 N_SHORT_c_23_n N_VGND_c_48_n 0.00240703f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_24 N_SHORT_c_27_n N_VGND_c_48_n 0.0273074f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_25 N_SHORT_c_22_n N_VGND_c_51_n 0.00376619f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_26 N_SHORT_c_23_n N_VGND_c_51_n 0.00472107f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_27 N_SHORT_c_24_n N_VGND_c_51_n 0.00472107f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_28 N_SHORT_c_25_n N_VGND_c_51_n 0.00472107f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_29 N_SHORT_c_26_n N_VGND_c_51_n 0.00449553f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_30 N_SHORT_c_22_n N_VGND_c_52_n 0.00399306f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_31 N_SHORT_c_23_n N_VGND_c_52_n 0.00495008f $X=1.02 $Y=0.995 $X2=0 $Y2=0
cc_32 N_SHORT_c_24_n N_VGND_c_52_n 0.00495008f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_33 N_SHORT_c_25_n N_VGND_c_52_n 0.00495008f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_34 N_SHORT_c_26_n N_VGND_c_52_n 0.00495008f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_35 N_SHORT_c_25_n N_VPWR_c_68_n 0.00230061f $X=1.74 $Y=0.995 $X2=0 $Y2=0
cc_36 N_SHORT_c_26_n N_VPWR_c_68_n 0.0106307f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_37 N_SHORT_c_27_n N_VPWR_c_68_n 0.0584087f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_38 N_SHORT_c_28_n N_VPWR_c_68_n 0.0144528f $X=2.1 $Y=1.16 $X2=0 $Y2=0
cc_39 N_VGND_c_51_n N_VPWR_c_68_n 0.0072329f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_40 N_VGND_c_52_n N_VPWR_c_68_n 0.0105274f $X=2.53 $Y=0 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__xnor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
M1000 Y a_27_297# a_560_47# VNB nshort w=650000u l=150000u
+  ad=3.38e+11p pd=3.64e+06u as=5.4925e+11p ps=5.59e+06u
M1001 VPWR a_27_297# Y VPB phighvt w=1e+06u l=150000u
+  ad=1.35e+12p pd=1.27e+07u as=5.75e+11p ps=5.15e+06u
M1002 a_474_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=8.1e+11p pd=7.62e+06u as=0p ps=0u
M1003 VPWR B a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=8.25e+11p ps=7.65e+06u
M1004 a_560_47# a_27_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_474_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=5.3625e+11p ps=5.55e+06u
M1008 a_27_47# B a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1009 a_27_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B a_560_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B a_474_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_560_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_560_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_474_297# B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_297# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A a_560_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


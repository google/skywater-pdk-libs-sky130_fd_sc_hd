* File: sky130_fd_sc_hd__o21bai_4.pex.spice
* Created: Tue Sep  1 19:22:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21BAI_4%B1_N 3 6 8 11 12 13
c27 12 0 1.91671e-19 $X=0.39 $Y=1.16
r28 11 14 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.16
+ $X2=0.402 $Y2=1.325
r29 11 13 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.16
+ $X2=0.402 $Y2=0.995
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.39
+ $Y=1.16 $X2=0.39 $Y2=1.16
r31 8 12 8.45022 $w=2.08e-07 $l=1.6e-07 $layer=LI1_cond $X=0.23 $Y=1.18 $X2=0.39
+ $Y2=1.18
r32 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.52 $Y=1.985
+ $X2=0.52 $Y2=1.325
r33 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.56 $X2=0.52
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%A_33_297# 1 2 9 13 15 17 20 22 24 27 29 31
+ 32 34 35 37 39 43 46 48 54 59 60 71
c95 71 0 2.68957e-19 $X=2.72 $Y=1.16
c96 48 0 1.77925e-19 $X=0.81 $Y=1.455
c97 32 0 1.56657e-19 $X=2.72 $Y=0.995
r98 70 71 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.3 $Y=1.16 $X2=2.72
+ $Y2=1.16
r99 69 70 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.2 $Y=1.16 $X2=2.3
+ $Y2=1.16
r100 66 67 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.78 $Y=1.16 $X2=1.88
+ $Y2=1.16
r101 65 66 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=1.16
+ $X2=1.78 $Y2=1.16
r102 64 65 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.36 $Y=1.16 $X2=1.46
+ $Y2=1.16
r103 55 69 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.05 $Y=1.16
+ $X2=2.2 $Y2=1.16
r104 55 67 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.05 $Y=1.16
+ $X2=1.88 $Y2=1.16
r105 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.05
+ $Y=1.16 $X2=2.05 $Y2=1.16
r106 52 64 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.03 $Y=1.16
+ $X2=1.36 $Y2=1.16
r107 52 61 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.03 $Y=1.16 $X2=0.94
+ $Y2=1.16
r108 51 54 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=1.03 $Y=1.18
+ $X2=2.05 $Y2=1.18
r109 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.16 $X2=1.03 $Y2=1.16
r110 49 60 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=1.18
+ $X2=0.81 $Y2=1.18
r111 49 51 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.895 $Y=1.18
+ $X2=1.03 $Y2=1.18
r112 47 60 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.81 $Y=1.285
+ $X2=0.81 $Y2=1.18
r113 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.81 $Y=1.285
+ $X2=0.81 $Y2=1.455
r114 46 60 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.81 $Y=1.075
+ $X2=0.81 $Y2=1.18
r115 46 59 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.81 $Y=1.075
+ $X2=0.81 $Y2=0.895
r116 41 59 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0.73
+ $X2=0.73 $Y2=0.895
r117 41 43 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.73 $Y=0.73
+ $X2=0.73 $Y2=0.39
r118 40 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=1.54
+ $X2=0.31 $Y2=1.54
r119 39 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.725 $Y=1.54
+ $X2=0.81 $Y2=1.455
r120 39 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.725 $Y=1.54
+ $X2=0.475 $Y2=1.54
r121 35 58 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.625
+ $X2=0.31 $Y2=1.54
r122 35 37 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.31 $Y=1.625
+ $X2=0.31 $Y2=2.3
r123 32 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=0.995
+ $X2=2.72 $Y2=1.16
r124 32 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.72 $Y=0.995
+ $X2=2.72 $Y2=0.56
r125 29 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=0.995
+ $X2=2.3 $Y2=1.16
r126 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.3 $Y=0.995
+ $X2=2.3 $Y2=0.56
r127 25 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.325
+ $X2=2.2 $Y2=1.16
r128 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.2 $Y=1.325
+ $X2=2.2 $Y2=1.985
r129 22 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.16
r130 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=0.56
r131 18 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.16
r132 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.985
r133 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.16
r134 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r135 11 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.16
r136 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.985
r137 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.325
+ $X2=0.94 $Y2=1.16
r138 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.94 $Y=1.325
+ $X2=0.94 $Y2=1.985
r139 2 58 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.485 $X2=0.31 $Y2=1.62
r140 2 37 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.485 $X2=0.31 $Y2=2.3
r141 1 43 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r85 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.25 $Y=1.16 $X2=4.4
+ $Y2=1.16
r86 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.25
+ $Y=1.16 $X2=4.25 $Y2=1.16
r87 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.98 $Y=1.16
+ $X2=4.25 $Y2=1.16
r88 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.56 $Y=1.16
+ $X2=3.98 $Y2=1.16
r89 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.23 $Y=1.16
+ $X2=3.56 $Y2=1.16
r90 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.23
+ $Y=1.16 $X2=3.23 $Y2=1.16
r91 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.14 $Y=1.16 $X2=3.23
+ $Y2=1.16
r92 29 40 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=4.25 $Y2=1.175
r93 29 35 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.23 $Y2=1.175
r94 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=1.325
+ $X2=4.4 $Y2=1.16
r95 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.4 $Y=1.325 $X2=4.4
+ $Y2=1.985
r96 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=0.995
+ $X2=4.4 $Y2=1.16
r97 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.4 $Y=0.995 $X2=4.4
+ $Y2=0.56
r98 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.325
+ $X2=3.98 $Y2=1.16
r99 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.98 $Y=1.325
+ $X2=3.98 $Y2=1.985
r100 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=1.16
r101 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=0.56
r102 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.325
+ $X2=3.56 $Y2=1.16
r103 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.56 $Y=1.325
+ $X2=3.56 $Y2=1.985
r104 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=0.995
+ $X2=3.56 $Y2=1.16
r105 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.56 $Y=0.995
+ $X2=3.56 $Y2=0.56
r106 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.325
+ $X2=3.14 $Y2=1.16
r107 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.14 $Y=1.325
+ $X2=3.14 $Y2=1.985
r108 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=0.995
+ $X2=3.14 $Y2=1.16
r109 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.14 $Y=0.995
+ $X2=3.14 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 31 32 33
+ 48
r79 46 48 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.9 $Y=1.16 $X2=6.08
+ $Y2=1.16
r80 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.9 $Y=1.16
+ $X2=5.9 $Y2=1.16
r81 44 46 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=5.66 $Y=1.16 $X2=5.9
+ $Y2=1.16
r82 43 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.24 $Y=1.16
+ $X2=5.66 $Y2=1.16
r83 41 43 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.88 $Y=1.16
+ $X2=5.24 $Y2=1.16
r84 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.88
+ $Y=1.16 $X2=4.88 $Y2=1.16
r85 38 41 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.82 $Y=1.16 $X2=4.88
+ $Y2=1.16
r86 32 33 13.6618 $w=3.78e-07 $l=3.75e-07 $layer=LI1_cond $X=6.21 $Y=1.18
+ $X2=6.585 $Y2=1.18
r87 32 47 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=6.21 $Y=1.18 $X2=5.9
+ $Y2=1.18
r88 31 47 32.2164 $w=2.08e-07 $l=6.1e-07 $layer=LI1_cond $X=5.29 $Y=1.18 $X2=5.9
+ $Y2=1.18
r89 31 42 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=5.29 $Y=1.18
+ $X2=4.88 $Y2=1.18
r90 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.08 $Y=1.325
+ $X2=6.08 $Y2=1.16
r91 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.08 $Y=1.325
+ $X2=6.08 $Y2=1.985
r92 22 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.08 $Y=0.995
+ $X2=6.08 $Y2=1.16
r93 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.08 $Y=0.995
+ $X2=6.08 $Y2=0.56
r94 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.66 $Y=1.325
+ $X2=5.66 $Y2=1.16
r95 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.66 $Y=1.325
+ $X2=5.66 $Y2=1.985
r96 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.66 $Y=0.995
+ $X2=5.66 $Y2=1.16
r97 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.66 $Y=0.995
+ $X2=5.66 $Y2=0.56
r98 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.325
+ $X2=5.24 $Y2=1.16
r99 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.24 $Y=1.325
+ $X2=5.24 $Y2=1.985
r100 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.16
r101 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r102 4 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.82 $Y=1.325
+ $X2=4.82 $Y2=1.16
r103 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.82 $Y=1.325
+ $X2=4.82 $Y2=1.985
r104 1 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=1.16
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%VPWR 1 2 3 4 5 20 24 28 32 34 38 40 41 42
+ 44 49 60 61 64 67 70 73
r98 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r99 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r100 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r101 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r102 61 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r103 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r104 58 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.995 $Y=2.72
+ $X2=5.87 $Y2=2.72
r105 58 60 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.995 $Y=2.72
+ $X2=6.67 $Y2=2.72
r106 57 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r107 57 71 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=2.53 $Y2=2.72
r108 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r109 54 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.535 $Y=2.72
+ $X2=2.41 $Y2=2.72
r110 54 56 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=2.535 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 53 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 53 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r114 50 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.695 $Y=2.72
+ $X2=1.57 $Y2=2.72
r115 50 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.695 $Y=2.72
+ $X2=2.07 $Y2=2.72
r116 49 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.41 $Y2=2.72
r117 49 52 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.07 $Y2=2.72
r118 48 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r119 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r121 45 64 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.75 $Y2=2.72
r122 45 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r123 44 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.57 $Y2=2.72
r124 44 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 42 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r126 40 56 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.905 $Y=2.72
+ $X2=4.83 $Y2=2.72
r127 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=2.72
+ $X2=5.03 $Y2=2.72
r128 36 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=2.635
+ $X2=5.87 $Y2=2.72
r129 36 38 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.87 $Y=2.635
+ $X2=5.87 $Y2=1.96
r130 35 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=2.72
+ $X2=5.03 $Y2=2.72
r131 34 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.745 $Y=2.72
+ $X2=5.87 $Y2=2.72
r132 34 35 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.745 $Y=2.72
+ $X2=5.155 $Y2=2.72
r133 30 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=2.635
+ $X2=5.03 $Y2=2.72
r134 30 32 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.03 $Y=2.635
+ $X2=5.03 $Y2=1.96
r135 26 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=2.635
+ $X2=2.41 $Y2=2.72
r136 26 28 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.41 $Y=2.635
+ $X2=2.41 $Y2=1.96
r137 22 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.635
+ $X2=1.57 $Y2=2.72
r138 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.57 $Y=2.635
+ $X2=1.57 $Y2=1.96
r139 18 64 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r140 18 20 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r141 5 38 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.735
+ $Y=1.485 $X2=5.87 $Y2=1.96
r142 4 32 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.485 $X2=5.03 $Y2=1.96
r143 3 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.485 $X2=2.41 $Y2=1.96
r144 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.435
+ $Y=1.485 $X2=1.57 $Y2=1.96
r145 1 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%Y 1 2 3 4 5 6 19 21 23 25 31 33 35 39 47 51
+ 53 54 60
r85 62 63 0.132898 $w=4.48e-07 $l=5e-09 $layer=LI1_cond $X=2.67 $Y=1.535
+ $X2=2.67 $Y2=1.54
r86 54 63 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=2.445 $Y=1.54
+ $X2=2.67 $Y2=1.54
r87 54 62 0.132898 $w=4.48e-07 $l=5e-09 $layer=LI1_cond $X=2.67 $Y=1.53 $X2=2.67
+ $Y2=1.535
r88 54 60 14.9447 $w=4.48e-07 $l=4.55e-07 $layer=LI1_cond $X=2.67 $Y=1.53
+ $X2=2.67 $Y2=1.075
r89 45 54 12.918 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.115 $Y=1.54
+ $X2=2.445 $Y2=1.54
r90 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.115 $Y=1.54
+ $X2=1.99 $Y2=1.54
r91 40 51 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=1.535
+ $X2=3.35 $Y2=1.535
r92 39 53 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.065 $Y=1.535
+ $X2=4.19 $Y2=1.535
r93 39 40 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=4.065 $Y=1.535
+ $X2=3.475 $Y2=1.535
r94 36 62 6.14847 $w=1.8e-07 $l=2.25e-07 $layer=LI1_cond $X=2.895 $Y=1.535
+ $X2=2.67 $Y2=1.535
r95 35 51 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=1.535
+ $X2=3.35 $Y2=1.535
r96 35 36 20.3333 $w=1.78e-07 $l=3.3e-07 $layer=LI1_cond $X=3.225 $Y=1.535
+ $X2=2.895 $Y2=1.535
r97 33 49 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.815 $X2=2.56
+ $Y2=0.73
r98 33 60 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.56 $Y=0.815
+ $X2=2.56 $Y2=1.075
r99 29 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=1.625
+ $X2=1.99 $Y2=1.54
r100 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.99 $Y=1.625
+ $X2=1.99 $Y2=2.3
r101 25 49 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.445 $Y=0.73
+ $X2=2.56 $Y2=0.73
r102 25 27 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.445 $Y=0.73
+ $X2=1.67 $Y2=0.73
r103 24 44 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.275 $Y=1.54
+ $X2=1.17 $Y2=1.54
r104 23 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.865 $Y=1.54
+ $X2=1.99 $Y2=1.54
r105 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.865 $Y=1.54
+ $X2=1.275 $Y2=1.54
r106 19 44 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=1.625
+ $X2=1.17 $Y2=1.54
r107 19 21 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=1.17 $Y=1.625
+ $X2=1.17 $Y2=2.3
r108 6 53 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.055
+ $Y=1.485 $X2=4.19 $Y2=1.62
r109 5 51 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.215
+ $Y=1.485 $X2=3.35 $Y2=1.62
r110 4 47 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.485 $X2=1.99 $Y2=1.62
r111 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.485 $X2=1.99 $Y2=2.3
r112 3 44 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.485 $X2=1.15 $Y2=1.62
r113 3 21 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.485 $X2=1.15 $Y2=2.3
r114 2 49 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.235 $X2=2.51 $Y2=0.73
r115 1 27 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%A_561_297# 1 2 3 4 5 18 20 21 24 26 28 29
+ 30 34 36 38 40 42 48
c65 18 0 7.72863e-20 $X=2.93 $Y=1.96
r66 38 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.29 $Y=1.625
+ $X2=6.29 $Y2=1.54
r67 38 40 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.29 $Y=1.625
+ $X2=6.29 $Y2=2.3
r68 37 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.575 $Y=1.54
+ $X2=5.45 $Y2=1.54
r69 36 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.165 $Y=1.54
+ $X2=6.29 $Y2=1.54
r70 36 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.165 $Y=1.54
+ $X2=5.575 $Y2=1.54
r71 32 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=1.625
+ $X2=5.45 $Y2=1.54
r72 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.45 $Y=1.625
+ $X2=5.45 $Y2=2.3
r73 31 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.735 $Y=1.54
+ $X2=4.61 $Y2=1.54
r74 30 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.325 $Y=1.54
+ $X2=5.45 $Y2=1.54
r75 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.325 $Y=1.54
+ $X2=4.735 $Y2=1.54
r76 29 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=2.295
+ $X2=4.61 $Y2=2.38
r77 28 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=1.625
+ $X2=4.61 $Y2=1.54
r78 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.61 $Y=1.625
+ $X2=4.61 $Y2=2.295
r79 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=2.38
+ $X2=3.77 $Y2=2.38
r80 26 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.485 $Y=2.38
+ $X2=4.61 $Y2=2.38
r81 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.485 $Y=2.38
+ $X2=3.895 $Y2=2.38
r82 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.295
+ $X2=3.77 $Y2=2.38
r83 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.77 $Y=2.295
+ $X2=3.77 $Y2=1.96
r84 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.645 $Y=2.38
+ $X2=3.77 $Y2=2.38
r85 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.645 $Y=2.38
+ $X2=3.055 $Y2=2.38
r86 16 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.915 $Y=2.295
+ $X2=3.055 $Y2=2.38
r87 16 18 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.915 $Y=2.295
+ $X2=2.915 $Y2=1.96
r88 5 50 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.155
+ $Y=1.485 $X2=6.29 $Y2=1.62
r89 5 40 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.155
+ $Y=1.485 $X2=6.29 $Y2=2.3
r90 4 48 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.485 $X2=5.45 $Y2=1.62
r91 4 34 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.485 $X2=5.45 $Y2=2.3
r92 3 46 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.61 $Y2=2.3
r93 3 44 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.61 $Y2=1.62
r94 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.635
+ $Y=1.485 $X2=3.77 $Y2=1.96
r95 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=2.93 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40
+ 41 43 44 46 47 48 67 68
r98 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r99 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r100 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r101 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r102 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r103 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r104 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r105 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r106 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r107 53 56 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.99
+ $Y2=0
r108 52 55 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.99
+ $Y2=0
r109 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r110 50 71 3.40825 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r111 50 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r112 48 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r113 48 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r114 46 64 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.785 $Y=0 $X2=5.75
+ $Y2=0
r115 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=0 $X2=5.87
+ $Y2=0
r116 45 67 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=5.955 $Y=0
+ $X2=6.67 $Y2=0
r117 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=0 $X2=5.87
+ $Y2=0
r118 43 61 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.945 $Y=0
+ $X2=4.83 $Y2=0
r119 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.03
+ $Y2=0
r120 42 64 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.115 $Y=0
+ $X2=5.75 $Y2=0
r121 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0 $X2=5.03
+ $Y2=0
r122 40 58 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.105 $Y=0
+ $X2=3.91 $Y2=0
r123 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.19
+ $Y2=0
r124 39 61 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.83 $Y2=0
r125 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.275 $Y=0 $X2=4.19
+ $Y2=0
r126 37 55 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=0
+ $X2=2.99 $Y2=0
r127 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.35
+ $Y2=0
r128 36 58 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.435 $Y=0
+ $X2=3.91 $Y2=0
r129 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.35
+ $Y2=0
r130 32 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=0.085
+ $X2=5.87 $Y2=0
r131 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.87 $Y=0.085
+ $X2=5.87 $Y2=0.39
r132 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r133 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.39
r134 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0
r135 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0.39
r136 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r137 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.39
r138 16 71 3.40825 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.197 $Y2=0
r139 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.31 $Y2=0.39
r140 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.735
+ $Y=0.235 $X2=5.87 $Y2=0.39
r141 4 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.895
+ $Y=0.235 $X2=5.03 $Y2=0.39
r142 3 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.055
+ $Y=0.235 $X2=4.19 $Y2=0.39
r143 2 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.235 $X2=3.35 $Y2=0.39
r144 1 18 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.31 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_4%A_225_47# 1 2 3 4 5 6 7 22 28 29 30 34 36
+ 40 42 46 48 52 58 59 60
c112 29 0 1.56657e-19 $X=2.97 $Y=0.725
r113 50 52 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.29 $Y=0.725
+ $X2=6.29 $Y2=0.39
r114 49 60 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.615 $Y=0.815
+ $X2=5.45 $Y2=0.815
r115 48 50 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.125 $Y=0.815
+ $X2=6.29 $Y2=0.725
r116 48 49 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.125 $Y=0.815
+ $X2=5.615 $Y2=0.815
r117 44 60 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.45 $Y=0.725
+ $X2=5.45 $Y2=0.815
r118 44 46 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.45 $Y=0.725
+ $X2=5.45 $Y2=0.39
r119 43 59 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.775 $Y=0.815
+ $X2=4.61 $Y2=0.815
r120 42 60 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=0.815
+ $X2=5.45 $Y2=0.815
r121 42 43 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.285 $Y=0.815
+ $X2=4.775 $Y2=0.815
r122 38 59 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.61 $Y=0.725
+ $X2=4.61 $Y2=0.815
r123 38 40 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.61 $Y=0.725
+ $X2=4.61 $Y2=0.39
r124 37 58 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=0.815
+ $X2=3.77 $Y2=0.815
r125 36 59 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0.815
+ $X2=4.61 $Y2=0.815
r126 36 37 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.445 $Y=0.815
+ $X2=3.935 $Y2=0.815
r127 32 58 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.77 $Y2=0.815
r128 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.77 $Y2=0.39
r129 31 57 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0.815
+ $X2=2.97 $Y2=0.815
r130 30 58 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=0.815
+ $X2=3.77 $Y2=0.815
r131 30 31 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.605 $Y=0.815
+ $X2=3.095 $Y2=0.815
r132 29 57 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.97 $Y=0.725 $X2=2.97
+ $Y2=0.815
r133 28 55 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=0.475
+ $X2=2.97 $Y2=0.39
r134 28 29 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.97 $Y=0.475
+ $X2=2.97 $Y2=0.725
r135 24 27 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.25 $Y=0.39
+ $X2=2.09 $Y2=0.39
r136 22 55 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=0.39
+ $X2=2.97 $Y2=0.39
r137 22 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.845 $Y=0.39
+ $X2=2.09 $Y2=0.39
r138 7 52 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.155
+ $Y=0.235 $X2=6.29 $Y2=0.39
r139 6 46 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.315
+ $Y=0.235 $X2=5.45 $Y2=0.39
r140 5 40 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.475
+ $Y=0.235 $X2=4.61 $Y2=0.39
r141 4 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.635
+ $Y=0.235 $X2=3.77 $Y2=0.39
r142 3 57 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.93 $Y2=0.73
r143 3 55 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.93 $Y2=0.39
r144 2 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.09 $Y2=0.39
r145 1 24 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.39
.ends


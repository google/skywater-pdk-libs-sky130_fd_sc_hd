* File: sky130_fd_sc_hd__o2bb2ai_1.spice
* Created: Tue Sep  1 19:24:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2bb2ai_1.pex.spice"
.subckt sky130_fd_sc_hd__o2bb2ai_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1008 A_112_47# N_A1_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.17875 PD=0.86 PS=1.85 NRD=9.228 NRS=1.836 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_A_112_297#_M1006_d N_A2_N_M1006_g A_112_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.2405 AS=0.06825 PD=2.04 PS=0.86 NRD=19.38 NRS=9.228 M=1 R=4.33333
+ SA=75000.6 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1000 N_A_394_47#_M1000_d N_A_112_297#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B2_M1003_g N_A_394_47#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1001 N_A_394_47#_M1001_d N_B1_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_112_297#_M1004_d N_A1_N_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A2_N_M1009_g N_A_112_297#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.42 AS=0.135 PD=1.84 PS=1.27 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_A_112_297#_M1007_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.42 PD=1.27 PS=1.84 NRD=0 NRS=14.7553 M=1 R=6.66667 SA=75001.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1005 A_478_297# N_B2_M1005_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g A_478_297# VPB PHIGHVT L=0.15 W=1 AD=0.275
+ AS=0.135 PD=2.55 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75002.4 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o2bb2ai_1.pxi.spice"
*
.ends
*
*

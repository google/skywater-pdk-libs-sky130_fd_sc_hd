* File: sky130_fd_sc_hd__decap_12.spice.pex
* Created: Thu Aug 27 14:13:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DECAP_12%VGND 1 9 10 11 12 14 22 34 37
r26 36 37 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r27 34 36 0.448529 $w=8.16e-07 $l=3e-08 $layer=LI1_cond $X=5.26 $Y=0.385
+ $X2=5.29 $Y2=0.385
r28 31 37 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=5.29
+ $Y2=0
r29 30 31 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r30 24 27 0.25811 $w=1.418e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.645
+ $X2=0.26 $Y2=0.645
r31 21 30 15.4006 $w=1.418e-06 $l=1.79e-06 $layer=LI1_cond $X=2.48 $Y=0.645
+ $X2=0.69 $Y2=0.645
r32 20 22 8.47369 $w=1.49e-06 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.87
+ $X2=2.645 $Y2=1.87
r33 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.48
+ $Y=1.29 $X2=2.48 $Y2=1.29
r34 17 30 1.11848 $w=1.418e-06 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=0.645
+ $X2=0.69 $Y2=0.645
r35 17 27 2.5811 $w=1.418e-06 $l=3e-07 $layer=LI1_cond $X=0.56 $Y=0.645 $X2=0.26
+ $Y2=0.645
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.56
+ $Y=1.29 $X2=0.56 $Y2=1.29
r37 14 20 19.2327 $w=1.49e-06 $l=5.8e-07 $layer=POLY_cond $X=1.9 $Y=1.87
+ $X2=2.48 $Y2=1.87
r38 14 16 44.4343 $w=1.49e-06 $l=1.34e-06 $layer=POLY_cond $X=1.9 $Y=1.87
+ $X2=0.56 $Y2=1.87
r39 12 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r40 12 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r41 11 21 2.97997 $w=1.418e-06 $l=3.40147e-07 $layer=LI1_cond $X=2.665 $Y=0.385
+ $X2=2.48 $Y2=0.645
r42 10 34 4.13877 $w=9.4e-07 $l=3e-07 $layer=LI1_cond $X=4.96 $Y=0.385 $X2=5.26
+ $Y2=0.385
r43 10 11 29.7862 $w=9.38e-07 $l=2.295e-06 $layer=LI1_cond $X=4.96 $Y=0.385
+ $X2=2.665 $Y2=0.385
r44 9 22 4.90531 $w=1.13e-06 $l=1.15e-07 $layer=POLY_cond $X=2.76 $Y=2.05
+ $X2=2.645 $Y2=2.05
r45 1 34 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=5.125 $Y=0.235
+ $X2=5.26 $Y2=0.475
r46 1 27 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__DECAP_12%VPWR 1 9 10 11 12 17 19 30 33
r25 32 33 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r26 30 32 0.212051 $w=1.726e-06 $l=3e-08 $layer=LI1_cond $X=5.26 $Y=1.915
+ $X2=5.29 $Y2=1.915
r27 23 26 0.323894 $w=1.13e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.175
+ $X2=0.26 $Y2=2.175
r28 20 30 2.26188 $w=1.726e-06 $l=3.2e-07 $layer=LI1_cond $X=4.94 $Y=1.915
+ $X2=5.26 $Y2=1.915
r29 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.94
+ $Y=1.11 $X2=4.94 $Y2=1.11
r30 16 20 13.5713 $w=1.726e-06 $l=1.92e-06 $layer=LI1_cond $X=3.02 $Y=1.915
+ $X2=4.94 $Y2=1.915
r31 15 19 84.3769 $w=1.17e-06 $l=1.92e-06 $layer=POLY_cond $X=3.02 $Y=0.69
+ $X2=4.94 $Y2=0.69
r32 15 17 12.167 $w=1.17e-06 $l=1.65e-07 $layer=POLY_cond $X=3.02 $Y=0.69
+ $X2=2.855 $Y2=0.69
r33 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.02
+ $Y=1.11 $X2=3.02 $Y2=1.11
r34 12 33 1.43978 $w=4.8e-07 $l=5.06e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=5.29 $Y2=2.72
r35 12 23 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r36 11 26 4.56277 $w=1.26e-06 $l=4.55e-07 $layer=LI1_cond $X=0.715 $Y=2.175
+ $X2=0.26 $Y2=2.175
r37 10 16 2.21943 $w=1.726e-06 $l=3.40147e-07 $layer=LI1_cond $X=2.835 $Y=2.175
+ $X2=3.02 $Y2=1.915
r38 10 11 20.527 $w=1.258e-06 $l=2.12e-06 $layer=LI1_cond $X=2.835 $Y=2.175
+ $X2=0.715 $Y2=2.175
r39 9 17 5.65309 $w=8.1e-07 $l=9.5e-08 $layer=POLY_cond $X=2.76 $Y=0.51
+ $X2=2.855 $Y2=0.51
r40 1 30 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.615 $X2=5.26 $Y2=1.83
r41 1 26 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends


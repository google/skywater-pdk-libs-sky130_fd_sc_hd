* File: sky130_fd_sc_hd__o221a_1.spice
* Created: Thu Aug 27 14:36:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o221a_1.spice.pex"
.subckt sky130_fd_sc_hd__o221a_1  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1011 N_A_149_47#_M1011_d N_C1_M1011_g N_A_51_297#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.099125 AS=0.2015 PD=0.955 PS=1.92 NRD=4.608 NRS=8.304 M=1
+ R=4.33333 SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_A_240_47#_M1007_d N_B1_M1007_g N_A_149_47#_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.099125 PD=0.92 PS=0.955 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_A_149_47#_M1006_d N_B2_M1006_g N_A_240_47#_M1007_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_240_47#_M1002_d N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_240_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_51_297#_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VPWR_M1009_d N_C1_M1009_g N_A_51_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.34 PD=1.33 PS=2.68 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75000.3
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1005 A_245_297# N_B1_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.165 PD=1.21 PS=1.33 NRD=9.8303 NRS=6.8753 M=1 R=6.66667 SA=75000.7
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1001 N_A_51_297#_M1001_d N_B2_M1001_g A_245_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.4125 AS=0.105 PD=1.825 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.1
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1010 A_512_297# N_A2_M1010_g N_A_51_297#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.4125 PD=1.21 PS=1.825 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75002.1
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_512_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.105 PD=1.33 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.4 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1008 N_X_M1008_d N_A_51_297#_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.165 PD=2.56 PS=1.33 NRD=2.9353 NRS=10.8153 M=1 R=6.66667
+ SA=75002.9 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_37 VNB 0 1.22672e-19 $X=0.145 $Y=-0.085
c_70 VPB 0 1.40821e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__o221a_1.spice.SKY130_FD_SC_HD__O221A_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__dfbbn_1.pxi.spice
* Created: Thu Aug 27 14:13:59 2020
* 
x_PM_SKY130_FD_SC_HD__DFBBN_1%CLK_N N_CLK_N_c_262_n N_CLK_N_c_257_n
+ N_CLK_N_M1033_g N_CLK_N_c_263_n N_CLK_N_M1011_g N_CLK_N_c_258_n
+ N_CLK_N_c_264_n CLK_N CLK_N N_CLK_N_c_260_n N_CLK_N_c_261_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%CLK_N
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_27_47# N_A_27_47#_M1033_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1013_g N_A_27_47#_M1000_g N_A_27_47#_M1021_g N_A_27_47#_c_303_n
+ N_A_27_47#_c_304_n N_A_27_47#_M1038_g N_A_27_47#_c_306_n N_A_27_47#_c_307_n
+ N_A_27_47#_M1001_g N_A_27_47#_M1022_g N_A_27_47#_c_550_p N_A_27_47#_c_308_n
+ N_A_27_47#_c_309_n N_A_27_47#_c_329_n N_A_27_47#_c_310_n N_A_27_47#_c_311_n
+ N_A_27_47#_c_330_n N_A_27_47#_c_331_n N_A_27_47#_c_332_n N_A_27_47#_c_312_n
+ N_A_27_47#_c_313_n N_A_27_47#_c_314_n N_A_27_47#_c_315_n N_A_27_47#_c_316_n
+ N_A_27_47#_c_317_n N_A_27_47#_c_318_n N_A_27_47#_c_319_n N_A_27_47#_c_320_n
+ N_A_27_47#_c_321_n N_A_27_47#_c_322_n N_A_27_47#_c_323_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DFBBN_1%D N_D_M1002_g N_D_M1017_g D D N_D_c_565_n
+ N_D_c_566_n PM_SKY130_FD_SC_HD__DFBBN_1%D
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_193_47# N_A_193_47#_M1013_d N_A_193_47#_M1000_d
+ N_A_193_47#_c_605_n N_A_193_47#_M1026_g N_A_193_47#_M1014_g
+ N_A_193_47#_M1034_g N_A_193_47#_c_606_n N_A_193_47#_c_607_n
+ N_A_193_47#_M1036_g N_A_193_47#_c_609_n N_A_193_47#_c_610_n
+ N_A_193_47#_c_617_n N_A_193_47#_c_618_n N_A_193_47#_c_619_n
+ N_A_193_47#_c_620_n N_A_193_47#_c_621_n N_A_193_47#_c_622_n
+ N_A_193_47#_c_623_n N_A_193_47#_c_624_n N_A_193_47#_c_625_n
+ N_A_193_47#_c_626_n N_A_193_47#_c_611_n PM_SKY130_FD_SC_HD__DFBBN_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_647_21# N_A_647_21#_M1035_d N_A_647_21#_M1004_d
+ N_A_647_21#_M1007_g N_A_647_21#_M1023_g N_A_647_21#_M1028_g
+ N_A_647_21#_c_808_n N_A_647_21#_M1019_g N_A_647_21#_c_817_n
+ N_A_647_21#_c_864_p N_A_647_21#_c_832_n N_A_647_21#_c_809_n
+ N_A_647_21#_c_810_n N_A_647_21#_c_811_n N_A_647_21#_c_819_n
+ N_A_647_21#_c_820_n N_A_647_21#_c_837_n N_A_647_21#_c_812_n
+ N_A_647_21#_c_813_n PM_SKY130_FD_SC_HD__DFBBN_1%A_647_21#
x_PM_SKY130_FD_SC_HD__DFBBN_1%SET_B N_SET_B_c_954_n N_SET_B_M1004_g
+ N_SET_B_M1016_g N_SET_B_M1009_g N_SET_B_c_958_n N_SET_B_M1012_g SET_B
+ N_SET_B_c_961_n N_SET_B_c_962_n N_SET_B_c_963_n N_SET_B_c_964_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%SET_B
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_473_413# N_A_473_413#_M1026_d
+ N_A_473_413#_M1021_d N_A_473_413#_M1035_g N_A_473_413#_M1024_g
+ N_A_473_413#_c_1097_n N_A_473_413#_c_1098_n N_A_473_413#_c_1092_n
+ N_A_473_413#_c_1087_n N_A_473_413#_c_1088_n N_A_473_413#_c_1089_n
+ N_A_473_413#_c_1090_n PM_SKY130_FD_SC_HD__DFBBN_1%A_473_413#
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_941_21# N_A_941_21#_M1015_s N_A_941_21#_M1029_s
+ N_A_941_21#_M1031_g N_A_941_21#_M1018_g N_A_941_21#_M1005_g
+ N_A_941_21#_M1032_g N_A_941_21#_c_1193_n N_A_941_21#_c_1194_n
+ N_A_941_21#_c_1204_n N_A_941_21#_c_1205_n N_A_941_21#_c_1195_n
+ N_A_941_21#_c_1196_n N_A_941_21#_c_1197_n N_A_941_21#_c_1198_n
+ N_A_941_21#_c_1199_n N_A_941_21#_c_1208_n N_A_941_21#_c_1209_n
+ N_A_941_21#_c_1210_n N_A_941_21#_c_1211_n N_A_941_21#_c_1200_n
+ N_A_941_21#_c_1201_n PM_SKY130_FD_SC_HD__DFBBN_1%A_941_21#
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_1415_315# N_A_1415_315#_M1025_d
+ N_A_1415_315#_M1012_d N_A_1415_315#_M1008_g N_A_1415_315#_M1020_g
+ N_A_1415_315#_c_1360_n N_A_1415_315#_M1030_g N_A_1415_315#_M1039_g
+ N_A_1415_315#_c_1361_n N_A_1415_315#_c_1362_n N_A_1415_315#_c_1363_n
+ N_A_1415_315#_c_1364_n N_A_1415_315#_c_1365_n N_A_1415_315#_M1010_g
+ N_A_1415_315#_c_1375_n N_A_1415_315#_M1006_g N_A_1415_315#_c_1366_n
+ N_A_1415_315#_c_1367_n N_A_1415_315#_c_1376_n N_A_1415_315#_c_1377_n
+ N_A_1415_315#_c_1378_n N_A_1415_315#_c_1379_n N_A_1415_315#_c_1380_n
+ N_A_1415_315#_c_1492_p N_A_1415_315#_c_1408_n N_A_1415_315#_c_1368_n
+ N_A_1415_315#_c_1382_n N_A_1415_315#_c_1383_n N_A_1415_315#_c_1384_n
+ N_A_1415_315#_c_1401_n N_A_1415_315#_c_1431_n N_A_1415_315#_c_1369_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%A_1415_315#
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_1256_413# N_A_1256_413#_M1001_d
+ N_A_1256_413#_M1034_d N_A_1256_413#_M1025_g N_A_1256_413#_M1003_g
+ N_A_1256_413#_c_1566_n N_A_1256_413#_c_1569_n N_A_1256_413#_c_1555_n
+ N_A_1256_413#_c_1561_n N_A_1256_413#_c_1556_n N_A_1256_413#_c_1557_n
+ N_A_1256_413#_c_1558_n N_A_1256_413#_c_1559_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%A_1256_413#
x_PM_SKY130_FD_SC_HD__DFBBN_1%RESET_B N_RESET_B_M1029_g N_RESET_B_M1015_g
+ RESET_B N_RESET_B_c_1668_n PM_SKY130_FD_SC_HD__DFBBN_1%RESET_B
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_2136_47# N_A_2136_47#_M1010_s
+ N_A_2136_47#_M1006_s N_A_2136_47#_M1027_g N_A_2136_47#_M1037_g
+ N_A_2136_47#_c_1705_n N_A_2136_47#_c_1711_n N_A_2136_47#_c_1706_n
+ N_A_2136_47#_c_1707_n N_A_2136_47#_c_1708_n N_A_2136_47#_c_1709_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%A_2136_47#
x_PM_SKY130_FD_SC_HD__DFBBN_1%VPWR N_VPWR_M1011_d N_VPWR_M1017_s N_VPWR_M1023_d
+ N_VPWR_M1018_d N_VPWR_M1008_d N_VPWR_M1005_d N_VPWR_M1029_d N_VPWR_M1006_d
+ N_VPWR_c_1760_n N_VPWR_c_1761_n N_VPWR_c_1762_n N_VPWR_c_1763_n
+ N_VPWR_c_1764_n N_VPWR_c_1765_n N_VPWR_c_1766_n N_VPWR_c_1767_n
+ N_VPWR_c_1768_n VPWR VPWR N_VPWR_c_1769_n N_VPWR_c_1770_n N_VPWR_c_1771_n
+ N_VPWR_c_1772_n N_VPWR_c_1773_n N_VPWR_c_1774_n N_VPWR_c_1775_n
+ N_VPWR_c_1759_n N_VPWR_c_1777_n N_VPWR_c_1778_n N_VPWR_c_1779_n
+ N_VPWR_c_1780_n N_VPWR_c_1781_n N_VPWR_c_1782_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%VPWR
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_381_47# N_A_381_47#_M1002_d N_A_381_47#_M1017_d
+ N_A_381_47#_c_1943_n N_A_381_47#_c_1944_n N_A_381_47#_c_1945_n
+ N_A_381_47#_c_1947_n N_A_381_47#_c_1948_n N_A_381_47#_c_1978_n
+ N_A_381_47#_c_1949_n PM_SKY130_FD_SC_HD__DFBBN_1%A_381_47#
x_PM_SKY130_FD_SC_HD__DFBBN_1%Q_N N_Q_N_M1030_d N_Q_N_M1039_d N_Q_N_c_2021_n
+ N_Q_N_c_2018_n Q_N Q_N Q_N N_Q_N_c_2020_n Q_N PM_SKY130_FD_SC_HD__DFBBN_1%Q_N
x_PM_SKY130_FD_SC_HD__DFBBN_1%Q N_Q_M1027_d N_Q_M1037_d N_Q_c_2049_n
+ N_Q_c_2052_n N_Q_c_2050_n Q Q Q PM_SKY130_FD_SC_HD__DFBBN_1%Q
x_PM_SKY130_FD_SC_HD__DFBBN_1%VGND N_VGND_M1033_d N_VGND_M1002_s N_VGND_M1007_d
+ N_VGND_M1019_s N_VGND_M1020_d N_VGND_M1015_d N_VGND_M1010_d N_VGND_c_2067_n
+ N_VGND_c_2068_n N_VGND_c_2069_n N_VGND_c_2070_n N_VGND_c_2071_n
+ N_VGND_c_2072_n N_VGND_c_2073_n N_VGND_c_2074_n N_VGND_c_2075_n
+ N_VGND_c_2076_n N_VGND_c_2077_n N_VGND_c_2078_n N_VGND_c_2079_n VGND VGND
+ N_VGND_c_2080_n N_VGND_c_2081_n N_VGND_c_2082_n N_VGND_c_2083_n
+ N_VGND_c_2084_n N_VGND_c_2085_n N_VGND_c_2086_n N_VGND_c_2087_n
+ N_VGND_c_2088_n N_VGND_c_2089_n PM_SKY130_FD_SC_HD__DFBBN_1%VGND
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_791_47# N_A_791_47#_M1016_d N_A_791_47#_M1031_d
+ N_A_791_47#_c_2257_n N_A_791_47#_c_2260_n N_A_791_47#_c_2267_n
+ PM_SKY130_FD_SC_HD__DFBBN_1%A_791_47#
x_PM_SKY130_FD_SC_HD__DFBBN_1%A_1555_47# N_A_1555_47#_M1009_d
+ N_A_1555_47#_M1032_d N_A_1555_47#_c_2292_n N_A_1555_47#_c_2288_n
+ N_A_1555_47#_c_2293_n PM_SKY130_FD_SC_HD__DFBBN_1%A_1555_47#
cc_1 VNB N_CLK_N_c_257_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_N_c_258_n 0.0233703f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK_N 0.0189188f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_N_c_260_n 0.0195341f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_CLK_N_c_261_n 0.0141411f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1013_g 0.0382826f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_303_n 0.0133397f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_27_47#_c_304_n 0.0047037f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_9 VNB N_A_27_47#_M1038_g 0.0197664f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_10 VNB N_A_27_47#_c_306_n 0.00878847f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_11 VNB N_A_27_47#_c_307_n 0.0179705f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_12 VNB N_A_27_47#_c_308_n 9.27212e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_309_n 0.00640562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_310_n 0.00137395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_311_n 0.027308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_312_n 0.0247224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_313_n 0.00419271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_314_n 0.0012554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_315_n 0.0207662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_316_n 0.00235584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_317_n 0.00293177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_318_n 0.00200585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_319_n 0.00104784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_320_n 0.0229463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_321_n 0.0249277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_322_n 0.00498131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_323_n 0.00672408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_D_M1002_g 0.0339092f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_29 VNB N_D_c_565_n 0.0258448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_D_c_566_n 0.00419137f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_31 VNB N_A_193_47#_c_605_n 0.0178504f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_32 VNB N_A_193_47#_c_606_n 0.0124337f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_33 VNB N_A_193_47#_c_607_n 0.00441338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_M1036_g 0.0460424f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_35 VNB N_A_193_47#_c_609_n 0.00411619f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_36 VNB N_A_193_47#_c_610_n 0.0303522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_611_n 0.0161622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_647_21#_M1007_g 0.0422736f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_39 VNB N_A_647_21#_c_808_n 0.0200445f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_40 VNB N_A_647_21#_c_809_n 0.00190301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_647_21#_c_810_n 0.00419895f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_42 VNB N_A_647_21#_c_811_n 0.0115295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_647_21#_c_812_n 0.00591507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_647_21#_c_813_n 0.0323382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_SET_B_c_954_n 0.0324673f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_46 VNB N_SET_B_M1004_g 0.00696335f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_47 VNB N_SET_B_M1016_g 0.0204057f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_48 VNB N_SET_B_M1009_g 0.0201994f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_49 VNB N_SET_B_c_958_n 0.0315063f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_50 VNB N_SET_B_M1012_g 0.00600733f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_51 VNB SET_B 0.00764108f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_52 VNB N_SET_B_c_961_n 0.0143319f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_53 VNB N_SET_B_c_962_n 0.00190663f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_54 VNB N_SET_B_c_963_n 0.00108341f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_55 VNB N_SET_B_c_964_n 0.00753532f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_56 VNB N_A_473_413#_M1035_g 0.0258405f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_57 VNB N_A_473_413#_c_1087_n 0.00430594f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_58 VNB N_A_473_413#_c_1088_n 0.00748589f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_59 VNB N_A_473_413#_c_1089_n 0.00392752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_473_413#_c_1090_n 0.0141708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_941_21#_M1031_g 0.0293266f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_62 VNB N_A_941_21#_M1032_g 0.0278383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_941_21#_c_1193_n 0.0112954f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_64 VNB N_A_941_21#_c_1194_n 0.00191901f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_65 VNB N_A_941_21#_c_1195_n 0.00262532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_941_21#_c_1196_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_941_21#_c_1197_n 0.0214041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_941_21#_c_1198_n 0.00250659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_941_21#_c_1199_n 0.00364137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_941_21#_c_1200_n 0.0186918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_941_21#_c_1201_n 3.26335e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1415_315#_M1020_g 0.043407f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_73 VNB N_A_1415_315#_c_1360_n 0.0204041f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_74 VNB N_A_1415_315#_c_1361_n 0.0582626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1415_315#_c_1362_n 0.0156851f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_76 VNB N_A_1415_315#_c_1363_n 0.00812918f $X=-0.19 $Y=-0.24 $X2=0.24
+ $Y2=1.235
cc_77 VNB N_A_1415_315#_c_1364_n 4.80417e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_78 VNB N_A_1415_315#_c_1365_n 0.0183894f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_79 VNB N_A_1415_315#_c_1366_n 0.0180366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1415_315#_c_1367_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1415_315#_c_1368_n 0.00319517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1415_315#_c_1369_n 0.00272728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1256_413#_M1025_g 0.0225426f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_84 VNB N_A_1256_413#_c_1555_n 0.0111717f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_85 VNB N_A_1256_413#_c_1556_n 0.0106187f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_86 VNB N_A_1256_413#_c_1557_n 4.9687e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1256_413#_c_1558_n 0.00200975f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_88 VNB N_A_1256_413#_c_1559_n 0.0197989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_RESET_B_M1015_g 0.0348161f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_90 VNB RESET_B 0.00351479f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_91 VNB N_RESET_B_c_1668_n 0.0292509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2136_47#_c_1705_n 0.0072656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_2136_47#_c_1706_n 0.00515122f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_94 VNB N_A_2136_47#_c_1707_n 0.025727f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_95 VNB N_A_2136_47#_c_1708_n 2.88662e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_96 VNB N_A_2136_47#_c_1709_n 0.0201038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VPWR_c_1759_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_381_47#_c_1943_n 0.00960564f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_99 VNB N_A_381_47#_c_1944_n 0.0043665f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_100 VNB N_A_381_47#_c_1945_n 0.00317304f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_101 VNB N_Q_N_c_2018_n 0.00377204f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_102 VNB Q_N 0.00140118f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_103 VNB N_Q_N_c_2020_n 0.00366681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_Q_c_2049_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_105 VNB N_Q_c_2050_n 0.0229373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB Q 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_107 VNB N_VGND_c_2067_n 4.08532e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_108 VNB N_VGND_c_2068_n 0.00537094f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_109 VNB N_VGND_c_2069_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2070_n 0.00606447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2071_n 0.00267847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2072_n 0.00476184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2073_n 0.002607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2074_n 0.0443368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2075_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2076_n 0.0381013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2077_n 0.00545594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2078_n 0.040336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2079_n 0.00491654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2080_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2081_n 0.0156788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2082_n 0.0529546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2083_n 0.0287938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2084_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2085_n 0.5617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2086_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2087_n 0.005552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2088_n 0.00462385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2089_n 0.00440183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VPB N_CLK_N_c_262_n 0.0118979f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_131 VPB N_CLK_N_c_263_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_132 VPB N_CLK_N_c_264_n 0.0238011f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_133 VPB CLK_N 0.0179925f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_134 VPB N_CLK_N_c_260_n 0.0100928f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_135 VPB N_A_27_47#_M1000_g 0.0363084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_136 VPB N_A_27_47#_M1021_g 0.045988f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_137 VPB N_A_27_47#_c_303_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_138 VPB N_A_27_47#_c_304_n 0.0032343f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_139 VPB N_A_27_47#_M1022_g 0.0215753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_329_n 0.00194467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_330_n 0.00383512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_331_n 0.0281213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_332_n 0.00354649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_317_n 0.00323841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_319_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_320_n 0.0117662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_323_n 3.29025e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_D_M1017_g 0.0559187f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_149 VPB N_D_c_565_n 0.00540326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_D_c_566_n 0.0069444f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_151 VPB N_A_193_47#_M1014_g 0.0215876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_193_47#_M1034_g 0.020906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_193_47#_c_606_n 0.0178865f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_154 VPB N_A_193_47#_c_607_n 0.00403646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_193_47#_c_609_n 0.00245106f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_156 VPB N_A_193_47#_c_617_n 0.00871552f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_157 VPB N_A_193_47#_c_618_n 0.00466989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_193_47#_c_619_n 0.00875464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_193_47#_c_620_n 0.00166205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_193_47#_c_621_n 0.00361682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_193_47#_c_622_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_193_47#_c_623_n 0.00575159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_193_47#_c_624_n 0.0283351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_193_47#_c_625_n 0.00471853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_193_47#_c_626_n 0.0125285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_193_47#_c_611_n 0.0175606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_647_21#_M1007_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_168 VPB N_A_647_21#_M1023_g 0.0210587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_169 VPB N_A_647_21#_M1028_g 0.0317411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_170 VPB N_A_647_21#_c_817_n 0.0055347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_647_21#_c_810_n 0.00619168f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_172 VPB N_A_647_21#_c_819_n 0.00575673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_647_21#_c_820_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_647_21#_c_813_n 0.00659461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_SET_B_M1004_g 0.0508831f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_176 VPB N_SET_B_M1012_g 0.0515333f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_177 VPB N_A_473_413#_M1024_g 0.0203673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_178 VPB N_A_473_413#_c_1092_n 0.0121994f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_179 VPB N_A_473_413#_c_1088_n 0.00789134f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_180 VPB N_A_473_413#_c_1089_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_473_413#_c_1090_n 0.0165426f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_941_21#_M1018_g 0.0205161f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_183 VPB N_A_941_21#_M1005_g 0.0207759f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_184 VPB N_A_941_21#_c_1204_n 0.00126237f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_185 VPB N_A_941_21#_c_1205_n 0.00527345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_941_21#_c_1196_n 0.00162652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_941_21#_c_1197_n 0.0228551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_941_21#_c_1208_n 0.0286431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_941_21#_c_1209_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_941_21#_c_1210_n 0.00737873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_941_21#_c_1211_n 0.00302735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_941_21#_c_1200_n 0.0212626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_941_21#_c_1201_n 0.00361185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1415_315#_M1008_g 0.0210257f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_195 VPB N_A_1415_315#_M1020_g 0.0159543f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_196 VPB N_A_1415_315#_M1039_g 0.0245523f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_197 VPB N_A_1415_315#_c_1362_n 0.00543649f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_198 VPB N_A_1415_315#_c_1364_n 0.0131679f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_199 VPB N_A_1415_315#_c_1375_n 0.0188717f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_200 VPB N_A_1415_315#_c_1376_n 0.0180742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1415_315#_c_1377_n 0.00426841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1415_315#_c_1378_n 0.0364062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1415_315#_c_1379_n 0.0034494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1415_315#_c_1380_n 8.78324e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1415_315#_c_1368_n 0.0032794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1415_315#_c_1382_n 0.00621558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_1415_315#_c_1383_n 0.00168728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_1415_315#_c_1384_n 2.32251e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_1415_315#_c_1369_n 2.41008e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_1256_413#_M1003_g 0.0224692f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_211 VPB N_A_1256_413#_c_1561_n 0.00609106f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.07
cc_212 VPB N_A_1256_413#_c_1556_n 0.00541384f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_213 VPB N_A_1256_413#_c_1557_n 7.48159e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_1256_413#_c_1558_n 0.00179991f $X=-0.19 $Y=1.305 $X2=0.26
+ $Y2=1.53
cc_215 VPB N_A_1256_413#_c_1559_n 0.0108842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_RESET_B_M1029_g 0.0248948f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_217 VPB RESET_B 7.97678e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_218 VPB N_RESET_B_c_1668_n 0.00965023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_2136_47#_M1037_g 0.0242905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_2136_47#_c_1711_n 0.0132505f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_221 VPB N_A_2136_47#_c_1706_n 0.00532263f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_222 VPB N_A_2136_47#_c_1707_n 0.00571877f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_223 VPB N_VPWR_c_1760_n 0.00105358f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_224 VPB N_VPWR_c_1761_n 0.00629486f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_225 VPB N_VPWR_c_1762_n 0.00313724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1763_n 0.00562862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1764_n 0.00350025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1765_n 0.0292737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1766_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1767_n 0.00407681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1768_n 0.0229981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1769_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1770_n 0.0155587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1771_n 0.0408432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1772_n 0.0591311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1773_n 0.0298382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1774_n 0.0293379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1775_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1759_n 0.0684784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1777_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1778_n 0.00555916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1779_n 0.00609488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1780_n 0.00929447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1781_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1782_n 0.00430944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_A_381_47#_c_1943_n 0.0098785f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_247 VPB N_A_381_47#_c_1947_n 0.00988091f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_248 VPB N_A_381_47#_c_1948_n 0.00333288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_A_381_47#_c_1949_n 0.00182829f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_250 VPB N_Q_N_c_2021_n 0.00137514f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_251 VPB N_Q_N_c_2018_n 0.00384084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_252 VPB Q_N 0.00760625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_Q_c_2052_n 0.00609566f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_254 VPB N_Q_c_2050_n 0.00768289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB Q 0.0337655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 N_CLK_N_c_257_n N_A_27_47#_M1013_g 0.0200656f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_257 CLK_N N_A_27_47#_M1013_g 3.13492e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_258 N_CLK_N_c_261_n N_A_27_47#_M1013_g 0.00499141f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_259 N_CLK_N_c_264_n N_A_27_47#_M1000_g 0.0275676f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_260 CLK_N N_A_27_47#_M1000_g 5.79634e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_261 N_CLK_N_c_260_n N_A_27_47#_M1000_g 0.00521293f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_262 N_CLK_N_c_257_n N_A_27_47#_c_308_n 0.00684762f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_263 N_CLK_N_c_258_n N_A_27_47#_c_308_n 0.00799602f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_264 CLK_N N_A_27_47#_c_308_n 0.00698378f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_265 N_CLK_N_c_258_n N_A_27_47#_c_309_n 0.00620138f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_266 CLK_N N_A_27_47#_c_309_n 0.0143701f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_267 N_CLK_N_c_260_n N_A_27_47#_c_309_n 2.99031e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_268 N_CLK_N_c_263_n N_A_27_47#_c_329_n 0.0129414f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_269 N_CLK_N_c_264_n N_A_27_47#_c_329_n 0.0013404f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_270 CLK_N N_A_27_47#_c_329_n 0.00690269f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_271 N_CLK_N_c_263_n N_A_27_47#_c_332_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_272 N_CLK_N_c_264_n N_A_27_47#_c_332_n 0.00374438f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_273 CLK_N N_A_27_47#_c_332_n 0.0153137f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_274 N_CLK_N_c_260_n N_A_27_47#_c_332_n 2.3617e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_275 N_CLK_N_c_258_n N_A_27_47#_c_313_n 0.0017102f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_276 N_CLK_N_c_261_n N_A_27_47#_c_313_n 0.00154323f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_277 N_CLK_N_c_258_n N_A_27_47#_c_317_n 0.00161727f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_278 N_CLK_N_c_264_n N_A_27_47#_c_317_n 0.00455491f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_279 CLK_N N_A_27_47#_c_317_n 0.0506358f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_280 N_CLK_N_c_260_n N_A_27_47#_c_317_n 0.0010036f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_281 N_CLK_N_c_261_n N_A_27_47#_c_317_n 0.0020643f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_282 CLK_N N_A_27_47#_c_320_n 0.00164115f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_283 N_CLK_N_c_260_n N_A_27_47#_c_320_n 0.0169859f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_284 N_CLK_N_c_263_n N_VPWR_c_1760_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_285 N_CLK_N_c_263_n N_VPWR_c_1769_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_286 N_CLK_N_c_263_n N_VPWR_c_1759_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_287 N_CLK_N_c_257_n N_VGND_c_2067_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_288 N_CLK_N_c_257_n N_VGND_c_2080_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_289 N_CLK_N_c_258_n N_VGND_c_2080_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_290 N_CLK_N_c_257_n N_VGND_c_2085_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_312_n N_D_M1002_g 0.00346149f $X=2.845 $Y=0.85 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_304_n N_D_M1017_g 0.0336995f $X=2.365 $Y=1.32 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_304_n N_D_c_565_n 0.00467503f $X=2.365 $Y=1.32 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_312_n N_D_c_565_n 0.00129446f $X=2.845 $Y=0.85 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_304_n N_D_c_566_n 0.00320876f $X=2.365 $Y=1.32 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_312_n N_D_c_566_n 0.0119589f $X=2.845 $Y=0.85 $X2=0 $Y2=0
cc_297 N_A_27_47#_M1038_g N_A_193_47#_c_605_n 0.00882622f $X=2.83 $Y=0.415 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_322_n N_A_193_47#_c_605_n 5.15019e-19 $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1021_g N_A_193_47#_M1014_g 0.0190567f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_330_n N_A_193_47#_c_606_n 0.00783754f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_331_n N_A_193_47#_c_606_n 0.021675f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_319_n N_A_193_47#_c_606_n 3.23054e-19 $X=6.21 $Y=1.19 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_323_n N_A_193_47#_c_606_n 0.0111119f $X=6.295 $Y=1.182 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_311_n N_A_193_47#_c_607_n 0.0173623f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_319_n N_A_193_47#_c_607_n 9.01357e-19 $X=6.21 $Y=1.19 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_323_n N_A_193_47#_c_607_n 0.00481144f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_307 N_A_27_47#_c_307_n N_A_193_47#_M1036_g 0.0130863f $X=6.32 $Y=0.705 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_310_n N_A_193_47#_M1036_g 0.00170335f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_311_n N_A_193_47#_M1036_g 0.0211332f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_323_n N_A_193_47#_M1036_g 0.00779497f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_M1021_g N_A_193_47#_c_609_n 0.00533691f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_303_n N_A_193_47#_c_609_n 0.010154f $X=2.755 $Y=1.32 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_304_n N_A_193_47#_c_609_n 0.0020394f $X=2.365 $Y=1.32 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1038_g N_A_193_47#_c_609_n 4.45841e-19 $X=2.83 $Y=0.415 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_312_n N_A_193_47#_c_609_n 0.017282f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_314_n N_A_193_47#_c_609_n 0.00934078f $X=3.027 $Y=1.12 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_318_n N_A_193_47#_c_609_n 4.74166e-19 $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_321_n N_A_193_47#_c_609_n 0.00674133f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_322_n N_A_193_47#_c_609_n 0.0210004f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_304_n N_A_193_47#_c_610_n 0.0220418f $X=2.365 $Y=1.32 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1038_g N_A_193_47#_c_610_n 0.0213475f $X=2.83 $Y=0.415 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_312_n N_A_193_47#_c_610_n 0.00483145f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_322_n N_A_193_47#_c_610_n 0.00153496f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1021_g N_A_193_47#_c_617_n 0.0069032f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1000_g N_A_193_47#_c_618_n 0.00459685f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_329_n N_A_193_47#_c_618_n 0.00562897f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_317_n N_A_193_47#_c_618_n 0.00113911f $X=0.695 $Y=0.85 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_303_n N_A_193_47#_c_619_n 3.83457e-19 $X=2.755 $Y=1.32 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_316_n N_A_193_47#_c_619_n 0.11126f $X=3.135 $Y=1.19 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_M1021_g N_A_193_47#_c_620_n 5.24592e-19 $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_M1022_g N_A_193_47#_c_621_n 0.00133927f $X=6.625 $Y=2.275
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_330_n N_A_193_47#_c_621_n 0.00483121f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_331_n N_A_193_47#_c_621_n 0.00219663f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_M1021_g N_A_193_47#_c_622_n 0.0174486f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_303_n N_A_193_47#_c_622_n 0.0212221f $X=2.755 $Y=1.32 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_322_n N_A_193_47#_c_622_n 3.18577e-19 $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_M1021_g N_A_193_47#_c_623_n 0.0103132f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_303_n N_A_193_47#_c_623_n 0.00654686f $X=2.755 $Y=1.32 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_322_n N_A_193_47#_c_623_n 0.00339609f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1022_g N_A_193_47#_c_624_n 0.0192968f $X=6.625 $Y=2.275 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_330_n N_A_193_47#_c_624_n 5.88448e-19 $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_331_n N_A_193_47#_c_624_n 0.0169266f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_315_n N_A_193_47#_c_624_n 2.37019e-19 $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_323_n N_A_193_47#_c_624_n 3.74988e-19 $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_M1022_g N_A_193_47#_c_625_n 6.52047e-19 $X=6.625 $Y=2.275
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_330_n N_A_193_47#_c_625_n 0.0168759f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_331_n N_A_193_47#_c_625_n 0.00153059f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_319_n N_A_193_47#_c_625_n 5.52451e-19 $X=6.21 $Y=1.19 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_323_n N_A_193_47#_c_625_n 0.00921846f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_330_n N_A_193_47#_c_626_n 0.00347329f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_M1013_g N_A_193_47#_c_611_n 0.0270893f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_308_n N_A_193_47#_c_611_n 0.0116433f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_329_n N_A_193_47#_c_611_n 0.0088687f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_312_n N_A_193_47#_c_611_n 0.0237208f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_313_n N_A_193_47#_c_611_n 0.00146306f $X=0.84 $Y=0.85 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_317_n N_A_193_47#_c_611_n 0.0704454f $X=0.695 $Y=0.85 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_M1038_g N_A_647_21#_M1007_g 0.0245694f $X=2.83 $Y=0.415 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_306_n N_A_647_21#_M1007_g 0.0105189f $X=2.83 $Y=1.245 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_315_n N_A_647_21#_M1007_g 7.74803e-19 $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_318_n N_A_647_21#_M1007_g 0.00642269f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_321_n N_A_647_21#_M1007_g 0.0200662f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_322_n N_A_647_21#_M1007_g 0.00189958f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_307_n N_A_647_21#_c_808_n 0.0170372f $X=6.32 $Y=0.705 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_310_n N_A_647_21#_c_808_n 0.00157071f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_311_n N_A_647_21#_c_808_n 0.0105048f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_315_n N_A_647_21#_c_817_n 0.00196084f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_315_n N_A_647_21#_c_832_n 0.00348372f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_315_n N_A_647_21#_c_809_n 0.00165548f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_315_n N_A_647_21#_c_810_n 0.016449f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_315_n N_A_647_21#_c_811_n 0.00907541f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_315_n N_A_647_21#_c_819_n 8.24776e-19 $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_315_n N_A_647_21#_c_837_n 6.83984e-19 $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_310_n N_A_647_21#_c_812_n 0.00700206f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_311_n N_A_647_21#_c_812_n 9.34624e-19 $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_315_n N_A_647_21#_c_812_n 0.015092f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_319_n N_A_647_21#_c_812_n 3.46518e-19 $X=6.21 $Y=1.19 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_323_n N_A_647_21#_c_812_n 0.00922241f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_315_n N_A_647_21#_c_813_n 0.00365485f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_323_n N_A_647_21#_c_813_n 0.00232132f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_315_n N_SET_B_c_954_n 0.00392015f $X=6.065 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_381 N_A_27_47#_c_315_n N_SET_B_M1004_g 0.0011704f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_315_n SET_B 0.00593372f $X=6.065 $Y=1.19 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_310_n N_SET_B_c_961_n 0.0170283f $X=6.32 $Y=0.87 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_311_n N_SET_B_c_961_n 0.00246584f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_315_n N_SET_B_c_961_n 0.158116f $X=6.065 $Y=1.19 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_319_n N_SET_B_c_961_n 0.0254613f $X=6.21 $Y=1.19 $X2=0 $Y2=0
cc_387 N_A_27_47#_c_323_n N_SET_B_c_961_n 0.00910371f $X=6.295 $Y=1.182 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_315_n N_SET_B_c_962_n 0.0265123f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_315_n N_A_473_413#_M1035_g 0.00188875f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_M1021_g N_A_473_413#_c_1097_n 0.00275336f $X=2.29 $Y=2.275
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_M1038_g N_A_473_413#_c_1098_n 0.00883573f $X=2.83 $Y=0.415
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_312_n N_A_473_413#_c_1098_n 0.00579266f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_318_n N_A_473_413#_c_1098_n 0.00257401f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_321_n N_A_473_413#_c_1098_n 5.24878e-19 $X=2.89 $Y=0.93
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_322_n N_A_473_413#_c_1098_n 0.0194937f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1021_g N_A_473_413#_c_1092_n 8.73767e-19 $X=2.29 $Y=2.275
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_316_n N_A_473_413#_c_1092_n 3.03433e-19 $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_M1038_g N_A_473_413#_c_1087_n 0.00119254f $X=2.83 $Y=0.415
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_306_n N_A_473_413#_c_1087_n 8.54957e-19 $X=2.83 $Y=1.245
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_315_n N_A_473_413#_c_1087_n 0.0145635f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_318_n N_A_473_413#_c_1087_n 0.0138897f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_321_n N_A_473_413#_c_1087_n 7.78235e-19 $X=2.89 $Y=0.93
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_322_n N_A_473_413#_c_1087_n 0.0244377f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_315_n N_A_473_413#_c_1088_n 0.0375702f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_306_n N_A_473_413#_c_1089_n 0.00268952f $X=2.83 $Y=1.245
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_315_n N_A_473_413#_c_1089_n 0.0109965f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_316_n N_A_473_413#_c_1089_n 0.00666557f $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_321_n N_A_473_413#_c_1089_n 5.70846e-19 $X=2.89 $Y=0.93
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_322_n N_A_473_413#_c_1089_n 0.0053097f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_c_315_n N_A_473_413#_c_1090_n 0.00386813f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_315_n N_A_941_21#_M1031_g 0.00150073f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_315_n N_A_941_21#_c_1196_n 0.0122882f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_315_n N_A_941_21#_c_1197_n 0.00603655f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_330_n N_A_941_21#_c_1208_n 0.0173527f $X=6.655 $Y=1.74 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_331_n N_A_941_21#_c_1208_n 0.00184742f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_315_n N_A_941_21#_c_1208_n 0.014133f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_319_n N_A_941_21#_c_1208_n 0.0261705f $X=6.21 $Y=1.19 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_323_n N_A_941_21#_c_1208_n 0.00750434f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_315_n N_A_941_21#_c_1209_n 0.0276968f $X=6.065 $Y=1.19 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_330_n N_A_941_21#_c_1210_n 0.00264766f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_315_n N_A_941_21#_c_1210_n 0.00618009f $X=6.065 $Y=1.19
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_330_n N_A_1415_315#_M1020_g 3.1988e-19 $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_M1022_g N_A_1415_315#_c_1378_n 0.0224334f $X=6.625 $Y=2.275
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_330_n N_A_1415_315#_c_1378_n 4.29767e-19 $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_331_n N_A_1415_315#_c_1378_n 0.0130101f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_M1022_g N_A_1256_413#_c_1566_n 0.00933665f $X=6.625 $Y=2.275
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_330_n N_A_1256_413#_c_1566_n 0.00676569f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_428 N_A_27_47#_c_331_n N_A_1256_413#_c_1566_n 0.0028948f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_307_n N_A_1256_413#_c_1569_n 0.00721774f $X=6.32 $Y=0.705
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_310_n N_A_1256_413#_c_1569_n 0.0046226f $X=6.32 $Y=0.87
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_311_n N_A_1256_413#_c_1569_n 9.76146e-19 $X=6.32 $Y=0.87
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_323_n N_A_1256_413#_c_1569_n 0.00311508f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_310_n N_A_1256_413#_c_1555_n 0.00957451f $X=6.32 $Y=0.87
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_319_n N_A_1256_413#_c_1555_n 6.68034e-19 $X=6.21 $Y=1.19
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_323_n N_A_1256_413#_c_1555_n 0.0105978f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_M1022_g N_A_1256_413#_c_1561_n 0.00635237f $X=6.625 $Y=2.275
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_330_n N_A_1256_413#_c_1561_n 0.0359924f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_331_n N_A_1256_413#_c_1561_n 0.00186193f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_330_n N_A_1256_413#_c_1557_n 0.00817073f $X=6.655 $Y=1.74
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_319_n N_A_1256_413#_c_1557_n 2.72722e-19 $X=6.21 $Y=1.19
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_323_n N_A_1256_413#_c_1557_n 0.00601065f $X=6.295 $Y=1.182
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_329_n N_VPWR_M1011_d 0.00167655f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_443 N_A_27_47#_M1000_g N_VPWR_c_1760_n 0.0082474f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_329_n N_VPWR_c_1760_n 0.0175536f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_445 N_A_27_47#_c_332_n N_VPWR_c_1760_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_446 N_A_27_47#_M1000_g N_VPWR_c_1761_n 0.00193825f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_M1021_g N_VPWR_c_1761_n 0.00113398f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_329_n N_VPWR_c_1769_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_332_n N_VPWR_c_1769_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_450 N_A_27_47#_M1000_g N_VPWR_c_1770_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_M1021_g N_VPWR_c_1771_n 0.00541732f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_M1022_g N_VPWR_c_1772_n 0.00367119f $X=6.625 $Y=2.275 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1000_g N_VPWR_c_1759_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_M1021_g N_VPWR_c_1759_n 0.00621511f $X=2.29 $Y=2.275 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_M1022_g N_VPWR_c_1759_n 0.00554407f $X=6.625 $Y=2.275 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_329_n N_VPWR_c_1759_n 0.00507261f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_332_n N_VPWR_c_1759_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_312_n N_A_381_47#_c_1943_n 0.0148981f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_312_n N_A_381_47#_c_1944_n 0.0207493f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_322_n N_A_381_47#_c_1944_n 0.00214915f $X=2.89 $Y=0.93 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_312_n N_A_381_47#_c_1945_n 0.00431455f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_462 N_A_27_47#_M1021_g N_A_381_47#_c_1947_n 0.00141699f $X=2.29 $Y=2.275
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_M1021_g N_A_381_47#_c_1949_n 0.00738444f $X=2.29 $Y=2.275
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_c_308_n N_VGND_M1033_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_465 N_A_27_47#_M1013_g N_VGND_c_2067_n 0.00777283f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_308_n N_VGND_c_2067_n 0.0158742f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_467 N_A_27_47#_c_313_n N_VGND_c_2067_n 0.00116283f $X=0.84 $Y=0.85 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_320_n N_VGND_c_2067_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1013_g N_VGND_c_2068_n 0.00305176f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_312_n N_VGND_c_2068_n 0.00132494f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_307_n N_VGND_c_2070_n 0.001573f $X=6.32 $Y=0.705 $X2=0 $Y2=0
cc_472 N_A_27_47#_M1038_g N_VGND_c_2074_n 0.00359964f $X=2.83 $Y=0.415 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_307_n N_VGND_c_2078_n 0.00387466f $X=6.32 $Y=0.705 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_310_n N_VGND_c_2078_n 0.00173925f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_311_n N_VGND_c_2078_n 2.14983e-19 $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_550_p N_VGND_c_2080_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_308_n N_VGND_c_2080_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_M1013_g N_VGND_c_2081_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_M1033_s N_VGND_c_2085_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_M1013_g N_VGND_c_2085_n 0.00581646f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_M1038_g N_VGND_c_2085_n 0.00559273f $X=2.83 $Y=0.415 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_307_n N_VGND_c_2085_n 0.00580109f $X=6.32 $Y=0.705 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_550_p N_VGND_c_2085_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_c_308_n N_VGND_c_2085_n 0.00526087f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_310_n N_VGND_c_2085_n 0.00154594f $X=6.32 $Y=0.87 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_312_n N_VGND_c_2085_n 0.0939486f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_313_n N_VGND_c_2085_n 0.0131302f $X=0.84 $Y=0.85 $X2=0 $Y2=0
cc_488 N_A_27_47#_c_318_n N_VGND_c_2085_n 0.0153531f $X=2.99 $Y=0.85 $X2=0 $Y2=0
cc_489 N_A_27_47#_c_322_n A_581_47# 0.00109904f $X=2.89 $Y=0.93 $X2=-0.19
+ $Y2=-0.24
cc_490 N_D_M1002_g N_A_193_47#_c_605_n 0.0212313f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_491 N_D_M1002_g N_A_193_47#_c_609_n 0.0012555f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_492 N_D_c_565_n N_A_193_47#_c_609_n 0.00106245f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_493 N_D_c_566_n N_A_193_47#_c_609_n 0.0453933f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_494 N_D_c_565_n N_A_193_47#_c_610_n 0.00136462f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_495 N_D_c_566_n N_A_193_47#_c_610_n 2.34518e-19 $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_496 N_D_c_566_n N_A_193_47#_c_617_n 0.00466646f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_497 N_D_M1017_g N_A_193_47#_c_618_n 4.11004e-19 $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_498 N_D_M1017_g N_A_193_47#_c_623_n 0.00106391f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_499 N_D_c_566_n N_A_193_47#_c_623_n 0.00408526f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_500 N_D_M1002_g N_A_193_47#_c_611_n 0.00369511f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_501 N_D_M1017_g N_A_193_47#_c_611_n 0.00452067f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_502 N_D_M1017_g N_VPWR_c_1761_n 0.0117356f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_503 N_D_M1017_g N_VPWR_c_1771_n 0.0035268f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_504 N_D_M1017_g N_VPWR_c_1759_n 0.0039725f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_505 N_D_M1002_g N_A_381_47#_c_1943_n 0.00537833f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_506 N_D_M1017_g N_A_381_47#_c_1943_n 0.00775166f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_507 N_D_c_565_n N_A_381_47#_c_1943_n 0.00753248f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_508 N_D_c_566_n N_A_381_47#_c_1943_n 0.0486094f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_509 N_D_M1002_g N_A_381_47#_c_1944_n 0.0125635f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_510 N_D_c_565_n N_A_381_47#_c_1944_n 0.0021626f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_511 N_D_c_566_n N_A_381_47#_c_1944_n 0.0246039f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_512 N_D_M1017_g N_A_381_47#_c_1947_n 0.0129489f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_513 N_D_c_565_n N_A_381_47#_c_1947_n 0.00167192f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_514 N_D_c_566_n N_A_381_47#_c_1947_n 0.0289371f $X=1.83 $Y=1.17 $X2=0 $Y2=0
cc_515 N_D_M1017_g N_A_381_47#_c_1949_n 0.00258776f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_516 N_D_M1002_g N_VGND_c_2068_n 0.00946079f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_517 N_D_M1002_g N_VGND_c_2074_n 0.00339367f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_518 N_D_M1002_g N_VGND_c_2085_n 0.00393034f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_519 N_A_193_47#_c_609_n N_A_647_21#_M1007_g 5.35023e-19 $X=2.41 $Y=0.87 $X2=0
+ $Y2=0
cc_520 N_A_193_47#_c_619_n N_A_647_21#_M1023_g 0.00197541f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_M1034_g N_A_647_21#_M1028_g 0.0164618f $X=6.205 $Y=2.275
+ $X2=0 $Y2=0
cc_522 N_A_193_47#_c_607_n N_A_647_21#_M1028_g 0.00557961f $X=6.28 $Y=1.32 $X2=0
+ $Y2=0
cc_523 N_A_193_47#_c_619_n N_A_647_21#_M1028_g 0.00750594f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_524 N_A_193_47#_c_624_n N_A_647_21#_M1028_g 0.00910409f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_525 N_A_193_47#_c_625_n N_A_647_21#_M1028_g 0.00264318f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_526 N_A_193_47#_c_619_n N_A_647_21#_c_817_n 0.0240118f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_c_619_n N_A_647_21#_c_832_n 0.0279846f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_528 N_A_193_47#_c_619_n N_A_647_21#_c_819_n 0.0141612f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_M1014_g N_A_647_21#_c_820_n 0.0161827f $X=2.71 $Y=2.275 $X2=0
+ $Y2=0
cc_530 N_A_193_47#_c_619_n N_A_647_21#_c_820_n 0.00193898f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_531 N_A_193_47#_c_622_n N_A_647_21#_c_820_n 0.00927772f $X=2.74 $Y=1.74 $X2=0
+ $Y2=0
cc_532 N_A_193_47#_c_619_n N_A_647_21#_c_837_n 0.00959465f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_533 N_A_193_47#_c_607_n N_A_647_21#_c_813_n 0.00268671f $X=6.28 $Y=1.32 $X2=0
+ $Y2=0
cc_534 N_A_193_47#_M1036_g N_SET_B_c_961_n 0.00575227f $X=6.74 $Y=0.415 $X2=0
+ $Y2=0
cc_535 N_A_193_47#_M1014_g N_A_473_413#_c_1097_n 0.0091014f $X=2.71 $Y=2.275
+ $X2=0 $Y2=0
cc_536 N_A_193_47#_c_617_n N_A_473_413#_c_1097_n 2.09728e-19 $X=2.385 $Y=1.87
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_c_619_n N_A_473_413#_c_1097_n 0.00506942f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_538 N_A_193_47#_c_620_n N_A_473_413#_c_1097_n 0.00303545f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_539 N_A_193_47#_c_622_n N_A_473_413#_c_1097_n 0.00186639f $X=2.74 $Y=1.74
+ $X2=0 $Y2=0
cc_540 N_A_193_47#_c_623_n N_A_473_413#_c_1097_n 0.0152514f $X=2.74 $Y=1.74
+ $X2=0 $Y2=0
cc_541 N_A_193_47#_c_609_n N_A_473_413#_c_1098_n 0.00620645f $X=2.41 $Y=0.87
+ $X2=0 $Y2=0
cc_542 N_A_193_47#_c_610_n N_A_473_413#_c_1098_n 8.57926e-19 $X=2.41 $Y=0.87
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_M1014_g N_A_473_413#_c_1092_n 0.00650943f $X=2.71 $Y=2.275
+ $X2=0 $Y2=0
cc_544 N_A_193_47#_c_609_n N_A_473_413#_c_1092_n 0.00666284f $X=2.41 $Y=0.87
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_619_n N_A_473_413#_c_1092_n 0.013911f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_620_n N_A_473_413#_c_1092_n 0.00149623f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_c_622_n N_A_473_413#_c_1092_n 0.00203066f $X=2.74 $Y=1.74
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_c_623_n N_A_473_413#_c_1092_n 0.0282877f $X=2.74 $Y=1.74
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_619_n N_A_473_413#_c_1088_n 0.00350894f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_550 N_A_193_47#_c_609_n N_A_473_413#_c_1089_n 0.00728915f $X=2.41 $Y=0.87
+ $X2=0 $Y2=0
cc_551 N_A_193_47#_c_619_n N_A_473_413#_c_1089_n 0.00456576f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_552 N_A_193_47#_c_619_n N_A_941_21#_M1018_g 0.00576309f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_553 N_A_193_47#_c_619_n N_A_941_21#_c_1196_n 0.00477237f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_554 N_A_193_47#_c_619_n N_A_941_21#_c_1197_n 3.78923e-19 $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_555 N_A_193_47#_c_606_n N_A_941_21#_c_1208_n 0.00389341f $X=6.665 $Y=1.32
+ $X2=0 $Y2=0
cc_556 N_A_193_47#_c_619_n N_A_941_21#_c_1208_n 0.0139809f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_557 N_A_193_47#_c_621_n N_A_941_21#_c_1208_n 0.0255925f $X=6.21 $Y=1.87 $X2=0
+ $Y2=0
cc_558 N_A_193_47#_c_624_n N_A_941_21#_c_1208_n 0.00183171f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_559 N_A_193_47#_c_625_n N_A_941_21#_c_1208_n 0.00622232f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_560 N_A_193_47#_c_626_n N_A_941_21#_c_1208_n 0.00371469f $X=6.145 $Y=1.575
+ $X2=0 $Y2=0
cc_561 N_A_193_47#_c_619_n N_A_941_21#_c_1209_n 0.0264578f $X=6.065 $Y=1.87
+ $X2=0 $Y2=0
cc_562 N_A_193_47#_c_624_n N_A_941_21#_c_1209_n 7.96394e-19 $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_563 N_A_193_47#_c_625_n N_A_941_21#_c_1209_n 0.00130051f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_564 N_A_193_47#_c_626_n N_A_941_21#_c_1209_n 7.27878e-19 $X=6.145 $Y=1.575
+ $X2=0 $Y2=0
cc_565 N_A_193_47#_c_619_n N_A_941_21#_c_1210_n 0.020032f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_566 N_A_193_47#_c_624_n N_A_941_21#_c_1210_n 6.45403e-19 $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_567 N_A_193_47#_c_625_n N_A_941_21#_c_1210_n 0.00461622f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_568 N_A_193_47#_c_626_n N_A_941_21#_c_1210_n 0.00148716f $X=6.145 $Y=1.575
+ $X2=0 $Y2=0
cc_569 N_A_193_47#_M1036_g N_A_1415_315#_M1020_g 0.0428021f $X=6.74 $Y=0.415
+ $X2=0 $Y2=0
cc_570 N_A_193_47#_M1034_g N_A_1256_413#_c_1566_n 0.00496872f $X=6.205 $Y=2.275
+ $X2=0 $Y2=0
cc_571 N_A_193_47#_c_621_n N_A_1256_413#_c_1566_n 0.00187313f $X=6.21 $Y=1.87
+ $X2=0 $Y2=0
cc_572 N_A_193_47#_c_625_n N_A_1256_413#_c_1566_n 0.00141396f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_573 N_A_193_47#_M1036_g N_A_1256_413#_c_1569_n 0.00963939f $X=6.74 $Y=0.415
+ $X2=0 $Y2=0
cc_574 N_A_193_47#_M1036_g N_A_1256_413#_c_1555_n 0.0106791f $X=6.74 $Y=0.415
+ $X2=0 $Y2=0
cc_575 N_A_193_47#_c_621_n N_A_1256_413#_c_1561_n 0.00214622f $X=6.21 $Y=1.87
+ $X2=0 $Y2=0
cc_576 N_A_193_47#_c_625_n N_A_1256_413#_c_1561_n 0.0013353f $X=6.145 $Y=1.74
+ $X2=0 $Y2=0
cc_577 N_A_193_47#_M1036_g N_A_1256_413#_c_1557_n 0.00154559f $X=6.74 $Y=0.415
+ $X2=0 $Y2=0
cc_578 N_A_193_47#_c_619_n N_VPWR_M1018_d 0.00670518f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_579 N_A_193_47#_c_611_n N_VPWR_c_1760_n 0.0127345f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_580 N_A_193_47#_c_617_n N_VPWR_c_1761_n 0.00179826f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_581 N_A_193_47#_c_611_n N_VPWR_c_1761_n 0.0243483f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_582 N_A_193_47#_c_619_n N_VPWR_c_1762_n 0.00160449f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_583 N_A_193_47#_c_619_n N_VPWR_c_1763_n 0.0137399f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_584 N_A_193_47#_c_611_n N_VPWR_c_1770_n 0.0156296f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_585 N_A_193_47#_M1014_g N_VPWR_c_1771_n 0.00367119f $X=2.71 $Y=2.275 $X2=0
+ $Y2=0
cc_586 N_A_193_47#_M1034_g N_VPWR_c_1772_n 0.00424681f $X=6.205 $Y=2.275 $X2=0
+ $Y2=0
cc_587 N_A_193_47#_c_625_n N_VPWR_c_1772_n 0.00254851f $X=6.145 $Y=1.74 $X2=0
+ $Y2=0
cc_588 N_A_193_47#_M1014_g N_VPWR_c_1759_n 0.00562272f $X=2.71 $Y=2.275 $X2=0
+ $Y2=0
cc_589 N_A_193_47#_M1034_g N_VPWR_c_1759_n 0.0061745f $X=6.205 $Y=2.275 $X2=0
+ $Y2=0
cc_590 N_A_193_47#_c_617_n N_VPWR_c_1759_n 0.0498118f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_591 N_A_193_47#_c_618_n N_VPWR_c_1759_n 0.0151864f $X=1.295 $Y=1.87 $X2=0
+ $Y2=0
cc_592 N_A_193_47#_c_619_n N_VPWR_c_1759_n 0.159156f $X=6.065 $Y=1.87 $X2=0
+ $Y2=0
cc_593 N_A_193_47#_c_620_n N_VPWR_c_1759_n 0.0160117f $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_594 N_A_193_47#_c_621_n N_VPWR_c_1759_n 0.0148451f $X=6.21 $Y=1.87 $X2=0
+ $Y2=0
cc_595 N_A_193_47#_c_623_n N_VPWR_c_1759_n 3.19863e-19 $X=2.74 $Y=1.74 $X2=0
+ $Y2=0
cc_596 N_A_193_47#_c_624_n N_VPWR_c_1759_n 3.05853e-19 $X=6.145 $Y=1.74 $X2=0
+ $Y2=0
cc_597 N_A_193_47#_c_625_n N_VPWR_c_1759_n 0.00131252f $X=6.145 $Y=1.74 $X2=0
+ $Y2=0
cc_598 N_A_193_47#_c_611_n N_VPWR_c_1759_n 0.00381175f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_599 N_A_193_47#_c_618_n N_A_381_47#_c_1943_n 0.00122075f $X=1.295 $Y=1.87
+ $X2=0 $Y2=0
cc_600 N_A_193_47#_c_611_n N_A_381_47#_c_1943_n 0.0733134f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_601 N_A_193_47#_c_605_n N_A_381_47#_c_1944_n 0.00218654f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_602 N_A_193_47#_c_609_n N_A_381_47#_c_1944_n 0.00812531f $X=2.41 $Y=0.87
+ $X2=0 $Y2=0
cc_603 N_A_193_47#_c_611_n N_A_381_47#_c_1945_n 0.015688f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_604 N_A_193_47#_c_617_n N_A_381_47#_c_1947_n 0.0308583f $X=2.385 $Y=1.87
+ $X2=0 $Y2=0
cc_605 N_A_193_47#_c_620_n N_A_381_47#_c_1947_n 7.06279e-19 $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_606 N_A_193_47#_c_623_n N_A_381_47#_c_1947_n 0.00962693f $X=2.74 $Y=1.74
+ $X2=0 $Y2=0
cc_607 N_A_193_47#_c_617_n N_A_381_47#_c_1948_n 0.0155963f $X=2.385 $Y=1.87
+ $X2=0 $Y2=0
cc_608 N_A_193_47#_c_618_n N_A_381_47#_c_1948_n 9.50689e-19 $X=1.295 $Y=1.87
+ $X2=0 $Y2=0
cc_609 N_A_193_47#_c_611_n N_A_381_47#_c_1948_n 0.0123978f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_610 N_A_193_47#_c_605_n N_A_381_47#_c_1978_n 0.00394877f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_611 N_A_193_47#_c_620_n N_A_381_47#_c_1949_n 8.71477e-19 $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_612 N_A_193_47#_c_619_n A_891_329# 0.00105375f $X=6.065 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_613 N_A_193_47#_c_619_n A_1112_329# 0.00532504f $X=6.065 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_614 N_A_193_47#_c_605_n N_VGND_c_2068_n 0.00121308f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_615 N_A_193_47#_c_611_n N_VGND_c_2068_n 0.00885393f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_616 N_A_193_47#_M1036_g N_VGND_c_2071_n 0.0012984f $X=6.74 $Y=0.415 $X2=0
+ $Y2=0
cc_617 N_A_193_47#_c_605_n N_VGND_c_2074_n 0.00531235f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_618 N_A_193_47#_c_609_n N_VGND_c_2074_n 0.00113905f $X=2.41 $Y=0.87 $X2=0
+ $Y2=0
cc_619 N_A_193_47#_M1036_g N_VGND_c_2078_n 0.00359964f $X=6.74 $Y=0.415 $X2=0
+ $Y2=0
cc_620 N_A_193_47#_c_611_n N_VGND_c_2081_n 0.00955835f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_621 N_A_193_47#_M1013_d N_VGND_c_2085_n 0.00217251f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_622 N_A_193_47#_c_605_n N_VGND_c_2085_n 0.00655518f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_623 N_A_193_47#_M1036_g N_VGND_c_2085_n 0.0053641f $X=6.74 $Y=0.415 $X2=0
+ $Y2=0
cc_624 N_A_193_47#_c_609_n N_VGND_c_2085_n 0.00118661f $X=2.41 $Y=0.87 $X2=0
+ $Y2=0
cc_625 N_A_193_47#_c_611_n N_VGND_c_2085_n 0.0038044f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_626 N_A_647_21#_M1007_g N_SET_B_c_954_n 0.0189927f $X=3.31 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_627 N_A_647_21#_M1007_g N_SET_B_M1004_g 0.0137896f $X=3.31 $Y=0.445 $X2=0
+ $Y2=0
cc_628 N_A_647_21#_M1023_g N_SET_B_M1004_g 0.0101628f $X=3.31 $Y=2.275 $X2=0
+ $Y2=0
cc_629 N_A_647_21#_c_817_n N_SET_B_M1004_g 0.0159332f $X=4.085 $Y=1.91 $X2=0
+ $Y2=0
cc_630 N_A_647_21#_c_864_p N_SET_B_M1004_g 0.00507112f $X=4.17 $Y=2.21 $X2=0
+ $Y2=0
cc_631 N_A_647_21#_c_819_n N_SET_B_M1004_g 0.00473578f $X=3.42 $Y=1.74 $X2=0
+ $Y2=0
cc_632 N_A_647_21#_c_820_n N_SET_B_M1004_g 0.020182f $X=3.42 $Y=1.74 $X2=0 $Y2=0
cc_633 N_A_647_21#_M1007_g N_SET_B_M1016_g 0.0145491f $X=3.31 $Y=0.445 $X2=0
+ $Y2=0
cc_634 N_A_647_21#_c_809_n N_SET_B_M1016_g 7.05788e-19 $X=4.6 $Y=1.065 $X2=0
+ $Y2=0
cc_635 N_A_647_21#_M1007_g SET_B 0.00110276f $X=3.31 $Y=0.445 $X2=0 $Y2=0
cc_636 N_A_647_21#_c_809_n SET_B 0.00825406f $X=4.6 $Y=1.065 $X2=0 $Y2=0
cc_637 N_A_647_21#_M1035_d N_SET_B_c_961_n 5.1491e-19 $X=4.435 $Y=0.235 $X2=0
+ $Y2=0
cc_638 N_A_647_21#_c_808_n N_SET_B_c_961_n 0.00519346f $X=5.72 $Y=0.985 $X2=0
+ $Y2=0
cc_639 N_A_647_21#_c_809_n N_SET_B_c_961_n 0.0208059f $X=4.6 $Y=1.065 $X2=0
+ $Y2=0
cc_640 N_A_647_21#_c_811_n N_SET_B_c_961_n 0.0211522f $X=5.495 $Y=0.98 $X2=0
+ $Y2=0
cc_641 N_A_647_21#_c_812_n N_SET_B_c_961_n 0.0109474f $X=5.66 $Y=0.98 $X2=0
+ $Y2=0
cc_642 N_A_647_21#_c_809_n N_SET_B_c_962_n 0.00230334f $X=4.6 $Y=1.065 $X2=0
+ $Y2=0
cc_643 N_A_647_21#_c_809_n N_A_473_413#_M1035_g 0.00718524f $X=4.6 $Y=1.065
+ $X2=0 $Y2=0
cc_644 N_A_647_21#_c_810_n N_A_473_413#_M1035_g 0.00191659f $X=4.6 $Y=1.785
+ $X2=0 $Y2=0
cc_645 N_A_647_21#_c_832_n N_A_473_413#_M1024_g 0.0126303f $X=4.515 $Y=1.91
+ $X2=0 $Y2=0
cc_646 N_A_647_21#_M1023_g N_A_473_413#_c_1097_n 0.00191115f $X=3.31 $Y=2.275
+ $X2=0 $Y2=0
cc_647 N_A_647_21#_M1007_g N_A_473_413#_c_1098_n 0.00854236f $X=3.31 $Y=0.445
+ $X2=0 $Y2=0
cc_648 N_A_647_21#_M1007_g N_A_473_413#_c_1092_n 0.0154362f $X=3.31 $Y=0.445
+ $X2=0 $Y2=0
cc_649 N_A_647_21#_c_819_n N_A_473_413#_c_1092_n 0.0330453f $X=3.42 $Y=1.74
+ $X2=0 $Y2=0
cc_650 N_A_647_21#_M1007_g N_A_473_413#_c_1087_n 0.0188177f $X=3.31 $Y=0.445
+ $X2=0 $Y2=0
cc_651 N_A_647_21#_c_817_n N_A_473_413#_c_1088_n 0.0141289f $X=4.085 $Y=1.91
+ $X2=0 $Y2=0
cc_652 N_A_647_21#_c_832_n N_A_473_413#_c_1088_n 0.00218253f $X=4.515 $Y=1.91
+ $X2=0 $Y2=0
cc_653 N_A_647_21#_c_810_n N_A_473_413#_c_1088_n 0.0246731f $X=4.6 $Y=1.785
+ $X2=0 $Y2=0
cc_654 N_A_647_21#_c_837_n N_A_473_413#_c_1088_n 0.00650509f $X=4.17 $Y=1.87
+ $X2=0 $Y2=0
cc_655 N_A_647_21#_M1007_g N_A_473_413#_c_1089_n 0.0109165f $X=3.31 $Y=0.445
+ $X2=0 $Y2=0
cc_656 N_A_647_21#_c_819_n N_A_473_413#_c_1089_n 0.0169843f $X=3.42 $Y=1.74
+ $X2=0 $Y2=0
cc_657 N_A_647_21#_c_820_n N_A_473_413#_c_1089_n 0.0011995f $X=3.42 $Y=1.74
+ $X2=0 $Y2=0
cc_658 N_A_647_21#_c_810_n N_A_473_413#_c_1090_n 0.0092978f $X=4.6 $Y=1.785
+ $X2=0 $Y2=0
cc_659 N_A_647_21#_c_837_n N_A_473_413#_c_1090_n 9.09922e-19 $X=4.17 $Y=1.87
+ $X2=0 $Y2=0
cc_660 N_A_647_21#_c_809_n N_A_941_21#_M1031_g 0.00955091f $X=4.6 $Y=1.065 $X2=0
+ $Y2=0
cc_661 N_A_647_21#_c_810_n N_A_941_21#_M1031_g 0.00587629f $X=4.6 $Y=1.785 $X2=0
+ $Y2=0
cc_662 N_A_647_21#_c_811_n N_A_941_21#_M1031_g 0.00930678f $X=5.495 $Y=0.98
+ $X2=0 $Y2=0
cc_663 N_A_647_21#_c_812_n N_A_941_21#_M1031_g 0.00136887f $X=5.66 $Y=0.98 $X2=0
+ $Y2=0
cc_664 N_A_647_21#_c_813_n N_A_941_21#_M1031_g 0.00197459f $X=5.66 $Y=1.15 $X2=0
+ $Y2=0
cc_665 N_A_647_21#_M1028_g N_A_941_21#_M1018_g 0.0153539f $X=5.485 $Y=2.065
+ $X2=0 $Y2=0
cc_666 N_A_647_21#_c_832_n N_A_941_21#_M1018_g 0.00219889f $X=4.515 $Y=1.91
+ $X2=0 $Y2=0
cc_667 N_A_647_21#_c_810_n N_A_941_21#_M1018_g 0.00171343f $X=4.6 $Y=1.785 $X2=0
+ $Y2=0
cc_668 N_A_647_21#_M1028_g N_A_941_21#_c_1196_n 2.86505e-19 $X=5.485 $Y=2.065
+ $X2=0 $Y2=0
cc_669 N_A_647_21#_c_810_n N_A_941_21#_c_1196_n 0.0309285f $X=4.6 $Y=1.785 $X2=0
+ $Y2=0
cc_670 N_A_647_21#_c_811_n N_A_941_21#_c_1196_n 0.0205705f $X=5.495 $Y=0.98
+ $X2=0 $Y2=0
cc_671 N_A_647_21#_c_813_n N_A_941_21#_c_1196_n 0.00382982f $X=5.66 $Y=1.15
+ $X2=0 $Y2=0
cc_672 N_A_647_21#_c_811_n N_A_941_21#_c_1197_n 0.00594187f $X=5.495 $Y=0.98
+ $X2=0 $Y2=0
cc_673 N_A_647_21#_c_812_n N_A_941_21#_c_1197_n 7.54142e-19 $X=5.66 $Y=0.98
+ $X2=0 $Y2=0
cc_674 N_A_647_21#_c_813_n N_A_941_21#_c_1197_n 0.0166765f $X=5.66 $Y=1.15 $X2=0
+ $Y2=0
cc_675 N_A_647_21#_c_812_n N_A_941_21#_c_1209_n 9.59092e-19 $X=5.66 $Y=0.98
+ $X2=0 $Y2=0
cc_676 N_A_647_21#_c_813_n N_A_941_21#_c_1209_n 0.00358318f $X=5.66 $Y=1.15
+ $X2=0 $Y2=0
cc_677 N_A_647_21#_M1028_g N_A_941_21#_c_1210_n 0.0143059f $X=5.485 $Y=2.065
+ $X2=0 $Y2=0
cc_678 N_A_647_21#_c_811_n N_A_941_21#_c_1210_n 0.00760725f $X=5.495 $Y=0.98
+ $X2=0 $Y2=0
cc_679 N_A_647_21#_c_812_n N_A_941_21#_c_1210_n 0.0207118f $X=5.66 $Y=0.98 $X2=0
+ $Y2=0
cc_680 N_A_647_21#_c_813_n N_A_941_21#_c_1210_n 0.00632961f $X=5.66 $Y=1.15
+ $X2=0 $Y2=0
cc_681 N_A_647_21#_M1028_g N_A_1256_413#_c_1566_n 7.04843e-19 $X=5.485 $Y=2.065
+ $X2=0 $Y2=0
cc_682 N_A_647_21#_c_808_n N_A_1256_413#_c_1569_n 6.8835e-19 $X=5.72 $Y=0.985
+ $X2=0 $Y2=0
cc_683 N_A_647_21#_M1023_g N_VPWR_c_1762_n 0.00326498f $X=3.31 $Y=2.275 $X2=0
+ $Y2=0
cc_684 N_A_647_21#_c_817_n N_VPWR_c_1762_n 0.0124698f $X=4.085 $Y=1.91 $X2=0
+ $Y2=0
cc_685 N_A_647_21#_c_864_p N_VPWR_c_1762_n 0.00820313f $X=4.17 $Y=2.21 $X2=0
+ $Y2=0
cc_686 N_A_647_21#_c_819_n N_VPWR_c_1762_n 0.0125544f $X=3.42 $Y=1.74 $X2=0
+ $Y2=0
cc_687 N_A_647_21#_c_820_n N_VPWR_c_1762_n 7.62241e-19 $X=3.42 $Y=1.74 $X2=0
+ $Y2=0
cc_688 N_A_647_21#_M1028_g N_VPWR_c_1763_n 0.0163458f $X=5.485 $Y=2.065 $X2=0
+ $Y2=0
cc_689 N_A_647_21#_c_832_n N_VPWR_c_1763_n 0.0048929f $X=4.515 $Y=1.91 $X2=0
+ $Y2=0
cc_690 N_A_647_21#_c_817_n N_VPWR_c_1765_n 0.00474052f $X=4.085 $Y=1.91 $X2=0
+ $Y2=0
cc_691 N_A_647_21#_c_864_p N_VPWR_c_1765_n 0.00725778f $X=4.17 $Y=2.21 $X2=0
+ $Y2=0
cc_692 N_A_647_21#_c_832_n N_VPWR_c_1765_n 0.00598455f $X=4.515 $Y=1.91 $X2=0
+ $Y2=0
cc_693 N_A_647_21#_M1023_g N_VPWR_c_1771_n 0.00535335f $X=3.31 $Y=2.275 $X2=0
+ $Y2=0
cc_694 N_A_647_21#_c_819_n N_VPWR_c_1771_n 0.00111392f $X=3.42 $Y=1.74 $X2=0
+ $Y2=0
cc_695 N_A_647_21#_M1028_g N_VPWR_c_1772_n 0.00585385f $X=5.485 $Y=2.065 $X2=0
+ $Y2=0
cc_696 N_A_647_21#_M1004_d N_VPWR_c_1759_n 0.0031612f $X=3.915 $Y=2.065 $X2=0
+ $Y2=0
cc_697 N_A_647_21#_M1023_g N_VPWR_c_1759_n 0.00664368f $X=3.31 $Y=2.275 $X2=0
+ $Y2=0
cc_698 N_A_647_21#_M1028_g N_VPWR_c_1759_n 0.00762825f $X=5.485 $Y=2.065 $X2=0
+ $Y2=0
cc_699 N_A_647_21#_c_817_n N_VPWR_c_1759_n 0.00386836f $X=4.085 $Y=1.91 $X2=0
+ $Y2=0
cc_700 N_A_647_21#_c_864_p N_VPWR_c_1759_n 0.0029026f $X=4.17 $Y=2.21 $X2=0
+ $Y2=0
cc_701 N_A_647_21#_c_832_n N_VPWR_c_1759_n 0.00505387f $X=4.515 $Y=1.91 $X2=0
+ $Y2=0
cc_702 N_A_647_21#_c_819_n N_VPWR_c_1759_n 0.00128163f $X=3.42 $Y=1.74 $X2=0
+ $Y2=0
cc_703 N_A_647_21#_c_832_n A_891_329# 0.00339576f $X=4.515 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_704 N_A_647_21#_c_810_n A_891_329# 0.00178287f $X=4.6 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_705 N_A_647_21#_M1007_g N_VGND_c_2069_n 0.00361232f $X=3.31 $Y=0.445 $X2=0
+ $Y2=0
cc_706 N_A_647_21#_c_808_n N_VGND_c_2070_n 0.0113057f $X=5.72 $Y=0.985 $X2=0
+ $Y2=0
cc_707 N_A_647_21#_c_811_n N_VGND_c_2070_n 0.00440912f $X=5.495 $Y=0.98 $X2=0
+ $Y2=0
cc_708 N_A_647_21#_c_812_n N_VGND_c_2070_n 0.00379129f $X=5.66 $Y=0.98 $X2=0
+ $Y2=0
cc_709 N_A_647_21#_c_813_n N_VGND_c_2070_n 8.52393e-19 $X=5.66 $Y=1.15 $X2=0
+ $Y2=0
cc_710 N_A_647_21#_M1007_g N_VGND_c_2074_n 0.0035977f $X=3.31 $Y=0.445 $X2=0
+ $Y2=0
cc_711 N_A_647_21#_c_808_n N_VGND_c_2078_n 0.0046653f $X=5.72 $Y=0.985 $X2=0
+ $Y2=0
cc_712 N_A_647_21#_M1035_d N_VGND_c_2085_n 0.00178362f $X=4.435 $Y=0.235 $X2=0
+ $Y2=0
cc_713 N_A_647_21#_M1007_g N_VGND_c_2085_n 0.00580574f $X=3.31 $Y=0.445 $X2=0
+ $Y2=0
cc_714 N_A_647_21#_c_808_n N_VGND_c_2085_n 0.00486196f $X=5.72 $Y=0.985 $X2=0
+ $Y2=0
cc_715 N_A_647_21#_M1035_d N_A_791_47#_c_2257_n 0.0030477f $X=4.435 $Y=0.235
+ $X2=0 $Y2=0
cc_716 N_A_647_21#_c_809_n N_A_791_47#_c_2257_n 0.0147704f $X=4.6 $Y=1.065 $X2=0
+ $Y2=0
cc_717 N_A_647_21#_c_811_n N_A_791_47#_c_2257_n 0.00259503f $X=5.495 $Y=0.98
+ $X2=0 $Y2=0
cc_718 N_A_647_21#_c_808_n N_A_791_47#_c_2260_n 0.00441801f $X=5.72 $Y=0.985
+ $X2=0 $Y2=0
cc_719 N_A_647_21#_c_811_n N_A_791_47#_c_2260_n 0.0106429f $X=5.495 $Y=0.98
+ $X2=0 $Y2=0
cc_720 N_SET_B_c_954_n N_A_473_413#_M1035_g 0.00619508f $X=3.84 $Y=1.145 $X2=0
+ $Y2=0
cc_721 N_SET_B_M1016_g N_A_473_413#_M1035_g 0.0197608f $X=3.88 $Y=0.445 $X2=0
+ $Y2=0
cc_722 SET_B N_A_473_413#_M1035_g 0.00183601f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_723 N_SET_B_c_961_n N_A_473_413#_M1035_g 0.00491921f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_962_n N_A_473_413#_M1035_g 0.00134231f $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_725 N_SET_B_M1004_g N_A_473_413#_M1024_g 0.0228864f $X=3.84 $Y=2.275 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_954_n N_A_473_413#_c_1087_n 0.00216489f $X=3.84 $Y=1.145 $X2=0
+ $Y2=0
cc_727 N_SET_B_M1004_g N_A_473_413#_c_1087_n 6.04572e-19 $X=3.84 $Y=2.275 $X2=0
+ $Y2=0
cc_728 N_SET_B_M1016_g N_A_473_413#_c_1087_n 0.00182721f $X=3.88 $Y=0.445 $X2=0
+ $Y2=0
cc_729 SET_B N_A_473_413#_c_1087_n 0.0244028f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_730 N_SET_B_c_962_n N_A_473_413#_c_1087_n 0.00111115f $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_731 N_SET_B_c_954_n N_A_473_413#_c_1088_n 0.00310411f $X=3.84 $Y=1.145 $X2=0
+ $Y2=0
cc_732 N_SET_B_M1004_g N_A_473_413#_c_1088_n 0.0131452f $X=3.84 $Y=2.275 $X2=0
+ $Y2=0
cc_733 SET_B N_A_473_413#_c_1088_n 0.0245807f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_734 N_SET_B_c_961_n N_A_473_413#_c_1088_n 0.00270886f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_962_n N_A_473_413#_c_1088_n 6.67689e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_SET_B_M1004_g N_A_473_413#_c_1089_n 5.20457e-19 $X=3.84 $Y=2.275 $X2=0
+ $Y2=0
cc_737 N_SET_B_M1004_g N_A_473_413#_c_1090_n 0.021088f $X=3.84 $Y=2.275 $X2=0
+ $Y2=0
cc_738 N_SET_B_c_961_n N_A_941_21#_M1031_g 0.00317213f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_739 N_SET_B_c_961_n N_A_941_21#_c_1196_n 5.29205e-19 $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_740 N_SET_B_M1012_g N_A_941_21#_c_1208_n 0.00589111f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_741 N_SET_B_c_961_n N_A_941_21#_c_1208_n 0.050802f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_742 N_SET_B_c_963_n N_A_941_21#_c_1208_n 0.0133806f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_743 N_SET_B_M1012_g N_A_1415_315#_M1008_g 0.0122611f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_744 N_SET_B_M1009_g N_A_1415_315#_M1020_g 0.0204909f $X=7.7 $Y=0.445 $X2=0
+ $Y2=0
cc_745 N_SET_B_c_958_n N_A_1415_315#_M1020_g 0.0230585f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_746 N_SET_B_M1012_g N_A_1415_315#_M1020_g 0.0124819f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_961_n N_A_1415_315#_M1020_g 0.00460114f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_748 N_SET_B_c_964_n N_A_1415_315#_M1020_g 0.00643702f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_749 N_SET_B_M1012_g N_A_1415_315#_c_1377_n 0.0071072f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_750 N_SET_B_M1012_g N_A_1415_315#_c_1378_n 0.0197578f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_751 N_SET_B_M1012_g N_A_1415_315#_c_1379_n 0.0139289f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_752 N_SET_B_c_964_n N_A_1415_315#_c_1368_n 0.00739337f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_753 N_SET_B_M1009_g N_A_1415_315#_c_1401_n 4.79271e-19 $X=7.7 $Y=0.445 $X2=0
+ $Y2=0
cc_754 N_SET_B_c_963_n N_A_1415_315#_c_1401_n 6.38044e-19 $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_755 N_SET_B_c_964_n N_A_1415_315#_c_1401_n 0.00396857f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_756 N_SET_B_M1009_g N_A_1256_413#_M1025_g 0.0215737f $X=7.7 $Y=0.445 $X2=0
+ $Y2=0
cc_757 N_SET_B_c_958_n N_A_1256_413#_M1025_g 0.00161465f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_758 N_SET_B_c_964_n N_A_1256_413#_M1025_g 0.00277477f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_759 N_SET_B_M1012_g N_A_1256_413#_M1003_g 0.0286249f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_760 N_SET_B_c_961_n N_A_1256_413#_c_1569_n 0.0088488f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_SET_B_c_961_n N_A_1256_413#_c_1555_n 0.0168353f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_762 N_SET_B_c_963_n N_A_1256_413#_c_1555_n 4.07638e-19 $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_763 N_SET_B_c_964_n N_A_1256_413#_c_1555_n 0.0207849f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_764 N_SET_B_M1012_g N_A_1256_413#_c_1561_n 6.40011e-19 $X=7.755 $Y=2.275
+ $X2=0 $Y2=0
cc_765 N_SET_B_c_958_n N_A_1256_413#_c_1556_n 0.00480597f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_766 N_SET_B_M1012_g N_A_1256_413#_c_1556_n 0.0118761f $X=7.755 $Y=2.275 $X2=0
+ $Y2=0
cc_767 N_SET_B_c_961_n N_A_1256_413#_c_1556_n 0.00529578f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_768 N_SET_B_c_963_n N_A_1256_413#_c_1556_n 9.47842e-19 $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_769 N_SET_B_c_964_n N_A_1256_413#_c_1556_n 0.0364733f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_770 N_SET_B_c_958_n N_A_1256_413#_c_1558_n 0.00112625f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_771 N_SET_B_c_958_n N_A_1256_413#_c_1559_n 0.0215562f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_772 N_SET_B_M1004_g N_VPWR_c_1762_n 0.0094739f $X=3.84 $Y=2.275 $X2=0 $Y2=0
cc_773 N_SET_B_M1004_g N_VPWR_c_1765_n 0.00373914f $X=3.84 $Y=2.275 $X2=0 $Y2=0
cc_774 N_SET_B_M1012_g N_VPWR_c_1768_n 0.00368415f $X=7.755 $Y=2.275 $X2=0 $Y2=0
cc_775 N_SET_B_M1004_g N_VPWR_c_1759_n 0.00439789f $X=3.84 $Y=2.275 $X2=0 $Y2=0
cc_776 N_SET_B_M1012_g N_VPWR_c_1759_n 0.00455672f $X=7.755 $Y=2.275 $X2=0 $Y2=0
cc_777 N_SET_B_M1012_g N_VPWR_c_1780_n 0.00881438f $X=7.755 $Y=2.275 $X2=0 $Y2=0
cc_778 N_SET_B_c_961_n N_VGND_M1019_s 0.00213341f $X=7.515 $Y=0.85 $X2=0 $Y2=0
cc_779 N_SET_B_c_954_n N_VGND_c_2069_n 8.58768e-19 $X=3.84 $Y=1.145 $X2=0 $Y2=0
cc_780 N_SET_B_M1016_g N_VGND_c_2069_n 0.00289978f $X=3.88 $Y=0.445 $X2=0 $Y2=0
cc_781 SET_B N_VGND_c_2069_n 0.010979f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_782 N_SET_B_c_961_n N_VGND_c_2070_n 0.00429522f $X=7.515 $Y=0.85 $X2=0 $Y2=0
cc_783 N_SET_B_M1009_g N_VGND_c_2071_n 0.002969f $X=7.7 $Y=0.445 $X2=0 $Y2=0
cc_784 N_SET_B_c_958_n N_VGND_c_2071_n 4.17175e-19 $X=7.755 $Y=1.18 $X2=0 $Y2=0
cc_785 N_SET_B_c_961_n N_VGND_c_2071_n 0.00204623f $X=7.515 $Y=0.85 $X2=0 $Y2=0
cc_786 N_SET_B_c_963_n N_VGND_c_2071_n 3.2427e-19 $X=7.66 $Y=0.85 $X2=0 $Y2=0
cc_787 N_SET_B_c_964_n N_VGND_c_2071_n 0.0159382f $X=7.66 $Y=0.85 $X2=0 $Y2=0
cc_788 N_SET_B_M1016_g N_VGND_c_2076_n 0.00422832f $X=3.88 $Y=0.445 $X2=0 $Y2=0
cc_789 SET_B N_VGND_c_2076_n 0.00221313f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_790 N_SET_B_M1009_g N_VGND_c_2082_n 0.00423333f $X=7.7 $Y=0.445 $X2=0 $Y2=0
cc_791 N_SET_B_c_964_n N_VGND_c_2082_n 0.00222084f $X=7.66 $Y=0.85 $X2=0 $Y2=0
cc_792 N_SET_B_M1016_g N_VGND_c_2085_n 0.00587817f $X=3.88 $Y=0.445 $X2=0 $Y2=0
cc_793 N_SET_B_M1009_g N_VGND_c_2085_n 0.00588395f $X=7.7 $Y=0.445 $X2=0 $Y2=0
cc_794 SET_B N_VGND_c_2085_n 0.00214053f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_795 N_SET_B_c_961_n N_VGND_c_2085_n 0.167605f $X=7.515 $Y=0.85 $X2=0 $Y2=0
cc_796 N_SET_B_c_962_n N_VGND_c_2085_n 0.0147327f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_797 N_SET_B_c_963_n N_VGND_c_2085_n 0.0141435f $X=7.66 $Y=0.85 $X2=0 $Y2=0
cc_798 N_SET_B_c_964_n N_VGND_c_2085_n 0.00190444f $X=7.66 $Y=0.85 $X2=0 $Y2=0
cc_799 N_SET_B_c_961_n N_A_791_47#_M1016_d 0.00182666f $X=7.515 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_800 N_SET_B_c_962_n N_A_791_47#_M1016_d 6.76077e-19 $X=4.055 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_801 N_SET_B_c_961_n N_A_791_47#_M1031_d 0.00215149f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_802 N_SET_B_c_961_n N_A_791_47#_c_2257_n 0.00555941f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_803 N_SET_B_c_961_n N_A_791_47#_c_2260_n 0.00234876f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_804 N_SET_B_M1016_g N_A_791_47#_c_2267_n 0.00335852f $X=3.88 $Y=0.445 $X2=0
+ $Y2=0
cc_805 SET_B N_A_791_47#_c_2267_n 0.00237046f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_806 N_SET_B_c_961_n N_A_791_47#_c_2267_n 0.00393563f $X=7.515 $Y=0.85 $X2=0
+ $Y2=0
cc_807 N_SET_B_c_962_n N_A_791_47#_c_2267_n 0.00215379f $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_808 N_SET_B_c_961_n A_1159_47# 0.00377207f $X=7.515 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_809 N_SET_B_M1009_g N_A_1555_47#_c_2288_n 0.00400944f $X=7.7 $Y=0.445 $X2=0
+ $Y2=0
cc_810 N_SET_B_c_963_n N_A_1555_47#_c_2288_n 2.64311e-19 $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_811 N_SET_B_c_964_n N_A_1555_47#_c_2288_n 0.00324102f $X=7.66 $Y=0.85 $X2=0
+ $Y2=0
cc_812 N_A_473_413#_M1035_g N_A_941_21#_M1031_g 0.030629f $X=4.36 $Y=0.555 $X2=0
+ $Y2=0
cc_813 N_A_473_413#_M1024_g N_A_941_21#_M1018_g 0.0493171f $X=4.38 $Y=2.065
+ $X2=0 $Y2=0
cc_814 N_A_473_413#_c_1090_n N_A_941_21#_c_1197_n 0.0167931f $X=4.26 $Y=1.32
+ $X2=0 $Y2=0
cc_815 N_A_473_413#_M1024_g N_VPWR_c_1762_n 0.00136797f $X=4.38 $Y=2.065 $X2=0
+ $Y2=0
cc_816 N_A_473_413#_M1024_g N_VPWR_c_1765_n 0.00432313f $X=4.38 $Y=2.065 $X2=0
+ $Y2=0
cc_817 N_A_473_413#_c_1097_n N_VPWR_c_1771_n 0.0377433f $X=2.995 $Y=2.335 $X2=0
+ $Y2=0
cc_818 N_A_473_413#_M1021_d N_VPWR_c_1759_n 0.00173085f $X=2.365 $Y=2.065 $X2=0
+ $Y2=0
cc_819 N_A_473_413#_M1024_g N_VPWR_c_1759_n 0.00600471f $X=4.38 $Y=2.065 $X2=0
+ $Y2=0
cc_820 N_A_473_413#_c_1097_n N_VPWR_c_1759_n 0.0132511f $X=2.995 $Y=2.335 $X2=0
+ $Y2=0
cc_821 N_A_473_413#_c_1097_n N_A_381_47#_c_1949_n 0.0112063f $X=2.995 $Y=2.335
+ $X2=0 $Y2=0
cc_822 N_A_473_413#_c_1097_n A_557_413# 0.00858887f $X=2.995 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_823 N_A_473_413#_c_1092_n A_557_413# 0.00579571f $X=3.08 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_824 N_A_473_413#_c_1098_n N_VGND_c_2074_n 0.0549341f $X=3.245 $Y=0.365 $X2=0
+ $Y2=0
cc_825 N_A_473_413#_M1035_g N_VGND_c_2076_n 0.00357877f $X=4.36 $Y=0.555 $X2=0
+ $Y2=0
cc_826 N_A_473_413#_M1026_d N_VGND_c_2085_n 0.00251173f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_827 N_A_473_413#_M1035_g N_VGND_c_2085_n 0.00536866f $X=4.36 $Y=0.555 $X2=0
+ $Y2=0
cc_828 N_A_473_413#_c_1098_n N_VGND_c_2085_n 0.0218827f $X=3.245 $Y=0.365 $X2=0
+ $Y2=0
cc_829 N_A_473_413#_c_1098_n A_581_47# 0.00568226f $X=3.245 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_830 N_A_473_413#_M1035_g N_A_791_47#_c_2257_n 0.00821062f $X=4.36 $Y=0.555
+ $X2=0 $Y2=0
cc_831 N_A_473_413#_c_1088_n N_A_791_47#_c_2267_n 0.00116076f $X=4.095 $Y=1.32
+ $X2=0 $Y2=0
cc_832 N_A_473_413#_c_1090_n N_A_791_47#_c_2267_n 5.81529e-19 $X=4.26 $Y=1.32
+ $X2=0 $Y2=0
cc_833 N_A_941_21#_c_1208_n N_A_1415_315#_M1020_g 0.00413345f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_834 N_A_941_21#_c_1208_n N_A_1415_315#_c_1377_n 0.015309f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_835 N_A_941_21#_c_1208_n N_A_1415_315#_c_1378_n 0.00935182f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_836 N_A_941_21#_c_1208_n N_A_1415_315#_c_1379_n 0.010417f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_837 N_A_941_21#_c_1208_n N_A_1415_315#_c_1408_n 0.0095166f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_838 N_A_941_21#_M1005_g N_A_1415_315#_c_1368_n 0.0116118f $X=8.645 $Y=2.065
+ $X2=0 $Y2=0
cc_839 N_A_941_21#_M1032_g N_A_1415_315#_c_1368_n 0.005494f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_840 N_A_941_21#_c_1194_n N_A_1415_315#_c_1368_n 0.00526859f $X=9.055 $Y=0.84
+ $X2=0 $Y2=0
cc_841 N_A_941_21#_c_1204_n N_A_1415_315#_c_1368_n 0.00845921f $X=9.055 $Y=1.66
+ $X2=0 $Y2=0
cc_842 N_A_941_21#_c_1198_n N_A_1415_315#_c_1368_n 0.0322778f $X=8.912 $Y=1.252
+ $X2=0 $Y2=0
cc_843 N_A_941_21#_c_1199_n N_A_1415_315#_c_1368_n 0.0105487f $X=8.912 $Y=1.11
+ $X2=0 $Y2=0
cc_844 N_A_941_21#_c_1208_n N_A_1415_315#_c_1368_n 0.0258804f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_845 N_A_941_21#_c_1211_n N_A_1415_315#_c_1368_n 5.93104e-19 $X=8.94 $Y=1.53
+ $X2=0 $Y2=0
cc_846 N_A_941_21#_c_1200_n N_A_1415_315#_c_1368_n 0.00728565f $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_847 N_A_941_21#_M1029_s N_A_1415_315#_c_1382_n 0.00494817f $X=9.25 $Y=1.505
+ $X2=0 $Y2=0
cc_848 N_A_941_21#_M1005_g N_A_1415_315#_c_1382_n 0.0100735f $X=8.645 $Y=2.065
+ $X2=0 $Y2=0
cc_849 N_A_941_21#_c_1204_n N_A_1415_315#_c_1382_n 0.0212769f $X=9.055 $Y=1.66
+ $X2=0 $Y2=0
cc_850 N_A_941_21#_c_1205_n N_A_1415_315#_c_1382_n 0.0322624f $X=9.375 $Y=1.66
+ $X2=0 $Y2=0
cc_851 N_A_941_21#_c_1208_n N_A_1415_315#_c_1382_n 0.00594443f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_852 N_A_941_21#_c_1211_n N_A_1415_315#_c_1382_n 0.00170464f $X=8.94 $Y=1.53
+ $X2=0 $Y2=0
cc_853 N_A_941_21#_c_1200_n N_A_1415_315#_c_1382_n 8.52182e-19 $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_854 N_A_941_21#_c_1205_n N_A_1415_315#_c_1383_n 0.00840283f $X=9.375 $Y=1.66
+ $X2=0 $Y2=0
cc_855 N_A_941_21#_c_1208_n N_A_1415_315#_c_1384_n 0.00453864f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_856 N_A_941_21#_M1032_g N_A_1415_315#_c_1401_n 0.00391303f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_857 N_A_941_21#_c_1194_n N_A_1415_315#_c_1401_n 0.00580837f $X=9.055 $Y=0.84
+ $X2=0 $Y2=0
cc_858 N_A_941_21#_c_1195_n N_A_1415_315#_c_1401_n 0.00249642f $X=9.39 $Y=0.43
+ $X2=0 $Y2=0
cc_859 N_A_941_21#_c_1208_n N_A_1415_315#_c_1401_n 3.49044e-19 $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_860 N_A_941_21#_M1005_g N_A_1415_315#_c_1431_n 0.00266575f $X=8.645 $Y=2.065
+ $X2=0 $Y2=0
cc_861 N_A_941_21#_M1032_g N_A_1256_413#_M1025_g 0.0300558f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_862 N_A_941_21#_M1005_g N_A_1256_413#_M1003_g 0.0452334f $X=8.645 $Y=2.065
+ $X2=0 $Y2=0
cc_863 N_A_941_21#_c_1208_n N_A_1256_413#_M1003_g 0.00852621f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_864 N_A_941_21#_c_1208_n N_A_1256_413#_c_1561_n 0.021932f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_865 N_A_941_21#_c_1208_n N_A_1256_413#_c_1556_n 0.0219758f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_866 N_A_941_21#_c_1208_n N_A_1256_413#_c_1558_n 0.00733551f $X=8.795 $Y=1.53
+ $X2=0 $Y2=0
cc_867 N_A_941_21#_c_1200_n N_A_1256_413#_c_1558_n 2.05377e-19 $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_868 N_A_941_21#_M1032_g N_A_1256_413#_c_1559_n 0.00446489f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_869 N_A_941_21#_c_1200_n N_A_1256_413#_c_1559_n 0.0452334f $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_870 N_A_941_21#_c_1205_n N_RESET_B_M1029_g 0.00360287f $X=9.375 $Y=1.66 $X2=0
+ $Y2=0
cc_871 N_A_941_21#_c_1211_n N_RESET_B_M1029_g 0.00260155f $X=8.94 $Y=1.53 $X2=0
+ $Y2=0
cc_872 N_A_941_21#_c_1200_n N_RESET_B_M1029_g 0.00242743f $X=8.855 $Y=1.32 $X2=0
+ $Y2=0
cc_873 N_A_941_21#_c_1201_n N_RESET_B_M1029_g 0.00312031f $X=8.855 $Y=1.32 $X2=0
+ $Y2=0
cc_874 N_A_941_21#_c_1193_n N_RESET_B_M1015_g 0.00676877f $X=9.265 $Y=0.84 $X2=0
+ $Y2=0
cc_875 N_A_941_21#_c_1195_n N_RESET_B_M1015_g 0.00291288f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_876 N_A_941_21#_c_1199_n N_RESET_B_M1015_g 0.00229156f $X=8.912 $Y=1.11 $X2=0
+ $Y2=0
cc_877 N_A_941_21#_c_1193_n RESET_B 0.0195128f $X=9.265 $Y=0.84 $X2=0 $Y2=0
cc_878 N_A_941_21#_c_1205_n RESET_B 0.0155567f $X=9.375 $Y=1.66 $X2=0 $Y2=0
cc_879 N_A_941_21#_c_1199_n RESET_B 0.0184648f $X=8.912 $Y=1.11 $X2=0 $Y2=0
cc_880 N_A_941_21#_c_1200_n RESET_B 5.44868e-19 $X=8.855 $Y=1.32 $X2=0 $Y2=0
cc_881 N_A_941_21#_M1032_g N_RESET_B_c_1668_n 0.00208799f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_882 N_A_941_21#_c_1193_n N_RESET_B_c_1668_n 0.00537728f $X=9.265 $Y=0.84
+ $X2=0 $Y2=0
cc_883 N_A_941_21#_c_1205_n N_RESET_B_c_1668_n 0.00527649f $X=9.375 $Y=1.66
+ $X2=0 $Y2=0
cc_884 N_A_941_21#_c_1199_n N_RESET_B_c_1668_n 0.0027306f $X=8.912 $Y=1.11 $X2=0
+ $Y2=0
cc_885 N_A_941_21#_c_1200_n N_RESET_B_c_1668_n 0.00881374f $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_886 N_A_941_21#_c_1201_n N_RESET_B_c_1668_n 4.73172e-19 $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_887 N_A_941_21#_c_1196_n N_VPWR_M1018_d 0.00297048f $X=5.02 $Y=1.32 $X2=0
+ $Y2=0
cc_888 N_A_941_21#_c_1210_n N_VPWR_M1018_d 0.00221014f $X=5.75 $Y=1.53 $X2=0
+ $Y2=0
cc_889 N_A_941_21#_c_1204_n N_VPWR_M1005_d 0.00308033f $X=9.055 $Y=1.66 $X2=0
+ $Y2=0
cc_890 N_A_941_21#_M1018_g N_VPWR_c_1763_n 0.00353361f $X=4.8 $Y=2.065 $X2=0
+ $Y2=0
cc_891 N_A_941_21#_c_1196_n N_VPWR_c_1763_n 0.011531f $X=5.02 $Y=1.32 $X2=0
+ $Y2=0
cc_892 N_A_941_21#_c_1197_n N_VPWR_c_1763_n 0.00111411f $X=5.02 $Y=1.32 $X2=0
+ $Y2=0
cc_893 N_A_941_21#_c_1210_n N_VPWR_c_1763_n 7.83548e-19 $X=5.75 $Y=1.53 $X2=0
+ $Y2=0
cc_894 N_A_941_21#_M1018_g N_VPWR_c_1765_n 0.00583607f $X=4.8 $Y=2.065 $X2=0
+ $Y2=0
cc_895 N_A_941_21#_M1005_g N_VPWR_c_1767_n 0.0140513f $X=8.645 $Y=2.065 $X2=0
+ $Y2=0
cc_896 N_A_941_21#_M1005_g N_VPWR_c_1768_n 0.00197639f $X=8.645 $Y=2.065 $X2=0
+ $Y2=0
cc_897 N_A_941_21#_M1018_g N_VPWR_c_1759_n 0.00670824f $X=4.8 $Y=2.065 $X2=0
+ $Y2=0
cc_898 N_A_941_21#_M1005_g N_VPWR_c_1759_n 0.00248516f $X=8.645 $Y=2.065 $X2=0
+ $Y2=0
cc_899 N_A_941_21#_c_1210_n A_1112_329# 0.00272182f $X=5.75 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_900 N_A_941_21#_M1031_g N_VGND_c_2070_n 0.00327939f $X=4.78 $Y=0.555 $X2=0
+ $Y2=0
cc_901 N_A_941_21#_c_1193_n N_VGND_c_2072_n 0.00333537f $X=9.265 $Y=0.84 $X2=0
+ $Y2=0
cc_902 N_A_941_21#_c_1195_n N_VGND_c_2072_n 0.00601533f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_903 N_A_941_21#_M1031_g N_VGND_c_2076_n 0.00357877f $X=4.78 $Y=0.555 $X2=0
+ $Y2=0
cc_904 N_A_941_21#_M1032_g N_VGND_c_2082_n 0.00357877f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_905 N_A_941_21#_c_1193_n N_VGND_c_2082_n 0.00300947f $X=9.265 $Y=0.84 $X2=0
+ $Y2=0
cc_906 N_A_941_21#_c_1194_n N_VGND_c_2082_n 0.00158839f $X=9.055 $Y=0.84 $X2=0
+ $Y2=0
cc_907 N_A_941_21#_c_1195_n N_VGND_c_2082_n 0.0135199f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_908 N_A_941_21#_M1015_s N_VGND_c_2085_n 0.00382354f $X=9.265 $Y=0.235 $X2=0
+ $Y2=0
cc_909 N_A_941_21#_M1031_g N_VGND_c_2085_n 0.00661646f $X=4.78 $Y=0.555 $X2=0
+ $Y2=0
cc_910 N_A_941_21#_M1032_g N_VGND_c_2085_n 0.00657948f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_911 N_A_941_21#_c_1193_n N_VGND_c_2085_n 0.00541125f $X=9.265 $Y=0.84 $X2=0
+ $Y2=0
cc_912 N_A_941_21#_c_1194_n N_VGND_c_2085_n 0.00302863f $X=9.055 $Y=0.84 $X2=0
+ $Y2=0
cc_913 N_A_941_21#_c_1195_n N_VGND_c_2085_n 0.00796608f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_914 N_A_941_21#_M1031_g N_A_791_47#_c_2257_n 0.0105472f $X=4.78 $Y=0.555
+ $X2=0 $Y2=0
cc_915 N_A_941_21#_c_1194_n N_A_1555_47#_M1032_d 0.0043423f $X=9.055 $Y=0.84
+ $X2=0 $Y2=0
cc_916 N_A_941_21#_M1032_g N_A_1555_47#_c_2292_n 0.0112959f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_917 N_A_941_21#_c_1194_n N_A_1555_47#_c_2293_n 0.00983417f $X=9.055 $Y=0.84
+ $X2=0 $Y2=0
cc_918 N_A_941_21#_c_1195_n N_A_1555_47#_c_2293_n 0.0151854f $X=9.39 $Y=0.43
+ $X2=0 $Y2=0
cc_919 N_A_941_21#_c_1198_n N_A_1555_47#_c_2293_n 0.00178436f $X=8.912 $Y=1.252
+ $X2=0 $Y2=0
cc_920 N_A_941_21#_c_1200_n N_A_1555_47#_c_2293_n 6.33841e-19 $X=8.855 $Y=1.32
+ $X2=0 $Y2=0
cc_921 N_A_1415_315#_c_1368_n N_A_1256_413#_M1025_g 0.00253508f $X=8.515
+ $Y=1.915 $X2=0 $Y2=0
cc_922 N_A_1415_315#_c_1401_n N_A_1256_413#_M1025_g 0.00857144f $X=8.45 $Y=0.75
+ $X2=0 $Y2=0
cc_923 N_A_1415_315#_c_1408_n N_A_1256_413#_M1003_g 0.0117409f $X=8.43 $Y=2
+ $X2=0 $Y2=0
cc_924 N_A_1415_315#_M1008_g N_A_1256_413#_c_1566_n 0.00437824f $X=7.15 $Y=2.275
+ $X2=0 $Y2=0
cc_925 N_A_1415_315#_M1020_g N_A_1256_413#_c_1569_n 0.0017146f $X=7.215 $Y=0.445
+ $X2=0 $Y2=0
cc_926 N_A_1415_315#_M1020_g N_A_1256_413#_c_1555_n 0.011896f $X=7.215 $Y=0.445
+ $X2=0 $Y2=0
cc_927 N_A_1415_315#_M1008_g N_A_1256_413#_c_1561_n 0.00792191f $X=7.15 $Y=2.275
+ $X2=0 $Y2=0
cc_928 N_A_1415_315#_M1020_g N_A_1256_413#_c_1561_n 0.00587016f $X=7.215
+ $Y=0.445 $X2=0 $Y2=0
cc_929 N_A_1415_315#_c_1377_n N_A_1256_413#_c_1561_n 0.0235931f $X=7.335 $Y=1.74
+ $X2=0 $Y2=0
cc_930 N_A_1415_315#_c_1378_n N_A_1256_413#_c_1561_n 0.00710752f $X=7.335
+ $Y=1.74 $X2=0 $Y2=0
cc_931 N_A_1415_315#_c_1380_n N_A_1256_413#_c_1561_n 0.0127349f $X=7.5 $Y=2
+ $X2=0 $Y2=0
cc_932 N_A_1415_315#_M1020_g N_A_1256_413#_c_1556_n 0.0114629f $X=7.215 $Y=0.445
+ $X2=0 $Y2=0
cc_933 N_A_1415_315#_c_1377_n N_A_1256_413#_c_1556_n 0.0154844f $X=7.335 $Y=1.74
+ $X2=0 $Y2=0
cc_934 N_A_1415_315#_c_1378_n N_A_1256_413#_c_1556_n 0.00327097f $X=7.335
+ $Y=1.74 $X2=0 $Y2=0
cc_935 N_A_1415_315#_c_1379_n N_A_1256_413#_c_1556_n 0.00638264f $X=7.94 $Y=2
+ $X2=0 $Y2=0
cc_936 N_A_1415_315#_c_1384_n N_A_1256_413#_c_1556_n 0.00164491f $X=8.025 $Y=2
+ $X2=0 $Y2=0
cc_937 N_A_1415_315#_c_1408_n N_A_1256_413#_c_1558_n 0.00157994f $X=8.43 $Y=2
+ $X2=0 $Y2=0
cc_938 N_A_1415_315#_c_1368_n N_A_1256_413#_c_1558_n 0.0240523f $X=8.515
+ $Y=1.915 $X2=0 $Y2=0
cc_939 N_A_1415_315#_c_1384_n N_A_1256_413#_c_1558_n 0.00106299f $X=8.025 $Y=2
+ $X2=0 $Y2=0
cc_940 N_A_1415_315#_c_1401_n N_A_1256_413#_c_1558_n 0.00240462f $X=8.45 $Y=0.75
+ $X2=0 $Y2=0
cc_941 N_A_1415_315#_c_1408_n N_A_1256_413#_c_1559_n 3.5483e-19 $X=8.43 $Y=2
+ $X2=0 $Y2=0
cc_942 N_A_1415_315#_c_1368_n N_A_1256_413#_c_1559_n 0.0130958f $X=8.515
+ $Y=1.915 $X2=0 $Y2=0
cc_943 N_A_1415_315#_c_1384_n N_A_1256_413#_c_1559_n 4.29792e-19 $X=8.025 $Y=2
+ $X2=0 $Y2=0
cc_944 N_A_1415_315#_M1039_g N_RESET_B_M1029_g 0.0287825f $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_945 N_A_1415_315#_c_1382_n N_RESET_B_M1029_g 0.0142369f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_946 N_A_1415_315#_c_1383_n N_RESET_B_M1029_g 0.00948427f $X=9.945 $Y=1.915
+ $X2=0 $Y2=0
cc_947 N_A_1415_315#_c_1360_n N_RESET_B_M1015_g 0.0198209f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_948 N_A_1415_315#_c_1362_n N_RESET_B_M1015_g 0.0189873f $X=10.175 $Y=1.16
+ $X2=0 $Y2=0
cc_949 N_A_1415_315#_c_1369_n N_RESET_B_M1015_g 0.00222119f $X=10.04 $Y=1.16
+ $X2=0 $Y2=0
cc_950 N_A_1415_315#_c_1362_n RESET_B 7.20757e-19 $X=10.175 $Y=1.16 $X2=0 $Y2=0
cc_951 N_A_1415_315#_c_1382_n RESET_B 0.0031078f $X=9.86 $Y=2 $X2=0 $Y2=0
cc_952 N_A_1415_315#_c_1369_n RESET_B 0.0193191f $X=10.04 $Y=1.16 $X2=0 $Y2=0
cc_953 N_A_1415_315#_M1039_g N_RESET_B_c_1668_n 6.94565e-19 $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_954 N_A_1415_315#_c_1383_n N_RESET_B_c_1668_n 4.34361e-19 $X=9.945 $Y=1.915
+ $X2=0 $Y2=0
cc_955 N_A_1415_315#_c_1369_n N_RESET_B_c_1668_n 7.06091e-19 $X=10.04 $Y=1.16
+ $X2=0 $Y2=0
cc_956 N_A_1415_315#_c_1364_n N_A_2136_47#_M1037_g 0.0046261f $X=10.89 $Y=1.535
+ $X2=0 $Y2=0
cc_957 N_A_1415_315#_c_1376_n N_A_2136_47#_M1037_g 0.0111659f $X=11.015 $Y=1.61
+ $X2=0 $Y2=0
cc_958 N_A_1415_315#_c_1360_n N_A_2136_47#_c_1705_n 0.00110305f $X=10.075
+ $Y=0.995 $X2=0 $Y2=0
cc_959 N_A_1415_315#_c_1363_n N_A_2136_47#_c_1705_n 0.00388761f $X=10.89
+ $Y=1.025 $X2=0 $Y2=0
cc_960 N_A_1415_315#_c_1365_n N_A_2136_47#_c_1705_n 0.00981326f $X=11.015
+ $Y=0.73 $X2=0 $Y2=0
cc_961 N_A_1415_315#_c_1366_n N_A_2136_47#_c_1705_n 0.00979941f $X=11.015
+ $Y=0.805 $X2=0 $Y2=0
cc_962 N_A_1415_315#_M1039_g N_A_2136_47#_c_1711_n 0.00166592f $X=10.075
+ $Y=1.985 $X2=0 $Y2=0
cc_963 N_A_1415_315#_c_1364_n N_A_2136_47#_c_1711_n 0.00715595f $X=10.89
+ $Y=1.535 $X2=0 $Y2=0
cc_964 N_A_1415_315#_c_1375_n N_A_2136_47#_c_1711_n 0.0108344f $X=11.015
+ $Y=1.685 $X2=0 $Y2=0
cc_965 N_A_1415_315#_c_1376_n N_A_2136_47#_c_1711_n 0.0101822f $X=11.015 $Y=1.61
+ $X2=0 $Y2=0
cc_966 N_A_1415_315#_c_1366_n N_A_2136_47#_c_1706_n 0.00368279f $X=11.015
+ $Y=0.805 $X2=0 $Y2=0
cc_967 N_A_1415_315#_c_1376_n N_A_2136_47#_c_1706_n 0.00324612f $X=11.015
+ $Y=1.61 $X2=0 $Y2=0
cc_968 N_A_1415_315#_c_1363_n N_A_2136_47#_c_1707_n 0.0131369f $X=10.89 $Y=1.025
+ $X2=0 $Y2=0
cc_969 N_A_1415_315#_c_1361_n N_A_2136_47#_c_1708_n 0.0133077f $X=10.815 $Y=1.16
+ $X2=0 $Y2=0
cc_970 N_A_1415_315#_c_1363_n N_A_2136_47#_c_1708_n 0.00116339f $X=10.89
+ $Y=1.025 $X2=0 $Y2=0
cc_971 N_A_1415_315#_c_1364_n N_A_2136_47#_c_1708_n 0.00115562f $X=10.89
+ $Y=1.535 $X2=0 $Y2=0
cc_972 N_A_1415_315#_c_1367_n N_A_2136_47#_c_1708_n 0.00732445f $X=10.89 $Y=1.16
+ $X2=0 $Y2=0
cc_973 N_A_1415_315#_c_1363_n N_A_2136_47#_c_1709_n 0.0025256f $X=10.89 $Y=1.025
+ $X2=0 $Y2=0
cc_974 N_A_1415_315#_c_1365_n N_A_2136_47#_c_1709_n 0.0159526f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_975 N_A_1415_315#_c_1379_n N_VPWR_M1008_d 0.00124767f $X=7.94 $Y=2 $X2=0
+ $Y2=0
cc_976 N_A_1415_315#_c_1380_n N_VPWR_M1008_d 0.00256616f $X=7.5 $Y=2 $X2=0 $Y2=0
cc_977 N_A_1415_315#_c_1382_n N_VPWR_M1005_d 0.00457725f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_978 N_A_1415_315#_c_1382_n N_VPWR_M1029_d 0.00750664f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_979 N_A_1415_315#_c_1383_n N_VPWR_M1029_d 0.00487804f $X=9.945 $Y=1.915 $X2=0
+ $Y2=0
cc_980 N_A_1415_315#_c_1375_n N_VPWR_c_1764_n 0.00446368f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_981 N_A_1415_315#_c_1492_p N_VPWR_c_1767_n 0.00381845f $X=8.025 $Y=2.21 $X2=0
+ $Y2=0
cc_982 N_A_1415_315#_c_1382_n N_VPWR_c_1767_n 0.0840218f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_983 N_A_1415_315#_c_1379_n N_VPWR_c_1768_n 0.00359839f $X=7.94 $Y=2 $X2=0
+ $Y2=0
cc_984 N_A_1415_315#_c_1492_p N_VPWR_c_1768_n 0.00725596f $X=8.025 $Y=2.21 $X2=0
+ $Y2=0
cc_985 N_A_1415_315#_c_1408_n N_VPWR_c_1768_n 0.00452819f $X=8.43 $Y=2 $X2=0
+ $Y2=0
cc_986 N_A_1415_315#_c_1382_n N_VPWR_c_1768_n 6.38179e-19 $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_987 N_A_1415_315#_c_1431_n N_VPWR_c_1768_n 0.00268434f $X=8.515 $Y=2 $X2=0
+ $Y2=0
cc_988 N_A_1415_315#_M1008_g N_VPWR_c_1772_n 0.00578102f $X=7.15 $Y=2.275 $X2=0
+ $Y2=0
cc_989 N_A_1415_315#_c_1380_n N_VPWR_c_1772_n 0.00103314f $X=7.5 $Y=2 $X2=0
+ $Y2=0
cc_990 N_A_1415_315#_M1039_g N_VPWR_c_1774_n 0.0046653f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_991 N_A_1415_315#_c_1375_n N_VPWR_c_1774_n 0.00464873f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_992 N_A_1415_315#_M1012_d N_VPWR_c_1759_n 0.00385648f $X=7.83 $Y=2.065 $X2=0
+ $Y2=0
cc_993 N_A_1415_315#_M1008_g N_VPWR_c_1759_n 0.0113228f $X=7.15 $Y=2.275 $X2=0
+ $Y2=0
cc_994 N_A_1415_315#_M1039_g N_VPWR_c_1759_n 0.00929621f $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_995 N_A_1415_315#_c_1375_n N_VPWR_c_1759_n 0.00924075f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_996 N_A_1415_315#_c_1378_n N_VPWR_c_1759_n 6.58877e-19 $X=7.335 $Y=1.74 $X2=0
+ $Y2=0
cc_997 N_A_1415_315#_c_1379_n N_VPWR_c_1759_n 0.00704318f $X=7.94 $Y=2 $X2=0
+ $Y2=0
cc_998 N_A_1415_315#_c_1380_n N_VPWR_c_1759_n 0.00300249f $X=7.5 $Y=2 $X2=0
+ $Y2=0
cc_999 N_A_1415_315#_c_1492_p N_VPWR_c_1759_n 0.00608739f $X=8.025 $Y=2.21 $X2=0
+ $Y2=0
cc_1000 N_A_1415_315#_c_1408_n N_VPWR_c_1759_n 0.00829558f $X=8.43 $Y=2 $X2=0
+ $Y2=0
cc_1001 N_A_1415_315#_c_1382_n N_VPWR_c_1759_n 0.00710897f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_1002 N_A_1415_315#_c_1431_n N_VPWR_c_1759_n 0.00494768f $X=8.515 $Y=2 $X2=0
+ $Y2=0
cc_1003 N_A_1415_315#_M1008_g N_VPWR_c_1780_n 0.00635699f $X=7.15 $Y=2.275 $X2=0
+ $Y2=0
cc_1004 N_A_1415_315#_c_1378_n N_VPWR_c_1780_n 7.54485e-19 $X=7.335 $Y=1.74
+ $X2=0 $Y2=0
cc_1005 N_A_1415_315#_c_1379_n N_VPWR_c_1780_n 0.0106677f $X=7.94 $Y=2 $X2=0
+ $Y2=0
cc_1006 N_A_1415_315#_c_1380_n N_VPWR_c_1780_n 0.0147832f $X=7.5 $Y=2 $X2=0
+ $Y2=0
cc_1007 N_A_1415_315#_c_1492_p N_VPWR_c_1780_n 0.00687131f $X=8.025 $Y=2.21
+ $X2=0 $Y2=0
cc_1008 N_A_1415_315#_M1039_g N_VPWR_c_1781_n 0.0100464f $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_1009 N_A_1415_315#_c_1382_n N_VPWR_c_1781_n 0.00915613f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_1010 N_A_1415_315#_c_1408_n A_1672_329# 3.91203e-19 $X=8.43 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1011 N_A_1415_315#_c_1368_n A_1672_329# 0.00296763f $X=8.515 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1012 N_A_1415_315#_c_1431_n A_1672_329# 0.00149905f $X=8.515 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1013 N_A_1415_315#_c_1361_n N_Q_N_c_2021_n 0.00383478f $X=10.815 $Y=1.16
+ $X2=0 $Y2=0
cc_1014 N_A_1415_315#_c_1375_n N_Q_N_c_2021_n 0.00131217f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_1015 N_A_1415_315#_c_1376_n N_Q_N_c_2021_n 5.75727e-19 $X=11.015 $Y=1.61
+ $X2=0 $Y2=0
cc_1016 N_A_1415_315#_c_1360_n N_Q_N_c_2018_n 0.00547914f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1017 N_A_1415_315#_M1039_g N_Q_N_c_2018_n 0.00269981f $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_1018 N_A_1415_315#_c_1361_n N_Q_N_c_2018_n 0.0206804f $X=10.815 $Y=1.16 $X2=0
+ $Y2=0
cc_1019 N_A_1415_315#_c_1362_n N_Q_N_c_2018_n 3.3844e-19 $X=10.175 $Y=1.16 $X2=0
+ $Y2=0
cc_1020 N_A_1415_315#_c_1364_n N_Q_N_c_2018_n 5.75727e-19 $X=10.89 $Y=1.535
+ $X2=0 $Y2=0
cc_1021 N_A_1415_315#_c_1366_n N_Q_N_c_2018_n 8.63605e-19 $X=11.015 $Y=0.805
+ $X2=0 $Y2=0
cc_1022 N_A_1415_315#_c_1383_n N_Q_N_c_2018_n 0.0126467f $X=9.945 $Y=1.915 $X2=0
+ $Y2=0
cc_1023 N_A_1415_315#_c_1369_n N_Q_N_c_2018_n 0.0224114f $X=10.04 $Y=1.16 $X2=0
+ $Y2=0
cc_1024 N_A_1415_315#_c_1361_n Q_N 0.00230535f $X=10.815 $Y=1.16 $X2=0 $Y2=0
cc_1025 N_A_1415_315#_c_1375_n Q_N 8.70693e-19 $X=11.015 $Y=1.685 $X2=0 $Y2=0
cc_1026 N_A_1415_315#_c_1365_n N_Q_N_c_2020_n 0.00104845f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_1027 N_A_1415_315#_M1020_g N_VGND_c_2071_n 0.0126997f $X=7.215 $Y=0.445 $X2=0
+ $Y2=0
cc_1028 N_A_1415_315#_c_1360_n N_VGND_c_2072_n 0.015252f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1029 N_A_1415_315#_c_1362_n N_VGND_c_2072_n 0.00200592f $X=10.175 $Y=1.16
+ $X2=0 $Y2=0
cc_1030 N_A_1415_315#_c_1369_n N_VGND_c_2072_n 0.0105583f $X=10.04 $Y=1.16 $X2=0
+ $Y2=0
cc_1031 N_A_1415_315#_c_1365_n N_VGND_c_2073_n 0.00418537f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_1032 N_A_1415_315#_M1020_g N_VGND_c_2078_n 0.00427505f $X=7.215 $Y=0.445
+ $X2=0 $Y2=0
cc_1033 N_A_1415_315#_c_1360_n N_VGND_c_2083_n 0.0046653f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1034 N_A_1415_315#_c_1365_n N_VGND_c_2083_n 0.00533769f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_1035 N_A_1415_315#_c_1366_n N_VGND_c_2083_n 2.84936e-19 $X=11.015 $Y=0.805
+ $X2=0 $Y2=0
cc_1036 N_A_1415_315#_M1025_d N_VGND_c_2085_n 0.00216833f $X=8.315 $Y=0.235
+ $X2=0 $Y2=0
cc_1037 N_A_1415_315#_M1020_g N_VGND_c_2085_n 0.00427939f $X=7.215 $Y=0.445
+ $X2=0 $Y2=0
cc_1038 N_A_1415_315#_c_1360_n N_VGND_c_2085_n 0.00934473f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1039 N_A_1415_315#_c_1365_n N_VGND_c_2085_n 0.0109143f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_1040 N_A_1415_315#_M1025_d N_A_1555_47#_c_2292_n 0.00339796f $X=8.315
+ $Y=0.235 $X2=0 $Y2=0
cc_1041 N_A_1415_315#_c_1401_n N_A_1555_47#_c_2292_n 0.0146622f $X=8.45 $Y=0.75
+ $X2=0 $Y2=0
cc_1042 N_A_1415_315#_M1020_g N_A_1555_47#_c_2288_n 2.56899e-19 $X=7.215
+ $Y=0.445 $X2=0 $Y2=0
cc_1043 N_A_1256_413#_M1003_g N_VPWR_c_1767_n 0.00231807f $X=8.285 $Y=2.065
+ $X2=0 $Y2=0
cc_1044 N_A_1256_413#_M1003_g N_VPWR_c_1768_n 0.00425094f $X=8.285 $Y=2.065
+ $X2=0 $Y2=0
cc_1045 N_A_1256_413#_c_1566_n N_VPWR_c_1772_n 0.0362326f $X=6.91 $Y=2.335 $X2=0
+ $Y2=0
cc_1046 N_A_1256_413#_M1034_d N_VPWR_c_1759_n 0.00205544f $X=6.28 $Y=2.065 $X2=0
+ $Y2=0
cc_1047 N_A_1256_413#_M1003_g N_VPWR_c_1759_n 0.00602674f $X=8.285 $Y=2.065
+ $X2=0 $Y2=0
cc_1048 N_A_1256_413#_c_1566_n N_VPWR_c_1759_n 0.0272569f $X=6.91 $Y=2.335 $X2=0
+ $Y2=0
cc_1049 N_A_1256_413#_M1003_g N_VPWR_c_1780_n 0.0013585f $X=8.285 $Y=2.065 $X2=0
+ $Y2=0
cc_1050 N_A_1256_413#_c_1566_n N_VPWR_c_1780_n 0.0105242f $X=6.91 $Y=2.335 $X2=0
+ $Y2=0
cc_1051 N_A_1256_413#_c_1566_n A_1340_413# 0.0071257f $X=6.91 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1052 N_A_1256_413#_c_1561_n A_1340_413# 0.00219581f $X=6.995 $Y=2.25
+ $X2=-0.19 $Y2=-0.24
cc_1053 N_A_1256_413#_c_1569_n N_VGND_c_2070_n 0.00536652f $X=6.91 $Y=0.365
+ $X2=0 $Y2=0
cc_1054 N_A_1256_413#_c_1569_n N_VGND_c_2071_n 0.0164982f $X=6.91 $Y=0.365 $X2=0
+ $Y2=0
cc_1055 N_A_1256_413#_c_1555_n N_VGND_c_2071_n 0.0043886f $X=6.995 $Y=1.235
+ $X2=0 $Y2=0
cc_1056 N_A_1256_413#_c_1569_n N_VGND_c_2078_n 0.0428541f $X=6.91 $Y=0.365 $X2=0
+ $Y2=0
cc_1057 N_A_1256_413#_M1025_g N_VGND_c_2082_n 0.00357877f $X=8.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1058 N_A_1256_413#_M1001_d N_VGND_c_2085_n 0.00177273f $X=6.395 $Y=0.235
+ $X2=0 $Y2=0
cc_1059 N_A_1256_413#_M1025_g N_VGND_c_2085_n 0.00559748f $X=8.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1060 N_A_1256_413#_c_1569_n N_VGND_c_2085_n 0.0129387f $X=6.91 $Y=0.365 $X2=0
+ $Y2=0
cc_1061 N_A_1256_413#_c_1569_n A_1363_47# 0.00516586f $X=6.91 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1062 N_A_1256_413#_c_1555_n A_1363_47# 0.00492562f $X=6.995 $Y=1.235
+ $X2=-0.19 $Y2=-0.24
cc_1063 N_A_1256_413#_M1025_g N_A_1555_47#_c_2292_n 0.00998936f $X=8.24 $Y=0.555
+ $X2=0 $Y2=0
cc_1064 N_A_1256_413#_c_1558_n N_A_1555_47#_c_2292_n 0.00271489f $X=8.175
+ $Y=1.24 $X2=0 $Y2=0
cc_1065 N_A_1256_413#_c_1559_n N_A_1555_47#_c_2292_n 2.62935e-19 $X=8.175
+ $Y=1.24 $X2=0 $Y2=0
cc_1066 N_A_1256_413#_M1025_g N_A_1555_47#_c_2288_n 0.00363416f $X=8.24 $Y=0.555
+ $X2=0 $Y2=0
cc_1067 N_A_1256_413#_c_1555_n N_A_1555_47#_c_2288_n 4.9689e-19 $X=6.995
+ $Y=1.235 $X2=0 $Y2=0
cc_1068 N_A_1256_413#_c_1558_n N_A_1555_47#_c_2288_n 0.00105031f $X=8.175
+ $Y=1.24 $X2=0 $Y2=0
cc_1069 N_RESET_B_M1029_g N_VPWR_c_1773_n 0.00655753f $X=9.59 $Y=1.825 $X2=0
+ $Y2=0
cc_1070 N_RESET_B_M1015_g N_VGND_c_2072_n 0.00472624f $X=9.6 $Y=0.445 $X2=0
+ $Y2=0
cc_1071 N_RESET_B_M1015_g N_VGND_c_2082_n 0.00585385f $X=9.6 $Y=0.445 $X2=0
+ $Y2=0
cc_1072 N_RESET_B_M1015_g N_VGND_c_2085_n 0.0120198f $X=9.6 $Y=0.445 $X2=0 $Y2=0
cc_1073 N_A_2136_47#_M1037_g N_VPWR_c_1764_n 0.0147189f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1074 N_A_2136_47#_c_1711_n N_VPWR_c_1764_n 0.0476506f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1075 N_A_2136_47#_c_1706_n N_VPWR_c_1764_n 0.010544f $X=11.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1076 N_A_2136_47#_c_1707_n N_VPWR_c_1764_n 0.00249491f $X=11.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1077 N_A_2136_47#_c_1711_n N_VPWR_c_1774_n 0.0169293f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1078 N_A_2136_47#_M1037_g N_VPWR_c_1775_n 0.0046653f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1079 N_A_2136_47#_M1037_g N_VPWR_c_1759_n 0.00895857f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1080 N_A_2136_47#_c_1711_n N_VPWR_c_1759_n 0.0115924f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1081 N_A_2136_47#_c_1711_n N_Q_N_c_2018_n 0.0871059f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1082 N_A_2136_47#_c_1708_n N_Q_N_c_2018_n 0.0251545f $X=10.817 $Y=1.16 $X2=0
+ $Y2=0
cc_1083 N_A_2136_47#_c_1705_n N_Q_N_c_2020_n 0.0590331f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1084 N_A_2136_47#_M1037_g N_Q_c_2052_n 0.00566837f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1085 N_A_2136_47#_c_1711_n N_Q_c_2052_n 0.0045901f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1086 N_A_2136_47#_M1037_g N_Q_c_2050_n 0.00488612f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1087 N_A_2136_47#_c_1706_n N_Q_c_2050_n 0.0266145f $X=11.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1088 N_A_2136_47#_c_1707_n N_Q_c_2050_n 0.00797367f $X=11.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1089 N_A_2136_47#_c_1709_n N_Q_c_2050_n 0.00640119f $X=11.422 $Y=0.995 $X2=0
+ $Y2=0
cc_1090 N_A_2136_47#_c_1705_n N_VGND_c_2073_n 0.0217483f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1091 N_A_2136_47#_c_1706_n N_VGND_c_2073_n 0.0105205f $X=11.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1092 N_A_2136_47#_c_1707_n N_VGND_c_2073_n 0.00246314f $X=11.41 $Y=1.16 $X2=0
+ $Y2=0
cc_1093 N_A_2136_47#_c_1709_n N_VGND_c_2073_n 0.00941229f $X=11.422 $Y=0.995
+ $X2=0 $Y2=0
cc_1094 N_A_2136_47#_c_1705_n N_VGND_c_2083_n 0.0199778f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1095 N_A_2136_47#_c_1709_n N_VGND_c_2084_n 0.0046653f $X=11.422 $Y=0.995
+ $X2=0 $Y2=0
cc_1096 N_A_2136_47#_M1010_s N_VGND_c_2085_n 0.00210122f $X=10.68 $Y=0.235 $X2=0
+ $Y2=0
cc_1097 N_A_2136_47#_c_1705_n N_VGND_c_2085_n 0.0118987f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1098 N_A_2136_47#_c_1709_n N_VGND_c_2085_n 0.00895857f $X=11.422 $Y=0.995
+ $X2=0 $Y2=0
cc_1099 N_VPWR_c_1759_n N_A_381_47#_M1017_d 0.00287829f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1761_n N_A_381_47#_c_1947_n 0.0127367f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1771_n N_A_381_47#_c_1947_n 0.00221328f $X=3.405 $Y=2.72 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1759_n N_A_381_47#_c_1947_n 0.00204441f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1103 N_VPWR_c_1761_n N_A_381_47#_c_1948_n 0.0116899f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1770_n N_A_381_47#_c_1948_n 3.86777e-19 $X=1.43 $Y=2.72 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1759_n N_A_381_47#_c_1948_n 7.1462e-19 $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1106 N_VPWR_c_1771_n N_A_381_47#_c_1949_n 0.0115924f $X=3.405 $Y=2.72 $X2=0
+ $Y2=0
cc_1107 N_VPWR_c_1759_n N_A_381_47#_c_1949_n 0.00307944f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1108 N_VPWR_c_1759_n A_557_413# 0.00355877f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1109 N_VPWR_c_1759_n A_891_329# 0.0026811f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1110 N_VPWR_c_1759_n A_1112_329# 0.00777501f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1111 N_VPWR_c_1759_n A_1340_413# 0.00305111f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1112 N_VPWR_c_1759_n A_1672_329# 0.00245039f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1113 N_VPWR_c_1759_n N_Q_N_M1039_d 0.00387172f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1764_n Q_N 0.00154465f $X=11.28 $Y=1.94 $X2=0 $Y2=0
cc_1115 N_VPWR_c_1774_n Q_N 0.0197934f $X=11.155 $Y=2.72 $X2=0 $Y2=0
cc_1116 N_VPWR_c_1759_n Q_N 0.0108988f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1117 N_VPWR_c_1759_n N_Q_M1037_d 0.00387172f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1118 N_VPWR_c_1775_n Q 0.018001f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1119 N_VPWR_c_1759_n Q 0.00993603f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1120 N_A_381_47#_c_1944_n N_VGND_M1002_s 0.00125196f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1121 N_A_381_47#_c_1945_n N_VGND_M1002_s 9.40198e-19 $X=1.575 $Y=0.73 $X2=0
+ $Y2=0
cc_1122 N_A_381_47#_c_1944_n N_VGND_c_2068_n 0.0106196f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1123 N_A_381_47#_c_1945_n N_VGND_c_2068_n 0.0115228f $X=1.575 $Y=0.73 $X2=0
+ $Y2=0
cc_1124 N_A_381_47#_c_1944_n N_VGND_c_2074_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1125 N_A_381_47#_c_1978_n N_VGND_c_2074_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1126 N_A_381_47#_c_1945_n N_VGND_c_2081_n 4.97798e-19 $X=1.575 $Y=0.73 $X2=0
+ $Y2=0
cc_1127 N_A_381_47#_M1002_d N_VGND_c_2085_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1128 N_A_381_47#_c_1944_n N_VGND_c_2085_n 0.00239595f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1129 N_A_381_47#_c_1945_n N_VGND_c_2085_n 8.52239e-19 $X=1.575 $Y=0.73 $X2=0
+ $Y2=0
cc_1130 N_A_381_47#_c_1978_n N_VGND_c_2085_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1131 N_Q_N_c_2018_n N_VGND_c_2072_n 0.00203781f $X=10.342 $Y=1.63 $X2=0 $Y2=0
cc_1132 N_Q_N_c_2020_n N_VGND_c_2083_n 0.0196011f $X=10.342 $Y=0.573 $X2=0 $Y2=0
cc_1133 N_Q_N_M1030_d N_VGND_c_2085_n 0.00387172f $X=10.15 $Y=0.235 $X2=0 $Y2=0
cc_1134 N_Q_N_c_2020_n N_VGND_c_2085_n 0.010859f $X=10.342 $Y=0.573 $X2=0 $Y2=0
cc_1135 Q N_VGND_c_2084_n 0.0179623f $X=11.645 $Y=0.425 $X2=0 $Y2=0
cc_1136 N_Q_M1027_d N_VGND_c_2085_n 0.00387172f $X=11.565 $Y=0.235 $X2=0 $Y2=0
cc_1137 Q N_VGND_c_2085_n 0.00992739f $X=11.645 $Y=0.425 $X2=0 $Y2=0
cc_1138 N_VGND_c_2085_n A_581_47# 0.0022723f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1139 N_VGND_c_2085_n N_A_791_47#_M1016_d 0.00214379f $X=11.73 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1140 N_VGND_c_2085_n N_A_791_47#_M1031_d 0.00204204f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1141 N_VGND_c_2070_n N_A_791_47#_c_2257_n 0.0112071f $X=5.51 $Y=0.38 $X2=0
+ $Y2=0
cc_1142 N_VGND_c_2076_n N_A_791_47#_c_2257_n 0.0113927f $X=5.325 $Y=0 $X2=0
+ $Y2=0
cc_1143 N_VGND_c_2085_n N_A_791_47#_c_2257_n 0.00305438f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1144 N_VGND_c_2070_n N_A_791_47#_c_2260_n 0.00235022f $X=5.51 $Y=0.38 $X2=0
+ $Y2=0
cc_1145 N_VGND_c_2076_n N_A_791_47#_c_2267_n 0.0540424f $X=5.325 $Y=0 $X2=0
+ $Y2=0
cc_1146 N_VGND_c_2085_n N_A_791_47#_c_2267_n 0.0159669f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1147 N_VGND_c_2085_n A_1159_47# 0.00617396f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1148 N_VGND_c_2085_n A_1363_47# 0.00261578f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1149 N_VGND_c_2085_n N_A_1555_47#_M1009_d 0.00307401f $X=11.73 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1150 N_VGND_c_2085_n N_A_1555_47#_M1032_d 0.00230679f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1151 N_VGND_c_2082_n N_A_1555_47#_c_2292_n 0.0382042f $X=9.725 $Y=0 $X2=0
+ $Y2=0
cc_1152 N_VGND_c_2085_n N_A_1555_47#_c_2292_n 0.0250101f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1153 N_VGND_c_2082_n N_A_1555_47#_c_2288_n 0.0199008f $X=9.725 $Y=0 $X2=0
+ $Y2=0
cc_1154 N_VGND_c_2085_n N_A_1555_47#_c_2288_n 0.0110702f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1155 N_VGND_c_2082_n N_A_1555_47#_c_2293_n 0.0110309f $X=9.725 $Y=0 $X2=0
+ $Y2=0
cc_1156 N_VGND_c_2085_n N_A_1555_47#_c_2293_n 0.0063548f $X=11.73 $Y=0 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.spice.pex
* Created: Thu Aug 27 14:26:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A 1 3 6 8 12 14
c28 12 0 1.86625e-19 $X=0.45 $Y=1.16
r29 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.45 $Y=1.16
+ $X2=0.66 $Y2=1.16
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.16 $X2=0.45 $Y2=1.16
r31 8 12 5.40943 $w=2.43e-07 $l=1.15e-07 $layer=LI1_cond $X=0.335 $Y=1.197
+ $X2=0.45 $Y2=1.197
r32 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.66 $Y=1.325
+ $X2=0.66 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.66 $Y=1.325 $X2=0.66
+ $Y2=1.985
r34 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.66 $Y=0.995
+ $X2=0.66 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.66 $Y=0.995 $X2=0.66
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_147_47# 1 2 7 9 12 14 16
+ 19 21 23 26 28 30 33 37 41 44 52 55 57 58 59 60 67
c125 60 0 1.86625e-19 $X=1.555 $Y=1.16
c126 58 0 1.68547e-19 $X=0.87 $Y=1.575
c127 26 0 7.39456e-20 $X=2.47 $Y=1.985
c128 14 0 1.6807e-19 $X=2.05 $Y=0.995
r129 66 67 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.47 $Y=1.16
+ $X2=2.89 $Y2=1.16
r130 63 64 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=2.05 $Y2=1.16
r131 60 63 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.555 $Y=1.16
+ $X2=1.63 $Y2=1.16
r132 57 58 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=1.66
+ $X2=0.87 $Y2=1.575
r133 53 66 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.1 $Y=1.16
+ $X2=2.47 $Y2=1.16
r134 53 64 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.1 $Y=1.16 $X2=2.05
+ $Y2=1.16
r135 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.1
+ $Y=1.16 $X2=2.1 $Y2=1.16
r136 50 60 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=1.08 $Y=1.16
+ $X2=1.555 $Y2=1.16
r137 49 52 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=1.08 $Y=1.175
+ $X2=2.1 $Y2=1.175
r138 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r139 47 59 2.15711 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=1.175
+ $X2=0.91 $Y2=1.175
r140 47 49 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=1.035 $Y=1.175
+ $X2=1.08 $Y2=1.175
r141 45 59 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=0.91 $Y=1.275 $X2=0.91
+ $Y2=1.175
r142 45 58 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=0.91 $Y=1.275
+ $X2=0.91 $Y2=1.575
r143 44 59 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=0.91 $Y=1.075 $X2=0.91
+ $Y2=1.175
r144 44 55 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=0.91 $Y=1.075
+ $X2=0.91 $Y2=0.815
r145 39 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.87 $Y=1.74 $X2=0.87
+ $Y2=1.66
r146 39 41 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=0.87 $Y=1.74 $X2=0.87
+ $Y2=2.34
r147 35 55 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=0.65
+ $X2=0.87 $Y2=0.815
r148 35 37 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.87 $Y=0.65
+ $X2=0.87 $Y2=0.39
r149 31 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=1.325
+ $X2=2.89 $Y2=1.16
r150 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.89 $Y=1.325
+ $X2=2.89 $Y2=1.985
r151 28 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=0.995
+ $X2=2.89 $Y2=1.16
r152 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.89 $Y=0.995
+ $X2=2.89 $Y2=0.56
r153 24 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.325
+ $X2=2.47 $Y2=1.16
r154 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.47 $Y=1.325
+ $X2=2.47 $Y2=1.985
r155 21 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=0.995
+ $X2=2.47 $Y2=1.16
r156 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.47 $Y=0.995
+ $X2=2.47 $Y2=0.56
r157 17 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.325
+ $X2=2.05 $Y2=1.16
r158 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.05 $Y=1.325
+ $X2=2.05 $Y2=1.985
r159 14 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=0.995
+ $X2=2.05 $Y2=1.16
r160 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.05 $Y=0.995
+ $X2=2.05 $Y2=0.56
r161 10 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.325
+ $X2=1.63 $Y2=1.16
r162 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.63 $Y=1.325
+ $X2=1.63 $Y2=1.985
r163 7 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=0.995
+ $X2=1.63 $Y2=1.16
r164 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.63 $Y=0.995
+ $X2=1.63 $Y2=0.56
r165 2 57 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=1.485 $X2=0.87 $Y2=1.66
r166 2 41 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=1.485 $X2=0.87 $Y2=2.34
r167 1 37 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.735
+ $Y=0.235 $X2=0.87 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%SLEEP 1 3 6 8 10 13 15 17
+ 20 22 24 27 29 40 41
r94 39 41 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.57 $Y2=1.16
r95 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r96 37 39 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=4.15 $Y=1.16 $X2=4.46
+ $Y2=1.16
r97 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.73 $Y=1.16
+ $X2=4.15 $Y2=1.16
r98 34 36 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.44 $Y=1.16
+ $X2=3.73 $Y2=1.16
r99 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r100 31 34 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=3.31 $Y=1.16
+ $X2=3.44 $Y2=1.16
r101 29 40 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=4.365 $Y=1.175
+ $X2=4.46 $Y2=1.175
r102 29 35 51.2955 $w=1.98e-07 $l=9.25e-07 $layer=LI1_cond $X=4.365 $Y=1.175
+ $X2=3.44 $Y2=1.175
r103 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.325
+ $X2=4.57 $Y2=1.16
r104 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.57 $Y=1.325
+ $X2=4.57 $Y2=1.985
r105 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=0.995
+ $X2=4.57 $Y2=1.16
r106 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.57 $Y=0.995
+ $X2=4.57 $Y2=0.56
r107 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.15 $Y=1.325
+ $X2=4.15 $Y2=1.16
r108 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.15 $Y=1.325
+ $X2=4.15 $Y2=1.985
r109 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.15 $Y=0.995
+ $X2=4.15 $Y2=1.16
r110 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.15 $Y=0.995
+ $X2=4.15 $Y2=0.56
r111 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.325
+ $X2=3.73 $Y2=1.16
r112 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.73 $Y=1.325
+ $X2=3.73 $Y2=1.985
r113 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=0.995
+ $X2=3.73 $Y2=1.16
r114 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.73 $Y=0.995
+ $X2=3.73 $Y2=0.56
r115 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.325
+ $X2=3.31 $Y2=1.16
r116 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.31 $Y=1.325
+ $X2=3.31 $Y2=1.985
r117 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.16
r118 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_341_47# 1 2 3 4 5 6 21 23
+ 25 28 30 32 35 37 39 42 44 46 49 51 53 55 58 60 63 67 69 73 75 79 84 85 86 91
+ 92 94 95 104 111 114
c220 104 0 1.60903e-20 $X=6.825 $Y=1.155
c221 95 0 1.41095e-19 $X=5.295 $Y=0.85
c222 60 0 1.6807e-19 $X=2.6 $Y=1.445
c223 55 0 1.22434e-19 $X=2.435 $Y=1.595
r224 103 104 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=6.395 $Y=1.155
+ $X2=6.825 $Y2=1.155
r225 102 103 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=5.965 $Y=1.155
+ $X2=6.395 $Y2=1.155
r226 101 102 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=5.535 $Y=1.155
+ $X2=5.965 $Y2=1.155
r227 98 101 21.5061 $w=5.1e-07 $l=2.05e-07 $layer=POLY_cond $X=5.33 $Y=1.155
+ $X2=5.535 $Y2=1.155
r228 98 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.16 $X2=5.33 $Y2=1.16
r229 95 99 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=5.302 $Y=0.85
+ $X2=5.302 $Y2=1.16
r230 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.295 $Y=0.85
+ $X2=5.295 $Y2=0.85
r231 91 94 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.15 $Y=0.85
+ $X2=5.295 $Y2=0.85
r232 91 92 2.51856 $w=1.4e-07 $l=2.035e-06 $layer=MET1_cond $X=5.15 $Y=0.85
+ $X2=3.115 $Y2=0.85
r233 89 114 6.74844 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.97 $Y=0.845
+ $X2=3.095 $Y2=0.845
r234 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.97 $Y=0.85
+ $X2=2.97 $Y2=0.85
r235 86 92 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=3 $Y=0.85
+ $X2=3.115 $Y2=0.85
r236 86 88 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=3 $Y=0.85 $X2=2.97
+ $Y2=0.85
r237 77 79 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.36 $Y=0.725
+ $X2=4.36 $Y2=0.39
r238 76 85 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0.815
+ $X2=3.52 $Y2=0.815
r239 75 77 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.195 $Y=0.815
+ $X2=4.36 $Y2=0.725
r240 75 76 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.195 $Y=0.815
+ $X2=3.685 $Y2=0.815
r241 71 85 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.52 $Y=0.725
+ $X2=3.52 $Y2=0.815
r242 71 73 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.52 $Y=0.725
+ $X2=3.52 $Y2=0.39
r243 69 85 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.52 $Y2=0.815
r244 69 114 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.095 $Y2=0.815
r245 65 84 5.99569 $w=2.5e-07 $l=1.85742e-07 $layer=LI1_cond $X=2.68 $Y=1.745
+ $X2=2.6 $Y2=1.595
r246 65 67 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.68 $Y=1.745
+ $X2=2.68 $Y2=1.96
r247 61 89 13.9254 $w=2.38e-07 $l=2.9e-07 $layer=LI1_cond $X=2.68 $Y=0.845
+ $X2=2.97 $Y2=0.845
r248 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.68 $Y=0.725
+ $X2=2.68 $Y2=0.39
r249 60 84 5.99569 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=2.6 $Y=1.445 $X2=2.6
+ $Y2=1.595
r250 59 61 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=2.6 $Y=0.845 $X2=2.68
+ $Y2=0.845
r251 59 111 8.66918 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=0.845
+ $X2=2.435 $Y2=0.845
r252 59 60 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.6 $Y=0.965
+ $X2=2.6 $Y2=1.445
r253 58 111 26.4949 $w=1.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.005 $Y=0.815
+ $X2=2.435 $Y2=0.815
r254 56 82 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.925 $Y=1.595
+ $X2=1.84 $Y2=1.595
r255 55 84 0.695019 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=1.595
+ $X2=2.6 $Y2=1.595
r256 55 56 19.5915 $w=2.98e-07 $l=5.1e-07 $layer=LI1_cond $X=2.435 $Y=1.595
+ $X2=1.925 $Y2=1.595
r257 51 82 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.84 $Y=1.745
+ $X2=1.84 $Y2=1.595
r258 51 53 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.84 $Y=1.745
+ $X2=1.84 $Y2=1.96
r259 47 58 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.84 $Y=0.725
+ $X2=2.005 $Y2=0.815
r260 47 49 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.84 $Y=0.725
+ $X2=1.84 $Y2=0.39
r261 44 104 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.825 $Y=1.41
+ $X2=6.825 $Y2=1.155
r262 44 46 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.825 $Y=1.41
+ $X2=6.825 $Y2=1.985
r263 40 104 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.825 $Y=0.9
+ $X2=6.825 $Y2=1.155
r264 40 42 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.825 $Y=0.9
+ $X2=6.825 $Y2=0.445
r265 37 103 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.395 $Y=1.41
+ $X2=6.395 $Y2=1.155
r266 37 39 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.395 $Y=1.41
+ $X2=6.395 $Y2=1.985
r267 33 103 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.395 $Y=0.9
+ $X2=6.395 $Y2=1.155
r268 33 35 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.395 $Y=0.9
+ $X2=6.395 $Y2=0.445
r269 30 102 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.965 $Y=1.41
+ $X2=5.965 $Y2=1.155
r270 30 32 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.965 $Y=1.41
+ $X2=5.965 $Y2=1.985
r271 26 102 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.965 $Y=0.9
+ $X2=5.965 $Y2=1.155
r272 26 28 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.965 $Y=0.9
+ $X2=5.965 $Y2=0.445
r273 23 101 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.535 $Y=1.41
+ $X2=5.535 $Y2=1.155
r274 23 25 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.535 $Y=1.41
+ $X2=5.535 $Y2=1.985
r275 19 101 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.535 $Y=0.9
+ $X2=5.535 $Y2=1.155
r276 19 21 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.535 $Y=0.9
+ $X2=5.535 $Y2=0.445
r277 6 84 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=1.485 $X2=2.68 $Y2=1.62
r278 6 67 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=1.485 $X2=2.68 $Y2=1.96
r279 5 82 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=1.485 $X2=1.84 $Y2=1.62
r280 5 53 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=1.485 $X2=1.84 $Y2=1.96
r281 4 79 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.225
+ $Y=0.235 $X2=4.36 $Y2=0.39
r282 3 73 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.52 $Y2=0.39
r283 2 63 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.545
+ $Y=0.235 $X2=2.68 $Y2=0.39
r284 1 49 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.705
+ $Y=0.235 $X2=1.84 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_1122_47# 1 2 3 4 15 19 23
+ 27 31 35 39 43 47 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119
+ 123 127 131 133 135 139 143 147 151 155 159 168 171 172
r336 168 169 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=12.565
+ $Y=1.16 $X2=12.565 $Y2=1.16
r337 165 168 235.098 $w=2.48e-07 $l=5.1e-06 $layer=LI1_cond $X=7.465 $Y=1.2
+ $X2=12.565 $Y2=1.2
r338 165 166 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=7.465
+ $Y=1.16 $X2=7.465 $Y2=1.16
r339 163 172 2.66945 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.74 $Y=1.2
+ $X2=6.615 $Y2=1.2
r340 163 165 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=6.74 $Y=1.2
+ $X2=7.465 $Y2=1.2
r341 159 161 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=6.61 $Y=1.615
+ $X2=6.61 $Y2=2.295
r342 157 172 3.44865 $w=1.9e-07 $l=1.27475e-07 $layer=LI1_cond $X=6.61 $Y=1.325
+ $X2=6.615 $Y2=1.2
r343 157 159 16.9282 $w=1.88e-07 $l=2.9e-07 $layer=LI1_cond $X=6.61 $Y=1.325
+ $X2=6.61 $Y2=1.615
r344 153 172 3.44865 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.615 $Y=1.075
+ $X2=6.615 $Y2=1.2
r345 153 155 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=6.615 $Y=1.075
+ $X2=6.615 $Y2=0.445
r346 152 171 0.681005 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=5.88 $Y=1.2
+ $X2=5.767 $Y2=1.2
r347 151 172 2.66945 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.49 $Y=1.2
+ $X2=6.615 $Y2=1.2
r348 151 152 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=6.49 $Y=1.2
+ $X2=5.88 $Y2=1.2
r349 147 149 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=5.75 $Y=1.62
+ $X2=5.75 $Y2=2.3
r350 145 171 6.01496 $w=2.07e-07 $l=1.33229e-07 $layer=LI1_cond $X=5.75 $Y=1.325
+ $X2=5.767 $Y2=1.2
r351 145 147 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=5.75 $Y=1.325
+ $X2=5.75 $Y2=1.62
r352 141 171 6.01496 $w=2.07e-07 $l=1.25e-07 $layer=LI1_cond $X=5.767 $Y=1.075
+ $X2=5.767 $Y2=1.2
r353 141 143 32.2684 $w=2.23e-07 $l=6.3e-07 $layer=LI1_cond $X=5.767 $Y=1.075
+ $X2=5.767 $Y2=0.445
r354 137 139 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.7 $Y=1.325
+ $X2=13.7 $Y2=1.985
r355 133 137 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=13.7 $Y=1.137
+ $X2=13.7 $Y2=1.325
r356 133 135 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=13.7 $Y=0.95
+ $X2=13.7 $Y2=0.445
r357 129 131 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.27 $Y=1.325
+ $X2=13.27 $Y2=1.985
r358 125 133 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=13.27 $Y=1.137
+ $X2=13.7 $Y2=1.137
r359 125 129 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=13.27 $Y=1.137
+ $X2=13.27 $Y2=1.325
r360 125 127 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=13.27 $Y=0.95
+ $X2=13.27 $Y2=0.445
r361 121 123 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.84 $Y=1.325
+ $X2=12.84 $Y2=1.985
r362 117 125 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=12.84 $Y=1.137
+ $X2=13.27 $Y2=1.137
r363 117 121 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=12.84 $Y=1.137
+ $X2=12.84 $Y2=1.325
r364 117 169 40.7846 $w=3.75e-07 $l=2.75e-07 $layer=POLY_cond $X=12.84 $Y=1.137
+ $X2=12.565 $Y2=1.137
r365 117 119 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=12.84 $Y=0.95
+ $X2=12.84 $Y2=0.445
r366 113 115 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.41 $Y=1.325
+ $X2=12.41 $Y2=1.985
r367 109 169 22.9877 $w=3.75e-07 $l=1.55e-07 $layer=POLY_cond $X=12.41 $Y=1.137
+ $X2=12.565 $Y2=1.137
r368 109 113 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=12.41 $Y=1.137
+ $X2=12.41 $Y2=1.325
r369 109 111 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=12.41 $Y=0.95
+ $X2=12.41 $Y2=0.445
r370 105 107 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.98 $Y=1.325
+ $X2=11.98 $Y2=1.985
r371 101 109 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=11.98 $Y=1.137
+ $X2=12.41 $Y2=1.137
r372 101 105 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=11.98 $Y=1.137
+ $X2=11.98 $Y2=1.325
r373 101 103 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.98 $Y=0.95
+ $X2=11.98 $Y2=0.445
r374 97 99 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.55 $Y=1.325
+ $X2=11.55 $Y2=1.985
r375 93 101 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=11.55 $Y=1.137
+ $X2=11.98 $Y2=1.137
r376 93 97 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=11.55 $Y=1.137
+ $X2=11.55 $Y2=1.325
r377 93 95 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.55 $Y=0.95
+ $X2=11.55 $Y2=0.445
r378 89 91 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.12 $Y=1.325
+ $X2=11.12 $Y2=1.985
r379 85 93 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=11.12 $Y=1.137
+ $X2=11.55 $Y2=1.137
r380 85 89 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=11.12 $Y=1.137
+ $X2=11.12 $Y2=1.325
r381 85 87 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.12 $Y=0.95
+ $X2=11.12 $Y2=0.445
r382 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.69 $Y=1.325
+ $X2=10.69 $Y2=1.985
r383 77 85 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=10.69 $Y=1.137
+ $X2=11.12 $Y2=1.137
r384 77 81 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=10.69 $Y=1.137
+ $X2=10.69 $Y2=1.325
r385 77 79 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=10.69 $Y=0.95
+ $X2=10.69 $Y2=0.445
r386 73 75 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.265 $Y=1.325
+ $X2=10.265 $Y2=1.985
r387 69 77 63.0308 $w=3.75e-07 $l=4.25e-07 $layer=POLY_cond $X=10.265 $Y=1.137
+ $X2=10.69 $Y2=1.137
r388 69 73 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=10.265 $Y=1.137
+ $X2=10.265 $Y2=1.325
r389 69 71 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=10.265 $Y=0.95
+ $X2=10.265 $Y2=0.445
r390 65 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.835 $Y=1.325
+ $X2=9.835 $Y2=1.985
r391 61 69 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=9.835 $Y=1.137
+ $X2=10.265 $Y2=1.137
r392 61 65 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=9.835 $Y=1.137
+ $X2=9.835 $Y2=1.325
r393 61 63 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.835 $Y=0.95
+ $X2=9.835 $Y2=0.445
r394 57 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.405 $Y=1.325
+ $X2=9.405 $Y2=1.985
r395 53 61 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=9.405 $Y=1.137
+ $X2=9.835 $Y2=1.137
r396 53 57 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=9.405 $Y=1.137
+ $X2=9.405 $Y2=1.325
r397 53 55 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.405 $Y=0.95
+ $X2=9.405 $Y2=0.445
r398 49 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.975 $Y=1.325
+ $X2=8.975 $Y2=1.985
r399 45 53 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=8.975 $Y=1.137
+ $X2=9.405 $Y2=1.137
r400 45 49 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.975 $Y=1.137
+ $X2=8.975 $Y2=1.325
r401 45 47 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.975 $Y=0.95
+ $X2=8.975 $Y2=0.445
r402 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.545 $Y=1.325
+ $X2=8.545 $Y2=1.985
r403 37 45 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=8.545 $Y=1.137
+ $X2=8.975 $Y2=1.137
r404 37 41 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.545 $Y=1.137
+ $X2=8.545 $Y2=1.325
r405 37 39 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.545 $Y=0.95
+ $X2=8.545 $Y2=0.445
r406 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.115 $Y=1.325
+ $X2=8.115 $Y2=1.985
r407 29 37 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=8.115 $Y=1.137
+ $X2=8.545 $Y2=1.137
r408 29 33 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.115 $Y=1.137
+ $X2=8.115 $Y2=1.325
r409 29 31 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.115 $Y=0.95
+ $X2=8.115 $Y2=0.445
r410 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.685 $Y=1.325
+ $X2=7.685 $Y2=1.985
r411 21 29 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=7.685 $Y=1.137
+ $X2=8.115 $Y2=1.137
r412 21 25 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=7.685 $Y=1.137
+ $X2=7.685 $Y2=1.325
r413 21 166 32.6277 $w=3.75e-07 $l=2.2e-07 $layer=POLY_cond $X=7.685 $Y=1.137
+ $X2=7.465 $Y2=1.137
r414 21 23 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.685 $Y=0.95
+ $X2=7.685 $Y2=0.445
r415 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.255 $Y=1.325
+ $X2=7.255 $Y2=1.985
r416 13 166 31.1446 $w=3.75e-07 $l=2.1e-07 $layer=POLY_cond $X=7.255 $Y=1.137
+ $X2=7.465 $Y2=1.137
r417 13 17 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=7.255 $Y=1.137
+ $X2=7.255 $Y2=1.325
r418 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.255 $Y=0.95
+ $X2=7.255 $Y2=0.445
r419 4 161 400 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=6.47
+ $Y=1.485 $X2=6.61 $Y2=2.295
r420 4 159 400 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_PDIFF $count=1 $X=6.47
+ $Y=1.485 $X2=6.61 $Y2=1.615
r421 3 149 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=5.61
+ $Y=1.485 $X2=5.75 $Y2=2.3
r422 3 147 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=5.61
+ $Y=1.485 $X2=5.75 $Y2=1.62
r423 2 155 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.47
+ $Y=0.235 $X2=6.61 $Y2=0.445
r424 1 143 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.235 $X2=5.75 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%VPWR 1 2 3 10 12 18 22 24
+ 26 31 41 42 48 51
c198 41 0 1.77237e-19 $X=14.03 $Y=2.72
r199 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r200 48 49 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r201 41 42 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=14.03
+ $Y=2.72 $X2=14.03 $Y2=2.72
r202 39 42 2.61778 $w=4.8e-07 $l=9.2e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=14.03 $Y2=2.72
r203 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r204 38 41 600.214 $w=1.68e-07 $l=9.2e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=14.03 $Y2=2.72
r205 38 39 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=4.83
+ $Y=2.72 $X2=4.83 $Y2=2.72
r206 36 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=2.72
+ $X2=4.36 $Y2=2.72
r207 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.525 $Y=2.72
+ $X2=4.83 $Y2=2.72
r208 35 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r209 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r210 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r211 32 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.56 $Y2=2.72
r212 32 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.91 $Y2=2.72
r213 31 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=4.36 $Y2=2.72
r214 31 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=3.91 $Y2=2.72
r215 30 49 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=3.45 $Y2=2.72
r216 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r217 27 45 5.39493 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.267 $Y2=2.72
r218 27 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.69 $Y2=2.72
r219 26 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.435 $Y=2.72
+ $X2=3.56 $Y2=2.72
r220 26 29 179.086 $w=1.68e-07 $l=2.745e-06 $layer=LI1_cond $X=3.435 $Y=2.72
+ $X2=0.69 $Y2=2.72
r221 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r222 24 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r223 20 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=2.635
+ $X2=4.36 $Y2=2.72
r224 20 22 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.36 $Y=2.635
+ $X2=4.36 $Y2=2
r225 16 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=2.635
+ $X2=3.56 $Y2=2.72
r226 16 18 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.56 $Y=2.635
+ $X2=3.56 $Y2=2
r227 12 15 19.3497 $w=4.03e-07 $l=6.8e-07 $layer=LI1_cond $X=0.332 $Y=1.66
+ $X2=0.332 $Y2=2.34
r228 10 45 3.01955 $w=4.05e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.332 $Y=2.635
+ $X2=0.267 $Y2=2.72
r229 10 15 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.332 $Y=2.635
+ $X2=0.332 $Y2=2.34
r230 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=1.485 $X2=4.36 $Y2=2
r231 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.385
+ $Y=1.485 $X2=3.52 $Y2=2
r232 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.485 $X2=0.45 $Y2=2.34
r233 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.485 $X2=0.45 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_255_297# 1 2 3 4 5 16 18
+ 20 24 26 28 29 30 34 36 38 40 44 50
c102 28 0 7.39456e-20 $X=3.1 $Y=1.665
c103 26 0 1.22434e-19 $X=2.935 $Y=2.38
r104 38 52 2.99957 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=4.835 $Y=1.665
+ $X2=4.835 $Y2=1.56
r105 38 40 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.835 $Y=1.665
+ $X2=4.835 $Y2=2.3
r106 37 50 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=1.56
+ $X2=3.94 $Y2=1.56
r107 36 52 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=4.695 $Y=1.56
+ $X2=4.835 $Y2=1.56
r108 36 37 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=4.695 $Y=1.56
+ $X2=4.025 $Y2=1.56
r109 32 50 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.94 $Y=1.665
+ $X2=3.94 $Y2=1.56
r110 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.94 $Y=1.665
+ $X2=3.94 $Y2=2.3
r111 31 46 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=1.56
+ $X2=3.1 $Y2=1.56
r112 30 50 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=1.56
+ $X2=3.94 $Y2=1.56
r113 30 31 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=3.855 $Y=1.56
+ $X2=3.265 $Y2=1.56
r114 29 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=2.295 $X2=3.1
+ $Y2=2.38
r115 28 46 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=3.1 $Y=1.665
+ $X2=3.1 $Y2=1.56
r116 28 29 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=3.1 $Y=1.665
+ $X2=3.1 $Y2=2.295
r117 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.38
+ $X2=2.26 $Y2=2.38
r118 26 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=2.38
+ $X2=3.1 $Y2=2.38
r119 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.935 $Y=2.38
+ $X2=2.425 $Y2=2.38
r120 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=2.295
+ $X2=2.26 $Y2=2.38
r121 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.26 $Y=2.295
+ $X2=2.26 $Y2=2.02
r122 21 43 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.585 $Y=2.38
+ $X2=1.395 $Y2=2.38
r123 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=2.38
+ $X2=2.26 $Y2=2.38
r124 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.095 $Y=2.38
+ $X2=1.585 $Y2=2.38
r125 16 43 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=2.295
+ $X2=1.395 $Y2=2.38
r126 16 18 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.395 $Y=2.295
+ $X2=1.395 $Y2=1.66
r127 5 52 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.485 $X2=4.78 $Y2=1.62
r128 5 40 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.485 $X2=4.78 $Y2=2.3
r129 4 50 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.485 $X2=3.94 $Y2=1.62
r130 4 34 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.485 $X2=3.94 $Y2=2.3
r131 3 48 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.485 $X2=3.1 $Y2=2.34
r132 3 46 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.485 $X2=3.1 $Y2=1.62
r133 2 24 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.125
+ $Y=1.485 $X2=2.26 $Y2=2.02
r134 1 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.485 $X2=1.42 $Y2=2.34
r135 1 18 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.485 $X2=1.42 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%KAPWR 1 2 3 4 5 6 7 8 9 10
+ 11 52 58 59 63 64 68 69 72 73 74 77 78 79 82 83 84 87 88 89 92 93 94 97 98 99
+ 102 103 104 107 108 111 117 123 161
c239 74 0 1.77237e-19 $X=8.03 $Y=2.21
c240 52 0 1.27506e-19 $X=13.78 $Y=2.24
c241 11 0 4.2343e-20 $X=13.775 $Y=1.485
r242 108 161 0.00921054 $w=2e-07 $l=1.2e-08 $layer=MET1_cond $X=0.252 $Y=2.24
+ $X2=0.24 $Y2=2.24
r243 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.925 $Y=2.21
+ $X2=13.925 $Y2=2.21
r244 101 104 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=13.045 $Y=2.21
+ $X2=13.19 $Y2=2.21
r245 101 103 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=13.045 $Y=2.21
+ $X2=12.9 $Y2=2.21
r246 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.045 $Y=2.21
+ $X2=13.045 $Y2=2.21
r247 99 103 0.429825 $w=2e-07 $l=5.6e-07 $layer=MET1_cond $X=12.34 $Y=2.24
+ $X2=12.9 $Y2=2.24
r248 96 99 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=12.195 $Y=2.21
+ $X2=12.34 $Y2=2.21
r249 96 98 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=12.195 $Y=2.21
+ $X2=12.05 $Y2=2.21
r250 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.195 $Y=2.21
+ $X2=12.195 $Y2=2.21
r251 94 98 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=11.485 $Y=2.24
+ $X2=12.05 $Y2=2.24
r252 91 94 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=11.34 $Y=2.21
+ $X2=11.485 $Y2=2.21
r253 91 93 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=11.34 $Y=2.21
+ $X2=11.195 $Y2=2.21
r254 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.34 $Y=2.21
+ $X2=11.34 $Y2=2.21
r255 89 93 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=10.625 $Y=2.24
+ $X2=11.195 $Y2=2.24
r256 86 89 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=10.48 $Y=2.21
+ $X2=10.625 $Y2=2.21
r257 86 88 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=10.48 $Y=2.21
+ $X2=10.335 $Y2=2.21
r258 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.48 $Y=2.21
+ $X2=10.48 $Y2=2.21
r259 84 88 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=9.77 $Y=2.24
+ $X2=10.335 $Y2=2.24
r260 81 84 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=9.625 $Y=2.21
+ $X2=9.77 $Y2=2.21
r261 81 83 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=9.625 $Y=2.21
+ $X2=9.48 $Y2=2.21
r262 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.625 $Y=2.21
+ $X2=9.625 $Y2=2.21
r263 79 83 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=8.91 $Y=2.24
+ $X2=9.48 $Y2=2.24
r264 76 79 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=8.765 $Y=2.21
+ $X2=8.91 $Y2=2.21
r265 76 78 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=8.765 $Y=2.21
+ $X2=8.62 $Y2=2.21
r266 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.765 $Y=2.21
+ $X2=8.765 $Y2=2.21
r267 74 78 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=8.03 $Y=2.24
+ $X2=8.62 $Y2=2.24
r268 71 74 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.885 $Y=2.21
+ $X2=8.03 $Y2=2.21
r269 71 73 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.885 $Y=2.21
+ $X2=7.74 $Y2=2.21
r270 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.885 $Y=2.21
+ $X2=7.885 $Y2=2.21
r271 69 73 0.429825 $w=2e-07 $l=5.6e-07 $layer=MET1_cond $X=7.18 $Y=2.24
+ $X2=7.74 $Y2=2.24
r272 67 123 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=7.04 $Y=2.21
+ $X2=7.04 $Y2=1.66
r273 66 69 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.035 $Y=2.21
+ $X2=7.18 $Y2=2.21
r274 66 68 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.035 $Y=2.21
+ $X2=6.89 $Y2=2.21
r275 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.035 $Y=2.21
+ $X2=7.035 $Y2=2.21
r276 64 68 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=6.325 $Y=2.24
+ $X2=6.89 $Y2=2.24
r277 62 117 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=6.18 $Y=2.21
+ $X2=6.18 $Y2=1.66
r278 61 64 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=6.18 $Y=2.21
+ $X2=6.325 $Y2=2.21
r279 61 63 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=6.18 $Y=2.21
+ $X2=6.035 $Y2=2.21
r280 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=2.21
+ $X2=6.18 $Y2=2.21
r281 59 63 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=5.465 $Y=2.24
+ $X2=6.035 $Y2=2.24
r282 58 108 3.77862 $w=2e-07 $l=4.923e-06 $layer=MET1_cond $X=5.175 $Y=2.24
+ $X2=0.252 $Y2=2.24
r283 57 111 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=5.32 $Y=2.21
+ $X2=5.32 $Y2=1.66
r284 56 59 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.32 $Y=2.21
+ $X2=5.465 $Y2=2.21
r285 56 58 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.32 $Y=2.21
+ $X2=5.175 $Y2=2.21
r286 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.32 $Y=2.21
+ $X2=5.32 $Y2=2.21
r287 52 106 0.0790316 $w=2.42e-07 $l=1.59295e-07 $layer=MET1_cond $X=13.78
+ $Y=2.24 $X2=13.925 $Y2=2.21
r288 52 104 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=13.78 $Y=2.24
+ $X2=13.19 $Y2=2.24
r289 11 107 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=13.775
+ $Y=1.485 $X2=13.915 $Y2=2.22
r290 10 102 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=12.915
+ $Y=1.485 $X2=13.055 $Y2=2.22
r291 9 97 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=12.055
+ $Y=1.485 $X2=12.195 $Y2=2.22
r292 8 92 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=11.195
+ $Y=1.485 $X2=11.335 $Y2=2.22
r293 7 87 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=10.34
+ $Y=1.485 $X2=10.48 $Y2=2.22
r294 6 82 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.62 $Y2=2.22
r295 5 77 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=8.62
+ $Y=1.485 $X2=8.76 $Y2=2.22
r296 4 72 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.485 $X2=7.9 $Y2=2.22
r297 3 67 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=1.485 $X2=7.04 $Y2=2.34
r298 3 123 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=1.485 $X2=7.04 $Y2=1.66
r299 2 62 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=1.485 $X2=6.18 $Y2=2.34
r300 2 117 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=1.485 $X2=6.18 $Y2=1.66
r301 1 57 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.485 $X2=5.32 $Y2=2.34
r302 1 111 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.485 $X2=5.32 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%X 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 51 55 56 57 61 65 67 71 75 77 81 85 87 91 95 97 101 105 107 111
+ 115 119 124 125 127 128 130 131 133 134 136 137 139 140 141 142 143 168 173
c300 141 0 1.18325e-19 $X=13.57 $Y=0.85
c301 16 0 1.27506e-19 $X=13.345 $Y=1.485
r302 171 173 0.603562 $w=1.516e-06 $l=7.5e-08 $layer=LI1_cond $X=13.285 $Y=1.615
+ $X2=13.285 $Y2=1.69
r303 158 168 0.966712 $w=1.516e-06 $l=2.33846e-07 $layer=LI1_cond $X=13.502
+ $Y=1.495 $X2=13.285 $Y2=1.53
r304 143 171 0.48285 $w=1.516e-06 $l=6e-08 $layer=LI1_cond $X=13.285 $Y=1.555
+ $X2=13.285 $Y2=1.615
r305 143 168 0.201187 $w=1.516e-06 $l=2.5e-08 $layer=LI1_cond $X=13.285 $Y=1.555
+ $X2=13.285 $Y2=1.53
r306 143 158 0.261803 $w=1.163e-06 $l=2.5e-08 $layer=LI1_cond $X=13.502 $Y=1.47
+ $X2=13.502 $Y2=1.495
r307 142 143 2.93219 $w=1.163e-06 $l=2.8e-07 $layer=LI1_cond $X=13.502 $Y=1.19
+ $X2=13.502 $Y2=1.47
r308 141 157 1.4003 $w=7.12e-07 $l=8.5e-08 $layer=LI1_cond $X=13.502 $Y=0.82
+ $X2=13.502 $Y2=0.905
r309 141 142 2.82747 $w=1.163e-06 $l=2.7e-07 $layer=LI1_cond $X=13.502 $Y=0.92
+ $X2=13.502 $Y2=1.19
r310 141 157 0.157082 $w=1.163e-06 $l=1.5e-08 $layer=LI1_cond $X=13.502 $Y=0.92
+ $X2=13.502 $Y2=0.905
r311 117 141 1.4003 $w=7.12e-07 $l=9.31128e-08 $layer=LI1_cond $X=13.485
+ $Y=0.735 $X2=13.502 $Y2=0.82
r312 117 119 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=13.485 $Y=0.735
+ $X2=13.485 $Y2=0.445
r313 116 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.745 $Y=0.82
+ $X2=12.615 $Y2=0.82
r314 115 141 6.76561 $w=1.7e-07 $l=5.82e-07 $layer=LI1_cond $X=12.92 $Y=0.82
+ $X2=13.502 $Y2=0.82
r315 115 116 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=12.92 $Y=0.82
+ $X2=12.745 $Y2=0.82
r316 109 140 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.615 $Y=0.735
+ $X2=12.615 $Y2=0.82
r317 109 111 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=12.615 $Y=0.735
+ $X2=12.615 $Y2=0.445
r318 108 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=11.885 $Y=1.615
+ $X2=11.755 $Y2=1.615
r319 107 171 12.2163 $w=2.4e-07 $l=8e-07 $layer=LI1_cond $X=12.485 $Y=1.615
+ $X2=13.285 $Y2=1.615
r320 107 108 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=12.485 $Y=1.615
+ $X2=11.885 $Y2=1.615
r321 106 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.885 $Y=0.82
+ $X2=11.755 $Y2=0.82
r322 105 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.485 $Y=0.82
+ $X2=12.615 $Y2=0.82
r323 105 106 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=12.485 $Y=0.82
+ $X2=11.885 $Y2=0.82
r324 99 137 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.755 $Y=0.735
+ $X2=11.755 $Y2=0.82
r325 99 101 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=11.755 $Y=0.735
+ $X2=11.755 $Y2=0.445
r326 98 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=11.025 $Y=1.615
+ $X2=10.895 $Y2=1.615
r327 97 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=11.625 $Y=1.615
+ $X2=11.755 $Y2=1.615
r328 97 98 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=11.625 $Y=1.615
+ $X2=11.025 $Y2=1.615
r329 96 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.025 $Y=0.82
+ $X2=10.895 $Y2=0.82
r330 95 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.625 $Y=0.82
+ $X2=11.755 $Y2=0.82
r331 95 96 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=11.625 $Y=0.82
+ $X2=11.025 $Y2=0.82
r332 89 134 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.895 $Y=0.735
+ $X2=10.895 $Y2=0.82
r333 89 91 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=10.895 $Y=0.735
+ $X2=10.895 $Y2=0.445
r334 88 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=10.18 $Y=1.615
+ $X2=10.05 $Y2=1.615
r335 87 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=10.765 $Y=1.615
+ $X2=10.895 $Y2=1.615
r336 87 88 28.0908 $w=2.38e-07 $l=5.85e-07 $layer=LI1_cond $X=10.765 $Y=1.615
+ $X2=10.18 $Y2=1.615
r337 86 131 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.18 $Y=0.82
+ $X2=10.042 $Y2=0.82
r338 85 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.765 $Y=0.82
+ $X2=10.895 $Y2=0.82
r339 85 86 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=10.765 $Y=0.82
+ $X2=10.18 $Y2=0.82
r340 79 131 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.042 $Y=0.735
+ $X2=10.042 $Y2=0.82
r341 79 81 12.153 $w=2.73e-07 $l=2.9e-07 $layer=LI1_cond $X=10.042 $Y=0.735
+ $X2=10.042 $Y2=0.445
r342 78 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=9.32 $Y=1.615
+ $X2=9.19 $Y2=1.615
r343 77 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=9.92 $Y=1.615
+ $X2=10.05 $Y2=1.615
r344 77 78 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=9.92 $Y=1.615
+ $X2=9.32 $Y2=1.615
r345 76 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.32 $Y=0.82
+ $X2=9.19 $Y2=0.82
r346 75 131 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=9.905 $Y=0.82
+ $X2=10.042 $Y2=0.82
r347 75 76 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.905 $Y=0.82
+ $X2=9.32 $Y2=0.82
r348 69 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.19 $Y=0.735
+ $X2=9.19 $Y2=0.82
r349 69 71 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=9.19 $Y=0.735
+ $X2=9.19 $Y2=0.445
r350 68 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=8.46 $Y=1.615
+ $X2=8.33 $Y2=1.615
r351 67 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=9.06 $Y=1.615
+ $X2=9.19 $Y2=1.615
r352 67 68 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=9.06 $Y=1.615
+ $X2=8.46 $Y2=1.615
r353 66 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.46 $Y=0.82
+ $X2=8.33 $Y2=0.82
r354 65 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.06 $Y=0.82
+ $X2=9.19 $Y2=0.82
r355 65 66 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=9.06 $Y=0.82 $X2=8.46
+ $Y2=0.82
r356 59 125 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=0.735
+ $X2=8.33 $Y2=0.82
r357 59 61 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=8.33 $Y=0.735
+ $X2=8.33 $Y2=0.445
r358 58 124 3.31033 $w=2.4e-07 $l=1.13e-07 $layer=LI1_cond $X=7.6 $Y=1.615
+ $X2=7.487 $Y2=1.615
r359 57 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=8.2 $Y=1.615
+ $X2=8.33 $Y2=1.615
r360 57 58 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=8.2 $Y=1.615 $X2=7.6
+ $Y2=1.615
r361 55 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.2 $Y=0.82
+ $X2=8.33 $Y2=0.82
r362 55 56 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.2 $Y=0.82 $X2=7.6
+ $Y2=0.82
r363 49 56 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.47 $Y=0.735
+ $X2=7.6 $Y2=0.82
r364 49 51 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=7.47 $Y=0.735
+ $X2=7.47 $Y2=0.445
r365 16 173 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=13.345
+ $Y=1.485 $X2=13.485 $Y2=1.69
r366 15 173 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=12.485
+ $Y=1.485 $X2=12.625 $Y2=1.69
r367 14 139 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=11.625
+ $Y=1.485 $X2=11.765 $Y2=1.69
r368 13 136 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=10.765
+ $Y=1.485 $X2=10.905 $Y2=1.69
r369 12 133 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=9.91
+ $Y=1.485 $X2=10.05 $Y2=1.69
r370 11 130 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=9.05
+ $Y=1.485 $X2=9.19 $Y2=1.69
r371 10 127 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=1.485 $X2=8.33 $Y2=1.69
r372 9 124 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=7.33
+ $Y=1.485 $X2=7.47 $Y2=1.69
r373 8 119 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.345
+ $Y=0.235 $X2=13.485 $Y2=0.445
r374 7 111 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.485
+ $Y=0.235 $X2=12.625 $Y2=0.445
r375 6 101 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.625
+ $Y=0.235 $X2=11.765 $Y2=0.445
r376 5 91 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.765
+ $Y=0.235 $X2=10.905 $Y2=0.445
r377 4 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.91
+ $Y=0.235 $X2=10.05 $Y2=0.445
r378 3 71 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.05
+ $Y=0.235 $X2=9.19 $Y2=0.445
r379 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.235 $X2=8.33 $Y2=0.445
r380 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.33
+ $Y=0.235 $X2=7.47 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%VGND 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 52 54 58 62 66 68 72 78 82 86 90 94 96 100 102 106 110
+ 114 116 118 121 122 124 125 126 127 129 130 132 133 135 136 137 138 140 141
+ 142 159 177 186 194 198 202 208 210 213 216 219 223 226
c257 202 0 1.60903e-20 $X=4.835 $Y=0.24
c258 159 0 1.41095e-19 $X=6.05 $Y=0
c259 140 0 7.59816e-20 $X=12.925 $Y=0
r260 222 223 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r261 219 220 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r262 216 217 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r263 214 217 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r264 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r265 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r266 207 208 9.83789 $w=6.48e-07 $l=1.3e-07 $layer=LI1_cond $X=5.32 $Y=0.24
+ $X2=5.45 $Y2=0.24
r267 204 207 0.552036 $w=6.48e-07 $l=3e-08 $layer=LI1_cond $X=5.29 $Y=0.24
+ $X2=5.32 $Y2=0.24
r268 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r269 202 204 8.37255 $w=6.48e-07 $l=4.55e-07 $layer=LI1_cond $X=4.835 $Y=0.24
+ $X2=5.29 $Y2=0.24
r270 201 205 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r271 200 202 0.092006 $w=6.48e-07 $l=5e-09 $layer=LI1_cond $X=4.83 $Y=0.24
+ $X2=4.835 $Y2=0.24
r272 200 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r273 197 200 0.92006 $w=6.48e-07 $l=5e-08 $layer=LI1_cond $X=4.78 $Y=0.24
+ $X2=4.83 $Y2=0.24
r274 197 198 9.00983 $w=6.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=0.24
+ $X2=4.695 $Y2=0.24
r275 194 195 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r276 191 226 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r277 189 223 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r278 188 189 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r279 186 222 4.35621 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=13.785 $Y=0
+ $X2=14.022 $Y2=0
r280 186 188 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=13.785 $Y=0
+ $X2=13.57 $Y2=0
r281 185 189 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.57 $Y2=0
r282 185 220 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r283 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r284 182 219 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.315 $Y=0
+ $X2=12.19 $Y2=0
r285 182 184 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.315 $Y=0
+ $X2=12.65 $Y2=0
r286 181 220 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r287 181 217 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r288 180 181 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r289 178 216 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.455 $Y=0
+ $X2=11.33 $Y2=0
r290 178 180 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.455 $Y=0
+ $X2=11.73 $Y2=0
r291 177 219 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.065 $Y=0
+ $X2=12.19 $Y2=0
r292 177 180 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.065 $Y=0
+ $X2=11.73 $Y2=0
r293 176 214 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r294 175 176 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r295 173 176 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r296 172 173 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r297 170 173 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r298 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r299 167 170 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r300 167 211 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r301 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r302 164 210 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.31 $Y=0 $X2=6.18
+ $Y2=0
r303 164 166 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.31 $Y=0
+ $X2=6.67 $Y2=0
r304 163 211 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r305 163 205 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r306 162 208 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.45
+ $Y2=0
r307 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r308 159 210 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.05 $Y=0 $X2=6.18
+ $Y2=0
r309 159 162 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.05 $Y=0 $X2=5.75
+ $Y2=0
r310 158 201 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r311 158 195 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r312 157 198 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.37 $Y=0
+ $X2=4.695 $Y2=0
r313 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r314 155 194 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=3.94 $Y2=0
r315 155 157 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=4.37 $Y2=0
r316 153 195 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r317 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r318 150 153 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r319 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r320 147 150 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r321 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r322 144 191 4.18769 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.267 $Y2=0
r323 144 146 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=1.15 $Y2=0
r324 142 147 0.260356 $w=4.8e-07 $l=9.15e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=1.15 $Y2=0
r325 142 226 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r326 140 184 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.925 $Y=0
+ $X2=12.65 $Y2=0
r327 140 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.925 $Y=0
+ $X2=13.055 $Y2=0
r328 139 188 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.185 $Y=0
+ $X2=13.57 $Y2=0
r329 139 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=13.185 $Y=0
+ $X2=13.055 $Y2=0
r330 137 175 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=9.49 $Y=0 $X2=9.43
+ $Y2=0
r331 137 138 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=9.49 $Y=0
+ $X2=9.612 $Y2=0
r332 135 172 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.63 $Y=0
+ $X2=8.51 $Y2=0
r333 135 136 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.63 $Y=0 $X2=8.76
+ $Y2=0
r334 134 175 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.89 $Y=0
+ $X2=9.43 $Y2=0
r335 134 136 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.89 $Y=0 $X2=8.76
+ $Y2=0
r336 132 169 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.77 $Y=0
+ $X2=7.59 $Y2=0
r337 132 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.9
+ $Y2=0
r338 131 172 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.03 $Y=0
+ $X2=8.51 $Y2=0
r339 131 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=7.9
+ $Y2=0
r340 129 166 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.91 $Y=0
+ $X2=6.67 $Y2=0
r341 129 130 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.91 $Y=0 $X2=7.04
+ $Y2=0
r342 128 169 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.17 $Y=0
+ $X2=7.59 $Y2=0
r343 128 130 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.04
+ $Y2=0
r344 126 152 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=0
+ $X2=2.99 $Y2=0
r345 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.1
+ $Y2=0
r346 124 149 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.175 $Y=0
+ $X2=2.07 $Y2=0
r347 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0
+ $X2=2.26 $Y2=0
r348 123 152 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.99 $Y2=0
r349 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.26 $Y2=0
r350 121 146 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.215 $Y=0
+ $X2=1.15 $Y2=0
r351 121 122 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.215 $Y=0
+ $X2=1.36 $Y2=0
r352 120 149 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.505 $Y=0
+ $X2=2.07 $Y2=0
r353 120 122 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.505 $Y=0
+ $X2=1.36 $Y2=0
r354 116 222 3.16147 $w=3e-07 $l=1.22327e-07 $layer=LI1_cond $X=13.935 $Y=0.085
+ $X2=14.022 $Y2=0
r355 116 118 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=13.935 $Y=0.085
+ $X2=13.935 $Y2=0.4
r356 112 141 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=13.055 $Y=0.085
+ $X2=13.055 $Y2=0
r357 112 114 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=13.055 $Y=0.085
+ $X2=13.055 $Y2=0.4
r358 108 219 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.19 $Y=0.085
+ $X2=12.19 $Y2=0
r359 108 110 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=12.19 $Y=0.085
+ $X2=12.19 $Y2=0.4
r360 104 216 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.33 $Y=0.085
+ $X2=11.33 $Y2=0
r361 104 106 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=11.33 $Y=0.085
+ $X2=11.33 $Y2=0.4
r362 103 213 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.472 $Y2=0
r363 102 216 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.205 $Y=0
+ $X2=11.33 $Y2=0
r364 102 103 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.205 $Y=0
+ $X2=10.595 $Y2=0
r365 98 213 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.472 $Y=0.085
+ $X2=10.472 $Y2=0
r366 98 100 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=10.472 $Y=0.085
+ $X2=10.472 $Y2=0.4
r367 97 138 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.612 $Y2=0
r368 96 213 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=10.35 $Y=0
+ $X2=10.472 $Y2=0
r369 96 97 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.35 $Y=0
+ $X2=9.735 $Y2=0
r370 92 138 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=9.612 $Y=0.085
+ $X2=9.612 $Y2=0
r371 92 94 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=9.612 $Y=0.085
+ $X2=9.612 $Y2=0.4
r372 88 136 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=0.085
+ $X2=8.76 $Y2=0
r373 88 90 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=8.76 $Y=0.085
+ $X2=8.76 $Y2=0.4
r374 84 133 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.085
+ $X2=7.9 $Y2=0
r375 84 86 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=7.9 $Y=0.085
+ $X2=7.9 $Y2=0.4
r376 80 130 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=0.085
+ $X2=7.04 $Y2=0
r377 80 82 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=7.04 $Y=0.085
+ $X2=7.04 $Y2=0.445
r378 76 210 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.18 $Y2=0
r379 76 78 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.18 $Y2=0.445
r380 70 194 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.94 $Y=0.085
+ $X2=3.94 $Y2=0
r381 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.94 $Y=0.085
+ $X2=3.94 $Y2=0.39
r382 69 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.1
+ $Y2=0
r383 68 194 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.94
+ $Y2=0
r384 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=3.185 $Y2=0
r385 64 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0
r386 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r387 60 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0
r388 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0.39
r389 56 122 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0
r390 56 58 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0.39
r391 52 191 3.25015 $w=2.9e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.39 $Y=0.085
+ $X2=0.267 $Y2=0
r392 52 54 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=0.39 $Y=0.085
+ $X2=0.39 $Y2=0.39
r393 17 118 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=13.775
+ $Y=0.235 $X2=13.915 $Y2=0.4
r394 16 114 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=12.915
+ $Y=0.235 $X2=13.055 $Y2=0.4
r395 15 110 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=12.055
+ $Y=0.235 $X2=12.195 $Y2=0.4
r396 14 106 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=11.195
+ $Y=0.235 $X2=11.335 $Y2=0.4
r397 13 100 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=10.34
+ $Y=0.235 $X2=10.48 $Y2=0.4
r398 12 94 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.48
+ $Y=0.235 $X2=9.62 $Y2=0.4
r399 11 90 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.62
+ $Y=0.235 $X2=8.76 $Y2=0.4
r400 10 86 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.76
+ $Y=0.235 $X2=7.9 $Y2=0.4
r401 9 82 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.235 $X2=7.04 $Y2=0.445
r402 8 78 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.235 $X2=6.18 $Y2=0.445
r403 7 207 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.195
+ $Y=0.235 $X2=5.32 $Y2=0.38
r404 6 197 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.645
+ $Y=0.235 $X2=4.78 $Y2=0.39
r405 5 72 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.235 $X2=3.94 $Y2=0.39
r406 4 66 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.965
+ $Y=0.235 $X2=3.1 $Y2=0.39
r407 3 62 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.235 $X2=2.26 $Y2=0.39
r408 2 58 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=1.295
+ $Y=0.235 $X2=1.42 $Y2=0.39
r409 1 54 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.315
+ $Y=0.235 $X2=0.45 $Y2=0.39
.ends


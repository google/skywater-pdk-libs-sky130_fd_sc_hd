* File: sky130_fd_sc_hd__mux2i_2.spice
* Created: Tue Sep  1 19:14:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2i_2.pex.spice"
.subckt sky130_fd_sc_hd__mux2i_2  VNB VPB S A0 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_S_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1004 N_A_193_47#_M1004_d N_S_M1004_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1009 N_A_193_47#_M1004_d N_S_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1008 N_A_361_47#_M1008_d N_A_27_47#_M1008_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_A_361_47#_M1008_d N_A_27_47#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_A0_M1002_g N_A_361_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_A0_M1005_g N_A_361_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.08775 PD=0.96 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1005_d N_A1_M1006_g N_A_193_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.089375 PD=0.96 PS=0.925 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1017 N_Y_M1017_d N_A1_M1017_g N_A_193_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.29575 AS=0.089375 PD=2.21 PS=0.925 NRD=35.076 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_S_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1010_d N_S_M1000_g N_A_193_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_S_M1001_g N_A_193_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1001_d N_A_27_47#_M1011_g N_A_361_297#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_27_47#_M1014_g N_A_361_297#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_193_297#_M1003_d N_A0_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_193_297#_M1003_d N_A0_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.155 PD=1.27 PS=1.31 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75000.6
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1012_s N_A1_M1007_g N_A_361_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.1375 PD=1.31 PS=1.275 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1015_d N_A1_M1015_g N_A_361_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.455 AS=0.1375 PD=2.91 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.4 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
c_43 VNB 0 1.34758e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__mux2i_2.pxi.spice"
*
.ends
*
*

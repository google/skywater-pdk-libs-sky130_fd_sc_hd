# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__lpflow_inputiso1n_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.735000 2.415000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.325000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.335000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.990000  1.495000 2.235000 1.665000 ;
      RECT 0.990000  1.665000 1.410000 1.915000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.495000  0.655000 2.235000 0.825000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.295000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1n_1
END LIBRARY

* File: sky130_fd_sc_hd__o22a_2.spice
* Created: Thu Aug 27 14:37:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o22a_2.pex.spice"
.subckt sky130_fd_sc_hd__o22a_2  VNB VPB B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_81_21#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1000_d N_A_81_21#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_81_21#_M1004_d N_B1_M1004_g N_A_301_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_301_47#_M1008_d N_B2_M1008_g N_A_81_21#_M1004_d VNB NSHORT L=0.15
+ W=0.65 AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_301_47#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_301_47#_M1009_d N_A1_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_81_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1001_d N_A_81_21#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.39 PD=1.27 PS=1.78 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75000.6
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1006 A_383_297# N_B1_M1006_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.39 PD=1.21 PS=1.78 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75001.6 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1007 N_A_81_21#_M1007_d N_B2_M1007_g A_383_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.235 AS=0.105 PD=1.47 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.9
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1003 A_579_297# N_A2_M1003_g N_A_81_21#_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.235 PD=1.21 PS=1.47 NRD=9.8303 NRS=38.3953 M=1 R=6.66667
+ SA=75002.5 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g A_579_297# VPB PHIGHVT L=0.15 W=1 AD=0.28
+ AS=0.105 PD=2.56 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.9 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__o22a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_isobufsrc_1.spice
* Created: Tue Sep  1 19:12:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_isobufsrc_1.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_isobufsrc_1  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_74_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_SLEEP_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.121799 PD=0.92 PS=1.19673 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_74_47#_M1004_g N_X_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_74_47#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0930507 AS=0.1092 PD=0.822254 PS=1.36 NRD=78.1105 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 A_265_297# N_SLEEP_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.221549 PD=1.21 PS=1.95775 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.4
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_74_47#_M1002_g A_265_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75000.8 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__lpflow_isobufsrc_1.pxi.spice"
*
.ends
*
*

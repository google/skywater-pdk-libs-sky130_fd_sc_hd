* File: sky130_fd_sc_hd__ebufn_8.pxi.spice
* Created: Thu Aug 27 14:19:40 2020
* 
x_PM_SKY130_FD_SC_HD__EBUFN_8%A N_A_c_156_n N_A_M1004_g N_A_M1019_g N_A_c_157_n
+ N_A_M1020_g N_A_M1036_g A A PM_SKY130_FD_SC_HD__EBUFN_8%A
x_PM_SKY130_FD_SC_HD__EBUFN_8%TE_B N_TE_B_c_205_n N_TE_B_M1031_g N_TE_B_M1025_g
+ N_TE_B_c_212_n N_TE_B_c_213_n N_TE_B_M1002_g N_TE_B_c_214_n N_TE_B_c_215_n
+ N_TE_B_M1008_g N_TE_B_c_216_n N_TE_B_c_217_n N_TE_B_M1011_g N_TE_B_c_218_n
+ N_TE_B_c_219_n N_TE_B_M1016_g N_TE_B_c_220_n N_TE_B_c_221_n N_TE_B_M1017_g
+ N_TE_B_c_222_n N_TE_B_c_223_n N_TE_B_M1022_g N_TE_B_c_224_n N_TE_B_c_225_n
+ N_TE_B_M1028_g N_TE_B_c_226_n N_TE_B_c_227_n N_TE_B_M1037_g N_TE_B_c_206_n
+ N_TE_B_c_207_n N_TE_B_c_230_n N_TE_B_c_231_n N_TE_B_c_232_n N_TE_B_c_233_n
+ N_TE_B_c_234_n N_TE_B_c_235_n N_TE_B_c_236_n N_TE_B_c_208_n N_TE_B_c_209_n
+ TE_B TE_B PM_SKY130_FD_SC_HD__EBUFN_8%TE_B
x_PM_SKY130_FD_SC_HD__EBUFN_8%A_301_47# N_A_301_47#_M1031_d N_A_301_47#_M1025_d
+ N_A_301_47#_c_377_n N_A_301_47#_M1000_g N_A_301_47#_c_378_n
+ N_A_301_47#_c_379_n N_A_301_47#_c_380_n N_A_301_47#_M1005_g
+ N_A_301_47#_c_381_n N_A_301_47#_c_382_n N_A_301_47#_M1007_g
+ N_A_301_47#_c_383_n N_A_301_47#_c_384_n N_A_301_47#_M1010_g
+ N_A_301_47#_c_385_n N_A_301_47#_c_386_n N_A_301_47#_M1012_g
+ N_A_301_47#_c_387_n N_A_301_47#_c_388_n N_A_301_47#_M1014_g
+ N_A_301_47#_c_389_n N_A_301_47#_c_390_n N_A_301_47#_M1015_g
+ N_A_301_47#_c_391_n N_A_301_47#_c_392_n N_A_301_47#_M1021_g
+ N_A_301_47#_c_393_n N_A_301_47#_c_394_n N_A_301_47#_c_395_n
+ N_A_301_47#_c_396_n N_A_301_47#_c_397_n N_A_301_47#_c_398_n
+ N_A_301_47#_c_402_n N_A_301_47#_c_399_n N_A_301_47#_c_400_n
+ N_A_301_47#_c_401_n N_A_301_47#_c_403_n N_A_301_47#_c_404_n
+ N_A_301_47#_c_440_n PM_SKY130_FD_SC_HD__EBUFN_8%A_301_47#
x_PM_SKY130_FD_SC_HD__EBUFN_8%A_116_47# N_A_116_47#_M1004_s N_A_116_47#_M1019_s
+ N_A_116_47#_M1001_g N_A_116_47#_M1003_g N_A_116_47#_M1006_g
+ N_A_116_47#_M1009_g N_A_116_47#_M1026_g N_A_116_47#_M1013_g
+ N_A_116_47#_M1027_g N_A_116_47#_M1018_g N_A_116_47#_M1029_g
+ N_A_116_47#_M1023_g N_A_116_47#_M1032_g N_A_116_47#_M1024_g
+ N_A_116_47#_M1033_g N_A_116_47#_M1030_g N_A_116_47#_M1034_g
+ N_A_116_47#_M1035_g N_A_116_47#_c_539_n N_A_116_47#_c_583_p
+ N_A_116_47#_c_540_n N_A_116_47#_c_541_n N_A_116_47#_c_552_n
+ N_A_116_47#_c_553_n N_A_116_47#_c_542_n N_A_116_47#_c_579_n
+ N_A_116_47#_c_543_n PM_SKY130_FD_SC_HD__EBUFN_8%A_116_47#
x_PM_SKY130_FD_SC_HD__EBUFN_8%VPWR N_VPWR_M1019_d N_VPWR_M1036_d N_VPWR_M1002_s
+ N_VPWR_M1011_s N_VPWR_M1017_s N_VPWR_M1028_s N_VPWR_c_675_n N_VPWR_c_676_n
+ N_VPWR_c_677_n N_VPWR_c_678_n N_VPWR_c_679_n N_VPWR_c_680_n N_VPWR_c_681_n
+ N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_684_n N_VPWR_c_685_n VPWR
+ N_VPWR_c_686_n N_VPWR_c_687_n N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_674_n
+ N_VPWR_c_691_n N_VPWR_c_692_n N_VPWR_c_693_n PM_SKY130_FD_SC_HD__EBUFN_8%VPWR
x_PM_SKY130_FD_SC_HD__EBUFN_8%A_407_309# N_A_407_309#_M1002_d
+ N_A_407_309#_M1008_d N_A_407_309#_M1016_d N_A_407_309#_M1022_d
+ N_A_407_309#_M1037_d N_A_407_309#_M1009_d N_A_407_309#_M1018_d
+ N_A_407_309#_M1024_d N_A_407_309#_M1035_d N_A_407_309#_c_811_n
+ N_A_407_309#_c_814_n N_A_407_309#_c_812_n N_A_407_309#_c_856_n
+ N_A_407_309#_c_818_n N_A_407_309#_c_863_n N_A_407_309#_c_821_n
+ N_A_407_309#_c_870_n N_A_407_309#_c_872_n N_A_407_309#_c_813_n
+ N_A_407_309#_c_824_n N_A_407_309#_c_825_n N_A_407_309#_c_826_n
+ N_A_407_309#_c_827_n PM_SKY130_FD_SC_HD__EBUFN_8%A_407_309#
x_PM_SKY130_FD_SC_HD__EBUFN_8%Z N_Z_M1001_d N_Z_M1026_d N_Z_M1029_d N_Z_M1033_d
+ N_Z_M1003_s N_Z_M1013_s N_Z_M1023_s N_Z_M1030_s N_Z_c_936_n Z Z Z Z Z Z Z Z Z
+ Z Z Z Z Z Z Z Z N_Z_c_906_n N_Z_c_903_n PM_SKY130_FD_SC_HD__EBUFN_8%Z
x_PM_SKY130_FD_SC_HD__EBUFN_8%VGND N_VGND_M1004_d N_VGND_M1020_d N_VGND_M1000_s
+ N_VGND_M1007_s N_VGND_M1012_s N_VGND_M1015_s N_VGND_c_1010_n N_VGND_c_1011_n
+ N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n
+ N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n
+ N_VGND_c_1020_n N_VGND_c_1021_n VGND N_VGND_c_1022_n N_VGND_c_1023_n
+ N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n
+ N_VGND_c_1028_n PM_SKY130_FD_SC_HD__EBUFN_8%VGND
x_PM_SKY130_FD_SC_HD__EBUFN_8%A_455_47# N_A_455_47#_M1000_d N_A_455_47#_M1005_d
+ N_A_455_47#_M1010_d N_A_455_47#_M1014_d N_A_455_47#_M1021_d
+ N_A_455_47#_M1006_s N_A_455_47#_M1027_s N_A_455_47#_M1032_s
+ N_A_455_47#_M1034_s N_A_455_47#_c_1144_n N_A_455_47#_c_1150_n
+ N_A_455_47#_c_1145_n N_A_455_47#_c_1223_n N_A_455_47#_c_1156_n
+ N_A_455_47#_c_1230_n N_A_455_47#_c_1160_n N_A_455_47#_c_1237_n
+ N_A_455_47#_c_1164_n N_A_455_47#_c_1146_n N_A_455_47#_c_1168_n
+ N_A_455_47#_c_1170_n N_A_455_47#_c_1172_n N_A_455_47#_c_1174_n
+ PM_SKY130_FD_SC_HD__EBUFN_8%A_455_47#
cc_1 VNB N_A_c_156_n 0.0211382f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=0.995
cc_2 VNB N_A_c_157_n 0.0509135f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.025
cc_3 VNB N_A_M1020_g 0.0173303f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.56
cc_4 VNB N_A_M1036_g 3.85873e-19 $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_5 VNB A 0.0148258f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_TE_B_c_205_n 0.0201327f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=0.995
cc_7 VNB N_TE_B_c_206_n 0.0249493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_TE_B_c_207_n 0.0201621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_TE_B_c_208_n 0.00186481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_TE_B_c_209_n 0.0169692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB TE_B 7.59431e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_301_47#_c_377_n 0.01763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_301_47#_c_378_n 0.00893548f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.56
cc_14 VNB N_A_301_47#_c_379_n 0.00752986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_301_47#_c_380_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.295
cc_16 VNB N_A_301_47#_c_381_n 0.00893472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_301_47#_c_382_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_18 VNB N_A_301_47#_c_383_n 0.00893548f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_19 VNB N_A_301_47#_c_384_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_20 VNB N_A_301_47#_c_385_n 0.00893472f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_21 VNB N_A_301_47#_c_386_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_301_47#_c_387_n 0.00893548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_301_47#_c_388_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_301_47#_c_389_n 0.00893472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_301_47#_c_390_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_301_47#_c_391_n 0.010572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_301_47#_c_392_n 0.0580155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_301_47#_c_393_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_301_47#_c_394_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_301_47#_c_395_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_301_47#_c_396_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_301_47#_c_397_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_301_47#_c_398_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_301_47#_c_399_n 0.00306725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_301_47#_c_400_n 0.0301483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_301_47#_c_401_n 0.0103832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_116_47#_M1001_g 0.0194198f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.56
cc_38 VNB N_A_116_47#_M1003_g 7.20486e-19 $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_39 VNB N_A_116_47#_M1006_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_40 VNB N_A_116_47#_M1009_g 3.77304e-19 $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_41 VNB N_A_116_47#_M1026_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_42 VNB N_A_116_47#_M1013_g 4.50174e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_116_47#_M1027_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_116_47#_M1018_g 4.50204e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_116_47#_M1029_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_116_47#_M1023_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_116_47#_M1032_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_116_47#_M1024_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_116_47#_M1033_g 0.0175011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_116_47#_M1030_g 4.49895e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_116_47#_M1034_g 0.0208147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_116_47#_M1035_g 4.89476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_116_47#_c_539_n 0.00161246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_116_47#_c_540_n 9.112e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_116_47#_c_541_n 0.00496447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_116_47#_c_542_n 3.01405e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_116_47#_c_543_n 0.128942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_674_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB Z 0.0224043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_Z_c_903_n 0.010637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1010_n 0.0106829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1011_n 0.0265872f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_63 VNB N_VGND_c_1012_n 0.00269826f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_64 VNB N_VGND_c_1013_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1014_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1015_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1016_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1017_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1018_n 0.0331239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1019_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1020_n 0.0110833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1021_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1022_n 0.0129098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1023_n 0.0110833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1024_n 0.0949418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1025_n 0.45679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1026_n 0.00516315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1027_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1028_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_455_47#_c_1144_n 0.00570911f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.53
cc_81 VNB N_A_455_47#_c_1145_n 0.00313518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_455_47#_c_1146_n 0.00882053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VPB N_A_M1019_g 0.0209796f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_84 VPB N_A_c_157_n 0.00948833f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.025
cc_85 VPB N_A_M1036_g 0.0193862f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_86 VPB A 0.0132012f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_87 VPB N_TE_B_M1025_g 0.0231272f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_88 VPB N_TE_B_c_212_n 0.0146714f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=0.56
cc_89 VPB N_TE_B_c_213_n 0.0172196f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.295
cc_90 VPB N_TE_B_c_214_n 0.0120194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_TE_B_c_215_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_92 VPB N_TE_B_c_216_n 0.0113042f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_93 VPB N_TE_B_c_217_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_94 VPB N_TE_B_c_218_n 0.0113042f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.16
cc_95 VPB N_TE_B_c_219_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_TE_B_c_220_n 0.0113042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_TE_B_c_221_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_TE_B_c_222_n 0.0113042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_TE_B_c_223_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_TE_B_c_224_n 0.0113042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_TE_B_c_225_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_TE_B_c_226_n 0.0238745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_TE_B_c_227_n 0.0172196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_TE_B_c_206_n 0.0143708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_TE_B_c_207_n 0.0127472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_TE_B_c_230_n 0.00612638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_TE_B_c_231_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_TE_B_c_232_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_TE_B_c_233_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_TE_B_c_234_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_TE_B_c_235_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_TE_B_c_236_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_TE_B_c_208_n 0.00186481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_TE_B_c_209_n 0.00494597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB TE_B 0.00111102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_301_47#_c_402_n 0.00893068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_301_47#_c_403_n 0.00156037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_301_47#_c_404_n 0.00259185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_116_47#_M1003_g 0.0267252f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_120 VPB N_A_116_47#_M1009_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_121 VPB N_A_116_47#_M1013_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_116_47#_M1018_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_116_47#_M1023_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_116_47#_M1024_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_116_47#_M1030_g 0.0191665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_116_47#_M1035_g 0.0230841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_116_47#_c_552_n 0.00212132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_116_47#_c_553_n 0.00213905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_116_47#_c_542_n 9.7779e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_675_n 0.010657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_676_n 0.0309481f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_132 VPB N_VPWR_c_677_n 0.00269826f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.16
cc_133 VPB N_VPWR_c_678_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_679_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_680_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_681_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_682_n 0.0110228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_683_n 0.00436274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_684_n 0.0110228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_685_n 0.00436274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_686_n 0.0128277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_687_n 0.0277448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_688_n 0.0110228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_689_n 0.100337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_674_n 0.0525071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_691_n 0.00517167f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_692_n 0.00436274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_693_n 0.00436274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_407_309#_c_811_n 0.00372278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_407_309#_c_812_n 0.00176412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_407_309#_c_813_n 0.0249987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB Z 0.00710692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB Z 0.0125296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_Z_c_906_n 0.0242819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 N_A_M1020_g N_TE_B_c_205_n 0.0217987f $X=0.925 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_M1036_g N_TE_B_M1025_g 0.0276113f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_c_157_n N_TE_B_c_208_n 0.00607751f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_158 N_A_M1020_g N_TE_B_c_208_n 5.64945e-19 $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A_M1036_g N_TE_B_c_208_n 5.61895e-19 $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1020_g N_TE_B_c_209_n 0.0214892f $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_161 N_A_M1020_g TE_B 0.008883f $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_M1036_g TE_B 0.00876899f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_M1036_g N_A_301_47#_c_402_n 4.44593e-19 $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1020_g N_A_301_47#_c_401_n 4.37219e-19 $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A_c_156_n N_A_116_47#_c_539_n 0.00371724f $X=0.505 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_M1020_g N_A_116_47#_c_539_n 0.00197811f $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_c_157_n N_A_116_47#_c_540_n 0.00540459f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_168 A N_A_116_47#_c_540_n 0.0345883f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A_c_157_n N_A_116_47#_c_541_n 0.0110937f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_170 N_A_c_157_n N_A_116_47#_c_552_n 0.00805321f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_171 A N_A_116_47#_c_552_n 0.0067549f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A_c_157_n N_A_116_47#_c_553_n 0.0109241f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_173 N_A_M1036_g N_A_116_47#_c_553_n 0.00375437f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_174 A N_VPWR_M1019_d 0.00400735f $X=0.145 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_175 N_A_M1019_g N_VPWR_c_676_n 0.0127975f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_c_157_n N_VPWR_c_676_n 0.00103558f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_177 N_A_M1036_g N_VPWR_c_676_n 6.68863e-19 $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_178 A N_VPWR_c_676_n 0.025872f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A_M1019_g N_VPWR_c_677_n 6.69841e-19 $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_M1036_g N_VPWR_c_677_n 0.0108177f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_M1019_g N_VPWR_c_686_n 0.00525069f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1036_g N_VPWR_c_686_n 0.0046653f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1019_g N_VPWR_c_674_n 0.00888907f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_M1036_g N_VPWR_c_674_n 0.00796766f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_c_156_n N_VGND_c_1011_n 0.0110579f $X=0.505 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_157_n N_VGND_c_1011_n 0.00195936f $X=0.925 $Y=1.025 $X2=0 $Y2=0
cc_187 N_A_M1020_g N_VGND_c_1011_n 6.39688e-19 $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_188 A N_VGND_c_1011_n 0.0276701f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_189 N_A_c_156_n N_VGND_c_1012_n 5.51156e-19 $X=0.505 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_M1020_g N_VGND_c_1012_n 0.00672509f $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_c_156_n N_VGND_c_1022_n 0.00525069f $X=0.505 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_M1020_g N_VGND_c_1022_n 0.0046653f $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_c_156_n N_VGND_c_1025_n 0.00888907f $X=0.505 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_M1020_g N_VGND_c_1025_n 0.00796766f $X=0.925 $Y=0.56 $X2=0 $Y2=0
cc_195 N_TE_B_c_231_n N_A_301_47#_c_378_n 0.0139594f $X=2.79 $Y=1.395 $X2=0
+ $Y2=0
cc_196 N_TE_B_c_214_n N_A_301_47#_c_379_n 0.0139594f $X=2.715 $Y=1.395 $X2=0
+ $Y2=0
cc_197 N_TE_B_c_207_n N_A_301_47#_c_379_n 0.00292154f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_198 N_TE_B_c_232_n N_A_301_47#_c_381_n 0.0139594f $X=3.21 $Y=1.395 $X2=0
+ $Y2=0
cc_199 N_TE_B_c_233_n N_A_301_47#_c_383_n 0.0139594f $X=3.63 $Y=1.395 $X2=0
+ $Y2=0
cc_200 N_TE_B_c_234_n N_A_301_47#_c_385_n 0.0139594f $X=4.05 $Y=1.395 $X2=0
+ $Y2=0
cc_201 N_TE_B_c_235_n N_A_301_47#_c_387_n 0.0139594f $X=4.47 $Y=1.395 $X2=0
+ $Y2=0
cc_202 N_TE_B_c_236_n N_A_301_47#_c_389_n 0.0139594f $X=4.89 $Y=1.395 $X2=0
+ $Y2=0
cc_203 N_TE_B_c_216_n N_A_301_47#_c_393_n 0.0139594f $X=3.135 $Y=1.395 $X2=0
+ $Y2=0
cc_204 N_TE_B_c_218_n N_A_301_47#_c_394_n 0.0139594f $X=3.555 $Y=1.395 $X2=0
+ $Y2=0
cc_205 N_TE_B_c_220_n N_A_301_47#_c_395_n 0.0139594f $X=3.975 $Y=1.395 $X2=0
+ $Y2=0
cc_206 N_TE_B_c_222_n N_A_301_47#_c_396_n 0.0139594f $X=4.395 $Y=1.395 $X2=0
+ $Y2=0
cc_207 N_TE_B_c_224_n N_A_301_47#_c_397_n 0.0139594f $X=4.815 $Y=1.395 $X2=0
+ $Y2=0
cc_208 N_TE_B_c_226_n N_A_301_47#_c_398_n 0.0139594f $X=5.235 $Y=1.395 $X2=0
+ $Y2=0
cc_209 N_TE_B_M1025_g N_A_301_47#_c_402_n 0.0103039f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_TE_B_c_213_n N_A_301_47#_c_402_n 0.00594189f $X=2.37 $Y=1.47 $X2=0
+ $Y2=0
cc_211 N_TE_B_c_205_n N_A_301_47#_c_399_n 0.00395306f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_TE_B_c_206_n N_A_301_47#_c_399_n 0.00909263f $X=1.92 $Y=1.232 $X2=0
+ $Y2=0
cc_213 N_TE_B_c_207_n N_A_301_47#_c_399_n 0.00229794f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_214 N_TE_B_c_208_n N_A_301_47#_c_399_n 0.00229846f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_215 TE_B N_A_301_47#_c_399_n 0.0078712f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_216 N_TE_B_c_212_n N_A_301_47#_c_400_n 0.0337992f $X=2.295 $Y=1.395 $X2=0
+ $Y2=0
cc_217 N_TE_B_c_207_n N_A_301_47#_c_400_n 0.012186f $X=2.07 $Y=1.232 $X2=0 $Y2=0
cc_218 N_TE_B_c_205_n N_A_301_47#_c_401_n 0.0127852f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_TE_B_c_206_n N_A_301_47#_c_401_n 0.00226063f $X=1.92 $Y=1.232 $X2=0
+ $Y2=0
cc_220 N_TE_B_M1025_g N_A_301_47#_c_403_n 0.00256246f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_TE_B_c_206_n N_A_301_47#_c_403_n 0.00228019f $X=1.92 $Y=1.232 $X2=0
+ $Y2=0
cc_222 N_TE_B_M1025_g N_A_301_47#_c_404_n 0.0018143f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_TE_B_c_213_n N_A_301_47#_c_404_n 9.88549e-19 $X=2.37 $Y=1.47 $X2=0
+ $Y2=0
cc_224 N_TE_B_c_206_n N_A_301_47#_c_404_n 0.00919668f $X=1.92 $Y=1.232 $X2=0
+ $Y2=0
cc_225 N_TE_B_c_207_n N_A_301_47#_c_404_n 0.00362194f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_226 N_TE_B_c_208_n N_A_301_47#_c_404_n 0.00370765f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_227 TE_B N_A_301_47#_c_404_n 0.0089926f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_228 N_TE_B_c_206_n N_A_301_47#_c_440_n 0.0142077f $X=1.92 $Y=1.232 $X2=0
+ $Y2=0
cc_229 N_TE_B_c_207_n N_A_301_47#_c_440_n 0.00445721f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_230 N_TE_B_c_208_n N_A_301_47#_c_440_n 0.0182328f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_231 TE_B N_A_116_47#_c_539_n 0.0202069f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_232 N_TE_B_c_208_n N_A_116_47#_c_540_n 0.0202069f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_233 N_TE_B_c_209_n N_A_116_47#_c_540_n 2.37905e-19 $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_234 N_TE_B_c_206_n N_A_116_47#_c_541_n 0.00162963f $X=1.92 $Y=1.232 $X2=0
+ $Y2=0
cc_235 N_TE_B_c_208_n N_A_116_47#_c_541_n 0.0436136f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_236 N_TE_B_c_209_n N_A_116_47#_c_541_n 0.00444123f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_237 N_TE_B_c_208_n N_A_116_47#_c_552_n 0.00237639f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_238 TE_B N_A_116_47#_c_553_n 0.0202069f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_239 TE_B N_VPWR_M1036_d 0.00388689f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_240 N_TE_B_M1025_g N_VPWR_c_677_n 0.00624081f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_241 N_TE_B_c_209_n N_VPWR_c_677_n 3.3572e-19 $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_242 TE_B N_VPWR_c_677_n 0.0235828f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_243 N_TE_B_c_213_n N_VPWR_c_678_n 0.00856801f $X=2.37 $Y=1.47 $X2=0 $Y2=0
cc_244 N_TE_B_c_215_n N_VPWR_c_678_n 0.00685342f $X=2.79 $Y=1.47 $X2=0 $Y2=0
cc_245 N_TE_B_c_217_n N_VPWR_c_678_n 5.14696e-19 $X=3.21 $Y=1.47 $X2=0 $Y2=0
cc_246 N_TE_B_c_215_n N_VPWR_c_679_n 5.14696e-19 $X=2.79 $Y=1.47 $X2=0 $Y2=0
cc_247 N_TE_B_c_217_n N_VPWR_c_679_n 0.00685342f $X=3.21 $Y=1.47 $X2=0 $Y2=0
cc_248 N_TE_B_c_219_n N_VPWR_c_679_n 0.00685342f $X=3.63 $Y=1.47 $X2=0 $Y2=0
cc_249 N_TE_B_c_221_n N_VPWR_c_679_n 5.14696e-19 $X=4.05 $Y=1.47 $X2=0 $Y2=0
cc_250 N_TE_B_c_219_n N_VPWR_c_680_n 5.14696e-19 $X=3.63 $Y=1.47 $X2=0 $Y2=0
cc_251 N_TE_B_c_221_n N_VPWR_c_680_n 0.00685342f $X=4.05 $Y=1.47 $X2=0 $Y2=0
cc_252 N_TE_B_c_223_n N_VPWR_c_680_n 0.00685342f $X=4.47 $Y=1.47 $X2=0 $Y2=0
cc_253 N_TE_B_c_225_n N_VPWR_c_680_n 5.14696e-19 $X=4.89 $Y=1.47 $X2=0 $Y2=0
cc_254 N_TE_B_c_223_n N_VPWR_c_681_n 5.14696e-19 $X=4.47 $Y=1.47 $X2=0 $Y2=0
cc_255 N_TE_B_c_225_n N_VPWR_c_681_n 0.00685342f $X=4.89 $Y=1.47 $X2=0 $Y2=0
cc_256 N_TE_B_c_227_n N_VPWR_c_681_n 0.00859487f $X=5.31 $Y=1.47 $X2=0 $Y2=0
cc_257 N_TE_B_c_219_n N_VPWR_c_682_n 0.00341689f $X=3.63 $Y=1.47 $X2=0 $Y2=0
cc_258 N_TE_B_c_221_n N_VPWR_c_682_n 0.00341689f $X=4.05 $Y=1.47 $X2=0 $Y2=0
cc_259 N_TE_B_c_223_n N_VPWR_c_684_n 0.00341689f $X=4.47 $Y=1.47 $X2=0 $Y2=0
cc_260 N_TE_B_c_225_n N_VPWR_c_684_n 0.00341689f $X=4.89 $Y=1.47 $X2=0 $Y2=0
cc_261 N_TE_B_M1025_g N_VPWR_c_687_n 0.00541359f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_262 N_TE_B_c_213_n N_VPWR_c_687_n 0.00341689f $X=2.37 $Y=1.47 $X2=0 $Y2=0
cc_263 N_TE_B_c_215_n N_VPWR_c_688_n 0.00341689f $X=2.79 $Y=1.47 $X2=0 $Y2=0
cc_264 N_TE_B_c_217_n N_VPWR_c_688_n 0.00341689f $X=3.21 $Y=1.47 $X2=0 $Y2=0
cc_265 N_TE_B_c_227_n N_VPWR_c_689_n 0.00341689f $X=5.31 $Y=1.47 $X2=0 $Y2=0
cc_266 N_TE_B_M1025_g N_VPWR_c_674_n 0.0111338f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_267 N_TE_B_c_213_n N_VPWR_c_674_n 0.00530897f $X=2.37 $Y=1.47 $X2=0 $Y2=0
cc_268 N_TE_B_c_215_n N_VPWR_c_674_n 0.0039829f $X=2.79 $Y=1.47 $X2=0 $Y2=0
cc_269 N_TE_B_c_217_n N_VPWR_c_674_n 0.0039829f $X=3.21 $Y=1.47 $X2=0 $Y2=0
cc_270 N_TE_B_c_219_n N_VPWR_c_674_n 0.0039829f $X=3.63 $Y=1.47 $X2=0 $Y2=0
cc_271 N_TE_B_c_221_n N_VPWR_c_674_n 0.0039829f $X=4.05 $Y=1.47 $X2=0 $Y2=0
cc_272 N_TE_B_c_223_n N_VPWR_c_674_n 0.0039829f $X=4.47 $Y=1.47 $X2=0 $Y2=0
cc_273 N_TE_B_c_225_n N_VPWR_c_674_n 0.0039829f $X=4.89 $Y=1.47 $X2=0 $Y2=0
cc_274 N_TE_B_c_227_n N_VPWR_c_674_n 0.00540327f $X=5.31 $Y=1.47 $X2=0 $Y2=0
cc_275 N_TE_B_c_213_n N_A_407_309#_c_814_n 0.0129586f $X=2.37 $Y=1.47 $X2=0
+ $Y2=0
cc_276 N_TE_B_c_214_n N_A_407_309#_c_814_n 3.62169e-19 $X=2.715 $Y=1.395 $X2=0
+ $Y2=0
cc_277 N_TE_B_c_215_n N_A_407_309#_c_814_n 0.0115215f $X=2.79 $Y=1.47 $X2=0
+ $Y2=0
cc_278 N_TE_B_c_207_n N_A_407_309#_c_812_n 0.00109405f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_279 N_TE_B_c_217_n N_A_407_309#_c_818_n 0.0115215f $X=3.21 $Y=1.47 $X2=0
+ $Y2=0
cc_280 N_TE_B_c_218_n N_A_407_309#_c_818_n 3.62169e-19 $X=3.555 $Y=1.395 $X2=0
+ $Y2=0
cc_281 N_TE_B_c_219_n N_A_407_309#_c_818_n 0.0115215f $X=3.63 $Y=1.47 $X2=0
+ $Y2=0
cc_282 N_TE_B_c_221_n N_A_407_309#_c_821_n 0.0115215f $X=4.05 $Y=1.47 $X2=0
+ $Y2=0
cc_283 N_TE_B_c_222_n N_A_407_309#_c_821_n 3.62169e-19 $X=4.395 $Y=1.395 $X2=0
+ $Y2=0
cc_284 N_TE_B_c_223_n N_A_407_309#_c_821_n 0.0115215f $X=4.47 $Y=1.47 $X2=0
+ $Y2=0
cc_285 N_TE_B_c_216_n N_A_407_309#_c_824_n 4.01342e-19 $X=3.135 $Y=1.395 $X2=0
+ $Y2=0
cc_286 N_TE_B_c_220_n N_A_407_309#_c_825_n 4.01342e-19 $X=3.975 $Y=1.395 $X2=0
+ $Y2=0
cc_287 N_TE_B_c_224_n N_A_407_309#_c_826_n 4.01342e-19 $X=4.815 $Y=1.395 $X2=0
+ $Y2=0
cc_288 N_TE_B_c_225_n N_A_407_309#_c_827_n 0.0115215f $X=4.89 $Y=1.47 $X2=0
+ $Y2=0
cc_289 N_TE_B_c_226_n N_A_407_309#_c_827_n 3.62169e-19 $X=5.235 $Y=1.395 $X2=0
+ $Y2=0
cc_290 N_TE_B_c_227_n N_A_407_309#_c_827_n 0.0136245f $X=5.31 $Y=1.47 $X2=0
+ $Y2=0
cc_291 N_TE_B_c_212_n N_Z_c_906_n 0.00664826f $X=2.295 $Y=1.395 $X2=0 $Y2=0
cc_292 N_TE_B_c_213_n N_Z_c_906_n 0.0136917f $X=2.37 $Y=1.47 $X2=0 $Y2=0
cc_293 N_TE_B_c_214_n N_Z_c_906_n 0.00442457f $X=2.715 $Y=1.395 $X2=0 $Y2=0
cc_294 N_TE_B_c_215_n N_Z_c_906_n 0.0115275f $X=2.79 $Y=1.47 $X2=0 $Y2=0
cc_295 N_TE_B_c_216_n N_Z_c_906_n 0.0043665f $X=3.135 $Y=1.395 $X2=0 $Y2=0
cc_296 N_TE_B_c_217_n N_Z_c_906_n 0.0115275f $X=3.21 $Y=1.47 $X2=0 $Y2=0
cc_297 N_TE_B_c_218_n N_Z_c_906_n 0.0043665f $X=3.555 $Y=1.395 $X2=0 $Y2=0
cc_298 N_TE_B_c_219_n N_Z_c_906_n 0.0115275f $X=3.63 $Y=1.47 $X2=0 $Y2=0
cc_299 N_TE_B_c_220_n N_Z_c_906_n 0.0043665f $X=3.975 $Y=1.395 $X2=0 $Y2=0
cc_300 N_TE_B_c_221_n N_Z_c_906_n 0.0115275f $X=4.05 $Y=1.47 $X2=0 $Y2=0
cc_301 N_TE_B_c_222_n N_Z_c_906_n 0.0043665f $X=4.395 $Y=1.395 $X2=0 $Y2=0
cc_302 N_TE_B_c_223_n N_Z_c_906_n 0.0115275f $X=4.47 $Y=1.47 $X2=0 $Y2=0
cc_303 N_TE_B_c_224_n N_Z_c_906_n 0.0043665f $X=4.815 $Y=1.395 $X2=0 $Y2=0
cc_304 N_TE_B_c_225_n N_Z_c_906_n 0.0115275f $X=4.89 $Y=1.47 $X2=0 $Y2=0
cc_305 N_TE_B_c_226_n N_Z_c_906_n 0.00643784f $X=5.235 $Y=1.395 $X2=0 $Y2=0
cc_306 N_TE_B_c_227_n N_Z_c_906_n 0.0146945f $X=5.31 $Y=1.47 $X2=0 $Y2=0
cc_307 N_TE_B_c_207_n N_Z_c_906_n 0.00279522f $X=2.07 $Y=1.232 $X2=0 $Y2=0
cc_308 N_TE_B_c_230_n N_Z_c_906_n 0.00156591f $X=2.37 $Y=1.395 $X2=0 $Y2=0
cc_309 N_TE_B_c_231_n N_Z_c_906_n 0.00146804f $X=2.79 $Y=1.395 $X2=0 $Y2=0
cc_310 N_TE_B_c_232_n N_Z_c_906_n 0.00146804f $X=3.21 $Y=1.395 $X2=0 $Y2=0
cc_311 N_TE_B_c_233_n N_Z_c_906_n 0.00146804f $X=3.63 $Y=1.395 $X2=0 $Y2=0
cc_312 N_TE_B_c_234_n N_Z_c_906_n 0.00146804f $X=4.05 $Y=1.395 $X2=0 $Y2=0
cc_313 N_TE_B_c_235_n N_Z_c_906_n 0.00146804f $X=4.47 $Y=1.395 $X2=0 $Y2=0
cc_314 N_TE_B_c_236_n N_Z_c_906_n 0.00146804f $X=4.89 $Y=1.395 $X2=0 $Y2=0
cc_315 TE_B N_VGND_M1020_d 0.00384013f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_316 N_TE_B_c_205_n N_VGND_c_1012_n 0.00409954f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_317 N_TE_B_c_209_n N_VGND_c_1012_n 3.24606e-19 $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_318 TE_B N_VGND_c_1012_n 0.0218659f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_319 N_TE_B_c_205_n N_VGND_c_1018_n 0.00541359f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_320 N_TE_B_c_205_n N_VGND_c_1025_n 0.0112237f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_321 TE_B N_VGND_c_1025_n 0.00173674f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_322 N_TE_B_c_205_n N_A_455_47#_c_1144_n 6.31784e-19 $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_TE_B_c_205_n N_A_455_47#_c_1145_n 3.46698e-19 $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_301_47#_c_392_n N_A_116_47#_M1001_g 0.0362291f $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_325 N_A_301_47#_c_392_n N_A_116_47#_c_541_n 7.53426e-19 $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_326 N_A_301_47#_c_400_n N_A_116_47#_c_541_n 0.16023f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_301_47#_c_401_n N_A_116_47#_c_541_n 0.0031471f $X=1.64 $Y=0.56 $X2=0
+ $Y2=0
cc_328 N_A_301_47#_c_403_n N_A_116_47#_c_541_n 0.00343878f $X=1.64 $Y=1.63 $X2=0
+ $Y2=0
cc_329 N_A_301_47#_c_440_n N_A_116_47#_c_541_n 0.0467388f $X=1.792 $Y=1.15 $X2=0
+ $Y2=0
cc_330 N_A_301_47#_c_400_n N_A_116_47#_c_542_n 2.36285e-19 $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_331 N_A_301_47#_c_392_n N_A_116_47#_c_579_n 4.24405e-19 $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_332 N_A_301_47#_c_400_n N_A_116_47#_c_579_n 0.0124827f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_A_301_47#_c_400_n N_A_116_47#_c_543_n 0.00100363f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_301_47#_c_402_n N_VPWR_c_687_n 0.0224721f $X=1.64 $Y=2.31 $X2=0 $Y2=0
cc_335 N_A_301_47#_M1025_d N_VPWR_c_674_n 0.00209319f $X=1.505 $Y=1.485 $X2=0
+ $Y2=0
cc_336 N_A_301_47#_c_402_n N_VPWR_c_674_n 0.013197f $X=1.64 $Y=2.31 $X2=0 $Y2=0
cc_337 N_A_301_47#_c_402_n N_A_407_309#_c_811_n 0.0327307f $X=1.64 $Y=2.31 $X2=0
+ $Y2=0
cc_338 N_A_301_47#_c_402_n N_A_407_309#_c_812_n 0.0151017f $X=1.64 $Y=2.31 $X2=0
+ $Y2=0
cc_339 N_A_301_47#_c_379_n N_Z_c_906_n 0.00214952f $X=2.685 $Y=1.035 $X2=0 $Y2=0
cc_340 N_A_301_47#_c_391_n N_Z_c_906_n 0.00101952f $X=5.475 $Y=1.035 $X2=0 $Y2=0
cc_341 N_A_301_47#_c_392_n N_Z_c_906_n 0.00780828f $X=5.55 $Y=0.96 $X2=0 $Y2=0
cc_342 N_A_301_47#_c_400_n N_Z_c_906_n 0.273878f $X=5.76 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_301_47#_c_404_n N_Z_c_906_n 0.0243711f $X=1.65 $Y=1.495 $X2=0 $Y2=0
cc_344 N_A_301_47#_c_377_n N_VGND_c_1013_n 0.00856801f $X=2.61 $Y=0.96 $X2=0
+ $Y2=0
cc_345 N_A_301_47#_c_380_n N_VGND_c_1013_n 0.00699289f $X=3.03 $Y=0.96 $X2=0
+ $Y2=0
cc_346 N_A_301_47#_c_382_n N_VGND_c_1013_n 6.07018e-19 $X=3.45 $Y=0.96 $X2=0
+ $Y2=0
cc_347 N_A_301_47#_c_380_n N_VGND_c_1014_n 6.07018e-19 $X=3.03 $Y=0.96 $X2=0
+ $Y2=0
cc_348 N_A_301_47#_c_382_n N_VGND_c_1014_n 0.00699289f $X=3.45 $Y=0.96 $X2=0
+ $Y2=0
cc_349 N_A_301_47#_c_384_n N_VGND_c_1014_n 0.00685342f $X=3.87 $Y=0.96 $X2=0
+ $Y2=0
cc_350 N_A_301_47#_c_386_n N_VGND_c_1014_n 5.54209e-19 $X=4.29 $Y=0.96 $X2=0
+ $Y2=0
cc_351 N_A_301_47#_c_384_n N_VGND_c_1015_n 0.00341689f $X=3.87 $Y=0.96 $X2=0
+ $Y2=0
cc_352 N_A_301_47#_c_386_n N_VGND_c_1015_n 0.00341689f $X=4.29 $Y=0.96 $X2=0
+ $Y2=0
cc_353 N_A_301_47#_c_384_n N_VGND_c_1016_n 5.54209e-19 $X=3.87 $Y=0.96 $X2=0
+ $Y2=0
cc_354 N_A_301_47#_c_386_n N_VGND_c_1016_n 0.00685342f $X=4.29 $Y=0.96 $X2=0
+ $Y2=0
cc_355 N_A_301_47#_c_388_n N_VGND_c_1016_n 0.00699289f $X=4.71 $Y=0.96 $X2=0
+ $Y2=0
cc_356 N_A_301_47#_c_390_n N_VGND_c_1016_n 6.07018e-19 $X=5.13 $Y=0.96 $X2=0
+ $Y2=0
cc_357 N_A_301_47#_c_388_n N_VGND_c_1017_n 6.07018e-19 $X=4.71 $Y=0.96 $X2=0
+ $Y2=0
cc_358 N_A_301_47#_c_390_n N_VGND_c_1017_n 0.00699289f $X=5.13 $Y=0.96 $X2=0
+ $Y2=0
cc_359 N_A_301_47#_c_392_n N_VGND_c_1017_n 0.00818769f $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_360 N_A_301_47#_c_377_n N_VGND_c_1018_n 0.00341689f $X=2.61 $Y=0.96 $X2=0
+ $Y2=0
cc_361 N_A_301_47#_c_401_n N_VGND_c_1018_n 0.0339167f $X=1.64 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_301_47#_c_380_n N_VGND_c_1020_n 0.00341689f $X=3.03 $Y=0.96 $X2=0
+ $Y2=0
cc_363 N_A_301_47#_c_382_n N_VGND_c_1020_n 0.00341689f $X=3.45 $Y=0.96 $X2=0
+ $Y2=0
cc_364 N_A_301_47#_c_388_n N_VGND_c_1023_n 0.00341689f $X=4.71 $Y=0.96 $X2=0
+ $Y2=0
cc_365 N_A_301_47#_c_390_n N_VGND_c_1023_n 0.00341689f $X=5.13 $Y=0.96 $X2=0
+ $Y2=0
cc_366 N_A_301_47#_c_392_n N_VGND_c_1024_n 0.00341689f $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_367 N_A_301_47#_M1031_d N_VGND_c_1025_n 0.00210122f $X=1.505 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_301_47#_c_377_n N_VGND_c_1025_n 0.00540327f $X=2.61 $Y=0.96 $X2=0
+ $Y2=0
cc_369 N_A_301_47#_c_380_n N_VGND_c_1025_n 0.0040262f $X=3.03 $Y=0.96 $X2=0
+ $Y2=0
cc_370 N_A_301_47#_c_382_n N_VGND_c_1025_n 0.0040262f $X=3.45 $Y=0.96 $X2=0
+ $Y2=0
cc_371 N_A_301_47#_c_384_n N_VGND_c_1025_n 0.0040262f $X=3.87 $Y=0.96 $X2=0
+ $Y2=0
cc_372 N_A_301_47#_c_386_n N_VGND_c_1025_n 0.0040262f $X=4.29 $Y=0.96 $X2=0
+ $Y2=0
cc_373 N_A_301_47#_c_388_n N_VGND_c_1025_n 0.0040262f $X=4.71 $Y=0.96 $X2=0
+ $Y2=0
cc_374 N_A_301_47#_c_390_n N_VGND_c_1025_n 0.0040262f $X=5.13 $Y=0.96 $X2=0
+ $Y2=0
cc_375 N_A_301_47#_c_392_n N_VGND_c_1025_n 0.00458661f $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_376 N_A_301_47#_c_401_n N_VGND_c_1025_n 0.0194095f $X=1.64 $Y=0.56 $X2=0
+ $Y2=0
cc_377 N_A_301_47#_c_401_n N_A_455_47#_c_1144_n 0.0343984f $X=1.64 $Y=0.56 $X2=0
+ $Y2=0
cc_378 N_A_301_47#_c_377_n N_A_455_47#_c_1150_n 0.0122782f $X=2.61 $Y=0.96 $X2=0
+ $Y2=0
cc_379 N_A_301_47#_c_378_n N_A_455_47#_c_1150_n 0.00186586f $X=2.955 $Y=1.035
+ $X2=0 $Y2=0
cc_380 N_A_301_47#_c_380_n N_A_455_47#_c_1150_n 0.0113204f $X=3.03 $Y=0.96 $X2=0
+ $Y2=0
cc_381 N_A_301_47#_c_400_n N_A_455_47#_c_1150_n 0.0379559f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_382 N_A_301_47#_c_400_n N_A_455_47#_c_1145_n 0.0254999f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_A_301_47#_c_401_n N_A_455_47#_c_1145_n 0.0181622f $X=1.64 $Y=0.56 $X2=0
+ $Y2=0
cc_384 N_A_301_47#_c_382_n N_A_455_47#_c_1156_n 0.0113204f $X=3.45 $Y=0.96 $X2=0
+ $Y2=0
cc_385 N_A_301_47#_c_383_n N_A_455_47#_c_1156_n 0.00186586f $X=3.795 $Y=1.035
+ $X2=0 $Y2=0
cc_386 N_A_301_47#_c_384_n N_A_455_47#_c_1156_n 0.0113204f $X=3.87 $Y=0.96 $X2=0
+ $Y2=0
cc_387 N_A_301_47#_c_400_n N_A_455_47#_c_1156_n 0.0377219f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_388 N_A_301_47#_c_386_n N_A_455_47#_c_1160_n 0.0113204f $X=4.29 $Y=0.96 $X2=0
+ $Y2=0
cc_389 N_A_301_47#_c_387_n N_A_455_47#_c_1160_n 0.00186586f $X=4.635 $Y=1.035
+ $X2=0 $Y2=0
cc_390 N_A_301_47#_c_388_n N_A_455_47#_c_1160_n 0.0113204f $X=4.71 $Y=0.96 $X2=0
+ $Y2=0
cc_391 N_A_301_47#_c_400_n N_A_455_47#_c_1160_n 0.0377219f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_A_301_47#_c_390_n N_A_455_47#_c_1164_n 0.0112683f $X=5.13 $Y=0.96 $X2=0
+ $Y2=0
cc_393 N_A_301_47#_c_391_n N_A_455_47#_c_1164_n 0.00186586f $X=5.475 $Y=1.035
+ $X2=0 $Y2=0
cc_394 N_A_301_47#_c_392_n N_A_455_47#_c_1164_n 0.0121329f $X=5.55 $Y=0.96 $X2=0
+ $Y2=0
cc_395 N_A_301_47#_c_400_n N_A_455_47#_c_1164_n 0.0377578f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_396 N_A_301_47#_c_381_n N_A_455_47#_c_1168_n 0.00193161f $X=3.375 $Y=1.035
+ $X2=0 $Y2=0
cc_397 N_A_301_47#_c_400_n N_A_455_47#_c_1168_n 0.0119538f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_398 N_A_301_47#_c_385_n N_A_455_47#_c_1170_n 0.00193392f $X=4.215 $Y=1.035
+ $X2=0 $Y2=0
cc_399 N_A_301_47#_c_400_n N_A_455_47#_c_1170_n 0.0119831f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_400 N_A_301_47#_c_389_n N_A_455_47#_c_1172_n 0.00193161f $X=5.055 $Y=1.035
+ $X2=0 $Y2=0
cc_401 N_A_301_47#_c_400_n N_A_455_47#_c_1172_n 0.0119538f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_402 N_A_301_47#_c_392_n N_A_455_47#_c_1174_n 0.00623981f $X=5.55 $Y=0.96
+ $X2=0 $Y2=0
cc_403 N_A_301_47#_c_400_n N_A_455_47#_c_1174_n 0.0180946f $X=5.76 $Y=1.16 $X2=0
+ $Y2=0
cc_404 N_A_116_47#_c_541_n N_VPWR_c_677_n 0.00123564f $X=6.52 $Y=1.19 $X2=0
+ $Y2=0
cc_405 N_A_116_47#_c_583_p N_VPWR_c_686_n 0.011928f $X=0.715 $Y=2.22 $X2=0 $Y2=0
cc_406 N_A_116_47#_M1003_g N_VPWR_c_689_n 0.00357877f $X=6.23 $Y=1.985 $X2=0
+ $Y2=0
cc_407 N_A_116_47#_M1009_g N_VPWR_c_689_n 0.00357877f $X=6.65 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_116_47#_M1013_g N_VPWR_c_689_n 0.00357877f $X=7.07 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_116_47#_M1018_g N_VPWR_c_689_n 0.00357877f $X=7.49 $Y=1.985 $X2=0
+ $Y2=0
cc_410 N_A_116_47#_M1023_g N_VPWR_c_689_n 0.00357877f $X=7.91 $Y=1.985 $X2=0
+ $Y2=0
cc_411 N_A_116_47#_M1024_g N_VPWR_c_689_n 0.00357877f $X=8.33 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A_116_47#_M1030_g N_VPWR_c_689_n 0.00357877f $X=8.75 $Y=1.985 $X2=0
+ $Y2=0
cc_413 N_A_116_47#_M1035_g N_VPWR_c_689_n 0.00357877f $X=9.17 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A_116_47#_M1019_s N_VPWR_c_674_n 0.00518834f $X=0.58 $Y=1.485 $X2=0
+ $Y2=0
cc_415 N_A_116_47#_M1003_g N_VPWR_c_674_n 0.00664112f $X=6.23 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A_116_47#_M1009_g N_VPWR_c_674_n 0.00522516f $X=6.65 $Y=1.985 $X2=0
+ $Y2=0
cc_417 N_A_116_47#_M1013_g N_VPWR_c_674_n 0.00522516f $X=7.07 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_A_116_47#_M1018_g N_VPWR_c_674_n 0.00522516f $X=7.49 $Y=1.985 $X2=0
+ $Y2=0
cc_419 N_A_116_47#_M1023_g N_VPWR_c_674_n 0.00522516f $X=7.91 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A_116_47#_M1024_g N_VPWR_c_674_n 0.00522516f $X=8.33 $Y=1.985 $X2=0
+ $Y2=0
cc_421 N_A_116_47#_M1030_g N_VPWR_c_674_n 0.00522516f $X=8.75 $Y=1.985 $X2=0
+ $Y2=0
cc_422 N_A_116_47#_M1035_g N_VPWR_c_674_n 0.00619805f $X=9.17 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A_116_47#_c_583_p N_VPWR_c_674_n 0.00704765f $X=0.715 $Y=2.22 $X2=0
+ $Y2=0
cc_424 N_A_116_47#_M1003_g N_A_407_309#_c_813_n 0.031735f $X=6.23 $Y=1.985 $X2=0
+ $Y2=0
cc_425 N_A_116_47#_M1009_g N_A_407_309#_c_813_n 0.017969f $X=6.65 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A_116_47#_M1013_g N_A_407_309#_c_813_n 0.0179753f $X=7.07 $Y=1.985
+ $X2=0 $Y2=0
cc_427 N_A_116_47#_M1018_g N_A_407_309#_c_813_n 0.0179753f $X=7.49 $Y=1.985
+ $X2=0 $Y2=0
cc_428 N_A_116_47#_M1023_g N_A_407_309#_c_813_n 0.0179753f $X=7.91 $Y=1.985
+ $X2=0 $Y2=0
cc_429 N_A_116_47#_M1024_g N_A_407_309#_c_813_n 0.0179753f $X=8.33 $Y=1.985
+ $X2=0 $Y2=0
cc_430 N_A_116_47#_M1030_g N_A_407_309#_c_813_n 0.0179753f $X=8.75 $Y=1.985
+ $X2=0 $Y2=0
cc_431 N_A_116_47#_M1035_g N_A_407_309#_c_813_n 0.0179753f $X=9.17 $Y=1.985
+ $X2=0 $Y2=0
cc_432 N_A_116_47#_M1001_g N_Z_c_936_n 0.00336436f $X=6.23 $Y=0.56 $X2=0 $Y2=0
cc_433 N_A_116_47#_M1006_g N_Z_c_936_n 0.010143f $X=6.65 $Y=0.56 $X2=0 $Y2=0
cc_434 N_A_116_47#_M1026_g N_Z_c_936_n 0.0102073f $X=7.07 $Y=0.56 $X2=0 $Y2=0
cc_435 N_A_116_47#_M1027_g N_Z_c_936_n 0.0102073f $X=7.49 $Y=0.56 $X2=0 $Y2=0
cc_436 N_A_116_47#_M1029_g N_Z_c_936_n 0.0102073f $X=7.91 $Y=0.56 $X2=0 $Y2=0
cc_437 N_A_116_47#_M1032_g N_Z_c_936_n 0.0102073f $X=8.33 $Y=0.56 $X2=0 $Y2=0
cc_438 N_A_116_47#_M1033_g N_Z_c_936_n 0.0102073f $X=8.75 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A_116_47#_M1034_g N_Z_c_936_n 0.0134794f $X=9.17 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A_116_47#_c_541_n N_Z_c_936_n 0.00151378f $X=6.52 $Y=1.19 $X2=0 $Y2=0
cc_441 N_A_116_47#_c_542_n N_Z_c_936_n 0.00191164f $X=6.665 $Y=1.19 $X2=0 $Y2=0
cc_442 N_A_116_47#_c_579_n N_Z_c_936_n 0.178269f $X=8.74 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_116_47#_c_543_n N_Z_c_936_n 0.0136691f $X=9.17 $Y=1.16 $X2=0 $Y2=0
cc_444 N_A_116_47#_M1034_g Z 0.0209399f $X=9.17 $Y=0.56 $X2=0 $Y2=0
cc_445 N_A_116_47#_c_579_n Z 0.0203821f $X=8.74 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_116_47#_M1003_g N_Z_c_906_n 0.0152137f $X=6.23 $Y=1.985 $X2=0 $Y2=0
cc_447 N_A_116_47#_M1009_g N_Z_c_906_n 0.0116539f $X=6.65 $Y=1.985 $X2=0 $Y2=0
cc_448 N_A_116_47#_M1013_g N_Z_c_906_n 0.0117437f $X=7.07 $Y=1.985 $X2=0 $Y2=0
cc_449 N_A_116_47#_M1018_g N_Z_c_906_n 0.0117437f $X=7.49 $Y=1.985 $X2=0 $Y2=0
cc_450 N_A_116_47#_M1023_g N_Z_c_906_n 0.0117437f $X=7.91 $Y=1.985 $X2=0 $Y2=0
cc_451 N_A_116_47#_M1024_g N_Z_c_906_n 0.0117437f $X=8.33 $Y=1.985 $X2=0 $Y2=0
cc_452 N_A_116_47#_M1030_g N_Z_c_906_n 0.0117437f $X=8.75 $Y=1.985 $X2=0 $Y2=0
cc_453 N_A_116_47#_M1035_g N_Z_c_906_n 0.0153674f $X=9.17 $Y=1.985 $X2=0 $Y2=0
cc_454 N_A_116_47#_c_541_n N_Z_c_906_n 0.0403215f $X=6.52 $Y=1.19 $X2=0 $Y2=0
cc_455 N_A_116_47#_c_542_n N_Z_c_906_n 0.0076828f $X=6.665 $Y=1.19 $X2=0 $Y2=0
cc_456 N_A_116_47#_c_579_n N_Z_c_906_n 0.218089f $X=8.74 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_116_47#_c_543_n N_Z_c_906_n 0.0140528f $X=9.17 $Y=1.16 $X2=0 $Y2=0
cc_458 N_A_116_47#_M1001_g N_VGND_c_1017_n 8.09705e-19 $X=6.23 $Y=0.56 $X2=0
+ $Y2=0
cc_459 N_A_116_47#_c_539_n N_VGND_c_1022_n 0.0102853f $X=0.715 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_116_47#_M1001_g N_VGND_c_1024_n 0.00357877f $X=6.23 $Y=0.56 $X2=0
+ $Y2=0
cc_461 N_A_116_47#_M1006_g N_VGND_c_1024_n 0.00357877f $X=6.65 $Y=0.56 $X2=0
+ $Y2=0
cc_462 N_A_116_47#_M1026_g N_VGND_c_1024_n 0.00357877f $X=7.07 $Y=0.56 $X2=0
+ $Y2=0
cc_463 N_A_116_47#_M1027_g N_VGND_c_1024_n 0.00357877f $X=7.49 $Y=0.56 $X2=0
+ $Y2=0
cc_464 N_A_116_47#_M1029_g N_VGND_c_1024_n 0.00357877f $X=7.91 $Y=0.56 $X2=0
+ $Y2=0
cc_465 N_A_116_47#_M1032_g N_VGND_c_1024_n 0.00357877f $X=8.33 $Y=0.56 $X2=0
+ $Y2=0
cc_466 N_A_116_47#_M1033_g N_VGND_c_1024_n 0.00357877f $X=8.75 $Y=0.56 $X2=0
+ $Y2=0
cc_467 N_A_116_47#_M1034_g N_VGND_c_1024_n 0.00357877f $X=9.17 $Y=0.56 $X2=0
+ $Y2=0
cc_468 N_A_116_47#_M1004_s N_VGND_c_1025_n 0.00519615f $X=0.58 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_A_116_47#_M1001_g N_VGND_c_1025_n 0.00582446f $X=6.23 $Y=0.56 $X2=0
+ $Y2=0
cc_470 N_A_116_47#_M1006_g N_VGND_c_1025_n 0.00522516f $X=6.65 $Y=0.56 $X2=0
+ $Y2=0
cc_471 N_A_116_47#_M1026_g N_VGND_c_1025_n 0.00522516f $X=7.07 $Y=0.56 $X2=0
+ $Y2=0
cc_472 N_A_116_47#_M1027_g N_VGND_c_1025_n 0.00522516f $X=7.49 $Y=0.56 $X2=0
+ $Y2=0
cc_473 N_A_116_47#_M1029_g N_VGND_c_1025_n 0.00522516f $X=7.91 $Y=0.56 $X2=0
+ $Y2=0
cc_474 N_A_116_47#_M1032_g N_VGND_c_1025_n 0.00522516f $X=8.33 $Y=0.56 $X2=0
+ $Y2=0
cc_475 N_A_116_47#_M1033_g N_VGND_c_1025_n 0.00522516f $X=8.75 $Y=0.56 $X2=0
+ $Y2=0
cc_476 N_A_116_47#_M1034_g N_VGND_c_1025_n 0.00619805f $X=9.17 $Y=0.56 $X2=0
+ $Y2=0
cc_477 N_A_116_47#_c_539_n N_VGND_c_1025_n 0.0069624f $X=0.715 $Y=0.445 $X2=0
+ $Y2=0
cc_478 N_A_116_47#_c_541_n N_A_455_47#_c_1150_n 0.00400213f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_479 N_A_116_47#_c_541_n N_A_455_47#_c_1145_n 0.00223802f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_480 N_A_116_47#_c_541_n N_A_455_47#_c_1156_n 0.00400213f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_481 N_A_116_47#_c_541_n N_A_455_47#_c_1160_n 0.00400213f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_482 N_A_116_47#_c_541_n N_A_455_47#_c_1164_n 0.00400213f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_483 N_A_116_47#_M1001_g N_A_455_47#_c_1146_n 0.0118535f $X=6.23 $Y=0.56 $X2=0
+ $Y2=0
cc_484 N_A_116_47#_M1006_g N_A_455_47#_c_1146_n 0.00809662f $X=6.65 $Y=0.56
+ $X2=0 $Y2=0
cc_485 N_A_116_47#_M1026_g N_A_455_47#_c_1146_n 0.00814603f $X=7.07 $Y=0.56
+ $X2=0 $Y2=0
cc_486 N_A_116_47#_M1027_g N_A_455_47#_c_1146_n 0.00814603f $X=7.49 $Y=0.56
+ $X2=0 $Y2=0
cc_487 N_A_116_47#_M1029_g N_A_455_47#_c_1146_n 0.00814603f $X=7.91 $Y=0.56
+ $X2=0 $Y2=0
cc_488 N_A_116_47#_M1032_g N_A_455_47#_c_1146_n 0.00814603f $X=8.33 $Y=0.56
+ $X2=0 $Y2=0
cc_489 N_A_116_47#_M1033_g N_A_455_47#_c_1146_n 0.00814603f $X=8.75 $Y=0.56
+ $X2=0 $Y2=0
cc_490 N_A_116_47#_M1034_g N_A_455_47#_c_1146_n 0.00814603f $X=9.17 $Y=0.56
+ $X2=0 $Y2=0
cc_491 N_A_116_47#_c_579_n N_A_455_47#_c_1146_n 0.0025603f $X=8.74 $Y=1.16 $X2=0
+ $Y2=0
cc_492 N_A_116_47#_c_541_n N_A_455_47#_c_1168_n 0.00114955f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_493 N_A_116_47#_c_541_n N_A_455_47#_c_1170_n 0.001153f $X=6.52 $Y=1.19 $X2=0
+ $Y2=0
cc_494 N_A_116_47#_c_541_n N_A_455_47#_c_1172_n 0.00114955f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_495 N_A_116_47#_c_541_n N_A_455_47#_c_1174_n 0.00699828f $X=6.52 $Y=1.19
+ $X2=0 $Y2=0
cc_496 N_VPWR_c_674_n N_A_407_309#_M1002_d 0.00227813f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_497 N_VPWR_c_674_n N_A_407_309#_M1008_d 0.00252188f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_674_n N_A_407_309#_M1016_d 0.00252188f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_674_n N_A_407_309#_M1022_d 0.00252188f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_674_n N_A_407_309#_M1037_d 0.00644954f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_674_n N_A_407_309#_M1009_d 0.00215227f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_674_n N_A_407_309#_M1018_d 0.00215227f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_674_n N_A_407_309#_M1024_d 0.00215227f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_674_n N_A_407_309#_M1035_d 0.00225742f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_687_n N_A_407_309#_c_811_n 0.0170644f $X=2.415 $Y=2.72 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_674_n N_A_407_309#_c_811_n 0.00950719f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_507 N_VPWR_M1002_s N_A_407_309#_c_814_n 0.0031354f $X=2.445 $Y=1.545 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_678_n N_A_407_309#_c_814_n 0.0160613f $X=2.58 $Y=2.36 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_687_n N_A_407_309#_c_814_n 0.0023303f $X=2.415 $Y=2.72 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_688_n N_A_407_309#_c_814_n 0.0023303f $X=3.255 $Y=2.72 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_674_n N_A_407_309#_c_814_n 0.00964389f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_688_n N_A_407_309#_c_856_n 0.0112554f $X=3.255 $Y=2.72 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_674_n N_A_407_309#_c_856_n 0.00644035f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_514 N_VPWR_M1011_s N_A_407_309#_c_818_n 0.0031354f $X=3.285 $Y=1.545 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_679_n N_A_407_309#_c_818_n 0.0160613f $X=3.42 $Y=2.36 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_682_n N_A_407_309#_c_818_n 0.0023303f $X=4.095 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_688_n N_A_407_309#_c_818_n 0.0023303f $X=3.255 $Y=2.72 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_674_n N_A_407_309#_c_818_n 0.00964389f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_682_n N_A_407_309#_c_863_n 0.0112554f $X=4.095 $Y=2.72 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_674_n N_A_407_309#_c_863_n 0.00644035f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_M1017_s N_A_407_309#_c_821_n 0.0031354f $X=4.125 $Y=1.545 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_680_n N_A_407_309#_c_821_n 0.0160613f $X=4.26 $Y=2.36 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_682_n N_A_407_309#_c_821_n 0.0023303f $X=4.095 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_684_n N_A_407_309#_c_821_n 0.0023303f $X=4.935 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_674_n N_A_407_309#_c_821_n 0.00964389f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_684_n N_A_407_309#_c_870_n 0.0112554f $X=4.935 $Y=2.72 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_674_n N_A_407_309#_c_870_n 0.00644035f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_689_n N_A_407_309#_c_872_n 0.251792f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_529 N_VPWR_c_674_n N_A_407_309#_c_872_n 0.152614f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_530 N_VPWR_M1028_s N_A_407_309#_c_827_n 0.0031354f $X=4.965 $Y=1.545 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_681_n N_A_407_309#_c_827_n 0.0160613f $X=5.1 $Y=2.36 $X2=0 $Y2=0
cc_532 N_VPWR_c_684_n N_A_407_309#_c_827_n 0.0023303f $X=4.935 $Y=2.72 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_689_n N_A_407_309#_c_827_n 0.0023303f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_674_n N_A_407_309#_c_827_n 0.00968468f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_674_n N_Z_M1003_s 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_536 N_VPWR_c_674_n N_Z_M1013_s 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_537 N_VPWR_c_674_n N_Z_M1023_s 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_538 N_VPWR_c_674_n N_Z_M1030_s 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_M1002_s N_Z_c_906_n 0.0016881f $X=2.445 $Y=1.545 $X2=0 $Y2=0
cc_540 N_VPWR_M1011_s N_Z_c_906_n 0.0016881f $X=3.285 $Y=1.545 $X2=0 $Y2=0
cc_541 N_VPWR_M1017_s N_Z_c_906_n 0.0016881f $X=4.125 $Y=1.545 $X2=0 $Y2=0
cc_542 N_VPWR_M1028_s N_Z_c_906_n 0.0016881f $X=4.965 $Y=1.545 $X2=0 $Y2=0
cc_543 N_A_407_309#_c_813_n N_Z_M1003_s 0.00316076f $X=9.38 $Y=2.02 $X2=0 $Y2=0
cc_544 N_A_407_309#_c_813_n N_Z_M1013_s 0.00316076f $X=9.38 $Y=2.02 $X2=0 $Y2=0
cc_545 N_A_407_309#_c_813_n N_Z_M1023_s 0.00316076f $X=9.38 $Y=2.02 $X2=0 $Y2=0
cc_546 N_A_407_309#_c_813_n N_Z_M1030_s 0.00316076f $X=9.38 $Y=2.02 $X2=0 $Y2=0
cc_547 N_A_407_309#_M1035_d Z 0.0035471f $X=9.245 $Y=1.485 $X2=0 $Y2=0
cc_548 N_A_407_309#_c_813_n Z 0.0222273f $X=9.38 $Y=2.02 $X2=0 $Y2=0
cc_549 N_A_407_309#_M1002_d N_Z_c_906_n 0.00251902f $X=2.035 $Y=1.545 $X2=0
+ $Y2=0
cc_550 N_A_407_309#_M1008_d N_Z_c_906_n 0.00168399f $X=2.865 $Y=1.545 $X2=0
+ $Y2=0
cc_551 N_A_407_309#_M1016_d N_Z_c_906_n 0.00168399f $X=3.705 $Y=1.545 $X2=0
+ $Y2=0
cc_552 N_A_407_309#_M1022_d N_Z_c_906_n 0.00168399f $X=4.545 $Y=1.545 $X2=0
+ $Y2=0
cc_553 N_A_407_309#_M1037_d N_Z_c_906_n 0.0125225f $X=5.385 $Y=1.545 $X2=0 $Y2=0
cc_554 N_A_407_309#_M1009_d N_Z_c_906_n 0.0016881f $X=6.725 $Y=1.485 $X2=0 $Y2=0
cc_555 N_A_407_309#_M1018_d N_Z_c_906_n 0.0016881f $X=7.565 $Y=1.485 $X2=0 $Y2=0
cc_556 N_A_407_309#_M1024_d N_Z_c_906_n 0.0016881f $X=8.405 $Y=1.485 $X2=0 $Y2=0
cc_557 N_A_407_309#_M1035_d N_Z_c_906_n 2.38066e-19 $X=9.245 $Y=1.485 $X2=0
+ $Y2=0
cc_558 N_A_407_309#_c_814_n N_Z_c_906_n 0.0329142f $X=2.915 $Y=1.98 $X2=0 $Y2=0
cc_559 N_A_407_309#_c_812_n N_Z_c_906_n 0.0203044f $X=2.245 $Y=1.98 $X2=0 $Y2=0
cc_560 N_A_407_309#_c_818_n N_Z_c_906_n 0.0329142f $X=3.755 $Y=1.98 $X2=0 $Y2=0
cc_561 N_A_407_309#_c_821_n N_Z_c_906_n 0.0329142f $X=4.595 $Y=1.98 $X2=0 $Y2=0
cc_562 N_A_407_309#_c_824_n N_Z_c_906_n 0.0129524f $X=3 $Y=1.98 $X2=0 $Y2=0
cc_563 N_A_407_309#_c_825_n N_Z_c_906_n 0.0129524f $X=3.84 $Y=1.98 $X2=0 $Y2=0
cc_564 N_A_407_309#_c_826_n N_Z_c_906_n 0.0129524f $X=4.68 $Y=1.98 $X2=0 $Y2=0
cc_565 N_A_407_309#_c_827_n N_Z_c_906_n 0.2711f $X=5.435 $Y=2.18 $X2=0 $Y2=0
cc_566 N_Z_M1001_d N_VGND_c_1025_n 0.00216833f $X=6.305 $Y=0.235 $X2=0 $Y2=0
cc_567 N_Z_M1026_d N_VGND_c_1025_n 0.00216833f $X=7.145 $Y=0.235 $X2=0 $Y2=0
cc_568 N_Z_M1029_d N_VGND_c_1025_n 0.00216833f $X=7.985 $Y=0.235 $X2=0 $Y2=0
cc_569 N_Z_M1033_d N_VGND_c_1025_n 0.00216833f $X=8.825 $Y=0.235 $X2=0 $Y2=0
cc_570 N_Z_c_936_n N_A_455_47#_M1006_s 0.0030582f $X=9.325 $Y=0.735 $X2=0 $Y2=0
cc_571 N_Z_c_936_n N_A_455_47#_M1027_s 0.00308199f $X=9.325 $Y=0.735 $X2=0 $Y2=0
cc_572 N_Z_c_936_n N_A_455_47#_M1032_s 0.00308199f $X=9.325 $Y=0.735 $X2=0 $Y2=0
cc_573 N_Z_c_936_n N_A_455_47#_M1034_s 6.34286e-19 $X=9.325 $Y=0.735 $X2=0 $Y2=0
cc_574 Z N_A_455_47#_M1034_s 4.96845e-19 $X=9.34 $Y=0.765 $X2=0 $Y2=0
cc_575 N_Z_c_903_n N_A_455_47#_M1034_s 0.00345418f $X=9.45 $Y=0.855 $X2=0 $Y2=0
cc_576 N_Z_M1001_d N_A_455_47#_c_1146_n 0.00305132f $X=6.305 $Y=0.235 $X2=0
+ $Y2=0
cc_577 N_Z_M1026_d N_A_455_47#_c_1146_n 0.00305132f $X=7.145 $Y=0.235 $X2=0
+ $Y2=0
cc_578 N_Z_M1029_d N_A_455_47#_c_1146_n 0.00305132f $X=7.985 $Y=0.235 $X2=0
+ $Y2=0
cc_579 N_Z_M1033_d N_A_455_47#_c_1146_n 0.00305132f $X=8.825 $Y=0.235 $X2=0
+ $Y2=0
cc_580 N_Z_c_936_n N_A_455_47#_c_1146_n 0.150263f $X=9.325 $Y=0.735 $X2=0 $Y2=0
cc_581 N_Z_c_903_n N_A_455_47#_c_1146_n 0.0194298f $X=9.45 $Y=0.855 $X2=0 $Y2=0
cc_582 N_Z_c_906_n N_A_455_47#_c_1174_n 0.00246104f $X=9.325 $Y=1.585 $X2=0
+ $Y2=0
cc_583 N_VGND_c_1025_n N_A_455_47#_M1000_d 0.00229009f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_584 N_VGND_c_1025_n N_A_455_47#_M1005_d 0.00255104f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_1025_n N_A_455_47#_M1010_d 0.00254582f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_1025_n N_A_455_47#_M1014_d 0.00255104f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_1025_n N_A_455_47#_M1021_d 0.00446531f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_1025_n N_A_455_47#_M1006_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_1025_n N_A_455_47#_M1027_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_1025_n N_A_455_47#_M1032_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_1025_n N_A_455_47#_M1034_s 0.00225742f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_1018_n N_A_455_47#_c_1144_n 0.0228093f $X=2.655 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_1025_n N_A_455_47#_c_1144_n 0.0125906f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_M1000_s N_A_455_47#_c_1150_n 0.00288179f $X=2.685 $Y=0.235 $X2=0
+ $Y2=0
cc_595 N_VGND_c_1013_n N_A_455_47#_c_1150_n 0.0162338f $X=2.82 $Y=0.36 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1018_n N_A_455_47#_c_1150_n 0.00234306f $X=2.655 $Y=0 $X2=0
+ $Y2=0
cc_597 N_VGND_c_1020_n N_A_455_47#_c_1150_n 0.00234306f $X=3.495 $Y=0 $X2=0
+ $Y2=0
cc_598 N_VGND_c_1025_n N_A_455_47#_c_1150_n 0.00978207f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_599 N_VGND_c_1020_n N_A_455_47#_c_1223_n 0.00998989f $X=3.495 $Y=0 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1025_n N_A_455_47#_c_1223_n 0.00637943f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_M1007_s N_A_455_47#_c_1156_n 0.00288179f $X=3.525 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_VGND_c_1014_n N_A_455_47#_c_1156_n 0.0162338f $X=3.66 $Y=0.36 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1015_n N_A_455_47#_c_1156_n 0.00234306f $X=4.335 $Y=0 $X2=0
+ $Y2=0
cc_604 N_VGND_c_1020_n N_A_455_47#_c_1156_n 0.00234306f $X=3.495 $Y=0 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1025_n N_A_455_47#_c_1156_n 0.00978207f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_c_1015_n N_A_455_47#_c_1230_n 0.0112958f $X=4.335 $Y=0 $X2=0 $Y2=0
cc_607 N_VGND_c_1025_n N_A_455_47#_c_1230_n 0.00644886f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_M1012_s N_A_455_47#_c_1160_n 0.00288179f $X=4.365 $Y=0.235 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1015_n N_A_455_47#_c_1160_n 0.00234306f $X=4.335 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1016_n N_A_455_47#_c_1160_n 0.0162338f $X=4.5 $Y=0.36 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1023_n N_A_455_47#_c_1160_n 0.00234306f $X=5.175 $Y=0 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1025_n N_A_455_47#_c_1160_n 0.00978207f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1023_n N_A_455_47#_c_1237_n 0.00998989f $X=5.175 $Y=0 $X2=0
+ $Y2=0
cc_614 N_VGND_c_1025_n N_A_455_47#_c_1237_n 0.00637943f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_M1015_s N_A_455_47#_c_1164_n 0.00292181f $X=5.205 $Y=0.235 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1017_n N_A_455_47#_c_1164_n 0.0162338f $X=5.34 $Y=0.36 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1023_n N_A_455_47#_c_1164_n 0.00234306f $X=5.175 $Y=0 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1024_n N_A_455_47#_c_1164_n 0.00234956f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1025_n N_A_455_47#_c_1164_n 0.00979243f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_620 N_VGND_c_1024_n N_A_455_47#_c_1146_n 0.193324f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_c_1025_n N_A_455_47#_c_1146_n 0.123597f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_c_1024_n N_A_455_47#_c_1174_n 0.0294126f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_c_1025_n N_A_455_47#_c_1174_n 0.0164292f $X=9.43 $Y=0 $X2=0 $Y2=0

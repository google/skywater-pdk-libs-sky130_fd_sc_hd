* File: sky130_fd_sc_hd__lpflow_isobufsrc_16.spice.pex
* Created: Thu Aug 27 14:25:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A 5 7 9 12 14 16 19 21 23 26 28
+ 30 33 36 37 45
r79 44 45 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.9 $Y=1.16 $X2=2.12
+ $Y2=1.16
r80 43 44 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.7 $Y=1.16 $X2=1.9
+ $Y2=1.16
r81 42 43 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.48 $Y=1.16 $X2=1.7
+ $Y2=1.16
r82 41 42 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.28 $Y=1.16 $X2=1.48
+ $Y2=1.16
r83 40 41 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.06 $Y=1.16
+ $X2=1.28 $Y2=1.16
r84 39 40 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.86 $Y=1.16 $X2=1.06
+ $Y2=1.16
r85 38 39 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.64 $Y=1.16
+ $X2=0.86 $Y2=1.16
r86 36 38 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.58 $Y=1.16 $X2=0.64
+ $Y2=1.16
r87 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r88 33 37 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.38 $Y=1.16 $X2=0.58
+ $Y2=1.16
r89 28 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.12 $Y=0.995
+ $X2=2.12 $Y2=1.16
r90 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.12 $Y=0.995
+ $X2=2.12 $Y2=0.56
r91 24 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=1.325
+ $X2=1.9 $Y2=1.16
r92 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.9 $Y=1.325 $X2=1.9
+ $Y2=1.985
r93 21 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=0.995
+ $X2=1.7 $Y2=1.16
r94 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.7 $Y=0.995 $X2=1.7
+ $Y2=0.56
r95 17 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=1.325
+ $X2=1.48 $Y2=1.16
r96 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.48 $Y=1.325
+ $X2=1.48 $Y2=1.985
r97 14 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.28 $Y=0.995
+ $X2=1.28 $Y2=1.16
r98 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.28 $Y=0.995
+ $X2=1.28 $Y2=0.56
r99 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.325
+ $X2=1.06 $Y2=1.16
r100 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.06 $Y=1.325
+ $X2=1.06 $Y2=1.985
r101 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.86 $Y=0.995
+ $X2=0.86 $Y2=1.16
r102 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.86 $Y=0.995
+ $X2=0.86 $Y2=0.56
r103 3 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.325
+ $X2=0.64 $Y2=1.16
r104 3 5 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.64 $Y=1.325
+ $X2=0.64 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A_143_297# 1 2 3 4 13 15 18 20
+ 22 25 27 29 32 34 36 39 41 43 46 48 50 53 55 57 60 62 64 67 69 71 74 76 78 81
+ 83 85 88 90 92 95 97 99 102 104 106 109 111 113 116 118 120 123 127 133 135
+ 136 139 145 152 156 157 161 180
r336 177 178 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.34 $Y=1.16
+ $X2=8.76 $Y2=1.16
r337 176 177 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7.92 $Y=1.16
+ $X2=8.34 $Y2=1.16
r338 175 176 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7.5 $Y=1.16
+ $X2=7.92 $Y2=1.16
r339 174 175 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7.08 $Y=1.16
+ $X2=7.5 $Y2=1.16
r340 173 174 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.66 $Y=1.16
+ $X2=7.08 $Y2=1.16
r341 172 173 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=6.66 $Y2=1.16
r342 171 172 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.82 $Y=1.16
+ $X2=6.24 $Y2=1.16
r343 170 171 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.4 $Y=1.16
+ $X2=5.82 $Y2=1.16
r344 169 170 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.98 $Y=1.16
+ $X2=5.4 $Y2=1.16
r345 168 169 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.98 $Y2=1.16
r346 167 168 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.14 $Y=1.16
+ $X2=4.56 $Y2=1.16
r347 166 167 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.72 $Y=1.16
+ $X2=4.14 $Y2=1.16
r348 165 166 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.3 $Y=1.16
+ $X2=3.72 $Y2=1.16
r349 158 160 8.64332 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=1.175
+ $X2=1.09 $Y2=1.175
r350 156 157 6.72958 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.85 $Y=1.62
+ $X2=0.85 $Y2=1.495
r351 153 180 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.09 $Y=1.16
+ $X2=9.18 $Y2=1.16
r352 153 178 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=9.09 $Y=1.16
+ $X2=8.76 $Y2=1.16
r353 152 153 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=9.09
+ $Y=1.16 $X2=9.09 $Y2=1.16
r354 150 165 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.97 $Y=1.16
+ $X2=3.3 $Y2=1.16
r355 150 162 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.97 $Y=1.16
+ $X2=2.88 $Y2=1.16
r356 149 152 323.221 $w=2.08e-07 $l=6.12e-06 $layer=LI1_cond $X=2.97 $Y=1.18
+ $X2=9.09 $Y2=1.18
r357 149 150 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=2.97
+ $Y=1.16 $X2=2.97 $Y2=1.16
r358 147 161 4.00838 $w=2.1e-07 $l=2.57488e-07 $layer=LI1_cond $X=2.035 $Y=1.18
+ $X2=1.78 $Y2=1.175
r359 147 149 49.381 $w=2.08e-07 $l=9.35e-07 $layer=LI1_cond $X=2.035 $Y=1.18
+ $X2=2.97 $Y2=1.18
r360 143 161 2.19032 $w=2.5e-07 $l=1.76635e-07 $layer=LI1_cond $X=1.91 $Y=1.065
+ $X2=1.78 $Y2=1.175
r361 143 145 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.91 $Y=1.065
+ $X2=1.91 $Y2=0.42
r362 139 141 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.69 $Y=1.62
+ $X2=1.69 $Y2=2.3
r363 137 161 2.19032 $w=3.3e-07 $l=1.48324e-07 $layer=LI1_cond $X=1.69 $Y=1.285
+ $X2=1.78 $Y2=1.175
r364 137 139 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=1.285
+ $X2=1.69 $Y2=1.62
r365 136 160 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.195 $Y=1.175
+ $X2=1.09 $Y2=1.175
r366 135 161 4.00838 $w=2.2e-07 $l=2.55e-07 $layer=LI1_cond $X=1.525 $Y=1.175
+ $X2=1.78 $Y2=1.175
r367 135 136 17.2866 $w=2.18e-07 $l=3.3e-07 $layer=LI1_cond $X=1.525 $Y=1.175
+ $X2=1.195 $Y2=1.175
r368 131 160 0.99856 $w=2.1e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=1.065
+ $X2=1.09 $Y2=1.175
r369 131 133 34.0649 $w=2.08e-07 $l=6.45e-07 $layer=LI1_cond $X=1.09 $Y=1.065
+ $X2=1.09 $Y2=0.42
r370 129 158 1.91462 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=0.925 $Y=1.285
+ $X2=0.925 $Y2=1.175
r371 129 157 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.925 $Y=1.285
+ $X2=0.925 $Y2=1.495
r372 125 156 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=0.85 $Y=1.66
+ $X2=0.85 $Y2=1.62
r373 125 127 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=0.85 $Y=1.66
+ $X2=0.85 $Y2=2.3
r374 121 180 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.18 $Y=1.325
+ $X2=9.18 $Y2=1.16
r375 121 123 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.18 $Y=1.325
+ $X2=9.18 $Y2=1.985
r376 118 180 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.18 $Y=0.995
+ $X2=9.18 $Y2=1.16
r377 118 120 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.18 $Y=0.995
+ $X2=9.18 $Y2=0.56
r378 114 178 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=1.325
+ $X2=8.76 $Y2=1.16
r379 114 116 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.76 $Y=1.325
+ $X2=8.76 $Y2=1.985
r380 111 178 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=0.995
+ $X2=8.76 $Y2=1.16
r381 111 113 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.76 $Y=0.995
+ $X2=8.76 $Y2=0.56
r382 107 177 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.34 $Y=1.325
+ $X2=8.34 $Y2=1.16
r383 107 109 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.34 $Y=1.325
+ $X2=8.34 $Y2=1.985
r384 104 177 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.34 $Y=0.995
+ $X2=8.34 $Y2=1.16
r385 104 106 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.34 $Y=0.995
+ $X2=8.34 $Y2=0.56
r386 100 176 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.92 $Y=1.325
+ $X2=7.92 $Y2=1.16
r387 100 102 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.92 $Y=1.325
+ $X2=7.92 $Y2=1.985
r388 97 176 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.92 $Y=0.995
+ $X2=7.92 $Y2=1.16
r389 97 99 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.92 $Y=0.995
+ $X2=7.92 $Y2=0.56
r390 93 175 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.5 $Y=1.325
+ $X2=7.5 $Y2=1.16
r391 93 95 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.5 $Y=1.325
+ $X2=7.5 $Y2=1.985
r392 90 175 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.5 $Y=0.995
+ $X2=7.5 $Y2=1.16
r393 90 92 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.5 $Y=0.995
+ $X2=7.5 $Y2=0.56
r394 86 174 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.08 $Y=1.325
+ $X2=7.08 $Y2=1.16
r395 86 88 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.08 $Y=1.325
+ $X2=7.08 $Y2=1.985
r396 83 174 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.08 $Y=0.995
+ $X2=7.08 $Y2=1.16
r397 83 85 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.08 $Y=0.995
+ $X2=7.08 $Y2=0.56
r398 79 173 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.325
+ $X2=6.66 $Y2=1.16
r399 79 81 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.66 $Y=1.325
+ $X2=6.66 $Y2=1.985
r400 76 173 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=0.995
+ $X2=6.66 $Y2=1.16
r401 76 78 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.66 $Y=0.995
+ $X2=6.66 $Y2=0.56
r402 72 172 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=1.325
+ $X2=6.24 $Y2=1.16
r403 72 74 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.24 $Y=1.325
+ $X2=6.24 $Y2=1.985
r404 69 172 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=0.995
+ $X2=6.24 $Y2=1.16
r405 69 71 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.24 $Y=0.995
+ $X2=6.24 $Y2=0.56
r406 65 171 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.82 $Y=1.325
+ $X2=5.82 $Y2=1.16
r407 65 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.82 $Y=1.325
+ $X2=5.82 $Y2=1.985
r408 62 171 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.82 $Y=0.995
+ $X2=5.82 $Y2=1.16
r409 62 64 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.82 $Y=0.995
+ $X2=5.82 $Y2=0.56
r410 58 170 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=1.325
+ $X2=5.4 $Y2=1.16
r411 58 60 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.4 $Y=1.325
+ $X2=5.4 $Y2=1.985
r412 55 170 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=0.995
+ $X2=5.4 $Y2=1.16
r413 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.4 $Y=0.995
+ $X2=5.4 $Y2=0.56
r414 51 169 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.98 $Y=1.325
+ $X2=4.98 $Y2=1.16
r415 51 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.98 $Y=1.325
+ $X2=4.98 $Y2=1.985
r416 48 169 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.98 $Y=0.995
+ $X2=4.98 $Y2=1.16
r417 48 50 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.98 $Y=0.995
+ $X2=4.98 $Y2=0.56
r418 44 168 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.56 $Y=1.325
+ $X2=4.56 $Y2=1.16
r419 44 46 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.56 $Y=1.325
+ $X2=4.56 $Y2=1.985
r420 41 168 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.56 $Y=0.995
+ $X2=4.56 $Y2=1.16
r421 41 43 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.56 $Y=0.995
+ $X2=4.56 $Y2=0.56
r422 37 167 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.325
+ $X2=4.14 $Y2=1.16
r423 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.14 $Y=1.325
+ $X2=4.14 $Y2=1.985
r424 34 167 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=0.995
+ $X2=4.14 $Y2=1.16
r425 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.14 $Y=0.995
+ $X2=4.14 $Y2=0.56
r426 30 166 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.325
+ $X2=3.72 $Y2=1.16
r427 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.72 $Y=1.325
+ $X2=3.72 $Y2=1.985
r428 27 166 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=0.995
+ $X2=3.72 $Y2=1.16
r429 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.72 $Y=0.995
+ $X2=3.72 $Y2=0.56
r430 23 165 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.325
+ $X2=3.3 $Y2=1.16
r431 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.3 $Y=1.325
+ $X2=3.3 $Y2=1.985
r432 20 165 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=0.995
+ $X2=3.3 $Y2=1.16
r433 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.3 $Y=0.995
+ $X2=3.3 $Y2=0.56
r434 16 162 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.325
+ $X2=2.88 $Y2=1.16
r435 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.88 $Y=1.325
+ $X2=2.88 $Y2=1.985
r436 13 162 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=0.995
+ $X2=2.88 $Y2=1.16
r437 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.88 $Y=0.995
+ $X2=2.88 $Y2=0.56
r438 4 141 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.485 $X2=1.69 $Y2=2.3
r439 4 139 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.485 $X2=1.69 $Y2=1.62
r440 3 156 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.485 $X2=0.85 $Y2=1.62
r441 3 127 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.485 $X2=0.85 $Y2=2.3
r442 2 145 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=1.775
+ $Y=0.235 $X2=1.91 $Y2=0.42
r443 1 133 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=0.235 $X2=1.07 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%SLEEP 1 3 6 8 10 13 15 17 20 22
+ 24 27 29 31 34 36 38 41 43 45 48 50 52 55 57 59 62 64 66 69 71 73 76 78 80 83
+ 85 87 90 92 94 97 99 101 104 106 108 111 113 119 137
r281 136 137 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=15.48 $Y=1.16
+ $X2=15.9 $Y2=1.16
r282 134 136 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=15.47 $Y=1.16
+ $X2=15.48 $Y2=1.16
r283 132 134 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=15.06 $Y=1.16
+ $X2=15.47 $Y2=1.16
r284 131 132 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=14.64 $Y=1.16
+ $X2=15.06 $Y2=1.16
r285 130 131 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=14.22 $Y=1.16
+ $X2=14.64 $Y2=1.16
r286 129 130 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=13.8 $Y=1.16
+ $X2=14.22 $Y2=1.16
r287 128 129 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=13.38 $Y=1.16
+ $X2=13.8 $Y2=1.16
r288 127 128 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.96 $Y=1.16
+ $X2=13.38 $Y2=1.16
r289 126 127 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.54 $Y=1.16
+ $X2=12.96 $Y2=1.16
r290 125 126 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.12 $Y=1.16
+ $X2=12.54 $Y2=1.16
r291 124 125 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.7 $Y=1.16
+ $X2=12.12 $Y2=1.16
r292 123 124 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.28 $Y=1.16
+ $X2=11.7 $Y2=1.16
r293 122 123 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=10.86 $Y=1.16
+ $X2=11.28 $Y2=1.16
r294 121 122 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=10.44 $Y=1.16
+ $X2=10.86 $Y2=1.16
r295 120 121 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=10.02 $Y=1.16
+ $X2=10.44 $Y2=1.16
r296 119 134 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=15.47
+ $Y=1.16 $X2=15.47 $Y2=1.16
r297 118 120 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=9.69 $Y=1.16
+ $X2=10.02 $Y2=1.16
r298 118 119 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=9.69
+ $Y=1.16 $X2=9.69 $Y2=1.16
r299 115 118 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.6 $Y=1.16
+ $X2=9.69 $Y2=1.16
r300 113 119 0.0590323 $w=6.198e-06 $l=3e-08 $layer=LI1_cond $X=12.55 $Y=1.19
+ $X2=12.55 $Y2=1.16
r301 109 137 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.9 $Y=1.325
+ $X2=15.9 $Y2=1.16
r302 109 111 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=15.9 $Y=1.325
+ $X2=15.9 $Y2=1.985
r303 106 137 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.9 $Y=0.995
+ $X2=15.9 $Y2=1.16
r304 106 108 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.9 $Y=0.995
+ $X2=15.9 $Y2=0.56
r305 102 136 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.48 $Y=1.325
+ $X2=15.48 $Y2=1.16
r306 102 104 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=15.48 $Y=1.325
+ $X2=15.48 $Y2=1.985
r307 99 136 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.48 $Y=0.995
+ $X2=15.48 $Y2=1.16
r308 99 101 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.48 $Y=0.995
+ $X2=15.48 $Y2=0.56
r309 95 132 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.06 $Y=1.325
+ $X2=15.06 $Y2=1.16
r310 95 97 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=15.06 $Y=1.325
+ $X2=15.06 $Y2=1.985
r311 92 132 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.06 $Y=0.995
+ $X2=15.06 $Y2=1.16
r312 92 94 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.06 $Y=0.995
+ $X2=15.06 $Y2=0.56
r313 88 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.64 $Y=1.325
+ $X2=14.64 $Y2=1.16
r314 88 90 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.64 $Y=1.325
+ $X2=14.64 $Y2=1.985
r315 85 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.64 $Y=0.995
+ $X2=14.64 $Y2=1.16
r316 85 87 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.64 $Y=0.995
+ $X2=14.64 $Y2=0.56
r317 81 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.22 $Y=1.325
+ $X2=14.22 $Y2=1.16
r318 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.22 $Y=1.325
+ $X2=14.22 $Y2=1.985
r319 78 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.22 $Y=0.995
+ $X2=14.22 $Y2=1.16
r320 78 80 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.22 $Y=0.995
+ $X2=14.22 $Y2=0.56
r321 74 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.8 $Y=1.325
+ $X2=13.8 $Y2=1.16
r322 74 76 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.8 $Y=1.325
+ $X2=13.8 $Y2=1.985
r323 71 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.8 $Y=0.995
+ $X2=13.8 $Y2=1.16
r324 71 73 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.8 $Y=0.995
+ $X2=13.8 $Y2=0.56
r325 67 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.38 $Y=1.325
+ $X2=13.38 $Y2=1.16
r326 67 69 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.38 $Y=1.325
+ $X2=13.38 $Y2=1.985
r327 64 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.38 $Y=0.995
+ $X2=13.38 $Y2=1.16
r328 64 66 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.38 $Y=0.995
+ $X2=13.38 $Y2=0.56
r329 60 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.96 $Y=1.325
+ $X2=12.96 $Y2=1.16
r330 60 62 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.96 $Y=1.325
+ $X2=12.96 $Y2=1.985
r331 57 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.96 $Y=0.995
+ $X2=12.96 $Y2=1.16
r332 57 59 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.96 $Y=0.995
+ $X2=12.96 $Y2=0.56
r333 53 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.54 $Y=1.325
+ $X2=12.54 $Y2=1.16
r334 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.54 $Y=1.325
+ $X2=12.54 $Y2=1.985
r335 50 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.54 $Y=0.995
+ $X2=12.54 $Y2=1.16
r336 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.54 $Y=0.995
+ $X2=12.54 $Y2=0.56
r337 46 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.12 $Y=1.325
+ $X2=12.12 $Y2=1.16
r338 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.12 $Y=1.325
+ $X2=12.12 $Y2=1.985
r339 43 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.12 $Y=0.995
+ $X2=12.12 $Y2=1.16
r340 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.12 $Y=0.995
+ $X2=12.12 $Y2=0.56
r341 39 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.7 $Y=1.325
+ $X2=11.7 $Y2=1.16
r342 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.7 $Y=1.325
+ $X2=11.7 $Y2=1.985
r343 36 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.7 $Y=0.995
+ $X2=11.7 $Y2=1.16
r344 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.7 $Y=0.995
+ $X2=11.7 $Y2=0.56
r345 32 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.28 $Y=1.325
+ $X2=11.28 $Y2=1.16
r346 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.28 $Y=1.325
+ $X2=11.28 $Y2=1.985
r347 29 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.28 $Y=0.995
+ $X2=11.28 $Y2=1.16
r348 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.28 $Y=0.995
+ $X2=11.28 $Y2=0.56
r349 25 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.86 $Y=1.325
+ $X2=10.86 $Y2=1.16
r350 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.86 $Y=1.325
+ $X2=10.86 $Y2=1.985
r351 22 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.86 $Y=0.995
+ $X2=10.86 $Y2=1.16
r352 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.86 $Y=0.995
+ $X2=10.86 $Y2=0.56
r353 18 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.44 $Y=1.325
+ $X2=10.44 $Y2=1.16
r354 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.44 $Y=1.325
+ $X2=10.44 $Y2=1.985
r355 15 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.44 $Y=0.995
+ $X2=10.44 $Y2=1.16
r356 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.44 $Y=0.995
+ $X2=10.44 $Y2=0.56
r357 11 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.02 $Y=1.325
+ $X2=10.02 $Y2=1.16
r358 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.02 $Y=1.325
+ $X2=10.02 $Y2=1.985
r359 8 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.02 $Y=0.995
+ $X2=10.02 $Y2=1.16
r360 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.02 $Y=0.995
+ $X2=10.02 $Y2=0.56
r361 4 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.6 $Y=1.325
+ $X2=9.6 $Y2=1.16
r362 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.6 $Y=1.325 $X2=9.6
+ $Y2=1.985
r363 1 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.6 $Y=0.995
+ $X2=9.6 $Y2=1.16
r364 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.6 $Y=0.995 $X2=9.6
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 36
+ 42 46 50 54 58 62 66 70 74 78 80 84 88 91 92 93 94 96 97 99 100 102 103 104
+ 105 106 115 133 143 144 147 150 153 156 159
r236 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r237 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r238 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r239 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r240 148 151 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r241 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r242 143 144 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r243 141 144 1.96334 $w=4.8e-07 $l=6.9e-06 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=16.33 $Y2=2.72
r244 141 160 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r245 140 143 450.16 $w=1.68e-07 $l=6.9e-06 $layer=LI1_cond $X=9.43 $Y=2.72
+ $X2=16.33 $Y2=2.72
r246 140 141 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r247 138 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.095 $Y=2.72
+ $X2=8.97 $Y2=2.72
r248 138 140 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.095 $Y=2.72
+ $X2=9.43 $Y2=2.72
r249 137 160 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r250 137 157 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r251 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r252 134 156 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.255 $Y=2.72
+ $X2=8.13 $Y2=2.72
r253 134 136 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.255 $Y=2.72
+ $X2=8.51 $Y2=2.72
r254 133 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.845 $Y=2.72
+ $X2=8.97 $Y2=2.72
r255 133 136 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.845 $Y=2.72
+ $X2=8.51 $Y2=2.72
r256 132 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r257 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r258 129 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r259 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r260 126 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r261 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r262 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r263 123 154 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r264 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r265 120 153 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.055 $Y=2.72
+ $X2=3.93 $Y2=2.72
r266 120 122 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.055 $Y=2.72
+ $X2=4.37 $Y2=2.72
r267 119 154 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r268 119 151 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r269 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r270 116 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.09 $Y2=2.72
r271 116 118 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.45 $Y2=2.72
r272 115 153 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.93 $Y2=2.72
r273 115 118 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.45 $Y2=2.72
r274 114 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r275 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r276 106 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r277 106 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r278 104 131 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.165 $Y=2.72
+ $X2=7.13 $Y2=2.72
r279 104 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.165 $Y=2.72
+ $X2=7.29 $Y2=2.72
r280 102 128 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.325 $Y=2.72
+ $X2=6.21 $Y2=2.72
r281 102 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.325 $Y=2.72
+ $X2=6.45 $Y2=2.72
r282 101 131 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=7.13 $Y2=2.72
r283 101 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.45 $Y2=2.72
r284 99 125 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.29 $Y2=2.72
r285 99 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.61 $Y2=2.72
r286 98 128 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=6.21 $Y2=2.72
r287 98 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.61 $Y2=2.72
r288 96 122 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.645 $Y=2.72
+ $X2=4.37 $Y2=2.72
r289 96 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.645 $Y=2.72
+ $X2=4.77 $Y2=2.72
r290 95 125 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=5.29 $Y2=2.72
r291 95 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.77 $Y2=2.72
r292 93 113 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.15 $Y2=2.72
r293 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.27 $Y2=2.72
r294 91 109 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.3 $Y=2.72 $X2=0.23
+ $Y2=2.72
r295 91 92 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.3 $Y=2.72
+ $X2=0.407 $Y2=2.72
r296 90 113 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=1.15 $Y2=2.72
r297 90 92 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.407 $Y2=2.72
r298 86 159 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=2.635
+ $X2=8.97 $Y2=2.72
r299 86 88 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.97 $Y=2.635
+ $X2=8.97 $Y2=2
r300 82 156 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.13 $Y=2.635
+ $X2=8.13 $Y2=2.72
r301 82 84 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.13 $Y=2.635
+ $X2=8.13 $Y2=2
r302 81 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.415 $Y=2.72
+ $X2=7.29 $Y2=2.72
r303 80 156 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.005 $Y=2.72
+ $X2=8.13 $Y2=2.72
r304 80 81 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.005 $Y=2.72
+ $X2=7.415 $Y2=2.72
r305 76 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.29 $Y=2.635
+ $X2=7.29 $Y2=2.72
r306 76 78 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.29 $Y=2.635
+ $X2=7.29 $Y2=2
r307 72 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=2.635
+ $X2=6.45 $Y2=2.72
r308 72 74 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.45 $Y=2.635
+ $X2=6.45 $Y2=2
r309 68 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.61 $Y=2.635
+ $X2=5.61 $Y2=2.72
r310 68 70 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=5.61 $Y=2.635
+ $X2=5.61 $Y2=2
r311 64 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=2.635
+ $X2=4.77 $Y2=2.72
r312 64 66 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.77 $Y=2.635
+ $X2=4.77 $Y2=2
r313 60 153 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=2.635
+ $X2=3.93 $Y2=2.72
r314 60 62 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.93 $Y=2.635
+ $X2=3.93 $Y2=2
r315 56 150 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=2.635
+ $X2=3.09 $Y2=2.72
r316 56 58 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.09 $Y=2.635
+ $X2=3.09 $Y2=2
r317 55 147 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.147 $Y2=2.72
r318 54 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=3.09 $Y2=2.72
r319 54 55 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.27 $Y2=2.72
r320 50 53 32.9269 $w=2.43e-07 $l=7e-07 $layer=LI1_cond $X=2.147 $Y=1.64
+ $X2=2.147 $Y2=2.34
r321 48 147 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.147 $Y=2.635
+ $X2=2.147 $Y2=2.72
r322 48 53 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=2.147 $Y=2.635
+ $X2=2.147 $Y2=2.34
r323 47 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.27 $Y2=2.72
r324 46 147 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.147 $Y2=2.72
r325 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.355 $Y2=2.72
r326 42 45 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.27 $Y=1.64 $X2=1.27
+ $Y2=2.34
r327 40 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2.72
r328 40 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2.34
r329 36 39 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=0.407 $Y=1.66
+ $X2=0.407 $Y2=2.34
r330 34 92 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.407 $Y=2.635
+ $X2=0.407 $Y2=2.72
r331 34 39 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.407 $Y=2.635
+ $X2=0.407 $Y2=2.34
r332 11 88 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.835
+ $Y=1.485 $X2=8.97 $Y2=2
r333 10 84 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.995
+ $Y=1.485 $X2=8.13 $Y2=2
r334 9 78 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.155
+ $Y=1.485 $X2=7.29 $Y2=2
r335 8 74 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.315
+ $Y=1.485 $X2=6.45 $Y2=2
r336 7 70 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.475
+ $Y=1.485 $X2=5.61 $Y2=2
r337 6 66 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.635
+ $Y=1.485 $X2=4.77 $Y2=2
r338 5 62 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.795
+ $Y=1.485 $X2=3.93 $Y2=2
r339 4 58 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.485 $X2=3.09 $Y2=2
r340 3 53 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.485 $X2=2.11 $Y2=2.34
r341 3 50 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.485 $X2=2.11 $Y2=1.64
r342 2 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.485 $X2=1.27 $Y2=2.34
r343 2 42 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.485 $X2=1.27 $Y2=1.64
r344 1 39 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.485 $X2=0.43 $Y2=2.34
r345 1 36 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.485 $X2=0.43 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A_505_297# 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 52 54 56 60 62 66 68 72 74 78 80 84 86 90 92 96 98 100
+ 101 102 106 108 112 114 118 120 124 126 130 132 136 138 142 144 148 153 155
+ 157 159 161 163 165 170 171 172 173 174 175 176
r215 146 148 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=16.11 $Y=2.295
+ $X2=16.11 $Y2=1.96
r216 145 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.395 $Y=2.38
+ $X2=15.27 $Y2=2.38
r217 144 146 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=15.985 $Y=2.38
+ $X2=16.11 $Y2=2.295
r218 144 145 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=15.985 $Y=2.38
+ $X2=15.395 $Y2=2.38
r219 140 176 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.27 $Y=2.295
+ $X2=15.27 $Y2=2.38
r220 140 142 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=15.27 $Y=2.295
+ $X2=15.27 $Y2=1.96
r221 139 175 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.555 $Y=2.38
+ $X2=14.43 $Y2=2.38
r222 138 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.145 $Y=2.38
+ $X2=15.27 $Y2=2.38
r223 138 139 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=15.145 $Y=2.38
+ $X2=14.555 $Y2=2.38
r224 134 175 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.43 $Y=2.295
+ $X2=14.43 $Y2=2.38
r225 134 136 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=14.43 $Y=2.295
+ $X2=14.43 $Y2=1.96
r226 133 174 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.715 $Y=2.38
+ $X2=13.59 $Y2=2.38
r227 132 175 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.305 $Y=2.38
+ $X2=14.43 $Y2=2.38
r228 132 133 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=14.305 $Y=2.38
+ $X2=13.715 $Y2=2.38
r229 128 174 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.59 $Y=2.295
+ $X2=13.59 $Y2=2.38
r230 128 130 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=13.59 $Y=2.295
+ $X2=13.59 $Y2=1.96
r231 127 173 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.875 $Y=2.38
+ $X2=12.75 $Y2=2.38
r232 126 174 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.465 $Y=2.38
+ $X2=13.59 $Y2=2.38
r233 126 127 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=13.465 $Y=2.38
+ $X2=12.875 $Y2=2.38
r234 122 173 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.75 $Y=2.295
+ $X2=12.75 $Y2=2.38
r235 122 124 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=12.75 $Y=2.295
+ $X2=12.75 $Y2=1.96
r236 121 172 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.035 $Y=2.38
+ $X2=11.91 $Y2=2.38
r237 120 173 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.625 $Y=2.38
+ $X2=12.75 $Y2=2.38
r238 120 121 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.625 $Y=2.38
+ $X2=12.035 $Y2=2.38
r239 116 172 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.91 $Y=2.295
+ $X2=11.91 $Y2=2.38
r240 116 118 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=11.91 $Y=2.295
+ $X2=11.91 $Y2=1.96
r241 115 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.195 $Y=2.38
+ $X2=11.07 $Y2=2.38
r242 114 172 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.785 $Y=2.38
+ $X2=11.91 $Y2=2.38
r243 114 115 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.785 $Y=2.38
+ $X2=11.195 $Y2=2.38
r244 110 171 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=2.295
+ $X2=11.07 $Y2=2.38
r245 110 112 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=11.07 $Y=2.295
+ $X2=11.07 $Y2=1.96
r246 109 170 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.355 $Y=2.38
+ $X2=10.23 $Y2=2.38
r247 108 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.945 $Y=2.38
+ $X2=11.07 $Y2=2.38
r248 108 109 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.945 $Y=2.38
+ $X2=10.355 $Y2=2.38
r249 104 170 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.23 $Y=2.295
+ $X2=10.23 $Y2=2.38
r250 104 106 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.23 $Y=2.295
+ $X2=10.23 $Y2=1.96
r251 103 169 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.515 $Y=2.38
+ $X2=9.39 $Y2=2.38
r252 102 170 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.105 $Y=2.38
+ $X2=10.23 $Y2=2.38
r253 102 103 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.105 $Y=2.38
+ $X2=9.515 $Y2=2.38
r254 101 169 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=2.295
+ $X2=9.39 $Y2=2.38
r255 100 167 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=9.39 $Y=1.665
+ $X2=9.39 $Y2=1.56
r256 100 101 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=9.39 $Y=1.665
+ $X2=9.39 $Y2=2.295
r257 99 165 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=8.675 $Y=1.56
+ $X2=8.55 $Y2=1.56
r258 98 167 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=9.265 $Y=1.56
+ $X2=9.39 $Y2=1.56
r259 98 99 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=9.265 $Y=1.56
+ $X2=8.675 $Y2=1.56
r260 94 165 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=8.55 $Y=1.665
+ $X2=8.55 $Y2=1.56
r261 94 96 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.55 $Y=1.665
+ $X2=8.55 $Y2=2.3
r262 93 163 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.835 $Y=1.56
+ $X2=7.71 $Y2=1.56
r263 92 165 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=8.425 $Y=1.56
+ $X2=8.55 $Y2=1.56
r264 92 93 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=8.425 $Y=1.56
+ $X2=7.835 $Y2=1.56
r265 88 163 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.71 $Y=1.665
+ $X2=7.71 $Y2=1.56
r266 88 90 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.71 $Y=1.665
+ $X2=7.71 $Y2=2.3
r267 87 161 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.995 $Y=1.56
+ $X2=6.87 $Y2=1.56
r268 86 163 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.585 $Y=1.56
+ $X2=7.71 $Y2=1.56
r269 86 87 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=7.585 $Y=1.56
+ $X2=6.995 $Y2=1.56
r270 82 161 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=6.87 $Y=1.665
+ $X2=6.87 $Y2=1.56
r271 82 84 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.87 $Y=1.665
+ $X2=6.87 $Y2=2.3
r272 81 159 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.155 $Y=1.56
+ $X2=6.03 $Y2=1.56
r273 80 161 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=6.745 $Y=1.56
+ $X2=6.87 $Y2=1.56
r274 80 81 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=6.745 $Y=1.56
+ $X2=6.155 $Y2=1.56
r275 76 159 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=6.03 $Y=1.665
+ $X2=6.03 $Y2=1.56
r276 76 78 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.03 $Y=1.665
+ $X2=6.03 $Y2=2.3
r277 75 157 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.315 $Y=1.56
+ $X2=5.19 $Y2=1.56
r278 74 159 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.905 $Y=1.56
+ $X2=6.03 $Y2=1.56
r279 74 75 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=5.905 $Y=1.56
+ $X2=5.315 $Y2=1.56
r280 70 157 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.19 $Y=1.665
+ $X2=5.19 $Y2=1.56
r281 70 72 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=5.19 $Y=1.665
+ $X2=5.19 $Y2=2.3
r282 69 155 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.475 $Y=1.56
+ $X2=4.35 $Y2=1.56
r283 68 157 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.065 $Y=1.56
+ $X2=5.19 $Y2=1.56
r284 68 69 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=5.065 $Y=1.56
+ $X2=4.475 $Y2=1.56
r285 64 155 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.35 $Y=1.665
+ $X2=4.35 $Y2=1.56
r286 64 66 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.35 $Y=1.665
+ $X2=4.35 $Y2=2.3
r287 63 153 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.635 $Y=1.56
+ $X2=3.51 $Y2=1.56
r288 62 155 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.225 $Y=1.56
+ $X2=4.35 $Y2=1.56
r289 62 63 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.225 $Y=1.56
+ $X2=3.635 $Y2=1.56
r290 58 153 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.51 $Y=1.665
+ $X2=3.51 $Y2=1.56
r291 58 60 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.51 $Y=1.665
+ $X2=3.51 $Y2=2.3
r292 57 151 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=2.795 $Y=1.56
+ $X2=2.635 $Y2=1.56
r293 56 153 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.385 $Y=1.56
+ $X2=3.51 $Y2=1.56
r294 56 57 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=3.385 $Y=1.56
+ $X2=2.795 $Y2=1.56
r295 52 151 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=1.56
r296 52 54 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=2.3
r297 17 148 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=15.975
+ $Y=1.485 $X2=16.11 $Y2=1.96
r298 16 142 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=15.135
+ $Y=1.485 $X2=15.27 $Y2=1.96
r299 15 136 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=14.295
+ $Y=1.485 $X2=14.43 $Y2=1.96
r300 14 130 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=13.455
+ $Y=1.485 $X2=13.59 $Y2=1.96
r301 13 124 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=12.615
+ $Y=1.485 $X2=12.75 $Y2=1.96
r302 12 118 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=11.775
+ $Y=1.485 $X2=11.91 $Y2=1.96
r303 11 112 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=10.935
+ $Y=1.485 $X2=11.07 $Y2=1.96
r304 10 106 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=10.095
+ $Y=1.485 $X2=10.23 $Y2=1.96
r305 9 169 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.255
+ $Y=1.485 $X2=9.39 $Y2=2.3
r306 9 167 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.255
+ $Y=1.485 $X2=9.39 $Y2=1.62
r307 8 165 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.415
+ $Y=1.485 $X2=8.55 $Y2=1.62
r308 8 96 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.415
+ $Y=1.485 $X2=8.55 $Y2=2.3
r309 7 163 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.485 $X2=7.71 $Y2=1.62
r310 7 90 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.485 $X2=7.71 $Y2=2.3
r311 6 161 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.485 $X2=6.87 $Y2=1.62
r312 6 84 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.485 $X2=6.87 $Y2=2.3
r313 5 159 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.895
+ $Y=1.485 $X2=6.03 $Y2=1.62
r314 5 78 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.895
+ $Y=1.485 $X2=6.03 $Y2=2.3
r315 4 157 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=1.485 $X2=5.19 $Y2=1.62
r316 4 72 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=1.485 $X2=5.19 $Y2=2.3
r317 3 155 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=1.485 $X2=4.35 $Y2=1.62
r318 3 66 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=1.485 $X2=4.35 $Y2=2.3
r319 2 153 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.485 $X2=3.51 $Y2=1.62
r320 2 60 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.485 $X2=3.51 $Y2=2.3
r321 1 151 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.67 $Y2=1.62
r322 1 54 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.67 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13
+ 14 15 16 17 18 19 20 21 22 23 24 75 77 78 81 83 87 89 93 95 99 101 105 107 111
+ 113 117 119 123 127 129 133 137 139 143 147 149 153 157 159 163 167 169 173
+ 177 179 183 187 189 193 197 198 199 200 201 202 203 204 206 207 209 210 212
+ 213 215 216 218 219 221 222 224 226 227
r467 227 230 2.15548 $w=4.52e-07 $l=1.64085e-07 $layer=LI1_cond $X=16.02 $Y=1.54
+ $X2=16.147 $Y2=1.455
r468 227 230 0.0913037 $w=6.53e-07 $l=5e-09 $layer=LI1_cond $X=16.147 $Y=1.45
+ $X2=16.147 $Y2=1.455
r469 225 227 9.9521 $w=6.53e-07 $l=5.45e-07 $layer=LI1_cond $X=16.147 $Y=0.905
+ $X2=16.147 $Y2=1.45
r470 225 226 2.10047 $w=4.92e-07 $l=1.86652e-07 $layer=LI1_cond $X=16.147
+ $Y=0.905 $X2=16 $Y2=0.815
r471 191 226 2.10047 $w=4.92e-07 $l=3.52136e-07 $layer=LI1_cond $X=15.69
+ $Y=0.725 $X2=16 $Y2=0.815
r472 191 193 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=15.69 $Y=0.725
+ $X2=15.69 $Y2=0.39
r473 190 222 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.015 $Y=0.815
+ $X2=14.85 $Y2=0.815
r474 189 226 5.1218 $w=1.8e-07 $l=4.75e-07 $layer=LI1_cond $X=15.525 $Y=0.815
+ $X2=16 $Y2=0.815
r475 189 190 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=15.525 $Y=0.815
+ $X2=15.015 $Y2=0.815
r476 188 224 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.975 $Y=1.54
+ $X2=14.85 $Y2=1.54
r477 187 227 5.01601 $w=1.7e-07 $l=4.55e-07 $layer=LI1_cond $X=15.565 $Y=1.54
+ $X2=16.02 $Y2=1.54
r478 187 188 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=15.565 $Y=1.54
+ $X2=14.975 $Y2=1.54
r479 181 222 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=14.85 $Y=0.725
+ $X2=14.85 $Y2=0.815
r480 181 183 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.85 $Y=0.725
+ $X2=14.85 $Y2=0.39
r481 180 219 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.175 $Y=0.815
+ $X2=14.01 $Y2=0.815
r482 179 222 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.685 $Y=0.815
+ $X2=14.85 $Y2=0.815
r483 179 180 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=14.685 $Y=0.815
+ $X2=14.175 $Y2=0.815
r484 178 221 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.135 $Y=1.54
+ $X2=14.01 $Y2=1.54
r485 177 224 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.725 $Y=1.54
+ $X2=14.85 $Y2=1.54
r486 177 178 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=14.725 $Y=1.54
+ $X2=14.135 $Y2=1.54
r487 171 219 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=14.01 $Y=0.725
+ $X2=14.01 $Y2=0.815
r488 171 173 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.01 $Y=0.725
+ $X2=14.01 $Y2=0.39
r489 170 216 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.335 $Y=0.815
+ $X2=13.17 $Y2=0.815
r490 169 219 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.845 $Y=0.815
+ $X2=14.01 $Y2=0.815
r491 169 170 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=13.845 $Y=0.815
+ $X2=13.335 $Y2=0.815
r492 168 218 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.295 $Y=1.54
+ $X2=13.17 $Y2=1.54
r493 167 221 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.885 $Y=1.54
+ $X2=14.01 $Y2=1.54
r494 167 168 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=13.885 $Y=1.54
+ $X2=13.295 $Y2=1.54
r495 161 216 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=13.17 $Y=0.725
+ $X2=13.17 $Y2=0.815
r496 161 163 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.17 $Y=0.725
+ $X2=13.17 $Y2=0.39
r497 160 213 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.495 $Y=0.815
+ $X2=12.33 $Y2=0.815
r498 159 216 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.005 $Y=0.815
+ $X2=13.17 $Y2=0.815
r499 159 160 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=13.005 $Y=0.815
+ $X2=12.495 $Y2=0.815
r500 158 215 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.455 $Y=1.54
+ $X2=12.33 $Y2=1.54
r501 157 218 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.045 $Y=1.54
+ $X2=13.17 $Y2=1.54
r502 157 158 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=13.045 $Y=1.54
+ $X2=12.455 $Y2=1.54
r503 151 213 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=12.33 $Y=0.725
+ $X2=12.33 $Y2=0.815
r504 151 153 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.33 $Y=0.725
+ $X2=12.33 $Y2=0.39
r505 150 210 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.655 $Y=0.815
+ $X2=11.49 $Y2=0.815
r506 149 213 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.165 $Y=0.815
+ $X2=12.33 $Y2=0.815
r507 149 150 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=12.165 $Y=0.815
+ $X2=11.655 $Y2=0.815
r508 148 212 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.615 $Y=1.54
+ $X2=11.49 $Y2=1.54
r509 147 215 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.205 $Y=1.54
+ $X2=12.33 $Y2=1.54
r510 147 148 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.205 $Y=1.54
+ $X2=11.615 $Y2=1.54
r511 141 210 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=11.49 $Y=0.725
+ $X2=11.49 $Y2=0.815
r512 141 143 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.49 $Y=0.725
+ $X2=11.49 $Y2=0.39
r513 140 207 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.815 $Y=0.815
+ $X2=10.65 $Y2=0.815
r514 139 210 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.325 $Y=0.815
+ $X2=11.49 $Y2=0.815
r515 139 140 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=11.325 $Y=0.815
+ $X2=10.815 $Y2=0.815
r516 138 209 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.775 $Y=1.54
+ $X2=10.65 $Y2=1.54
r517 137 212 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.365 $Y=1.54
+ $X2=11.49 $Y2=1.54
r518 137 138 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.365 $Y=1.54
+ $X2=10.775 $Y2=1.54
r519 131 207 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=10.65 $Y=0.725
+ $X2=10.65 $Y2=0.815
r520 131 133 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.65 $Y=0.725
+ $X2=10.65 $Y2=0.39
r521 130 204 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.975 $Y=0.815
+ $X2=9.81 $Y2=0.815
r522 129 207 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=0.815
+ $X2=10.65 $Y2=0.815
r523 129 130 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=10.485 $Y=0.815
+ $X2=9.975 $Y2=0.815
r524 128 206 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.935 $Y=1.54
+ $X2=9.81 $Y2=1.54
r525 127 209 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.525 $Y=1.54
+ $X2=10.65 $Y2=1.54
r526 127 128 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.525 $Y=1.54
+ $X2=9.935 $Y2=1.54
r527 121 204 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=9.81 $Y=0.725
+ $X2=9.81 $Y2=0.815
r528 121 123 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.81 $Y=0.725
+ $X2=9.81 $Y2=0.39
r529 120 203 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.135 $Y=0.815
+ $X2=8.97 $Y2=0.815
r530 119 204 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.645 $Y=0.815
+ $X2=9.81 $Y2=0.815
r531 119 120 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=9.645 $Y=0.815
+ $X2=9.135 $Y2=0.815
r532 115 203 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.97 $Y=0.725
+ $X2=8.97 $Y2=0.815
r533 115 117 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.97 $Y=0.725
+ $X2=8.97 $Y2=0.39
r534 114 202 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.295 $Y=0.815
+ $X2=8.13 $Y2=0.815
r535 113 203 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.805 $Y=0.815
+ $X2=8.97 $Y2=0.815
r536 113 114 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=8.805 $Y=0.815
+ $X2=8.295 $Y2=0.815
r537 109 202 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.13 $Y=0.725
+ $X2=8.13 $Y2=0.815
r538 109 111 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.13 $Y=0.725
+ $X2=8.13 $Y2=0.39
r539 108 201 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=0.815
+ $X2=7.29 $Y2=0.815
r540 107 202 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.965 $Y=0.815
+ $X2=8.13 $Y2=0.815
r541 107 108 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.965 $Y=0.815
+ $X2=7.455 $Y2=0.815
r542 103 201 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.29 $Y=0.725
+ $X2=7.29 $Y2=0.815
r543 103 105 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.29 $Y=0.725
+ $X2=7.29 $Y2=0.39
r544 102 200 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.615 $Y=0.815
+ $X2=6.45 $Y2=0.815
r545 101 201 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=0.815
+ $X2=7.29 $Y2=0.815
r546 101 102 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.125 $Y=0.815
+ $X2=6.615 $Y2=0.815
r547 97 200 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.45 $Y=0.725
+ $X2=6.45 $Y2=0.815
r548 97 99 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.45 $Y=0.725
+ $X2=6.45 $Y2=0.39
r549 96 199 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0.815
+ $X2=5.61 $Y2=0.815
r550 95 200 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.285 $Y=0.815
+ $X2=6.45 $Y2=0.815
r551 95 96 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.285 $Y=0.815
+ $X2=5.775 $Y2=0.815
r552 91 199 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.61 $Y=0.725
+ $X2=5.61 $Y2=0.815
r553 91 93 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.61 $Y=0.725
+ $X2=5.61 $Y2=0.39
r554 90 198 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=0.815
+ $X2=4.77 $Y2=0.815
r555 89 199 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.445 $Y=0.815
+ $X2=5.61 $Y2=0.815
r556 89 90 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.445 $Y=0.815
+ $X2=4.935 $Y2=0.815
r557 85 198 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.77 $Y=0.725
+ $X2=4.77 $Y2=0.815
r558 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.77 $Y=0.725
+ $X2=4.77 $Y2=0.39
r559 84 197 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0.815
+ $X2=3.93 $Y2=0.815
r560 83 198 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=0.815
+ $X2=4.77 $Y2=0.815
r561 83 84 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.605 $Y=0.815
+ $X2=4.095 $Y2=0.815
r562 79 197 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.93 $Y=0.725
+ $X2=3.93 $Y2=0.815
r563 79 81 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.93 $Y=0.725
+ $X2=3.93 $Y2=0.39
r564 77 197 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0.815
+ $X2=3.93 $Y2=0.815
r565 77 78 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.765 $Y=0.815
+ $X2=3.255 $Y2=0.815
r566 73 78 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.09 $Y=0.725
+ $X2=3.255 $Y2=0.815
r567 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.09 $Y=0.725
+ $X2=3.09 $Y2=0.39
r568 24 227 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=15.555
+ $Y=1.485 $X2=15.69 $Y2=1.62
r569 23 224 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=14.715
+ $Y=1.485 $X2=14.85 $Y2=1.62
r570 22 221 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=13.875
+ $Y=1.485 $X2=14.01 $Y2=1.62
r571 21 218 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=13.035
+ $Y=1.485 $X2=13.17 $Y2=1.62
r572 20 215 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=12.195
+ $Y=1.485 $X2=12.33 $Y2=1.62
r573 19 212 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=11.355
+ $Y=1.485 $X2=11.49 $Y2=1.62
r574 18 209 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=10.515
+ $Y=1.485 $X2=10.65 $Y2=1.62
r575 17 206 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=9.675
+ $Y=1.485 $X2=9.81 $Y2=1.62
r576 16 193 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=15.555
+ $Y=0.235 $X2=15.69 $Y2=0.39
r577 15 183 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=14.715
+ $Y=0.235 $X2=14.85 $Y2=0.39
r578 14 173 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=13.875
+ $Y=0.235 $X2=14.01 $Y2=0.39
r579 13 163 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=13.035
+ $Y=0.235 $X2=13.17 $Y2=0.39
r580 12 153 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=12.195
+ $Y=0.235 $X2=12.33 $Y2=0.39
r581 11 143 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=11.355
+ $Y=0.235 $X2=11.49 $Y2=0.39
r582 10 133 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.515
+ $Y=0.235 $X2=10.65 $Y2=0.39
r583 9 123 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.675
+ $Y=0.235 $X2=9.81 $Y2=0.39
r584 8 117 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.835
+ $Y=0.235 $X2=8.97 $Y2=0.39
r585 7 111 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.995
+ $Y=0.235 $X2=8.13 $Y2=0.39
r586 6 105 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.155
+ $Y=0.235 $X2=7.29 $Y2=0.39
r587 5 99 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.315
+ $Y=0.235 $X2=6.45 $Y2=0.39
r588 4 93 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.475
+ $Y=0.235 $X2=5.61 $Y2=0.39
r589 3 87 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.635
+ $Y=0.235 $X2=4.77 $Y2=0.39
r590 2 81 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.795
+ $Y=0.235 $X2=3.93 $Y2=0.39
r591 1 75 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.955
+ $Y=0.235 $X2=3.09 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 18 19 60 64 68 70 74 78 82 86 90 94 96 100 104 108 112 116 120
+ 122 126 130 134 136 138 141 142 144 145 147 148 150 151 153 154 155 156 158
+ 159 161 162 164 165 167 168 169 170 172 173 175 176 177 179 188 231 236 239
+ 242 245 248 252
r315 251 252 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r316 248 249 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r317 245 246 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r318 242 243 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r319 240 243 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r320 239 240 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r321 236 237 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r322 234 252 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=16.33 $Y2=0
r323 233 234 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r324 231 251 4.01862 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=16.025 $Y=0
+ $X2=16.292 $Y2=0
r325 231 233 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=16.025 $Y=0
+ $X2=15.87 $Y2=0
r326 230 234 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.95 $Y=0
+ $X2=15.87 $Y2=0
r327 229 230 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r328 227 230 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=14.95 $Y2=0
r329 227 249 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=13.57 $Y2=0
r330 226 227 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r331 224 248 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.675 $Y=0
+ $X2=13.59 $Y2=0
r332 224 226 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.675 $Y=0
+ $X2=14.03 $Y2=0
r333 223 249 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.57 $Y2=0
r334 222 223 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r335 220 223 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.65 $Y2=0
r336 219 220 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r337 217 220 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r338 216 217 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r339 214 217 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r340 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r341 211 214 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r342 211 246 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=8.51 $Y2=0
r343 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r344 208 245 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.635 $Y=0
+ $X2=8.55 $Y2=0
r345 208 210 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.635 $Y=0
+ $X2=8.97 $Y2=0
r346 207 246 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r347 206 207 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r348 204 207 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r349 203 204 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r350 201 204 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r351 200 201 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r352 198 201 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r353 197 198 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r354 195 198 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r355 195 243 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=3.45 $Y2=0
r356 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r357 192 242 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=3.51 $Y2=0
r358 192 194 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=3.91 $Y2=0
r359 191 240 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.53 $Y2=0
r360 190 191 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r361 188 239 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.48 $Y2=0
r362 188 190 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.07 $Y2=0
r363 187 191 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r364 187 237 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r365 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r366 184 236 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0
+ $X2=0.65 $Y2=0
r367 184 186 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0
+ $X2=1.15 $Y2=0
r368 179 236 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.65 $Y2=0
r369 179 181 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.23 $Y2=0
r370 177 237 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r371 177 181 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r372 175 229 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=15.185 $Y=0
+ $X2=14.95 $Y2=0
r373 175 176 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.185 $Y=0
+ $X2=15.27 $Y2=0
r374 174 233 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=15.355 $Y=0
+ $X2=15.87 $Y2=0
r375 174 176 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.355 $Y=0
+ $X2=15.27 $Y2=0
r376 172 226 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=14.345 $Y=0
+ $X2=14.03 $Y2=0
r377 172 173 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.345 $Y=0
+ $X2=14.43 $Y2=0
r378 171 229 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=14.515 $Y=0
+ $X2=14.95 $Y2=0
r379 171 173 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.515 $Y=0
+ $X2=14.43 $Y2=0
r380 169 222 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=12.665 $Y=0
+ $X2=12.65 $Y2=0
r381 169 170 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.665 $Y=0
+ $X2=12.75 $Y2=0
r382 167 219 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=11.73 $Y2=0
r383 167 168 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=11.91 $Y2=0
r384 166 222 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=11.995 $Y=0
+ $X2=12.65 $Y2=0
r385 166 168 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.995 $Y=0
+ $X2=11.91 $Y2=0
r386 164 216 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=10.81 $Y2=0
r387 164 165 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=11.07 $Y2=0
r388 163 219 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=11.73 $Y2=0
r389 163 165 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=11.07 $Y2=0
r390 161 213 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=9.89 $Y2=0
r391 161 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=10.23 $Y2=0
r392 160 216 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.81 $Y2=0
r393 160 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.23 $Y2=0
r394 158 210 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=8.97 $Y2=0
r395 158 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=9.39 $Y2=0
r396 157 213 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.475 $Y=0
+ $X2=9.89 $Y2=0
r397 157 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.475 $Y=0
+ $X2=9.39 $Y2=0
r398 155 206 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.59 $Y2=0
r399 155 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.71 $Y2=0
r400 153 203 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.785 $Y=0
+ $X2=6.67 $Y2=0
r401 153 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.785 $Y=0
+ $X2=6.87 $Y2=0
r402 152 206 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.955 $Y=0
+ $X2=7.59 $Y2=0
r403 152 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0
+ $X2=6.87 $Y2=0
r404 150 200 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=5.75 $Y2=0
r405 150 151 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=6.03 $Y2=0
r406 149 203 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.115 $Y=0
+ $X2=6.67 $Y2=0
r407 149 151 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=0
+ $X2=6.03 $Y2=0
r408 147 197 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.105 $Y=0
+ $X2=4.83 $Y2=0
r409 147 148 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=0
+ $X2=5.19 $Y2=0
r410 146 200 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.275 $Y=0
+ $X2=5.75 $Y2=0
r411 146 148 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.275 $Y=0
+ $X2=5.19 $Y2=0
r412 144 194 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.265 $Y=0
+ $X2=3.91 $Y2=0
r413 144 145 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=0
+ $X2=4.35 $Y2=0
r414 143 197 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.83 $Y2=0
r415 143 145 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.35 $Y2=0
r416 141 186 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.365 $Y=0
+ $X2=1.15 $Y2=0
r417 141 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.365 $Y=0
+ $X2=1.49 $Y2=0
r418 140 190 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=2.07 $Y2=0
r419 140 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=1.49 $Y2=0
r420 136 251 3.26607 $w=2.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=16.16 $Y=0.085
+ $X2=16.292 $Y2=0
r421 136 138 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=16.16 $Y=0.085
+ $X2=16.16 $Y2=0.39
r422 132 176 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.27 $Y=0.085
+ $X2=15.27 $Y2=0
r423 132 134 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=15.27 $Y=0.085
+ $X2=15.27 $Y2=0.39
r424 128 173 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.43 $Y=0.085
+ $X2=14.43 $Y2=0
r425 128 130 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.43 $Y=0.085
+ $X2=14.43 $Y2=0.39
r426 124 248 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.59 $Y=0.085
+ $X2=13.59 $Y2=0
r427 124 126 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.59 $Y=0.085
+ $X2=13.59 $Y2=0.39
r428 123 170 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.835 $Y=0
+ $X2=12.75 $Y2=0
r429 122 248 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.505 $Y=0
+ $X2=13.59 $Y2=0
r430 122 123 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.505 $Y=0
+ $X2=12.835 $Y2=0
r431 118 170 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.75 $Y=0.085
+ $X2=12.75 $Y2=0
r432 118 120 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=12.75 $Y=0.085
+ $X2=12.75 $Y2=0.39
r433 114 168 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.91 $Y=0.085
+ $X2=11.91 $Y2=0
r434 114 116 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.91 $Y=0.085
+ $X2=11.91 $Y2=0.39
r435 110 165 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=0.085
+ $X2=11.07 $Y2=0
r436 110 112 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.07 $Y=0.085
+ $X2=11.07 $Y2=0.39
r437 106 162 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.23 $Y=0.085
+ $X2=10.23 $Y2=0
r438 106 108 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.23 $Y=0.085
+ $X2=10.23 $Y2=0.39
r439 102 159 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=0.085
+ $X2=9.39 $Y2=0
r440 102 104 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.39 $Y=0.085
+ $X2=9.39 $Y2=0.39
r441 98 245 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.55 $Y=0.085
+ $X2=8.55 $Y2=0
r442 98 100 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.55 $Y=0.085
+ $X2=8.55 $Y2=0.39
r443 97 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.795 $Y=0 $X2=7.71
+ $Y2=0
r444 96 245 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=0 $X2=8.55
+ $Y2=0
r445 96 97 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.465 $Y=0
+ $X2=7.795 $Y2=0
r446 92 156 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.71 $Y=0.085
+ $X2=7.71 $Y2=0
r447 92 94 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.71 $Y=0.085
+ $X2=7.71 $Y2=0.39
r448 88 154 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.87 $Y=0.085
+ $X2=6.87 $Y2=0
r449 88 90 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.87 $Y=0.085
+ $X2=6.87 $Y2=0.39
r450 84 151 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0
r451 84 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0.39
r452 80 148 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0
r453 80 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0.39
r454 76 145 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.35 $Y=0.085
+ $X2=4.35 $Y2=0
r455 76 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.35 $Y=0.085
+ $X2=4.35 $Y2=0.39
r456 72 242 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.51 $Y=0.085
+ $X2=3.51 $Y2=0
r457 72 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.51 $Y=0.085
+ $X2=3.51 $Y2=0.39
r458 71 239 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=2.48 $Y2=0
r459 70 242 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.51
+ $Y2=0
r460 70 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.425 $Y=0
+ $X2=2.755 $Y2=0
r461 66 239 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0
r462 66 68 6.6328 $w=5.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0.39
r463 62 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=0.085
+ $X2=1.49 $Y2=0
r464 62 64 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=1.49 $Y=0.085
+ $X2=1.49 $Y2=0.39
r465 58 236 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.085
+ $X2=0.65 $Y2=0
r466 58 60 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.65 $Y=0.085
+ $X2=0.65 $Y2=0.39
r467 19 138 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=15.975
+ $Y=0.235 $X2=16.11 $Y2=0.39
r468 18 134 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=15.135
+ $Y=0.235 $X2=15.27 $Y2=0.39
r469 17 130 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=14.295
+ $Y=0.235 $X2=14.43 $Y2=0.39
r470 16 126 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=13.455
+ $Y=0.235 $X2=13.59 $Y2=0.39
r471 15 120 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=12.615
+ $Y=0.235 $X2=12.75 $Y2=0.39
r472 14 116 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=11.775
+ $Y=0.235 $X2=11.91 $Y2=0.39
r473 13 112 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.935
+ $Y=0.235 $X2=11.07 $Y2=0.39
r474 12 108 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.095
+ $Y=0.235 $X2=10.23 $Y2=0.39
r475 11 104 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.255
+ $Y=0.235 $X2=9.39 $Y2=0.39
r476 10 100 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.415
+ $Y=0.235 $X2=8.55 $Y2=0.39
r477 9 94 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.575
+ $Y=0.235 $X2=7.71 $Y2=0.39
r478 8 90 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.735
+ $Y=0.235 $X2=6.87 $Y2=0.39
r479 7 86 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.895
+ $Y=0.235 $X2=6.03 $Y2=0.39
r480 6 82 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.19 $Y2=0.39
r481 5 78 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.235 $X2=4.35 $Y2=0.39
r482 4 74 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.235 $X2=3.51 $Y2=0.39
r483 3 68 45.5 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_NDIFF $count=4 $X=2.195
+ $Y=0.235 $X2=2.67 $Y2=0.39
r484 2 64 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.355
+ $Y=0.235 $X2=1.49 $Y2=0.39
r485 1 60 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.525
+ $Y=0.235 $X2=0.65 $Y2=0.39
.ends


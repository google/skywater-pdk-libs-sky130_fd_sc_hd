* File: sky130_fd_sc_hd__and2b_1.spice
* Created: Thu Aug 27 14:07:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and2b_1.pex.spice"
.subckt sky130_fd_sc_hd__and2b_1  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_A_27_413#_M1007_d N_A_N_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_297_47# N_A_27_413#_M1001_g N_A_207_413#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1092 PD=0.66 PS=1.36 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g A_297_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0795252 AS=0.0504 PD=0.777196 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_207_413#_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.123075 PD=1.82 PS=1.2028 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_413#_M1003_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0714 AS=0.1092 PD=0.76 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1004 N_A_207_413#_M1004_d N_A_27_413#_M1004_g N_VPWR_M1003_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0609 AS=0.0714 PD=0.71 PS=0.76 NRD=2.3443 NRS=30.4759 M=1
+ R=2.8 SA=75000.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_207_413#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.134814 AS=0.0609 PD=1.0293 PS=0.71 NRD=21.0987 NRS=2.3443 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_207_413#_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.320986 PD=2.52 PS=2.4507 NRD=0 NRS=14.7553 M=1 R=6.66667
+ SA=75000.9 SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__and2b_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__xnor3_4.pxi.spice
* Created: Thu Aug 27 14:49:35 2020
* 
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_101_21# N_A_101_21#_M1024_d N_A_101_21#_M1011_d
+ N_A_101_21#_c_171_n N_A_101_21#_M1010_g N_A_101_21#_M1001_g
+ N_A_101_21#_c_172_n N_A_101_21#_M1015_g N_A_101_21#_M1002_g
+ N_A_101_21#_c_173_n N_A_101_21#_M1022_g N_A_101_21#_M1005_g
+ N_A_101_21#_c_174_n N_A_101_21#_M1027_g N_A_101_21#_M1014_g
+ N_A_101_21#_c_175_n N_A_101_21#_c_184_n N_A_101_21#_c_191_p
+ N_A_101_21#_c_196_p N_A_101_21#_c_224_p N_A_101_21#_c_176_n
+ N_A_101_21#_c_185_n N_A_101_21#_c_177_n N_A_101_21#_c_186_n
+ N_A_101_21#_c_187_n N_A_101_21#_c_178_n N_A_101_21#_c_200_p
+ N_A_101_21#_c_179_n PM_SKY130_FD_SC_HD__XNOR3_4%A_101_21#
x_PM_SKY130_FD_SC_HD__XNOR3_4%C N_C_c_306_n N_C_M1016_g N_C_c_311_n N_C_M1025_g
+ N_C_M1011_g N_C_c_307_n N_C_M1024_g N_C_c_308_n N_C_c_309_n N_C_c_310_n C
+ PM_SKY130_FD_SC_HD__XNOR3_4%C
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_492_93# N_A_492_93#_M1016_d N_A_492_93#_M1025_d
+ N_A_492_93#_c_374_n N_A_492_93#_M1026_g N_A_492_93#_M1020_g
+ N_A_492_93#_c_384_n N_A_492_93#_c_370_n N_A_492_93#_c_376_n
+ N_A_492_93#_c_377_n N_A_492_93#_c_378_n N_A_492_93#_c_371_n
+ N_A_492_93#_c_372_n N_A_492_93#_c_373_n PM_SKY130_FD_SC_HD__XNOR3_4%A_492_93#
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_1011_297# N_A_1011_297#_M1003_d
+ N_A_1011_297#_M1000_d N_A_1011_297#_M1021_g N_A_1011_297#_M1019_g
+ N_A_1011_297#_c_446_n N_A_1011_297#_M1008_g N_A_1011_297#_c_448_n
+ N_A_1011_297#_M1006_g N_A_1011_297#_c_449_n N_A_1011_297#_c_450_n
+ N_A_1011_297#_c_463_n N_A_1011_297#_c_451_n N_A_1011_297#_c_452_n
+ N_A_1011_297#_c_467_p N_A_1011_297#_c_453_n N_A_1011_297#_c_454_n
+ N_A_1011_297#_c_455_n N_A_1011_297#_c_456_n N_A_1011_297#_c_457_n
+ N_A_1011_297#_c_458_n PM_SKY130_FD_SC_HD__XNOR3_4%A_1011_297#
x_PM_SKY130_FD_SC_HD__XNOR3_4%B N_B_M1000_g N_B_M1003_g N_B_c_616_n N_B_c_617_n
+ N_B_M1007_g N_B_M1018_g N_B_c_626_n N_B_c_627_n N_B_M1023_g N_B_M1013_g
+ N_B_c_620_n N_B_c_621_n N_B_c_622_n N_B_c_631_n B N_B_c_623_n
+ PM_SKY130_FD_SC_HD__XNOR3_4%B
x_PM_SKY130_FD_SC_HD__XNOR3_4%A N_A_M1004_g N_A_M1017_g A N_A_c_735_n
+ N_A_c_736_n N_A_c_737_n PM_SKY130_FD_SC_HD__XNOR3_4%A
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_1117_297# N_A_1117_297#_M1007_s
+ N_A_1117_297#_M1006_d N_A_1117_297#_M1018_s N_A_1117_297#_M1008_d
+ N_A_1117_297#_c_779_n N_A_1117_297#_M1009_g N_A_1117_297#_M1012_g
+ N_A_1117_297#_c_780_n N_A_1117_297#_c_789_n N_A_1117_297#_c_781_n
+ N_A_1117_297#_c_782_n N_A_1117_297#_c_783_n N_A_1117_297#_c_791_n
+ N_A_1117_297#_c_784_n N_A_1117_297#_c_802_n N_A_1117_297#_c_785_n
+ N_A_1117_297#_c_786_n N_A_1117_297#_c_815_n N_A_1117_297#_c_816_n
+ PM_SKY130_FD_SC_HD__XNOR3_4%A_1117_297#
x_PM_SKY130_FD_SC_HD__XNOR3_4%VPWR N_VPWR_M1001_d N_VPWR_M1002_d N_VPWR_M1014_d
+ N_VPWR_M1000_s N_VPWR_M1017_d N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_917_n
+ N_VPWR_c_918_n N_VPWR_c_919_n N_VPWR_c_920_n N_VPWR_c_921_n N_VPWR_c_922_n
+ VPWR N_VPWR_c_923_n N_VPWR_c_924_n N_VPWR_c_925_n N_VPWR_c_926_n
+ N_VPWR_c_914_n N_VPWR_c_928_n N_VPWR_c_929_n N_VPWR_c_930_n N_VPWR_c_931_n
+ PM_SKY130_FD_SC_HD__XNOR3_4%VPWR
x_PM_SKY130_FD_SC_HD__XNOR3_4%X N_X_M1010_s N_X_M1022_s N_X_M1001_s N_X_M1005_s
+ N_X_c_1028_n N_X_c_1033_n N_X_c_1036_n N_X_c_1037_n N_X_c_1039_n N_X_c_1029_n
+ X N_X_c_1049_n PM_SKY130_FD_SC_HD__XNOR3_4%X
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_607_325# N_A_607_325#_M1020_d
+ N_A_607_325#_M1007_d N_A_607_325#_M1011_s N_A_607_325#_M1013_d
+ N_A_607_325#_c_1073_n N_A_607_325#_c_1067_n N_A_607_325#_c_1068_n
+ N_A_607_325#_c_1069_n N_A_607_325#_c_1075_n N_A_607_325#_c_1076_n
+ N_A_607_325#_c_1077_n N_A_607_325#_c_1078_n N_A_607_325#_c_1070_n
+ N_A_607_325#_c_1080_n N_A_607_325#_c_1116_n N_A_607_325#_c_1071_n
+ N_A_607_325#_c_1081_n N_A_607_325#_c_1072_n N_A_607_325#_c_1082_n
+ PM_SKY130_FD_SC_HD__XNOR3_4%A_607_325#
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_631_49# N_A_631_49#_M1024_s N_A_631_49#_M1023_d
+ N_A_631_49#_M1026_d N_A_631_49#_M1018_d N_A_631_49#_c_1228_n
+ N_A_631_49#_c_1216_n N_A_631_49#_c_1220_n N_A_631_49#_c_1257_n
+ N_A_631_49#_c_1221_n N_A_631_49#_c_1217_n N_A_631_49#_c_1329_p
+ N_A_631_49#_c_1218_n N_A_631_49#_c_1268_n N_A_631_49#_c_1288_n
+ N_A_631_49#_c_1223_n N_A_631_49#_c_1224_n N_A_631_49#_c_1225_n
+ N_A_631_49#_c_1226_n PM_SKY130_FD_SC_HD__XNOR3_4%A_631_49#
x_PM_SKY130_FD_SC_HD__XNOR3_4%A_1382_49# N_A_1382_49#_M1021_d
+ N_A_1382_49#_M1009_d N_A_1382_49#_M1019_d N_A_1382_49#_M1012_d
+ N_A_1382_49#_c_1345_n N_A_1382_49#_c_1357_n N_A_1382_49#_c_1349_n
+ N_A_1382_49#_c_1346_n N_A_1382_49#_c_1358_n N_A_1382_49#_c_1351_n
+ N_A_1382_49#_c_1347_n PM_SKY130_FD_SC_HD__XNOR3_4%A_1382_49#
x_PM_SKY130_FD_SC_HD__XNOR3_4%VGND N_VGND_M1010_d N_VGND_M1015_d N_VGND_M1027_d
+ N_VGND_M1003_s N_VGND_M1004_d N_VGND_c_1412_n N_VGND_c_1413_n N_VGND_c_1414_n
+ N_VGND_c_1415_n N_VGND_c_1416_n N_VGND_c_1417_n N_VGND_c_1418_n
+ N_VGND_c_1419_n N_VGND_c_1420_n N_VGND_c_1421_n N_VGND_c_1422_n
+ N_VGND_c_1423_n VGND N_VGND_c_1424_n N_VGND_c_1425_n N_VGND_c_1426_n
+ N_VGND_c_1427_n N_VGND_c_1428_n PM_SKY130_FD_SC_HD__XNOR3_4%VGND
cc_1 VNB N_A_101_21#_c_171_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_2 VNB N_A_101_21#_c_172_n 0.0160643f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.995
cc_3 VNB N_A_101_21#_c_173_n 0.0156266f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A_101_21#_c_174_n 0.0177713f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.995
cc_5 VNB N_A_101_21#_c_175_n 0.00105375f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.325
cc_6 VNB N_A_101_21#_c_176_n 0.00130544f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.695
cc_7 VNB N_A_101_21#_c_177_n 0.00178848f $X=-0.19 $Y=-0.24 $X2=2.485 $Y2=0.34
cc_8 VNB N_A_101_21#_c_178_n 0.0875417f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.16
cc_9 VNB N_A_101_21#_c_179_n 0.0170299f $X=-0.19 $Y=-0.24 $X2=3.45 $Y2=0.355
cc_10 VNB N_C_c_306_n 0.0195625f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=0.245
cc_11 VNB N_C_c_307_n 0.0212338f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_12 VNB N_C_c_308_n 0.010198f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_13 VNB N_C_c_309_n 0.0524249f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_14 VNB N_C_c_310_n 0.0123066f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.325
cc_15 VNB N_A_492_93#_c_370_n 0.00248343f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_16 VNB N_A_492_93#_c_371_n 0.00272073f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.995
cc_17 VNB N_A_492_93#_c_372_n 0.0221323f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.56
cc_18 VNB N_A_492_93#_c_373_n 0.0204272f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.985
cc_19 VNB N_A_1011_297#_M1021_g 0.0355486f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.56
cc_20 VNB N_A_1011_297#_c_446_n 0.0259644f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_21 VNB N_A_1011_297#_M1008_g 0.00127227f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.325
cc_22 VNB N_A_1011_297#_c_448_n 0.018065f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_23 VNB N_A_1011_297#_c_449_n 0.028835f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_24 VNB N_A_1011_297#_c_450_n 0.0140975f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_25 VNB N_A_1011_297#_c_451_n 0.00225945f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.325
cc_26 VNB N_A_1011_297#_c_452_n 0.00811041f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=0.78
cc_27 VNB N_A_1011_297#_c_453_n 0.0124845f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.96
cc_28 VNB N_A_1011_297#_c_454_n 6.17105e-19 $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=1.96
cc_29 VNB N_A_1011_297#_c_455_n 0.00274249f $X=-0.19 $Y=-0.24 $X2=2.6 $Y2=2.32
cc_30 VNB N_A_1011_297#_c_456_n 9.00189e-19 $X=-0.19 $Y=-0.24 $X2=3.645 $Y2=2.32
cc_31 VNB N_A_1011_297#_c_457_n 0.00544296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_1011_297#_c_458_n 0.0025002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_B_M1000_g 0.00411376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_B_M1003_g 0.0298518f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_35 VNB N_B_c_616_n 0.0515784f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.56
cc_36 VNB N_B_c_617_n 0.0170865f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.325
cc_37 VNB N_B_M1007_g 0.0285028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_B_M1018_g 0.00419882f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_39 VNB N_B_c_620_n 0.00493002f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.325
cc_40 VNB N_B_c_621_n 7.60368e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_B_c_622_n 0.0267383f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.325
cc_42 VNB N_B_c_623_n 0.0206335f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.425
cc_43 VNB N_A_c_735_n 0.0201493f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_44 VNB N_A_c_736_n 0.00393727f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_45 VNB N_A_c_737_n 0.0173356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1117_297#_c_779_n 0.0193901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1117_297#_c_780_n 0.00629819f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_48 VNB N_A_1117_297#_c_781_n 0.00264442f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.995
cc_49 VNB N_A_1117_297#_c_782_n 0.00179065f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.56
cc_50 VNB N_A_1117_297#_c_783_n 0.00347802f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.56
cc_51 VNB N_A_1117_297#_c_784_n 0.0235243f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.875
cc_52 VNB N_A_1117_297#_c_785_n 0.00204812f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=0.78
cc_53 VNB N_A_1117_297#_c_786_n 0.00464641f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.425
cc_54 VNB N_VPWR_c_914_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_X_c_1028_n 8.69283e-19 $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_56 VNB N_X_c_1029_n 8.39623e-19 $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.56
cc_57 VNB N_A_607_325#_c_1067_n 0.0106968f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.325
cc_58 VNB N_A_607_325#_c_1068_n 0.0134262f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.56
cc_59 VNB N_A_607_325#_c_1069_n 0.00277812f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.325
cc_60 VNB N_A_607_325#_c_1070_n 0.00223184f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.985
cc_61 VNB N_A_607_325#_c_1071_n 0.0103649f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=2.045
cc_62 VNB N_A_607_325#_c_1072_n 2.56766e-19 $X=-0.19 $Y=-0.24 $X2=2.485 $Y2=0.34
cc_63 VNB N_A_631_49#_c_1216_n 0.00886805f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_64 VNB N_A_631_49#_c_1217_n 0.00928634f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.325
cc_65 VNB N_A_631_49#_c_1218_n 0.00533463f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.56
cc_66 VNB N_A_1382_49#_c_1345_n 0.00783929f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_67 VNB N_A_1382_49#_c_1346_n 0.0307334f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.985
cc_68 VNB N_A_1382_49#_c_1347_n 0.0135316f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.875
cc_69 VNB N_VGND_c_1412_n 0.00419749f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_70 VNB N_VGND_c_1413_n 0.0194124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1414_n 0.00358658f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.325
cc_72 VNB N_VGND_c_1415_n 0.00226837f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.995
cc_73 VNB N_VGND_c_1416_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.985
cc_74 VNB N_VGND_c_1417_n 0.00468014f $X=-0.19 $Y=-0.24 $X2=2 $Y2=1.875
cc_75 VNB N_VGND_c_1418_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=0.78
cc_76 VNB N_VGND_c_1419_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.96
cc_77 VNB N_VGND_c_1420_n 0.0641689f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.425
cc_78 VNB N_VGND_c_1421_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.695
cc_79 VNB N_VGND_c_1422_n 0.0989889f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=2.235
cc_80 VNB N_VGND_c_1423_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=3.45 $Y2=0.34
cc_81 VNB N_VGND_c_1424_n 0.0159673f $X=-0.19 $Y=-0.24 $X2=1.982 $Y2=0.78
cc_82 VNB N_VGND_c_1425_n 0.0189867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1426_n 0.485372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1427_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1428_n 0.00353728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VPB N_A_101_21#_M1001_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_87 VPB N_A_101_21#_M1002_g 0.0181656f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_88 VPB N_A_101_21#_M1005_g 0.0181651f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.985
cc_89 VPB N_A_101_21#_M1014_g 0.0201602f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.985
cc_90 VPB N_A_101_21#_c_184_n 0.00152367f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.875
cc_91 VPB N_A_101_21#_c_185_n 0.00374454f $X=-0.19 $Y=1.305 $X2=2.515 $Y2=2.235
cc_92 VPB N_A_101_21#_c_186_n 0.00112766f $X=-0.19 $Y=1.305 $X2=2.6 $Y2=2.32
cc_93 VPB N_A_101_21#_c_187_n 0.0124058f $X=-0.19 $Y=1.305 $X2=3.645 $Y2=2.32
cc_94 VPB N_A_101_21#_c_178_n 0.0173651f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.16
cc_95 VPB N_C_c_311_n 0.0330326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_C_M1011_g 0.0323158f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.56
cc_97 VPB N_C_c_308_n 6.57939e-19 $X=-0.19 $Y=1.305 $X2=1 $Y2=0.56
cc_98 VPB N_C_c_309_n 0.0203296f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.56
cc_99 VPB N_C_c_310_n 0.00463557f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.325
cc_100 VPB N_A_492_93#_c_374_n 0.0261747f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=0.995
cc_101 VPB N_A_492_93#_c_370_n 0.00436454f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_102 VPB N_A_492_93#_c_376_n 0.0098968f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_492_93#_c_377_n 0.00173389f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_104 VPB N_A_492_93#_c_378_n 0.00184072f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.325
cc_105 VPB N_A_492_93#_c_371_n 2.68098e-19 $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.995
cc_106 VPB N_A_492_93#_c_372_n 0.00492238f $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.56
cc_107 VPB N_A_1011_297#_M1019_g 0.0247955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_1011_297#_M1008_g 0.0307087f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.325
cc_109 VPB N_A_1011_297#_c_449_n 0.0104529f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_110 VPB N_A_1011_297#_c_450_n 9.09516e-19 $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_111 VPB N_A_1011_297#_c_463_n 0.00806131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_1011_297#_c_458_n 0.00297191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_B_M1000_g 0.026301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_B_M1018_g 0.0236166f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_115 VPB N_B_c_626_n 0.110395f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_116 VPB N_B_c_627_n 0.0129123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_B_M1013_g 0.0314866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_B_c_621_n 9.25804e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_B_c_622_n 0.00514585f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.325
cc_120 VPB N_B_c_631_n 0.00168086f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=0.78
cc_121 VPB B 0.00780431f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=0.78
cc_122 VPB N_A_M1017_g 0.0197671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_c_735_n 0.00439035f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_124 VPB N_A_c_736_n 0.00141167f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_125 VPB N_A_1117_297#_M1012_g 0.0211416f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_126 VPB N_A_1117_297#_c_780_n 0.00271943f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_127 VPB N_A_1117_297#_c_789_n 0.00177722f $X=-0.19 $Y=1.305 $X2=1.45
+ $Y2=1.325
cc_128 VPB N_A_1117_297#_c_783_n 2.70069e-19 $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.56
cc_129 VPB N_A_1117_297#_c_791_n 0.0015591f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.325
cc_130 VPB N_A_1117_297#_c_784_n 0.004813f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.875
cc_131 VPB N_VPWR_c_915_n 0.00417382f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_132 VPB N_VPWR_c_916_n 0.0184034f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_133 VPB N_VPWR_c_917_n 0.00355058f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.985
cc_134 VPB N_VPWR_c_918_n 0.00675868f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.985
cc_135 VPB N_VPWR_c_919_n 0.00735011f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.875
cc_136 VPB N_VPWR_c_920_n 4.89207e-19 $X=-0.19 $Y=1.305 $X2=2.085 $Y2=1.96
cc_137 VPB N_VPWR_c_921_n 0.0112126f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=0.695
cc_138 VPB N_VPWR_c_922_n 0.00324402f $X=-0.19 $Y=1.305 $X2=2.515 $Y2=2.045
cc_139 VPB N_VPWR_c_923_n 0.0158681f $X=-0.19 $Y=1.305 $X2=3.645 $Y2=2.32
cc_140 VPB N_VPWR_c_924_n 0.0588598f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.16
cc_141 VPB N_VPWR_c_925_n 0.0887437f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=1.16
cc_142 VPB N_VPWR_c_926_n 0.0150434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_914_n 0.075831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_928_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_929_n 0.00517014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_930_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_931_n 0.00442675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_X_c_1029_n 0.00197606f $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.56
cc_149 VPB N_A_607_325#_c_1073_n 0.0110088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_607_325#_c_1069_n 0.00797136f $X=-0.19 $Y=1.305 $X2=1.45
+ $Y2=1.325
cc_151 VPB N_A_607_325#_c_1075_n 0.00296005f $X=-0.19 $Y=1.305 $X2=1.45
+ $Y2=1.985
cc_152 VPB N_A_607_325#_c_1076_n 0.00292375f $X=-0.19 $Y=1.305 $X2=1.85
+ $Y2=0.995
cc_153 VPB N_A_607_325#_c_1077_n 0.0105963f $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.56
cc_154 VPB N_A_607_325#_c_1078_n 0.00172555f $X=-0.19 $Y=1.305 $X2=1.85 $Y2=0.56
cc_155 VPB N_A_607_325#_c_1070_n 0.00149669f $X=-0.19 $Y=1.305 $X2=1.87
+ $Y2=1.985
cc_156 VPB N_A_607_325#_c_1080_n 0.0238947f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.325
cc_157 VPB N_A_607_325#_c_1081_n 3.60787e-19 $X=-0.19 $Y=1.305 $X2=3.45 $Y2=0.34
cc_158 VPB N_A_607_325#_c_1082_n 2.94232e-19 $X=-0.19 $Y=1.305 $X2=3.645
+ $Y2=2.32
cc_159 VPB N_A_631_49#_c_1216_n 0.00146756f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.56
cc_160 VPB N_A_631_49#_c_1220_n 0.00267409f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.325
cc_161 VPB N_A_631_49#_c_1221_n 6.69494e-19 $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.995
cc_162 VPB N_A_631_49#_c_1217_n 0.00210227f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.325
cc_163 VPB N_A_631_49#_c_1223_n 0.0147143f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.325
cc_164 VPB N_A_631_49#_c_1224_n 0.00333347f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.875
cc_165 VPB N_A_631_49#_c_1225_n 0.00870609f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.96
cc_166 VPB N_A_631_49#_c_1226_n 0.0014424f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=0.695
cc_167 VPB N_A_1382_49#_c_1345_n 0.00467504f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.56
cc_168 VPB N_A_1382_49#_c_1349_n 0.0147295f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_169 VPB N_A_1382_49#_c_1346_n 0.0229143f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.985
cc_170 VPB N_A_1382_49#_c_1351_n 0.0100871f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.325
cc_171 N_A_101_21#_c_174_n N_C_c_306_n 0.0147807f $X=1.85 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_172 N_A_101_21#_c_175_n N_C_c_306_n 0.00125959f $X=2 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_101_21#_c_191_p N_C_c_306_n 0.0117768f $X=2.315 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_101_21#_c_176_n N_C_c_306_n 0.0101804f $X=2.4 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_101_21#_c_177_n N_C_c_306_n 0.00609264f $X=2.485 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_101_21#_M1014_g N_C_c_311_n 0.0268586f $X=1.87 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_101_21#_c_184_n N_C_c_311_n 0.00650163f $X=2 $Y=1.875 $X2=0 $Y2=0
cc_178 N_A_101_21#_c_196_p N_C_c_311_n 0.0125297f $X=2.43 $Y=1.96 $X2=0 $Y2=0
cc_179 N_A_101_21#_c_185_n N_C_c_311_n 0.00658715f $X=2.515 $Y=2.235 $X2=0 $Y2=0
cc_180 N_A_101_21#_c_186_n N_C_c_311_n 0.00614426f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_181 N_A_101_21#_c_187_n N_C_M1011_g 0.0100647f $X=3.645 $Y=2.32 $X2=0 $Y2=0
cc_182 N_A_101_21#_c_200_p N_C_c_307_n 0.00628162f $X=3.72 $Y=0.37 $X2=0 $Y2=0
cc_183 N_A_101_21#_c_179_n N_C_c_307_n 0.00499109f $X=3.45 $Y=0.355 $X2=0 $Y2=0
cc_184 N_A_101_21#_c_175_n N_C_c_308_n 0.00157017f $X=2 $Y=1.325 $X2=0 $Y2=0
cc_185 N_A_101_21#_c_178_n N_C_c_308_n 0.0240529f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_101_21#_c_179_n N_C_c_309_n 0.00982945f $X=3.45 $Y=0.355 $X2=0 $Y2=0
cc_187 N_A_101_21#_c_179_n C 0.00344638f $X=3.45 $Y=0.355 $X2=0 $Y2=0
cc_188 N_A_101_21#_c_196_p N_A_492_93#_M1025_d 0.00409968f $X=2.43 $Y=1.96 $X2=0
+ $Y2=0
cc_189 N_A_101_21#_c_185_n N_A_492_93#_M1025_d 0.00259246f $X=2.515 $Y=2.235
+ $X2=0 $Y2=0
cc_190 N_A_101_21#_c_187_n N_A_492_93#_c_374_n 0.0118274f $X=3.645 $Y=2.32 $X2=0
+ $Y2=0
cc_191 N_A_101_21#_c_184_n N_A_492_93#_c_384_n 0.010447f $X=2 $Y=1.875 $X2=0
+ $Y2=0
cc_192 N_A_101_21#_c_191_p N_A_492_93#_c_384_n 0.00345572f $X=2.315 $Y=0.78
+ $X2=0 $Y2=0
cc_193 N_A_101_21#_c_196_p N_A_492_93#_c_384_n 0.0165826f $X=2.43 $Y=1.96 $X2=0
+ $Y2=0
cc_194 N_A_101_21#_c_187_n N_A_492_93#_c_384_n 0.00176797f $X=3.645 $Y=2.32
+ $X2=0 $Y2=0
cc_195 N_A_101_21#_c_175_n N_A_492_93#_c_370_n 0.0125392f $X=2 $Y=1.325 $X2=0
+ $Y2=0
cc_196 N_A_101_21#_c_184_n N_A_492_93#_c_370_n 0.00659166f $X=2 $Y=1.875 $X2=0
+ $Y2=0
cc_197 N_A_101_21#_c_178_n N_A_492_93#_c_370_n 7.97535e-19 $X=1.965 $Y=1.16
+ $X2=0 $Y2=0
cc_198 N_A_101_21#_c_179_n N_A_492_93#_c_370_n 0.0130244f $X=3.45 $Y=0.355 $X2=0
+ $Y2=0
cc_199 N_A_101_21#_M1011_d N_A_492_93#_c_376_n 0.00757366f $X=3.51 $Y=1.625
+ $X2=0 $Y2=0
cc_200 N_A_101_21#_c_187_n N_A_492_93#_c_376_n 0.0039224f $X=3.645 $Y=2.32 $X2=0
+ $Y2=0
cc_201 N_A_101_21#_M1011_d N_A_492_93#_c_377_n 5.89264e-19 $X=3.51 $Y=1.625
+ $X2=0 $Y2=0
cc_202 N_A_101_21#_c_187_n N_A_492_93#_c_378_n 0.00633062f $X=3.645 $Y=2.32
+ $X2=0 $Y2=0
cc_203 N_A_101_21#_c_200_p N_A_492_93#_c_373_n 0.00356056f $X=3.72 $Y=0.37 $X2=0
+ $Y2=0
cc_204 N_A_101_21#_c_184_n N_VPWR_M1014_d 0.00437587f $X=2 $Y=1.875 $X2=0 $Y2=0
cc_205 N_A_101_21#_c_196_p N_VPWR_M1014_d 0.00778804f $X=2.43 $Y=1.96 $X2=0
+ $Y2=0
cc_206 N_A_101_21#_c_224_p N_VPWR_M1014_d 8.79014e-19 $X=2.085 $Y=1.96 $X2=0
+ $Y2=0
cc_207 N_A_101_21#_M1001_g N_VPWR_c_915_n 0.00316354f $X=0.58 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_101_21#_M1001_g N_VPWR_c_916_n 0.00542953f $X=0.58 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_101_21#_M1002_g N_VPWR_c_916_n 0.00542953f $X=1 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_101_21#_M1002_g N_VPWR_c_917_n 0.00150929f $X=1 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_101_21#_M1005_g N_VPWR_c_917_n 0.00403828f $X=1.45 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_101_21#_c_178_n N_VPWR_c_917_n 0.00287436f $X=1.965 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A_101_21#_M1005_g N_VPWR_c_918_n 4.92168e-19 $X=1.45 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_101_21#_M1014_g N_VPWR_c_918_n 0.00842366f $X=1.87 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_101_21#_c_196_p N_VPWR_c_918_n 0.0126548f $X=2.43 $Y=1.96 $X2=0 $Y2=0
cc_216 N_A_101_21#_c_224_p N_VPWR_c_918_n 0.00931978f $X=2.085 $Y=1.96 $X2=0
+ $Y2=0
cc_217 N_A_101_21#_c_185_n N_VPWR_c_918_n 0.00141608f $X=2.515 $Y=2.235 $X2=0
+ $Y2=0
cc_218 N_A_101_21#_c_186_n N_VPWR_c_918_n 0.0136738f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_219 N_A_101_21#_M1005_g N_VPWR_c_923_n 0.00495816f $X=1.45 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_101_21#_M1014_g N_VPWR_c_923_n 0.0046653f $X=1.87 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_101_21#_c_196_p N_VPWR_c_924_n 0.00232824f $X=2.43 $Y=1.96 $X2=0
+ $Y2=0
cc_222 N_A_101_21#_c_186_n N_VPWR_c_924_n 0.00857493f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_223 N_A_101_21#_c_187_n N_VPWR_c_924_n 0.0575132f $X=3.645 $Y=2.32 $X2=0
+ $Y2=0
cc_224 N_A_101_21#_M1001_g N_VPWR_c_914_n 0.0105485f $X=0.58 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_101_21#_M1002_g N_VPWR_c_914_n 0.00958191f $X=1 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_101_21#_M1005_g N_VPWR_c_914_n 0.0085449f $X=1.45 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_101_21#_M1014_g N_VPWR_c_914_n 0.00789179f $X=1.87 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_101_21#_c_196_p N_VPWR_c_914_n 0.00552493f $X=2.43 $Y=1.96 $X2=0
+ $Y2=0
cc_229 N_A_101_21#_c_224_p N_VPWR_c_914_n 7.79838e-19 $X=2.085 $Y=1.96 $X2=0
+ $Y2=0
cc_230 N_A_101_21#_c_186_n N_VPWR_c_914_n 0.00627734f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_231 N_A_101_21#_c_187_n N_VPWR_c_914_n 0.0456534f $X=3.645 $Y=2.32 $X2=0
+ $Y2=0
cc_232 N_A_101_21#_c_171_n N_X_c_1028_n 0.0174388f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_101_21#_c_172_n N_X_c_1028_n 0.00193928f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_101_21#_M1001_g N_X_c_1033_n 0.0195882f $X=0.58 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_101_21#_M1002_g N_X_c_1033_n 0.0148433f $X=1 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_101_21#_M1005_g N_X_c_1033_n 7.32103e-19 $X=1.45 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_101_21#_c_178_n N_X_c_1036_n 0.0513174f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_101_21#_c_172_n N_X_c_1037_n 2.55752e-19 $X=1 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_101_21#_c_173_n N_X_c_1037_n 0.00640074f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_101_21#_c_178_n N_X_c_1039_n 0.0334941f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_101_21#_c_172_n N_X_c_1029_n 6.20832e-19 $X=1 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_101_21#_M1002_g N_X_c_1029_n 5.35663e-19 $X=1 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_101_21#_c_173_n N_X_c_1029_n 0.00560877f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_101_21#_M1005_g N_X_c_1029_n 0.00569082f $X=1.45 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_101_21#_c_174_n N_X_c_1029_n 0.00118116f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_101_21#_M1014_g N_X_c_1029_n 0.00114867f $X=1.87 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_101_21#_c_175_n N_X_c_1029_n 0.0363044f $X=2 $Y=1.325 $X2=0 $Y2=0
cc_248 N_A_101_21#_c_184_n N_X_c_1029_n 0.0139297f $X=2 $Y=1.875 $X2=0 $Y2=0
cc_249 N_A_101_21#_c_178_n N_X_c_1029_n 0.0165705f $X=1.965 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_101_21#_M1005_g N_X_c_1049_n 0.0115506f $X=1.45 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A_101_21#_c_187_n N_A_607_325#_M1011_s 0.00705836f $X=3.645 $Y=2.32
+ $X2=0 $Y2=0
cc_252 N_A_101_21#_M1011_d N_A_607_325#_c_1073_n 0.00468683f $X=3.51 $Y=1.625
+ $X2=0 $Y2=0
cc_253 N_A_101_21#_c_196_p N_A_607_325#_c_1073_n 0.00832414f $X=2.43 $Y=1.96
+ $X2=0 $Y2=0
cc_254 N_A_101_21#_c_185_n N_A_607_325#_c_1073_n 9.41079e-19 $X=2.515 $Y=2.235
+ $X2=0 $Y2=0
cc_255 N_A_101_21#_c_187_n N_A_607_325#_c_1073_n 0.0537701f $X=3.645 $Y=2.32
+ $X2=0 $Y2=0
cc_256 N_A_101_21#_c_179_n N_A_631_49#_M1024_s 0.0050721f $X=3.45 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_257 N_A_101_21#_M1024_d N_A_631_49#_c_1228_n 0.00636386f $X=3.575 $Y=0.245
+ $X2=0 $Y2=0
cc_258 N_A_101_21#_c_200_p N_A_631_49#_c_1218_n 0.0217348f $X=3.72 $Y=0.37 $X2=0
+ $Y2=0
cc_259 N_A_101_21#_c_179_n N_A_631_49#_c_1218_n 0.0164657f $X=3.45 $Y=0.355
+ $X2=0 $Y2=0
cc_260 N_A_101_21#_c_175_n N_VGND_M1027_d 0.00139163f $X=2 $Y=1.325 $X2=0 $Y2=0
cc_261 N_A_101_21#_c_191_p N_VGND_M1027_d 0.00877172f $X=2.315 $Y=0.78 $X2=0
+ $Y2=0
cc_262 N_A_101_21#_c_171_n N_VGND_c_1412_n 0.00565425f $X=0.58 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A_101_21#_c_171_n N_VGND_c_1413_n 0.00545968f $X=0.58 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_101_21#_c_172_n N_VGND_c_1413_n 0.00585385f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_101_21#_c_172_n N_VGND_c_1414_n 0.00202947f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_101_21#_c_173_n N_VGND_c_1414_n 0.00386709f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_101_21#_c_178_n N_VGND_c_1414_n 0.00221658f $X=1.965 $Y=1.16 $X2=0
+ $Y2=0
cc_268 N_A_101_21#_c_173_n N_VGND_c_1415_n 8.65536e-19 $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_101_21#_c_174_n N_VGND_c_1415_n 0.00935425f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A_101_21#_c_175_n N_VGND_c_1415_n 0.0104852f $X=2 $Y=1.325 $X2=0 $Y2=0
cc_271 N_A_101_21#_c_191_p N_VGND_c_1415_n 0.0045481f $X=2.315 $Y=0.78 $X2=0
+ $Y2=0
cc_272 N_A_101_21#_c_176_n N_VGND_c_1415_n 0.00720258f $X=2.4 $Y=0.695 $X2=0
+ $Y2=0
cc_273 N_A_101_21#_c_177_n N_VGND_c_1415_n 0.0140928f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_274 N_A_101_21#_c_178_n N_VGND_c_1415_n 5.56374e-19 $X=1.965 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_101_21#_c_191_p N_VGND_c_1420_n 0.00219715f $X=2.315 $Y=0.78 $X2=0
+ $Y2=0
cc_276 N_A_101_21#_c_177_n N_VGND_c_1420_n 0.0120884f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_277 N_A_101_21#_c_179_n N_VGND_c_1420_n 0.0844231f $X=3.45 $Y=0.355 $X2=0
+ $Y2=0
cc_278 N_A_101_21#_c_173_n N_VGND_c_1424_n 0.00531141f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_101_21#_c_174_n N_VGND_c_1424_n 0.0046653f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_101_21#_c_171_n N_VGND_c_1426_n 0.010718f $X=0.58 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_101_21#_c_172_n N_VGND_c_1426_n 0.010716f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_101_21#_c_173_n N_VGND_c_1426_n 0.00931445f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_101_21#_c_174_n N_VGND_c_1426_n 0.00796766f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_101_21#_c_175_n N_VGND_c_1426_n 7.88478e-19 $X=2 $Y=1.325 $X2=0 $Y2=0
cc_285 N_A_101_21#_c_191_p N_VGND_c_1426_n 0.00486078f $X=2.315 $Y=0.78 $X2=0
+ $Y2=0
cc_286 N_A_101_21#_c_177_n N_VGND_c_1426_n 0.00652842f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_287 N_A_101_21#_c_179_n N_VGND_c_1426_n 0.0514035f $X=3.45 $Y=0.355 $X2=0
+ $Y2=0
cc_288 N_C_M1011_g N_A_492_93#_c_374_n 0.037701f $X=3.435 $Y=2.045 $X2=0 $Y2=0
cc_289 N_C_c_310_n N_A_492_93#_c_374_n 0.00128239f $X=3.467 $Y=1.175 $X2=0 $Y2=0
cc_290 N_C_c_311_n N_A_492_93#_c_384_n 0.00939901f $X=2.385 $Y=1.325 $X2=0 $Y2=0
cc_291 N_C_c_309_n N_A_492_93#_c_384_n 0.00376155f $X=3.36 $Y=1.16 $X2=0 $Y2=0
cc_292 N_C_c_306_n N_A_492_93#_c_370_n 0.0047097f $X=2.385 $Y=0.995 $X2=0 $Y2=0
cc_293 N_C_c_311_n N_A_492_93#_c_370_n 0.00386891f $X=2.385 $Y=1.325 $X2=0 $Y2=0
cc_294 N_C_c_307_n N_A_492_93#_c_370_n 0.00249399f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C_c_309_n N_A_492_93#_c_370_n 0.0260984f $X=3.36 $Y=1.16 $X2=0 $Y2=0
cc_296 N_C_c_310_n N_A_492_93#_c_370_n 0.00491617f $X=3.467 $Y=1.175 $X2=0 $Y2=0
cc_297 C N_A_492_93#_c_370_n 0.0186011f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_298 N_C_M1011_g N_A_492_93#_c_376_n 0.0131528f $X=3.435 $Y=2.045 $X2=0 $Y2=0
cc_299 N_C_c_309_n N_A_492_93#_c_376_n 0.0121053f $X=3.36 $Y=1.16 $X2=0 $Y2=0
cc_300 N_C_c_310_n N_A_492_93#_c_376_n 0.00194181f $X=3.467 $Y=1.175 $X2=0 $Y2=0
cc_301 C N_A_492_93#_c_376_n 0.0348885f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_302 N_C_M1011_g N_A_492_93#_c_377_n 0.00357789f $X=3.435 $Y=2.045 $X2=0 $Y2=0
cc_303 N_C_c_310_n N_A_492_93#_c_377_n 6.37129e-19 $X=3.467 $Y=1.175 $X2=0 $Y2=0
cc_304 N_C_c_310_n N_A_492_93#_c_371_n 0.00344688f $X=3.467 $Y=1.175 $X2=0 $Y2=0
cc_305 C N_A_492_93#_c_371_n 0.0203401f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_306 N_C_c_310_n N_A_492_93#_c_372_n 0.0218135f $X=3.467 $Y=1.175 $X2=0 $Y2=0
cc_307 C N_A_492_93#_c_372_n 2.69217e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_308 N_C_c_307_n N_A_492_93#_c_373_n 0.0255134f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_309 N_C_c_311_n N_VPWR_c_918_n 0.00191684f $X=2.385 $Y=1.325 $X2=0 $Y2=0
cc_310 N_C_c_311_n N_VPWR_c_924_n 0.00403219f $X=2.385 $Y=1.325 $X2=0 $Y2=0
cc_311 N_C_M1011_g N_VPWR_c_924_n 0.00356303f $X=3.435 $Y=2.045 $X2=0 $Y2=0
cc_312 N_C_c_311_n N_VPWR_c_914_n 0.00522107f $X=2.385 $Y=1.325 $X2=0 $Y2=0
cc_313 N_C_M1011_g N_VPWR_c_914_n 0.00707416f $X=3.435 $Y=2.045 $X2=0 $Y2=0
cc_314 N_C_c_311_n N_A_607_325#_c_1073_n 9.60045e-19 $X=2.385 $Y=1.325 $X2=0
+ $Y2=0
cc_315 N_C_M1011_g N_A_607_325#_c_1073_n 0.00880042f $X=3.435 $Y=2.045 $X2=0
+ $Y2=0
cc_316 N_C_c_307_n N_A_631_49#_c_1228_n 0.00557156f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_317 C N_A_631_49#_c_1228_n 0.00255562f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_318 N_C_c_307_n N_A_631_49#_c_1218_n 0.00640201f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_319 N_C_c_309_n N_A_631_49#_c_1218_n 0.0055213f $X=3.36 $Y=1.16 $X2=0 $Y2=0
cc_320 C N_A_631_49#_c_1218_n 0.0287341f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_321 N_C_c_306_n N_VGND_c_1415_n 0.00130576f $X=2.385 $Y=0.995 $X2=0 $Y2=0
cc_322 N_C_c_306_n N_VGND_c_1420_n 8.79444e-19 $X=2.385 $Y=0.995 $X2=0 $Y2=0
cc_323 N_C_c_307_n N_VGND_c_1420_n 0.00357877f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_324 N_C_c_307_n N_VGND_c_1426_n 0.00671982f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_492_93#_c_374_n N_VPWR_c_919_n 0.0062797f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_326 N_A_492_93#_c_374_n N_VPWR_c_924_n 0.00338202f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_327 N_A_492_93#_c_374_n N_VPWR_c_914_n 0.00503145f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_328 N_A_492_93#_c_376_n N_A_607_325#_M1011_s 0.00362749f $X=3.73 $Y=1.62
+ $X2=0 $Y2=0
cc_329 N_A_492_93#_c_374_n N_A_607_325#_c_1073_n 0.01487f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_330 N_A_492_93#_c_376_n N_A_607_325#_c_1073_n 0.0523983f $X=3.73 $Y=1.62
+ $X2=0 $Y2=0
cc_331 N_A_492_93#_c_371_n N_A_607_325#_c_1073_n 0.00267573f $X=3.92 $Y=1.16
+ $X2=0 $Y2=0
cc_332 N_A_492_93#_c_372_n N_A_607_325#_c_1073_n 0.00101141f $X=3.92 $Y=1.16
+ $X2=0 $Y2=0
cc_333 N_A_492_93#_c_373_n N_A_607_325#_c_1068_n 0.00496015f $X=3.92 $Y=0.995
+ $X2=0 $Y2=0
cc_334 N_A_492_93#_c_374_n N_A_607_325#_c_1069_n 0.00456667f $X=3.92 $Y=1.325
+ $X2=0 $Y2=0
cc_335 N_A_492_93#_c_371_n N_A_631_49#_c_1228_n 0.0159681f $X=3.92 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_492_93#_c_372_n N_A_631_49#_c_1228_n 0.00169817f $X=3.92 $Y=1.16
+ $X2=0 $Y2=0
cc_337 N_A_492_93#_c_373_n N_A_631_49#_c_1228_n 0.0135605f $X=3.92 $Y=0.995
+ $X2=0 $Y2=0
cc_338 N_A_492_93#_c_374_n N_A_631_49#_c_1216_n 9.82177e-19 $X=3.92 $Y=1.325
+ $X2=0 $Y2=0
cc_339 N_A_492_93#_c_377_n N_A_631_49#_c_1216_n 0.00244972f $X=3.815 $Y=1.535
+ $X2=0 $Y2=0
cc_340 N_A_492_93#_c_371_n N_A_631_49#_c_1216_n 0.0244326f $X=3.92 $Y=1.16 $X2=0
+ $Y2=0
cc_341 N_A_492_93#_c_372_n N_A_631_49#_c_1216_n 0.00755993f $X=3.92 $Y=1.16
+ $X2=0 $Y2=0
cc_342 N_A_492_93#_c_373_n N_A_631_49#_c_1216_n 0.00577619f $X=3.92 $Y=0.995
+ $X2=0 $Y2=0
cc_343 N_A_492_93#_c_370_n N_A_631_49#_c_1218_n 0.0151382f $X=2.74 $Y=0.76 $X2=0
+ $Y2=0
cc_344 N_A_492_93#_c_373_n N_A_631_49#_c_1218_n 3.80178e-19 $X=3.92 $Y=0.995
+ $X2=0 $Y2=0
cc_345 N_A_492_93#_c_376_n N_A_631_49#_c_1224_n 5.8448e-19 $X=3.73 $Y=1.62 $X2=0
+ $Y2=0
cc_346 N_A_492_93#_c_377_n N_A_631_49#_c_1224_n 6.69003e-19 $X=3.815 $Y=1.535
+ $X2=0 $Y2=0
cc_347 N_A_492_93#_c_374_n N_A_631_49#_c_1225_n 0.006802f $X=3.92 $Y=1.325 $X2=0
+ $Y2=0
cc_348 N_A_492_93#_c_376_n N_A_631_49#_c_1225_n 0.0128201f $X=3.73 $Y=1.62 $X2=0
+ $Y2=0
cc_349 N_A_492_93#_c_377_n N_A_631_49#_c_1225_n 0.00775472f $X=3.815 $Y=1.535
+ $X2=0 $Y2=0
cc_350 N_A_492_93#_c_373_n N_VGND_c_1420_n 0.00414846f $X=3.92 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_492_93#_c_373_n N_VGND_c_1426_n 0.00723015f $X=3.92 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_1011_297#_c_463_n N_B_M1000_g 0.00527651f $X=5.325 $Y=1.58 $X2=0
+ $Y2=0
cc_353 N_A_1011_297#_c_458_n N_B_M1000_g 0.00474255f $X=5.36 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_1011_297#_c_467_p N_B_M1003_g 0.00371061f $X=5.435 $Y=0.85 $X2=0
+ $Y2=0
cc_355 N_A_1011_297#_c_458_n N_B_M1003_g 0.0140872f $X=5.36 $Y=0.74 $X2=0 $Y2=0
cc_356 N_A_1011_297#_c_452_n N_B_c_616_n 0.00436054f $X=6.525 $Y=0.85 $X2=0
+ $Y2=0
cc_357 N_A_1011_297#_c_458_n N_B_c_616_n 0.0122528f $X=5.36 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A_1011_297#_c_463_n N_B_c_617_n 0.00356061f $X=5.325 $Y=1.58 $X2=0
+ $Y2=0
cc_359 N_A_1011_297#_c_458_n N_B_c_617_n 0.00332114f $X=5.36 $Y=0.74 $X2=0 $Y2=0
cc_360 N_A_1011_297#_M1021_g N_B_M1007_g 0.0115983f $X=6.835 $Y=0.455 $X2=0
+ $Y2=0
cc_361 N_A_1011_297#_c_449_n N_B_M1007_g 0.0209917f $X=6.76 $Y=1.16 $X2=0 $Y2=0
cc_362 N_A_1011_297#_c_451_n N_B_M1007_g 0.00168544f $X=6.65 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_1011_297#_c_452_n N_B_M1007_g 6.73737e-19 $X=6.525 $Y=0.85 $X2=0
+ $Y2=0
cc_364 N_A_1011_297#_c_454_n N_B_M1007_g 6.65705e-19 $X=6.815 $Y=0.85 $X2=0
+ $Y2=0
cc_365 N_A_1011_297#_c_455_n N_B_M1007_g 0.0011633f $X=6.67 $Y=0.85 $X2=0 $Y2=0
cc_366 N_A_1011_297#_M1019_g N_B_M1018_g 0.0139116f $X=6.835 $Y=1.805 $X2=0
+ $Y2=0
cc_367 N_A_1011_297#_M1019_g N_B_c_626_n 0.00881703f $X=6.835 $Y=1.805 $X2=0
+ $Y2=0
cc_368 N_A_1011_297#_M1008_g N_B_M1013_g 0.0403239f $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_369 N_A_1011_297#_c_446_n N_B_c_621_n 0.00114568f $X=8.225 $Y=1.28 $X2=0
+ $Y2=0
cc_370 N_A_1011_297#_c_453_n N_B_c_621_n 0.00555012f $X=7.905 $Y=0.85 $X2=0
+ $Y2=0
cc_371 N_A_1011_297#_c_457_n N_B_c_621_n 0.0211354f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_372 N_A_1011_297#_c_446_n N_B_c_622_n 0.0189136f $X=8.225 $Y=1.28 $X2=0 $Y2=0
cc_373 N_A_1011_297#_c_450_n N_B_c_622_n 0.00771227f $X=6.835 $Y=1.16 $X2=0
+ $Y2=0
cc_374 N_A_1011_297#_c_453_n N_B_c_622_n 0.00134545f $X=7.905 $Y=0.85 $X2=0
+ $Y2=0
cc_375 N_A_1011_297#_c_457_n N_B_c_622_n 0.00169113f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_376 N_A_1011_297#_c_446_n B 8.1069e-19 $X=8.225 $Y=1.28 $X2=0 $Y2=0
cc_377 N_A_1011_297#_M1008_g B 0.00593518f $X=8.225 $Y=2.065 $X2=0 $Y2=0
cc_378 N_A_1011_297#_c_453_n B 0.00414594f $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_379 N_A_1011_297#_c_456_n B 0.00235209f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_380 N_A_1011_297#_c_457_n B 0.0183366f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_381 N_A_1011_297#_M1021_g N_B_c_623_n 0.00771227f $X=6.835 $Y=0.455 $X2=0
+ $Y2=0
cc_382 N_A_1011_297#_c_446_n N_B_c_623_n 0.00163786f $X=8.225 $Y=1.28 $X2=0
+ $Y2=0
cc_383 N_A_1011_297#_c_448_n N_B_c_623_n 0.0180222f $X=8.23 $Y=0.945 $X2=0 $Y2=0
cc_384 N_A_1011_297#_c_453_n N_B_c_623_n 0.00749482f $X=7.905 $Y=0.85 $X2=0
+ $Y2=0
cc_385 N_A_1011_297#_c_456_n N_B_c_623_n 0.00142159f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_386 N_A_1011_297#_c_457_n N_B_c_623_n 0.00206701f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_387 N_A_1011_297#_M1008_g N_A_M1017_g 0.0404776f $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_388 N_A_1011_297#_c_446_n N_A_c_735_n 0.0176934f $X=8.225 $Y=1.28 $X2=0 $Y2=0
cc_389 N_A_1011_297#_M1008_g N_A_c_735_n 0.00255062f $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_390 N_A_1011_297#_c_457_n N_A_c_735_n 7.00021e-19 $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_391 N_A_1011_297#_c_446_n N_A_c_736_n 0.00129629f $X=8.225 $Y=1.28 $X2=0
+ $Y2=0
cc_392 N_A_1011_297#_M1008_g N_A_c_736_n 5.31842e-19 $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_393 N_A_1011_297#_c_457_n N_A_c_736_n 0.016109f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_394 N_A_1011_297#_c_448_n N_A_c_737_n 0.0225442f $X=8.23 $Y=0.945 $X2=0 $Y2=0
cc_395 N_A_1011_297#_c_457_n N_A_c_737_n 2.68453e-19 $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_396 N_A_1011_297#_c_452_n N_A_1117_297#_M1007_s 8.53241e-19 $X=6.525 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_397 N_A_1011_297#_c_463_n N_A_1117_297#_c_780_n 0.0192437f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_398 N_A_1011_297#_c_452_n N_A_1117_297#_c_780_n 0.0124002f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_399 N_A_1011_297#_c_467_p N_A_1117_297#_c_780_n 6.57905e-19 $X=5.435 $Y=0.85
+ $X2=0 $Y2=0
cc_400 N_A_1011_297#_c_458_n N_A_1117_297#_c_780_n 0.0595696f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_401 N_A_1011_297#_M1008_g N_A_1117_297#_c_789_n 0.00235326f $X=8.225 $Y=2.065
+ $X2=0 $Y2=0
cc_402 N_A_1011_297#_c_448_n N_A_1117_297#_c_782_n 0.00164439f $X=8.23 $Y=0.945
+ $X2=0 $Y2=0
cc_403 N_A_1011_297#_c_456_n N_A_1117_297#_c_782_n 0.00485657f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_1011_297#_c_457_n N_A_1117_297#_c_782_n 0.00616889f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_405 N_A_1011_297#_M1021_g N_A_1117_297#_c_802_n 0.00602131f $X=6.835 $Y=0.455
+ $X2=0 $Y2=0
cc_406 N_A_1011_297#_c_448_n N_A_1117_297#_c_802_n 0.00716191f $X=8.23 $Y=0.945
+ $X2=0 $Y2=0
cc_407 N_A_1011_297#_c_451_n N_A_1117_297#_c_802_n 3.69046e-19 $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_408 N_A_1011_297#_c_452_n N_A_1117_297#_c_802_n 0.0490335f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_409 N_A_1011_297#_c_453_n N_A_1117_297#_c_802_n 0.0873524f $X=7.905 $Y=0.85
+ $X2=0 $Y2=0
cc_410 N_A_1011_297#_c_454_n N_A_1117_297#_c_802_n 0.0265516f $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_411 N_A_1011_297#_c_455_n N_A_1117_297#_c_802_n 0.00311774f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_412 N_A_1011_297#_c_456_n N_A_1117_297#_c_802_n 0.0265508f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_413 N_A_1011_297#_c_457_n N_A_1117_297#_c_802_n 0.00472786f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_414 N_A_1011_297#_c_452_n N_A_1117_297#_c_785_n 0.0261258f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_415 N_A_1011_297#_c_458_n N_A_1117_297#_c_785_n 0.00680928f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_416 N_A_1011_297#_c_452_n N_A_1117_297#_c_786_n 0.00110657f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_1011_297#_c_458_n N_A_1117_297#_c_786_n 0.0113597f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_418 N_A_1011_297#_c_448_n N_A_1117_297#_c_815_n 0.00153367f $X=8.23 $Y=0.945
+ $X2=0 $Y2=0
cc_419 N_A_1011_297#_c_448_n N_A_1117_297#_c_816_n 0.0077529f $X=8.23 $Y=0.945
+ $X2=0 $Y2=0
cc_420 N_A_1011_297#_M1008_g N_VPWR_c_920_n 0.00128985f $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_421 N_A_1011_297#_M1008_g N_VPWR_c_925_n 0.00362032f $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_422 N_A_1011_297#_M1000_d N_VPWR_c_914_n 0.00294931f $X=5.055 $Y=1.485 $X2=0
+ $Y2=0
cc_423 N_A_1011_297#_M1008_g N_VPWR_c_914_n 0.00570414f $X=8.225 $Y=2.065 $X2=0
+ $Y2=0
cc_424 N_A_1011_297#_c_452_n N_A_607_325#_M1007_d 0.00134889f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_425 N_A_1011_297#_c_454_n N_A_607_325#_M1007_d 5.4759e-19 $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_426 N_A_1011_297#_c_455_n N_A_607_325#_M1007_d 0.00561877f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_427 N_A_1011_297#_c_467_p N_A_607_325#_c_1068_n 0.00245527f $X=5.435 $Y=0.85
+ $X2=0 $Y2=0
cc_428 N_A_1011_297#_c_458_n N_A_607_325#_c_1068_n 0.00390808f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_429 N_A_1011_297#_c_463_n N_A_607_325#_c_1069_n 0.0142896f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_430 N_A_1011_297#_c_458_n N_A_607_325#_c_1069_n 0.00993319f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_431 N_A_1011_297#_M1000_d N_A_607_325#_c_1075_n 0.00549845f $X=5.055 $Y=1.485
+ $X2=0 $Y2=0
cc_432 N_A_1011_297#_c_463_n N_A_607_325#_c_1075_n 0.025068f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_433 N_A_1011_297#_M1000_d N_A_607_325#_c_1076_n 0.00296992f $X=5.055 $Y=1.485
+ $X2=0 $Y2=0
cc_434 N_A_1011_297#_M1000_d N_A_607_325#_c_1078_n 0.00287797f $X=5.055 $Y=1.485
+ $X2=0 $Y2=0
cc_435 N_A_1011_297#_M1019_g N_A_607_325#_c_1070_n 0.0017846f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_436 N_A_1011_297#_c_449_n N_A_607_325#_c_1070_n 7.1162e-19 $X=6.76 $Y=1.16
+ $X2=0 $Y2=0
cc_437 N_A_1011_297#_c_451_n N_A_607_325#_c_1070_n 0.0190267f $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_438 N_A_1011_297#_c_452_n N_A_607_325#_c_1070_n 0.00612761f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_439 N_A_1011_297#_c_454_n N_A_607_325#_c_1070_n 0.00109225f $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_440 N_A_1011_297#_c_455_n N_A_607_325#_c_1070_n 0.00299076f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_441 N_A_1011_297#_M1019_g N_A_607_325#_c_1080_n 0.00215111f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_442 N_A_1011_297#_M1008_g N_A_607_325#_c_1080_n 0.00693683f $X=8.225 $Y=2.065
+ $X2=0 $Y2=0
cc_443 N_A_1011_297#_M1021_g N_A_607_325#_c_1116_n 0.002299f $X=6.835 $Y=0.455
+ $X2=0 $Y2=0
cc_444 N_A_1011_297#_c_455_n N_A_607_325#_c_1116_n 0.00180873f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_445 N_A_1011_297#_c_458_n N_A_607_325#_c_1071_n 0.0066474f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_446 N_A_1011_297#_c_449_n N_A_607_325#_c_1072_n 2.22283e-19 $X=6.76 $Y=1.16
+ $X2=0 $Y2=0
cc_447 N_A_1011_297#_c_451_n N_A_607_325#_c_1072_n 0.00299453f $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_448 N_A_1011_297#_c_452_n N_A_607_325#_c_1072_n 0.0153691f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_449 N_A_1011_297#_c_454_n N_A_607_325#_c_1072_n 0.00134329f $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_450 N_A_1011_297#_c_455_n N_A_607_325#_c_1072_n 0.0140693f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_451 N_A_1011_297#_c_453_n N_A_631_49#_M1023_d 0.00109392f $X=7.905 $Y=0.85
+ $X2=0 $Y2=0
cc_452 N_A_1011_297#_c_456_n N_A_631_49#_M1023_d 7.4435e-19 $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_453 N_A_1011_297#_c_457_n N_A_631_49#_M1023_d 0.00406077f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_454 N_A_1011_297#_c_449_n N_A_631_49#_c_1220_n 0.00881942f $X=6.76 $Y=1.16
+ $X2=0 $Y2=0
cc_455 N_A_1011_297#_c_451_n N_A_631_49#_c_1220_n 0.0271004f $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_456 N_A_1011_297#_c_452_n N_A_631_49#_c_1220_n 5.63647e-19 $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_457 N_A_1011_297#_M1019_g N_A_631_49#_c_1257_n 0.00366596f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_458 N_A_1011_297#_M1019_g N_A_631_49#_c_1221_n 0.0155406f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_459 N_A_1011_297#_c_449_n N_A_631_49#_c_1221_n 7.42472e-19 $X=6.76 $Y=1.16
+ $X2=0 $Y2=0
cc_460 N_A_1011_297#_c_451_n N_A_631_49#_c_1221_n 0.00152864f $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_461 N_A_1011_297#_c_453_n N_A_631_49#_c_1221_n 0.00288457f $X=7.905 $Y=0.85
+ $X2=0 $Y2=0
cc_462 N_A_1011_297#_c_454_n N_A_631_49#_c_1221_n 6.69145e-19 $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_463 N_A_1011_297#_M1021_g N_A_631_49#_c_1217_n 0.0170866f $X=6.835 $Y=0.455
+ $X2=0 $Y2=0
cc_464 N_A_1011_297#_c_451_n N_A_631_49#_c_1217_n 0.0210201f $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_465 N_A_1011_297#_c_453_n N_A_631_49#_c_1217_n 0.0170211f $X=7.905 $Y=0.85
+ $X2=0 $Y2=0
cc_466 N_A_1011_297#_c_454_n N_A_631_49#_c_1217_n 0.00240264f $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_467 N_A_1011_297#_c_455_n N_A_631_49#_c_1217_n 0.0233531f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_468 N_A_1011_297#_c_448_n N_A_631_49#_c_1268_n 0.00328526f $X=8.23 $Y=0.945
+ $X2=0 $Y2=0
cc_469 N_A_1011_297#_c_453_n N_A_631_49#_c_1268_n 0.00149151f $X=7.905 $Y=0.85
+ $X2=0 $Y2=0
cc_470 N_A_1011_297#_c_456_n N_A_631_49#_c_1268_n 3.55136e-19 $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_471 N_A_1011_297#_c_457_n N_A_631_49#_c_1268_n 0.00528249f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_472 N_A_1011_297#_c_463_n N_A_631_49#_c_1223_n 0.0241272f $X=5.325 $Y=1.58
+ $X2=0 $Y2=0
cc_473 N_A_1011_297#_c_451_n N_A_631_49#_c_1223_n 8.40027e-19 $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_474 N_A_1011_297#_c_452_n N_A_631_49#_c_1223_n 0.0483077f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_475 N_A_1011_297#_c_467_p N_A_631_49#_c_1223_n 0.0124731f $X=5.435 $Y=0.85
+ $X2=0 $Y2=0
cc_476 N_A_1011_297#_c_458_n N_A_631_49#_c_1223_n 0.00191712f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_477 N_A_1011_297#_M1019_g N_A_631_49#_c_1226_n 0.00414368f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_478 N_A_1011_297#_c_449_n N_A_631_49#_c_1226_n 0.00431105f $X=6.76 $Y=1.16
+ $X2=0 $Y2=0
cc_479 N_A_1011_297#_c_451_n N_A_631_49#_c_1226_n 0.00243787f $X=6.65 $Y=0.995
+ $X2=0 $Y2=0
cc_480 N_A_1011_297#_c_454_n N_A_631_49#_c_1226_n 0.0153734f $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_481 N_A_1011_297#_c_453_n N_A_1382_49#_M1021_d 0.00166227f $X=7.905 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_482 N_A_1011_297#_M1019_g N_A_1382_49#_c_1345_n 0.00785518f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_483 N_A_1011_297#_c_453_n N_A_1382_49#_c_1345_n 0.0179438f $X=7.905 $Y=0.85
+ $X2=0 $Y2=0
cc_484 N_A_1011_297#_c_456_n N_A_1382_49#_c_1345_n 0.00214961f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_485 N_A_1011_297#_c_457_n N_A_1382_49#_c_1345_n 0.00583126f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_486 N_A_1011_297#_M1019_g N_A_1382_49#_c_1357_n 0.00421122f $X=6.835 $Y=1.805
+ $X2=0 $Y2=0
cc_487 N_A_1011_297#_M1008_g N_A_1382_49#_c_1358_n 0.0138456f $X=8.225 $Y=2.065
+ $X2=0 $Y2=0
cc_488 N_A_1011_297#_c_457_n N_A_1382_49#_c_1358_n 0.00161448f $X=8.05 $Y=0.85
+ $X2=0 $Y2=0
cc_489 N_A_1011_297#_c_467_p N_VGND_c_1416_n 0.0038492f $X=5.435 $Y=0.85 $X2=0
+ $Y2=0
cc_490 N_A_1011_297#_M1021_g N_VGND_c_1422_n 0.00575161f $X=6.835 $Y=0.455 $X2=0
+ $Y2=0
cc_491 N_A_1011_297#_c_448_n N_VGND_c_1422_n 0.00585385f $X=8.23 $Y=0.945 $X2=0
+ $Y2=0
cc_492 N_A_1011_297#_c_455_n N_VGND_c_1422_n 0.00308387f $X=6.67 $Y=0.85 $X2=0
+ $Y2=0
cc_493 N_A_1011_297#_c_457_n N_VGND_c_1422_n 7.70543e-19 $X=8.05 $Y=0.85 $X2=0
+ $Y2=0
cc_494 N_A_1011_297#_c_458_n N_VGND_c_1422_n 0.0072215f $X=5.36 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A_1011_297#_M1003_d N_VGND_c_1426_n 0.00197536f $X=5.225 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_A_1011_297#_M1021_g N_VGND_c_1426_n 0.00662684f $X=6.835 $Y=0.455 $X2=0
+ $Y2=0
cc_497 N_A_1011_297#_c_448_n N_VGND_c_1426_n 0.00607914f $X=8.23 $Y=0.945 $X2=0
+ $Y2=0
cc_498 N_A_1011_297#_c_452_n N_VGND_c_1426_n 0.00895484f $X=6.525 $Y=0.85 $X2=0
+ $Y2=0
cc_499 N_A_1011_297#_c_467_p N_VGND_c_1426_n 0.0148686f $X=5.435 $Y=0.85 $X2=0
+ $Y2=0
cc_500 N_A_1011_297#_c_458_n N_VGND_c_1426_n 0.00376573f $X=5.36 $Y=0.74 $X2=0
+ $Y2=0
cc_501 B N_A_M1017_g 2.12214e-19 $X=7.965 $Y=1.445 $X2=0 $Y2=0
cc_502 N_B_c_621_n N_A_c_736_n 0.00135728f $X=7.69 $Y=1.16 $X2=0 $Y2=0
cc_503 N_B_M1000_g N_A_1117_297#_c_780_n 0.00403038f $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_504 N_B_M1003_g N_A_1117_297#_c_780_n 0.00120589f $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_505 N_B_c_616_n N_A_1117_297#_c_780_n 0.0145602f $X=6.005 $Y=1.16 $X2=0 $Y2=0
cc_506 N_B_M1007_g N_A_1117_297#_c_780_n 0.00392248f $X=6.08 $Y=0.565 $X2=0
+ $Y2=0
cc_507 N_B_M1018_g N_A_1117_297#_c_780_n 0.00549757f $X=6.08 $Y=1.905 $X2=0
+ $Y2=0
cc_508 B N_A_1117_297#_c_789_n 0.0103993f $X=7.965 $Y=1.445 $X2=0 $Y2=0
cc_509 N_B_M1007_g N_A_1117_297#_c_802_n 0.00167912f $X=6.08 $Y=0.565 $X2=0
+ $Y2=0
cc_510 N_B_c_623_n N_A_1117_297#_c_802_n 0.00325031f $X=7.69 $Y=0.995 $X2=0
+ $Y2=0
cc_511 N_B_M1003_g N_A_1117_297#_c_785_n 4.212e-19 $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_512 N_B_M1007_g N_A_1117_297#_c_785_n 9.44608e-19 $X=6.08 $Y=0.565 $X2=0
+ $Y2=0
cc_513 N_B_M1003_g N_A_1117_297#_c_786_n 0.00330428f $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_514 N_B_c_616_n N_A_1117_297#_c_786_n 0.00222258f $X=6.005 $Y=1.16 $X2=0
+ $Y2=0
cc_515 N_B_M1007_g N_A_1117_297#_c_786_n 0.00459791f $X=6.08 $Y=0.565 $X2=0
+ $Y2=0
cc_516 N_B_M1000_g N_VPWR_c_919_n 0.0112156f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_517 N_B_M1000_g N_VPWR_c_925_n 0.00341689f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_518 N_B_c_627_n N_VPWR_c_925_n 0.0380719f $X=6.155 $Y=2.54 $X2=0 $Y2=0
cc_519 N_B_M1000_g N_VPWR_c_914_n 0.00540327f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_520 N_B_c_626_n N_VPWR_c_914_n 0.0390811f $X=7.635 $Y=2.54 $X2=0 $Y2=0
cc_521 N_B_c_627_n N_VPWR_c_914_n 0.00592494f $X=6.155 $Y=2.54 $X2=0 $Y2=0
cc_522 N_B_M1003_g N_A_607_325#_c_1068_n 0.0032688f $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_523 N_B_c_617_n N_A_607_325#_c_1069_n 0.0176593f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_524 N_B_M1000_g N_A_607_325#_c_1075_n 0.0157597f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_525 N_B_M1000_g N_A_607_325#_c_1076_n 0.00631689f $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_526 N_B_M1018_g N_A_607_325#_c_1076_n 9.10003e-19 $X=6.08 $Y=1.905 $X2=0
+ $Y2=0
cc_527 N_B_M1000_g N_A_607_325#_c_1078_n 0.00361658f $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_528 N_B_c_616_n N_A_607_325#_c_1070_n 0.00258995f $X=6.005 $Y=1.16 $X2=0
+ $Y2=0
cc_529 N_B_M1007_g N_A_607_325#_c_1070_n 0.0066461f $X=6.08 $Y=0.565 $X2=0 $Y2=0
cc_530 N_B_M1018_g N_A_607_325#_c_1070_n 0.0375937f $X=6.08 $Y=1.905 $X2=0 $Y2=0
cc_531 N_B_c_620_n N_A_607_325#_c_1070_n 0.00263255f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_532 N_B_M1018_g N_A_607_325#_c_1080_n 0.00536892f $X=6.08 $Y=1.905 $X2=0
+ $Y2=0
cc_533 N_B_c_626_n N_A_607_325#_c_1080_n 0.0277284f $X=7.635 $Y=2.54 $X2=0 $Y2=0
cc_534 N_B_M1013_g N_A_607_325#_c_1080_n 0.0122992f $X=7.71 $Y=1.965 $X2=0 $Y2=0
cc_535 N_B_M1007_g N_A_607_325#_c_1116_n 5.19748e-19 $X=6.08 $Y=0.565 $X2=0
+ $Y2=0
cc_536 N_B_M1003_g N_A_607_325#_c_1071_n 9.36944e-19 $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_537 N_B_c_617_n N_A_607_325#_c_1071_n 0.00379336f $X=5.225 $Y=1.16 $X2=0
+ $Y2=0
cc_538 N_B_M1007_g N_A_607_325#_c_1072_n 0.0110389f $X=6.08 $Y=0.565 $X2=0 $Y2=0
cc_539 N_B_M1018_g N_A_607_325#_c_1082_n 0.00739846f $X=6.08 $Y=1.905 $X2=0
+ $Y2=0
cc_540 N_B_c_617_n N_A_631_49#_c_1216_n 4.44674e-19 $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_541 N_B_M1018_g N_A_631_49#_c_1220_n 0.00133974f $X=6.08 $Y=1.905 $X2=0 $Y2=0
cc_542 N_B_M1018_g N_A_631_49#_c_1257_n 0.00404484f $X=6.08 $Y=1.905 $X2=0 $Y2=0
cc_543 N_B_c_623_n N_A_631_49#_c_1217_n 0.0026019f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_544 N_B_c_621_n N_A_631_49#_c_1268_n 0.00216976f $X=7.69 $Y=1.16 $X2=0 $Y2=0
cc_545 N_B_c_622_n N_A_631_49#_c_1268_n 0.00134398f $X=7.69 $Y=1.16 $X2=0 $Y2=0
cc_546 N_B_c_623_n N_A_631_49#_c_1268_n 0.00498906f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_547 N_B_c_623_n N_A_631_49#_c_1288_n 0.00521263f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_548 N_B_M1000_g N_A_631_49#_c_1223_n 0.0049882f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_549 N_B_c_616_n N_A_631_49#_c_1223_n 0.0041572f $X=6.005 $Y=1.16 $X2=0 $Y2=0
cc_550 N_B_M1018_g N_A_631_49#_c_1223_n 0.00263877f $X=6.08 $Y=1.905 $X2=0 $Y2=0
cc_551 N_B_M1018_g N_A_631_49#_c_1226_n 4.43803e-19 $X=6.08 $Y=1.905 $X2=0 $Y2=0
cc_552 N_B_M1013_g N_A_1382_49#_c_1345_n 0.0107026f $X=7.71 $Y=1.965 $X2=0 $Y2=0
cc_553 N_B_c_621_n N_A_1382_49#_c_1345_n 0.0325983f $X=7.69 $Y=1.16 $X2=0 $Y2=0
cc_554 N_B_c_631_n N_A_1382_49#_c_1345_n 0.0141708f $X=7.775 $Y=1.53 $X2=0 $Y2=0
cc_555 N_B_c_623_n N_A_1382_49#_c_1345_n 0.0103225f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_556 N_B_M1013_g N_A_1382_49#_c_1358_n 0.0096343f $X=7.71 $Y=1.965 $X2=0 $Y2=0
cc_557 N_B_c_622_n N_A_1382_49#_c_1358_n 0.00103367f $X=7.69 $Y=1.16 $X2=0 $Y2=0
cc_558 N_B_c_631_n N_A_1382_49#_c_1358_n 0.00720786f $X=7.775 $Y=1.53 $X2=0
+ $Y2=0
cc_559 B N_A_1382_49#_c_1358_n 0.0164129f $X=7.965 $Y=1.445 $X2=0 $Y2=0
cc_560 N_B_M1003_g N_VGND_c_1416_n 0.00438629f $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_561 N_B_c_617_n N_VGND_c_1416_n 0.0053187f $X=5.225 $Y=1.16 $X2=0 $Y2=0
cc_562 N_B_M1003_g N_VGND_c_1422_n 0.00560495f $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_563 N_B_M1007_g N_VGND_c_1422_n 0.00414252f $X=6.08 $Y=0.565 $X2=0 $Y2=0
cc_564 N_B_c_623_n N_VGND_c_1422_n 0.00357877f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_565 N_B_M1003_g N_VGND_c_1426_n 0.0107857f $X=5.15 $Y=0.56 $X2=0 $Y2=0
cc_566 N_B_M1007_g N_VGND_c_1426_n 0.00707108f $X=6.08 $Y=0.565 $X2=0 $Y2=0
cc_567 N_B_c_623_n N_VGND_c_1426_n 0.00596272f $X=7.69 $Y=0.995 $X2=0 $Y2=0
cc_568 N_A_c_737_n N_A_1117_297#_c_779_n 0.0247826f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_569 N_A_M1017_g N_A_1117_297#_M1012_g 0.0453081f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_570 N_A_M1017_g N_A_1117_297#_c_789_n 0.00974519f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_571 N_A_c_735_n N_A_1117_297#_c_789_n 0.00302292f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_572 N_A_c_736_n N_A_1117_297#_c_789_n 0.0269201f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_573 N_A_c_736_n N_A_1117_297#_c_781_n 0.0106752f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_574 N_A_c_737_n N_A_1117_297#_c_781_n 0.00845772f $X=8.66 $Y=0.995 $X2=0
+ $Y2=0
cc_575 N_A_c_735_n N_A_1117_297#_c_782_n 0.00357599f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_576 N_A_c_736_n N_A_1117_297#_c_782_n 0.0204454f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_577 N_A_c_737_n N_A_1117_297#_c_782_n 0.00178341f $X=8.66 $Y=0.995 $X2=0
+ $Y2=0
cc_578 N_A_c_735_n N_A_1117_297#_c_783_n 7.09491e-19 $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_579 N_A_c_736_n N_A_1117_297#_c_783_n 0.0206309f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_580 N_A_c_737_n N_A_1117_297#_c_783_n 0.00347974f $X=8.66 $Y=0.995 $X2=0
+ $Y2=0
cc_581 N_A_M1017_g N_A_1117_297#_c_791_n 0.00333575f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_582 N_A_c_735_n N_A_1117_297#_c_784_n 0.0211645f $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_583 N_A_c_736_n N_A_1117_297#_c_784_n 8.25692e-19 $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_584 N_A_c_736_n N_A_1117_297#_c_815_n 9.51454e-19 $X=8.65 $Y=1.16 $X2=0 $Y2=0
cc_585 N_A_c_737_n N_A_1117_297#_c_816_n 0.00774108f $X=8.66 $Y=0.995 $X2=0
+ $Y2=0
cc_586 N_A_M1017_g N_VPWR_c_920_n 0.00873272f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_587 N_A_M1017_g N_VPWR_c_925_n 0.00337001f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_588 N_A_M1017_g N_VPWR_c_914_n 0.00417888f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_589 N_A_M1017_g N_A_607_325#_c_1080_n 0.00145186f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_590 N_A_M1017_g N_A_1382_49#_c_1358_n 0.0121115f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_591 N_A_M1017_g N_A_1382_49#_c_1351_n 3.59394e-19 $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_592 N_A_c_737_n N_VGND_c_1417_n 0.00268723f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_593 N_A_c_737_n N_VGND_c_1422_n 0.0042601f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_594 N_A_c_737_n N_VGND_c_1426_n 0.00602447f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_595 N_A_1117_297#_c_789_n N_VPWR_M1017_d 0.00452045f $X=9.005 $Y=1.6 $X2=0
+ $Y2=0
cc_596 N_A_1117_297#_M1012_g N_VPWR_c_920_n 0.00837913f $X=9.15 $Y=1.985 $X2=0
+ $Y2=0
cc_597 N_A_1117_297#_M1012_g N_VPWR_c_926_n 0.00322931f $X=9.15 $Y=1.985 $X2=0
+ $Y2=0
cc_598 N_A_1117_297#_M1008_d N_VPWR_c_914_n 0.00382772f $X=8.3 $Y=1.645 $X2=0
+ $Y2=0
cc_599 N_A_1117_297#_M1012_g N_VPWR_c_914_n 0.00475509f $X=9.15 $Y=1.985 $X2=0
+ $Y2=0
cc_600 N_A_1117_297#_c_802_n N_A_607_325#_M1007_d 0.00511495f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_601 N_A_1117_297#_c_780_n N_A_607_325#_c_1075_n 0.0132911f $X=5.71 $Y=1.94
+ $X2=0 $Y2=0
cc_602 N_A_1117_297#_c_780_n N_A_607_325#_c_1076_n 0.00274773f $X=5.71 $Y=1.94
+ $X2=0 $Y2=0
cc_603 N_A_1117_297#_M1018_s N_A_607_325#_c_1077_n 0.00987712f $X=5.585 $Y=1.485
+ $X2=0 $Y2=0
cc_604 N_A_1117_297#_c_780_n N_A_607_325#_c_1077_n 0.0128549f $X=5.71 $Y=1.94
+ $X2=0 $Y2=0
cc_605 N_A_1117_297#_c_780_n N_A_607_325#_c_1070_n 0.0675782f $X=5.71 $Y=1.94
+ $X2=0 $Y2=0
cc_606 N_A_1117_297#_M1008_d N_A_607_325#_c_1080_n 0.00239642f $X=8.3 $Y=1.645
+ $X2=0 $Y2=0
cc_607 N_A_1117_297#_c_802_n N_A_607_325#_c_1116_n 0.0121742f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_608 N_A_1117_297#_c_785_n N_A_607_325#_c_1116_n 0.00146594f $X=5.895 $Y=0.51
+ $X2=0 $Y2=0
cc_609 N_A_1117_297#_c_786_n N_A_607_325#_c_1116_n 0.0093757f $X=5.75 $Y=0.51
+ $X2=0 $Y2=0
cc_610 N_A_1117_297#_c_780_n N_A_607_325#_c_1072_n 0.0121907f $X=5.71 $Y=1.94
+ $X2=0 $Y2=0
cc_611 N_A_1117_297#_c_802_n N_A_607_325#_c_1072_n 0.00296668f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_612 N_A_1117_297#_c_786_n N_A_607_325#_c_1072_n 0.00198934f $X=5.75 $Y=0.51
+ $X2=0 $Y2=0
cc_613 N_A_1117_297#_c_802_n N_A_631_49#_M1023_d 0.00332817f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_614 N_A_1117_297#_c_802_n N_A_631_49#_c_1217_n 0.0145685f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_615 N_A_1117_297#_c_802_n N_A_631_49#_c_1268_n 0.0145995f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_616 N_A_1117_297#_c_815_n N_A_631_49#_c_1268_n 0.00126391f $X=8.51 $Y=0.51
+ $X2=0 $Y2=0
cc_617 N_A_1117_297#_c_816_n N_A_631_49#_c_1268_n 0.00765914f $X=8.51 $Y=0.51
+ $X2=0 $Y2=0
cc_618 N_A_1117_297#_c_802_n N_A_631_49#_c_1288_n 0.0119237f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_619 N_A_1117_297#_M1018_s N_A_631_49#_c_1223_n 0.00802537f $X=5.585 $Y=1.485
+ $X2=0 $Y2=0
cc_620 N_A_1117_297#_c_780_n N_A_631_49#_c_1223_n 0.0183124f $X=5.71 $Y=1.94
+ $X2=0 $Y2=0
cc_621 N_A_1117_297#_c_802_n N_A_1382_49#_M1021_d 0.00653094f $X=8.365 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_622 N_A_1117_297#_c_802_n N_A_1382_49#_c_1345_n 0.00162336f $X=8.365 $Y=0.51
+ $X2=0 $Y2=0
cc_623 N_A_1117_297#_c_779_n N_A_1382_49#_c_1346_n 0.00964261f $X=9.15 $Y=0.995
+ $X2=0 $Y2=0
cc_624 N_A_1117_297#_M1012_g N_A_1382_49#_c_1346_n 0.0113295f $X=9.15 $Y=1.985
+ $X2=0 $Y2=0
cc_625 N_A_1117_297#_c_789_n N_A_1382_49#_c_1346_n 0.0130585f $X=9.005 $Y=1.6
+ $X2=0 $Y2=0
cc_626 N_A_1117_297#_c_783_n N_A_1382_49#_c_1346_n 0.040001f $X=9.09 $Y=1.325
+ $X2=0 $Y2=0
cc_627 N_A_1117_297#_c_791_n N_A_1382_49#_c_1346_n 0.00963537f $X=9.09 $Y=1.495
+ $X2=0 $Y2=0
cc_628 N_A_1117_297#_c_784_n N_A_1382_49#_c_1346_n 0.00752814f $X=9.15 $Y=1.16
+ $X2=0 $Y2=0
cc_629 N_A_1117_297#_M1008_d N_A_1382_49#_c_1358_n 0.00689243f $X=8.3 $Y=1.645
+ $X2=0 $Y2=0
cc_630 N_A_1117_297#_M1012_g N_A_1382_49#_c_1358_n 0.00253441f $X=9.15 $Y=1.985
+ $X2=0 $Y2=0
cc_631 N_A_1117_297#_c_789_n N_A_1382_49#_c_1358_n 0.0324094f $X=9.005 $Y=1.6
+ $X2=0 $Y2=0
cc_632 N_A_1117_297#_M1012_g N_A_1382_49#_c_1351_n 0.0090064f $X=9.15 $Y=1.985
+ $X2=0 $Y2=0
cc_633 N_A_1117_297#_c_789_n N_A_1382_49#_c_1351_n 0.00661258f $X=9.005 $Y=1.6
+ $X2=0 $Y2=0
cc_634 N_A_1117_297#_c_783_n N_A_1382_49#_c_1351_n 0.00152532f $X=9.09 $Y=1.325
+ $X2=0 $Y2=0
cc_635 N_A_1117_297#_c_784_n N_A_1382_49#_c_1351_n 7.17833e-19 $X=9.15 $Y=1.16
+ $X2=0 $Y2=0
cc_636 N_A_1117_297#_c_784_n N_A_1382_49#_c_1347_n 2.03932e-19 $X=9.15 $Y=1.16
+ $X2=0 $Y2=0
cc_637 N_A_1117_297#_c_815_n N_A_1382_49#_c_1347_n 4.91816e-19 $X=8.51 $Y=0.51
+ $X2=0 $Y2=0
cc_638 N_A_1117_297#_c_781_n N_VGND_M1004_d 0.00147467f $X=9.005 $Y=0.82 $X2=0
+ $Y2=0
cc_639 N_A_1117_297#_c_785_n N_VGND_c_1416_n 7.58969e-19 $X=5.895 $Y=0.51 $X2=0
+ $Y2=0
cc_640 N_A_1117_297#_c_779_n N_VGND_c_1417_n 0.00268723f $X=9.15 $Y=0.995 $X2=0
+ $Y2=0
cc_641 N_A_1117_297#_c_781_n N_VGND_c_1417_n 0.0111874f $X=9.005 $Y=0.82 $X2=0
+ $Y2=0
cc_642 N_A_1117_297#_c_783_n N_VGND_c_1417_n 0.00112709f $X=9.09 $Y=1.325 $X2=0
+ $Y2=0
cc_643 N_A_1117_297#_c_815_n N_VGND_c_1417_n 0.00115239f $X=8.51 $Y=0.51 $X2=0
+ $Y2=0
cc_644 N_A_1117_297#_c_781_n N_VGND_c_1422_n 0.00193763f $X=9.005 $Y=0.82 $X2=0
+ $Y2=0
cc_645 N_A_1117_297#_c_802_n N_VGND_c_1422_n 0.00504557f $X=8.365 $Y=0.51 $X2=0
+ $Y2=0
cc_646 N_A_1117_297#_c_785_n N_VGND_c_1422_n 2.9688e-19 $X=5.895 $Y=0.51 $X2=0
+ $Y2=0
cc_647 N_A_1117_297#_c_786_n N_VGND_c_1422_n 0.0244659f $X=5.75 $Y=0.51 $X2=0
+ $Y2=0
cc_648 N_A_1117_297#_c_815_n N_VGND_c_1422_n 3.63685e-19 $X=8.51 $Y=0.51 $X2=0
+ $Y2=0
cc_649 N_A_1117_297#_c_816_n N_VGND_c_1422_n 0.0143515f $X=8.51 $Y=0.51 $X2=0
+ $Y2=0
cc_650 N_A_1117_297#_c_779_n N_VGND_c_1425_n 0.00487842f $X=9.15 $Y=0.995 $X2=0
+ $Y2=0
cc_651 N_A_1117_297#_c_783_n N_VGND_c_1425_n 0.00181647f $X=9.09 $Y=1.325 $X2=0
+ $Y2=0
cc_652 N_A_1117_297#_M1006_d N_VGND_c_1426_n 0.00190368f $X=8.305 $Y=0.235 $X2=0
+ $Y2=0
cc_653 N_A_1117_297#_c_779_n N_VGND_c_1426_n 0.00845884f $X=9.15 $Y=0.995 $X2=0
+ $Y2=0
cc_654 N_A_1117_297#_c_781_n N_VGND_c_1426_n 0.00437041f $X=9.005 $Y=0.82 $X2=0
+ $Y2=0
cc_655 N_A_1117_297#_c_783_n N_VGND_c_1426_n 0.00372241f $X=9.09 $Y=1.325 $X2=0
+ $Y2=0
cc_656 N_A_1117_297#_c_802_n N_VGND_c_1426_n 0.215402f $X=8.365 $Y=0.51 $X2=0
+ $Y2=0
cc_657 N_A_1117_297#_c_785_n N_VGND_c_1426_n 0.028616f $X=5.895 $Y=0.51 $X2=0
+ $Y2=0
cc_658 N_A_1117_297#_c_786_n N_VGND_c_1426_n 0.00387583f $X=5.75 $Y=0.51 $X2=0
+ $Y2=0
cc_659 N_A_1117_297#_c_815_n N_VGND_c_1426_n 0.0285254f $X=8.51 $Y=0.51 $X2=0
+ $Y2=0
cc_660 N_A_1117_297#_c_816_n N_VGND_c_1426_n 0.00348354f $X=8.51 $Y=0.51 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_914_n N_X_M1001_s 0.00217524f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_662 N_VPWR_c_914_n N_X_M1005_s 0.0038878f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_663 N_VPWR_c_916_n N_X_c_1033_n 0.0150775f $X=1.125 $Y=2.72 $X2=0 $Y2=0
cc_664 N_VPWR_c_914_n N_X_c_1033_n 0.0119688f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_665 N_VPWR_c_917_n N_X_c_1036_n 0.0136043f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_666 N_VPWR_c_917_n N_X_c_1029_n 0.0062286f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_667 N_VPWR_c_917_n N_X_c_1049_n 0.0644832f $X=1.21 $Y=1.66 $X2=0 $Y2=0
cc_668 N_VPWR_c_923_n N_X_c_1049_n 0.0171953f $X=1.915 $Y=2.72 $X2=0 $Y2=0
cc_669 N_VPWR_c_914_n N_X_c_1049_n 0.010364f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_670 N_VPWR_c_914_n N_A_607_325#_M1013_d 0.00233026f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_919_n N_A_607_325#_c_1073_n 0.00147971f $X=4.77 $Y=2.32 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_924_n N_A_607_325#_c_1073_n 0.0114434f $X=4.605 $Y=2.72 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_914_n N_A_607_325#_c_1073_n 0.0210414f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_674 N_VPWR_M1000_s N_A_607_325#_c_1069_n 0.00637486f $X=4.645 $Y=2.175 $X2=0
+ $Y2=0
cc_675 N_VPWR_M1000_s N_A_607_325#_c_1075_n 0.00130442f $X=4.645 $Y=2.175 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_919_n N_A_607_325#_c_1075_n 0.00607843f $X=4.77 $Y=2.32 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_925_n N_A_607_325#_c_1075_n 0.00503515f $X=8.775 $Y=2.72 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_914_n N_A_607_325#_c_1075_n 0.00935628f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_919_n N_A_607_325#_c_1076_n 0.00173147f $X=4.77 $Y=2.32 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_925_n N_A_607_325#_c_1077_n 0.0300226f $X=8.775 $Y=2.72 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_914_n N_A_607_325#_c_1077_n 0.0193106f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_919_n N_A_607_325#_c_1078_n 0.00833535f $X=4.77 $Y=2.32 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_925_n N_A_607_325#_c_1078_n 0.0105925f $X=8.775 $Y=2.72 $X2=0
+ $Y2=0
cc_684 N_VPWR_c_914_n N_A_607_325#_c_1078_n 0.00644598f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_685 N_VPWR_c_920_n N_A_607_325#_c_1080_n 0.00704283f $X=8.94 $Y=2.36 $X2=0
+ $Y2=0
cc_686 N_VPWR_c_925_n N_A_607_325#_c_1080_n 0.12359f $X=8.775 $Y=2.72 $X2=0
+ $Y2=0
cc_687 N_VPWR_c_914_n N_A_607_325#_c_1080_n 0.07455f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_688 N_VPWR_M1000_s N_A_607_325#_c_1081_n 0.00224421f $X=4.645 $Y=2.175 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_919_n N_A_607_325#_c_1081_n 0.0144069f $X=4.77 $Y=2.32 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_914_n N_A_607_325#_c_1081_n 8.22076e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_925_n N_A_607_325#_c_1082_n 0.0103171f $X=8.775 $Y=2.72 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_914_n N_A_607_325#_c_1082_n 0.00587148f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_693 N_VPWR_M1000_s N_A_631_49#_c_1223_n 0.00100785f $X=4.645 $Y=2.175 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_914_n N_A_1382_49#_M1012_d 0.00248304f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_926_n N_A_1382_49#_c_1349_n 0.0197307f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_914_n N_A_1382_49#_c_1349_n 0.0111012f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_697 N_VPWR_M1017_d N_A_1382_49#_c_1358_n 0.00343874f $X=8.805 $Y=1.485 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_920_n N_A_1382_49#_c_1358_n 0.0162117f $X=8.94 $Y=2.36 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_925_n N_A_1382_49#_c_1358_n 0.00690051f $X=8.775 $Y=2.72 $X2=0
+ $Y2=0
cc_700 N_VPWR_c_914_n N_A_1382_49#_c_1358_n 0.0144976f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_926_n N_A_1382_49#_c_1351_n 0.00258024f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_914_n N_A_1382_49#_c_1351_n 0.00441029f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_703 N_X_c_1028_n N_VGND_c_1413_n 0.00854925f $X=0.79 $Y=0.56 $X2=0 $Y2=0
cc_704 N_X_c_1036_n N_VGND_c_1414_n 0.00981162f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_705 N_X_c_1037_n N_VGND_c_1414_n 0.0279087f $X=1.64 $Y=0.56 $X2=0 $Y2=0
cc_706 N_X_c_1037_n N_VGND_c_1424_n 0.00984675f $X=1.64 $Y=0.56 $X2=0 $Y2=0
cc_707 N_X_M1010_s N_VGND_c_1426_n 0.00405614f $X=0.655 $Y=0.235 $X2=0 $Y2=0
cc_708 N_X_M1022_s N_VGND_c_1426_n 0.00401728f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_709 N_X_c_1028_n N_VGND_c_1426_n 0.00878408f $X=0.79 $Y=0.56 $X2=0 $Y2=0
cc_710 N_X_c_1037_n N_VGND_c_1426_n 0.00925029f $X=1.64 $Y=0.56 $X2=0 $Y2=0
cc_711 N_A_607_325#_c_1073_n N_A_631_49#_M1026_d 0.0117309f $X=4.625 $Y=1.98
+ $X2=0 $Y2=0
cc_712 N_A_607_325#_c_1080_n N_A_631_49#_M1018_d 0.00884079f $X=8.005 $Y=2.36
+ $X2=0 $Y2=0
cc_713 N_A_607_325#_M1020_d N_A_631_49#_c_1228_n 0.0100433f $X=4.015 $Y=0.245
+ $X2=0 $Y2=0
cc_714 N_A_607_325#_c_1067_n N_A_631_49#_c_1228_n 0.0200889f $X=4.515 $Y=0.37
+ $X2=0 $Y2=0
cc_715 N_A_607_325#_c_1068_n N_A_631_49#_c_1228_n 0.0140571f $X=4.6 $Y=1.035
+ $X2=0 $Y2=0
cc_716 N_A_607_325#_M1020_d N_A_631_49#_c_1216_n 0.00292468f $X=4.015 $Y=0.245
+ $X2=0 $Y2=0
cc_717 N_A_607_325#_c_1068_n N_A_631_49#_c_1216_n 0.0179157f $X=4.6 $Y=1.035
+ $X2=0 $Y2=0
cc_718 N_A_607_325#_c_1069_n N_A_631_49#_c_1216_n 0.00902524f $X=4.71 $Y=1.895
+ $X2=0 $Y2=0
cc_719 N_A_607_325#_c_1071_n N_A_631_49#_c_1216_n 0.0132103f $X=4.71 $Y=1.12
+ $X2=0 $Y2=0
cc_720 N_A_607_325#_c_1070_n N_A_631_49#_c_1220_n 0.0111917f $X=6.05 $Y=2.275
+ $X2=0 $Y2=0
cc_721 N_A_607_325#_c_1072_n N_A_631_49#_c_1220_n 2.53366e-19 $X=6.05 $Y=0.772
+ $X2=0 $Y2=0
cc_722 N_A_607_325#_c_1070_n N_A_631_49#_c_1257_n 0.0308675f $X=6.05 $Y=2.275
+ $X2=0 $Y2=0
cc_723 N_A_607_325#_c_1080_n N_A_631_49#_c_1257_n 0.0235166f $X=8.005 $Y=2.36
+ $X2=0 $Y2=0
cc_724 N_A_607_325#_c_1080_n N_A_631_49#_c_1221_n 0.00873322f $X=8.005 $Y=2.36
+ $X2=0 $Y2=0
cc_725 N_A_607_325#_c_1116_n N_A_631_49#_c_1217_n 0.00284845f $X=6.29 $Y=0.545
+ $X2=0 $Y2=0
cc_726 N_A_607_325#_c_1073_n N_A_631_49#_c_1223_n 0.00437461f $X=4.625 $Y=1.98
+ $X2=0 $Y2=0
cc_727 N_A_607_325#_c_1069_n N_A_631_49#_c_1223_n 0.0161183f $X=4.71 $Y=1.895
+ $X2=0 $Y2=0
cc_728 N_A_607_325#_c_1075_n N_A_631_49#_c_1223_n 0.0108524f $X=5.27 $Y=1.98
+ $X2=0 $Y2=0
cc_729 N_A_607_325#_c_1070_n N_A_631_49#_c_1223_n 0.0191401f $X=6.05 $Y=2.275
+ $X2=0 $Y2=0
cc_730 N_A_607_325#_c_1071_n N_A_631_49#_c_1223_n 0.0052436f $X=4.71 $Y=1.12
+ $X2=0 $Y2=0
cc_731 N_A_607_325#_c_1072_n N_A_631_49#_c_1223_n 3.36438e-19 $X=6.05 $Y=0.772
+ $X2=0 $Y2=0
cc_732 N_A_607_325#_c_1073_n N_A_631_49#_c_1224_n 0.00415423f $X=4.625 $Y=1.98
+ $X2=0 $Y2=0
cc_733 N_A_607_325#_c_1069_n N_A_631_49#_c_1224_n 0.00275249f $X=4.71 $Y=1.895
+ $X2=0 $Y2=0
cc_734 N_A_607_325#_c_1073_n N_A_631_49#_c_1225_n 0.0251846f $X=4.625 $Y=1.98
+ $X2=0 $Y2=0
cc_735 N_A_607_325#_c_1069_n N_A_631_49#_c_1225_n 0.0231767f $X=4.71 $Y=1.895
+ $X2=0 $Y2=0
cc_736 N_A_607_325#_c_1070_n N_A_631_49#_c_1226_n 0.00132955f $X=6.05 $Y=2.275
+ $X2=0 $Y2=0
cc_737 N_A_607_325#_c_1080_n N_A_1382_49#_M1019_d 0.0055303f $X=8.005 $Y=2.36
+ $X2=0 $Y2=0
cc_738 N_A_607_325#_c_1080_n N_A_1382_49#_c_1357_n 0.0129278f $X=8.005 $Y=2.36
+ $X2=0 $Y2=0
cc_739 N_A_607_325#_M1013_d N_A_1382_49#_c_1358_n 0.00612338f $X=7.785 $Y=1.645
+ $X2=0 $Y2=0
cc_740 N_A_607_325#_c_1080_n N_A_1382_49#_c_1358_n 0.0467387f $X=8.005 $Y=2.36
+ $X2=0 $Y2=0
cc_741 N_A_607_325#_c_1067_n N_VGND_c_1416_n 0.014042f $X=4.515 $Y=0.37 $X2=0
+ $Y2=0
cc_742 N_A_607_325#_c_1068_n N_VGND_c_1416_n 0.0298884f $X=4.6 $Y=1.035 $X2=0
+ $Y2=0
cc_743 N_A_607_325#_c_1067_n N_VGND_c_1420_n 0.0344776f $X=4.515 $Y=0.37 $X2=0
+ $Y2=0
cc_744 N_A_607_325#_c_1116_n N_VGND_c_1422_n 0.00800682f $X=6.29 $Y=0.545 $X2=0
+ $Y2=0
cc_745 N_A_607_325#_c_1072_n N_VGND_c_1422_n 0.00224548f $X=6.05 $Y=0.772 $X2=0
+ $Y2=0
cc_746 N_A_607_325#_c_1067_n N_VGND_c_1426_n 0.0232692f $X=4.515 $Y=0.37 $X2=0
+ $Y2=0
cc_747 N_A_607_325#_c_1116_n N_VGND_c_1426_n 0.0018012f $X=6.29 $Y=0.545 $X2=0
+ $Y2=0
cc_748 N_A_631_49#_c_1217_n N_A_1382_49#_M1021_d 0.00729398f $X=7.01 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_749 N_A_631_49#_c_1329_p N_A_1382_49#_M1021_d 0.0024562f $X=7.095 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_750 N_A_631_49#_c_1288_n N_A_1382_49#_M1021_d 0.0107136f $X=7.605 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_751 N_A_631_49#_c_1221_n N_A_1382_49#_M1019_d 0.00414782f $X=6.925 $Y=1.53
+ $X2=0 $Y2=0
cc_752 N_A_631_49#_c_1257_n N_A_1382_49#_c_1345_n 0.00487817f $X=6.49 $Y=1.62
+ $X2=0 $Y2=0
cc_753 N_A_631_49#_c_1221_n N_A_1382_49#_c_1345_n 0.0134336f $X=6.925 $Y=1.53
+ $X2=0 $Y2=0
cc_754 N_A_631_49#_c_1217_n N_A_1382_49#_c_1345_n 0.0622566f $X=7.01 $Y=1.445
+ $X2=0 $Y2=0
cc_755 N_A_631_49#_c_1288_n N_A_1382_49#_c_1345_n 0.0106102f $X=7.605 $Y=0.36
+ $X2=0 $Y2=0
cc_756 N_A_631_49#_c_1226_n N_A_1382_49#_c_1345_n 0.0013871f $X=6.67 $Y=1.53
+ $X2=0 $Y2=0
cc_757 N_A_631_49#_c_1223_n N_VGND_c_1416_n 0.00553699f $X=6.525 $Y=1.53 $X2=0
+ $Y2=0
cc_758 N_A_631_49#_c_1228_n N_VGND_c_1420_n 0.00257941f $X=4.175 $Y=0.71 $X2=0
+ $Y2=0
cc_759 N_A_631_49#_c_1329_p N_VGND_c_1422_n 0.0104913f $X=7.095 $Y=0.34 $X2=0
+ $Y2=0
cc_760 N_A_631_49#_c_1288_n N_VGND_c_1422_n 0.0586043f $X=7.605 $Y=0.36 $X2=0
+ $Y2=0
cc_761 N_A_631_49#_M1023_d N_VGND_c_1426_n 0.00184103f $X=7.705 $Y=0.245 $X2=0
+ $Y2=0
cc_762 N_A_631_49#_c_1329_p N_VGND_c_1426_n 0.00184693f $X=7.095 $Y=0.34 $X2=0
+ $Y2=0
cc_763 N_A_631_49#_c_1218_n N_VGND_c_1426_n 0.00606683f $X=3.505 $Y=0.765 $X2=0
+ $Y2=0
cc_764 N_A_631_49#_c_1288_n N_VGND_c_1426_n 0.0092581f $X=7.605 $Y=0.36 $X2=0
+ $Y2=0
cc_765 N_A_1382_49#_c_1347_n N_VGND_c_1425_n 0.0197576f $X=9.49 $Y=0.42 $X2=0
+ $Y2=0
cc_766 N_A_1382_49#_M1009_d N_VGND_c_1426_n 0.00399944f $X=9.225 $Y=0.235 $X2=0
+ $Y2=0
cc_767 N_A_1382_49#_c_1347_n N_VGND_c_1426_n 0.0113402f $X=9.49 $Y=0.42 $X2=0
+ $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o31a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 1.055000 5.470000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.265000 1.055000 4.970000 1.360000 ;
        RECT 4.680000 1.360000 4.970000 1.530000 ;
        RECT 4.680000 1.530000 6.355000 1.700000 ;
        RECT 5.640000 1.055000 6.355000 1.530000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 1.055000 4.095000 1.360000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 1.055000 3.575000 1.355000 ;
        RECT 2.780000 1.355000 3.150000 1.695000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 1.765000 0.885000 ;
        RECT 0.085000 0.885000 0.735000 1.460000 ;
        RECT 0.085000 1.460000 1.750000 1.665000 ;
        RECT 0.680000 0.255000 0.895000 0.655000 ;
        RECT 0.680000 0.655000 1.765000 0.715000 ;
        RECT 0.680000 1.665000 0.895000 2.465000 ;
        RECT 1.565000 0.255000 1.765000 0.655000 ;
        RECT 1.565000 1.665000 1.750000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.085000  0.085000 0.510000 0.545000 ;
        RECT 1.065000  0.085000 1.395000 0.485000 ;
        RECT 1.935000  0.085000 2.250000 0.885000 ;
        RECT 3.760000  0.085000 4.090000 0.445000 ;
        RECT 4.600000  0.085000 4.930000 0.445000 ;
        RECT 5.440000  0.085000 5.770000 0.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.085000 1.835000 0.510000 2.635000 ;
        RECT 1.065000 1.835000 1.395000 2.635000 ;
        RECT 1.920000 1.460000 2.250000 2.635000 ;
        RECT 2.780000 2.240000 3.110000 2.635000 ;
        RECT 5.020000 2.240000 5.350000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.905000 1.055000 2.610000 1.290000 ;
      RECT 2.440000 0.255000 3.570000 0.465000 ;
      RECT 2.440000 0.635000 3.210000 0.885000 ;
      RECT 2.440000 0.885000 2.610000 1.055000 ;
      RECT 2.440000 1.290000 2.610000 1.870000 ;
      RECT 2.440000 1.870000 4.090000 2.070000 ;
      RECT 2.440000 2.070000 2.610000 2.465000 ;
      RECT 3.320000 1.530000 4.510000 1.700000 ;
      RECT 3.380000 0.465000 3.570000 0.635000 ;
      RECT 3.380000 0.635000 6.355000 0.885000 ;
      RECT 3.760000 2.070000 4.090000 2.465000 ;
      RECT 4.260000 0.255000 4.430000 0.635000 ;
      RECT 4.260000 1.700000 4.510000 2.465000 ;
      RECT 4.680000 1.870000 5.720000 2.070000 ;
      RECT 4.680000 2.070000 4.850000 2.465000 ;
      RECT 5.100000 0.255000 5.270000 0.635000 ;
      RECT 5.520000 2.070000 5.720000 2.465000 ;
      RECT 5.890000 1.870000 6.355000 2.465000 ;
      RECT 5.940000 0.255000 6.355000 0.635000 ;
    LAYER mcon ;
      RECT 4.285000 2.125000 4.455000 2.295000 ;
      RECT 6.125000 2.125000 6.295000 2.295000 ;
    LAYER met1 ;
      RECT 4.225000 2.095000 4.515000 2.140000 ;
      RECT 4.225000 2.140000 6.355000 2.280000 ;
      RECT 4.225000 2.280000 4.515000 2.325000 ;
      RECT 6.065000 2.095000 6.355000 2.140000 ;
      RECT 6.065000 2.280000 6.355000 2.325000 ;
  END
END sky130_fd_sc_hd__o31a_4
END LIBRARY

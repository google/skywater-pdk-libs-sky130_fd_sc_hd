* File: sky130_fd_sc_hd__nor4_1.pex.spice
* Created: Tue Sep  1 19:18:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4_1%D 1 3 6 8 9 16
c30 6 0 1.88106e-19 $X=0.47 $Y=1.985
r31 13 16 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.25 $Y=1.16
+ $X2=0.47 $Y2=1.16
r32 8 9 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.21 $Y=1.16 $X2=0.21
+ $Y2=0.85
r33 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r34 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r35 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r36 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_1%C 3 7 10 11 13 17 22
c46 22 0 1.88106e-19 $X=1.157 $Y=1.615
c47 11 0 7.80018e-20 $X=0.93 $Y=1.16
r48 13 22 0.388182 $w=1.98e-07 $l=7e-09 $layer=LI1_cond $X=1.15 $Y=1.515
+ $X2=1.157 $Y2=1.515
r49 13 22 0.10027 $w=8.33e-07 $l=7e-09 $layer=LI1_cond $X=1.15 $Y=2.032
+ $X2=1.157 $Y2=2.032
r50 11 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=0.93 $Y2=1.325
r51 11 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=0.93 $Y2=0.995
r52 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.16 $X2=0.93 $Y2=1.16
r53 8 13 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=1.515
+ $X2=1.15 $Y2=1.515
r54 8 10 12.7771 $w=2.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.96 $Y=1.415
+ $X2=0.96 $Y2=1.16
r55 7 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.985 $Y=0.56
+ $X2=0.985 $Y2=0.995
r56 3 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.88 $Y=1.985
+ $X2=0.88 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_1%B 1 3 6 10 13 15
c41 15 0 7.80018e-20 $X=1.61 $Y=1.87
c42 10 0 1.93867e-19 $X=1.41 $Y=1.16
r43 13 15 30.0115 $w=2.38e-07 $l=6.25e-07 $layer=LI1_cond $X=1.575 $Y=1.245
+ $X2=1.575 $Y2=1.87
r44 9 13 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=1.16
+ $X2=1.575 $Y2=1.16
r45 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.16 $X2=1.41 $Y2=1.16
r46 4 10 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r47 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325 $X2=1.41
+ $Y2=1.985
r48 1 10 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_1%A 1 3 6 8 13
c28 8 0 1.75897e-19 $X=2.07 $Y=0.85
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r30 10 13 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=2.06 $Y2=1.16
r31 8 14 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.085 $Y=0.85
+ $X2=2.085 $Y2=1.16
r32 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=1.985
r34 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.995 $X2=1.83
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_1%Y 1 2 3 10 11 12 18 24 28
c48 24 0 1.93867e-19 $X=1.62 $Y=0.55
r49 28 33 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.34
r50 24 26 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.55
+ $X2=1.62 $Y2=0.74
r51 21 22 7.701 $w=3.01e-07 $l=1.9e-07 $layer=LI1_cond $X=0.682 $Y=0.55
+ $X2=0.682 $Y2=0.74
r52 15 28 18.7487 $w=3.33e-07 $l=5.45e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.21
r53 15 18 21.7251 $w=1.68e-07 $l=3.33e-07 $layer=LI1_cond $X=0.257 $Y=1.58
+ $X2=0.59 $Y2=1.58
r54 13 22 4.08057 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.86 $Y=0.74
+ $X2=0.682 $Y2=0.74
r55 12 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0.74
+ $X2=1.62 $Y2=0.74
r56 12 13 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.535 $Y=0.74
+ $X2=0.86 $Y2=0.74
r57 11 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.59 $Y=1.495
+ $X2=0.59 $Y2=1.58
r58 10 22 5.73711 $w=3.01e-07 $l=1.27609e-07 $layer=LI1_cond $X=0.59 $Y=0.825
+ $X2=0.682 $Y2=0.74
r59 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.59 $Y=0.825
+ $X2=0.59 $Y2=1.495
r60 3 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r61 3 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r62 2 24 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.55
r63 1 21 182 $w=1.7e-07 $l=4.14337e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.775 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_1%VPWR 1 4 6 8 10 20
r27 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r28 17 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 12 16 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 10 19 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.127 $Y2=2.72
r32 10 16 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r33 8 17 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r35 4 19 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.085 $Y=2.635
+ $X2=2.127 $Y2=2.72
r36 4 6 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=2.085 $Y=2.635
+ $X2=2.085 $Y2=2
r37 1 6 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4_1%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
c43 18 0 1.75897e-19 $X=2.04 $Y=0.085
r44 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r45 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r46 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r47 33 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r48 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r49 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r50 30 32 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r51 29 41 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.087
+ $Y2=0
r52 29 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r53 28 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r54 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r55 25 35 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r56 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r57 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r58 24 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r59 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r60 22 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r61 18 41 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.087 $Y2=0
r62 18 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.39
r63 14 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r64 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r65 10 35 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r66 10 12 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.39
r67 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.39
r68 2 16 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.235 $X2=1.2 $Y2=0.39
r69 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__decap_6.spice
* Created: Tue Sep  1 19:02:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__decap_6.pex.spice"
.subckt sky130_fd_sc_hd__decap_6  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_VPWR_M1001_g N_VGND_M1001_s VNB NSHORT L=1.97 W=0.55
+ AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 M=1 R=0.279188 SA=984999
+ SB=984999 A=1.0835 P=5.04 MULT=1
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=1.97 W=0.87
+ AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 M=1 R=0.441624 SA=984999
+ SB=984999 A=1.7139 P=5.68 MULT=1
DX2_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__decap_6.pxi.spice"
*
.ends
*
*

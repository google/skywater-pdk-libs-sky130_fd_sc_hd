* File: sky130_fd_sc_hd__nor3_1.pxi.spice
* Created: Thu Aug 27 14:31:59 2020
* 
x_PM_SKY130_FD_SC_HD__NOR3_1%C N_C_c_37_n N_C_M1005_g N_C_M1004_g C N_C_c_39_n
+ PM_SKY130_FD_SC_HD__NOR3_1%C
x_PM_SKY130_FD_SC_HD__NOR3_1%B N_B_c_64_n N_B_M1002_g N_B_M1001_g N_B_c_65_n
+ N_B_c_66_n B B PM_SKY130_FD_SC_HD__NOR3_1%B
x_PM_SKY130_FD_SC_HD__NOR3_1%A N_A_c_103_n N_A_M1003_g N_A_M1000_g A A A
+ N_A_c_105_n PM_SKY130_FD_SC_HD__NOR3_1%A
x_PM_SKY130_FD_SC_HD__NOR3_1%Y N_Y_M1005_s N_Y_M1002_d N_Y_M1004_s N_Y_c_144_n
+ N_Y_c_146_n N_Y_c_167_n N_Y_c_158_n N_Y_c_139_n N_Y_c_140_n N_Y_c_164_n Y
+ N_Y_c_142_n N_Y_c_143_n Y PM_SKY130_FD_SC_HD__NOR3_1%Y
x_PM_SKY130_FD_SC_HD__NOR3_1%VPWR N_VPWR_M1000_d N_VPWR_c_206_n N_VPWR_c_207_n
+ VPWR N_VPWR_c_208_n N_VPWR_c_205_n PM_SKY130_FD_SC_HD__NOR3_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR3_1%VGND N_VGND_M1005_d N_VGND_M1003_d N_VGND_c_227_n
+ N_VGND_c_228_n N_VGND_c_229_n VGND N_VGND_c_230_n N_VGND_c_231_n
+ N_VGND_c_232_n N_VGND_c_233_n PM_SKY130_FD_SC_HD__NOR3_1%VGND
cc_1 VNB N_C_c_37_n 0.0219513f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB C 0.0143803f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_c_39_n 0.0355062f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B_c_64_n 0.0161955f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_B_c_65_n 0.00329554f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_6 VNB N_B_c_66_n 0.0200302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_c_103_n 0.0178908f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB A 0.0261988f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_9 VNB N_A_c_105_n 0.0368307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_139_n 0.00287947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_140_n 0.017363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_205_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_227_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_228_n 0.0119223f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_15 VNB N_VGND_c_229_n 0.012566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_230_n 0.0149052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_231_n 0.0115543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_232_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_233_n 0.123624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VPB N_C_M1004_g 0.0262632f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_21 VPB C 0.00356082f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_22 VPB N_C_c_39_n 0.00949799f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_23 VPB N_B_M1001_g 0.0181868f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_24 VPB N_B_c_65_n 5.65188e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_25 VPB N_B_c_66_n 0.00517728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB B 0.0019548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_M1000_g 0.0213063f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_28 VPB A 0.0158577f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_29 VPB N_A_c_105_n 0.0121657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_Y_c_139_n 0.00130071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_Y_c_142_n 0.00753565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_Y_c_143_n 0.030912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_206_n 0.0110025f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_34 VPB N_VPWR_c_207_n 0.0328657f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_35 VPB N_VPWR_c_208_n 0.0379439f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_36 VPB N_VPWR_c_205_n 0.0430082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 N_C_c_37_n N_B_c_64_n 0.0255041f $X=0.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_38 N_C_M1004_g N_B_M1001_g 0.0569056f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_39 C N_B_c_65_n 0.0264046f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_40 N_C_c_39_n N_B_c_65_n 0.0024723f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_41 C N_B_c_66_n 2.5326e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_42 N_C_c_39_n N_B_c_66_n 0.0207204f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_43 N_C_M1004_g B 0.00618236f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_44 N_C_c_37_n N_Y_c_144_n 0.0143828f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_45 C N_Y_c_144_n 0.00396858f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_46 N_C_M1004_g N_Y_c_146_n 0.0101518f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_47 C N_Y_c_140_n 0.0202418f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_48 N_C_c_39_n N_Y_c_140_n 0.00164655f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_49 N_C_M1004_g N_Y_c_142_n 7.32439e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_50 N_C_M1004_g N_Y_c_143_n 0.0107635f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_51 C N_Y_c_143_n 0.0251629f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_52 N_C_c_39_n N_Y_c_143_n 0.00196424f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_53 N_C_M1004_g N_VPWR_c_208_n 0.00360959f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_54 N_C_M1004_g N_VPWR_c_205_n 0.00621123f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_55 N_C_c_37_n N_VGND_c_227_n 0.0127917f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_56 N_C_c_37_n N_VGND_c_230_n 0.00341689f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_57 N_C_c_37_n N_VGND_c_233_n 0.0050171f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_58 N_B_c_64_n N_A_c_103_n 0.0228932f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_59 N_B_M1001_g N_A_M1000_g 0.0526224f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_60 B N_A_M1000_g 3.80691e-19 $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_61 N_B_c_65_n N_A_c_105_n 3.1445e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B_c_66_n N_A_c_105_n 0.0202376f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_63 N_B_c_64_n N_Y_c_144_n 0.0103948f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_64 N_B_c_65_n N_Y_c_144_n 0.0256654f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_65 N_B_c_66_n N_Y_c_144_n 0.00122018f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_66 N_B_M1001_g N_Y_c_146_n 0.0133463f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_67 B N_Y_c_146_n 0.00853825f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_68 N_B_c_66_n N_Y_c_158_n 2.29104e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B_c_64_n N_Y_c_139_n 0.00343469f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B_M1001_g N_Y_c_139_n 0.00117375f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_71 N_B_c_65_n N_Y_c_139_n 0.0250399f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B_c_66_n N_Y_c_139_n 0.00190138f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_73 B N_Y_c_139_n 0.00782711f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_74 N_B_c_66_n N_Y_c_164_n 5.26998e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B_M1001_g N_Y_c_143_n 0.00121251f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_76 B A_109_297# 0.00294271f $X=0.61 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_77 N_B_M1001_g N_VPWR_c_208_n 0.00361001f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B_M1001_g N_VPWR_c_205_n 0.00532425f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B_c_64_n N_VGND_c_227_n 0.00772378f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B_c_64_n N_VGND_c_229_n 8.32923e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_64_n N_VGND_c_231_n 0.00341689f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_82 N_B_c_64_n N_VGND_c_233_n 0.00405445f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_Y_c_146_n 0.00163992f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1000_g N_Y_c_167_n 0.00756125f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_c_103_n N_Y_c_158_n 0.00520611f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_86 A N_Y_c_158_n 0.0138064f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_87 N_A_c_103_n N_Y_c_139_n 0.00335527f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_M1000_g N_Y_c_139_n 0.0036243f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_89 A N_Y_c_139_n 0.048235f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_c_105_n N_Y_c_139_n 0.00829361f $X=1.57 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_M1000_g N_Y_c_164_n 0.00768989f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_92 A N_Y_c_164_n 0.012862f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_93 A N_VPWR_M1000_d 0.00456601f $X=1.53 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_94 N_A_M1000_g N_VPWR_c_207_n 0.00456315f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_95 A N_VPWR_c_207_n 0.0240802f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_96 N_A_c_105_n N_VPWR_c_207_n 0.00230035f $X=1.57 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_M1000_g N_VPWR_c_208_n 0.00585385f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_M1000_g N_VPWR_c_205_n 0.0116482f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_99 A N_VGND_M1003_d 0.00488309f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A_c_103_n N_VGND_c_227_n 8.32923e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_101 A N_VGND_c_228_n 0.00134855f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_102 N_A_c_103_n N_VGND_c_229_n 0.0098809f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_103 A N_VGND_c_229_n 0.0169195f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A_c_105_n N_VGND_c_229_n 0.00288712f $X=1.57 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_c_103_n N_VGND_c_231_n 0.00382526f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_c_103_n N_VGND_c_233_n 0.00538868f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_107 A N_VGND_c_233_n 0.00305454f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_108 N_Y_c_146_n A_109_297# 0.00357801f $X=1 $Y=2.365 $X2=-0.19 $Y2=-0.24
cc_109 N_Y_c_146_n A_193_297# 0.0034556f $X=1 $Y=2.365 $X2=-0.19 $Y2=-0.24
cc_110 N_Y_c_167_n A_193_297# 0.00926926f $X=1.085 $Y=2.28 $X2=-0.19 $Y2=-0.24
cc_111 N_Y_c_139_n A_193_297# 2.02674e-19 $X=1.23 $Y=1.495 $X2=-0.19 $Y2=-0.24
cc_112 N_Y_c_164_n A_193_297# 0.0035673f $X=1.23 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_113 N_Y_c_146_n N_VPWR_c_208_n 0.0391903f $X=1 $Y=2.365 $X2=0 $Y2=0
cc_114 N_Y_c_142_n N_VPWR_c_208_n 0.019625f $X=0.257 $Y=2.28 $X2=0 $Y2=0
cc_115 N_Y_M1004_s N_VPWR_c_205_n 0.00209863f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_116 N_Y_c_146_n N_VPWR_c_205_n 0.0264778f $X=1 $Y=2.365 $X2=0 $Y2=0
cc_117 N_Y_c_142_n N_VPWR_c_205_n 0.0125934f $X=0.257 $Y=2.28 $X2=0 $Y2=0
cc_118 N_Y_c_144_n N_VGND_M1005_d 0.00323154f $X=1.015 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_119 N_Y_c_144_n N_VGND_c_227_n 0.0160613f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_120 N_Y_c_144_n N_VGND_c_230_n 0.00232396f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_121 N_Y_c_140_n N_VGND_c_230_n 0.00928504f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_122 N_Y_c_144_n N_VGND_c_231_n 0.00232396f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_123 N_Y_c_158_n N_VGND_c_231_n 0.00790924f $X=1.23 $Y=0.825 $X2=0 $Y2=0
cc_124 N_Y_M1005_s N_VGND_c_233_n 0.0024189f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_125 N_Y_M1002_d N_VGND_c_233_n 0.00266592f $X=0.965 $Y=0.235 $X2=0 $Y2=0
cc_126 N_Y_c_144_n N_VGND_c_233_n 0.00971098f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_127 N_Y_c_158_n N_VGND_c_233_n 0.00944761f $X=1.23 $Y=0.825 $X2=0 $Y2=0
cc_128 N_Y_c_140_n N_VGND_c_233_n 0.00892296f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_129 A_109_297# N_VPWR_c_205_n 0.00217425f $X=0.545 $Y=1.485 $X2=0.712
+ $Y2=1.53
cc_130 A_193_297# N_VPWR_c_205_n 0.00442896f $X=0.965 $Y=1.485 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__and2_0.pex.spice
* Created: Tue Sep  1 18:56:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND2_0%A 2 5 9 11 12 15 16
r34 15 17 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.397 $Y=1.375
+ $X2=0.397 $Y2=1.21
r35 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.345
+ $Y=1.375 $X2=0.345 $Y2=1.375
r36 12 16 16.5351 $w=3.43e-07 $l=4.95e-07 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=1.375
r37 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.54 $Y=2.275
+ $X2=0.54 $Y2=1.88
r38 5 17 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.54 $Y=0.445
+ $X2=0.54 $Y2=1.21
r39 2 11 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.397 $Y=1.663
+ $X2=0.397 $Y2=1.88
r40 1 15 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=0.397 $Y=1.427
+ $X2=0.397 $Y2=1.375
r41 1 2 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=0.397 $Y=1.427
+ $X2=0.397 $Y2=1.663
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_0%B 3 7 9 10 14
c35 3 0 1.70382e-19 $X=0.9 $Y=0.445
r36 14 17 92.4199 $w=4.45e-07 $l=5.3e-07 $layer=POLY_cond $X=1.047 $Y=1.18
+ $X2=1.047 $Y2=1.71
r37 14 16 43.0534 $w=4.45e-07 $l=1.35e-07 $layer=POLY_cond $X=1.047 $Y=1.18
+ $X2=1.047 $Y2=1.045
r38 9 10 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.105 $Y=1.18
+ $X2=1.105 $Y2=1.53
r39 9 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.105
+ $Y=1.18 $X2=1.105 $Y2=1.18
r40 7 17 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.98 $Y=2.275
+ $X2=0.98 $Y2=1.71
r41 3 16 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.9 $Y=0.445 $X2=0.9
+ $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_0%A_40_47# 1 2 9 12 15 16 18 21 25 29 30 35 37
+ 38
r72 37 38 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.732 $Y=2.3
+ $X2=0.732 $Y2=2.135
r73 34 35 4.15858 $w=2.53e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.822
+ $X2=0.77 $Y2=0.822
r74 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=0.93 $X2=1.615 $Y2=0.93
r75 27 29 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.615 $Y=0.91
+ $X2=1.615 $Y2=0.93
r76 25 27 7.21882 $w=2.15e-07 $l=2.12238e-07 $layer=LI1_cond $X=1.45 $Y=0.802
+ $X2=1.615 $Y2=0.91
r77 25 35 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=1.45 $Y=0.802
+ $X2=0.77 $Y2=0.802
r78 23 34 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.685 $Y=0.95
+ $X2=0.685 $Y2=0.822
r79 23 38 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=0.685 $Y=0.95
+ $X2=0.685 $Y2=2.135
r80 19 34 15.7275 $w=2.53e-07 $l=3.48e-07 $layer=LI1_cond $X=0.337 $Y=0.822
+ $X2=0.685 $Y2=0.822
r81 19 21 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=0.337 $Y=0.695
+ $X2=0.337 $Y2=0.445
r82 17 30 55.6971 $w=3.45e-07 $l=3.33e-07 $layer=POLY_cond $X=1.652 $Y=1.263
+ $X2=1.652 $Y2=0.93
r83 17 18 47.5363 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=1.652 $Y=1.263
+ $X2=1.652 $Y2=1.435
r84 16 30 2.50888 $w=3.45e-07 $l=1.5e-08 $layer=POLY_cond $X=1.652 $Y=0.915
+ $X2=1.652 $Y2=0.93
r85 15 16 43.8566 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=1.63 $Y=0.765
+ $X2=1.63 $Y2=0.915
r86 12 18 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.75 $Y=2.165
+ $X2=1.75 $Y2=1.435
r87 9 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.51 $Y=0.445
+ $X2=1.51 $Y2=0.765
r88 2 37 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=2.065 $X2=0.765 $Y2=2.3
r89 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.325 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_0%VPWR 1 2 7 9 11 15 17 21 22 28
r34 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 22 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 19 28 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.62 $Y=2.72
+ $X2=1.365 $Y2=2.72
r38 19 21 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.62 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r40 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r41 13 28 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=2.635
+ $X2=1.365 $Y2=2.72
r42 13 15 14.8923 $w=5.08e-07 $l=6.35e-07 $layer=LI1_cond $X=1.365 $Y=2.635
+ $X2=1.365 $Y2=2
r43 12 25 4.1216 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=2.72
+ $X2=0.215 $Y2=2.72
r44 11 28 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.11 $Y=2.72
+ $X2=1.365 $Y2=2.72
r45 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.11 $Y=2.72
+ $X2=0.43 $Y2=2.72
r46 7 25 3.16309 $w=2.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.295 $Y=2.635
+ $X2=0.215 $Y2=2.72
r47 7 9 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=2.635
+ $X2=0.295 $Y2=2.34
r48 2 15 200 $w=1.7e-07 $l=5.01448e-07 $layer=licon1_PDIFF $count=3 $X=1.055
+ $Y=2.065 $X2=1.525 $Y2=2
r49 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=2.065 $X2=0.325 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_0%X 1 2 7 13 16 17
c19 7 0 1.70382e-19 $X=1.95 $Y=0.39
r20 16 17 6.09834 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=2.002 $Y=2
+ $X2=2.002 $Y2=1.835
r21 13 16 5.69442 $w=4.23e-07 $l=2.1e-07 $layer=LI1_cond $X=2.002 $Y=2.21
+ $X2=2.002 $Y2=2
r22 11 17 56.9698 $w=2.63e-07 $l=1.31e-06 $layer=LI1_cond $X=2.082 $Y=0.525
+ $X2=2.082 $Y2=1.835
r23 7 11 6.81727 $w=2.7e-07 $l=1.89855e-07 $layer=LI1_cond $X=1.95 $Y=0.39
+ $X2=2.082 $Y2=0.525
r24 7 9 9.60369 $w=2.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.95 $Y=0.39
+ $X2=1.725 $Y2=0.39
r25 2 16 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.845 $X2=1.965 $Y2=2
r26 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.725 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_0%VGND 1 4 6 13 14 18
r26 18 21 9.42908 $w=4.38e-07 $l=3.6e-07 $layer=LI1_cond $X=1.17 $Y=0 $X2=1.17
+ $Y2=0.36
r27 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r28 14 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r29 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r30 11 18 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.17
+ $Y2=0
r31 11 13 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=2.07
+ $Y2=0
r32 9 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r33 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r34 6 18 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.17
+ $Y2=0
r35 6 8 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.69
+ $Y2=0
r36 4 9 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r37 1 21 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=1.18 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__o22ai_4.pxi.spice
* Created: Thu Aug 27 14:38:06 2020
* 
x_PM_SKY130_FD_SC_HD__O22AI_4%A1 N_A1_c_105_n N_A1_M1013_g N_A1_M1002_g
+ N_A1_c_106_n N_A1_M1017_g N_A1_M1005_g N_A1_c_107_n N_A1_M1023_g N_A1_M1009_g
+ N_A1_c_108_n N_A1_M1027_g N_A1_M1015_g N_A1_c_118_n N_A1_c_119_n N_A1_c_109_n
+ N_A1_c_121_n N_A1_c_110_n N_A1_c_111_n A1 N_A1_c_113_n
+ PM_SKY130_FD_SC_HD__O22AI_4%A1
x_PM_SKY130_FD_SC_HD__O22AI_4%A2 N_A2_c_237_n N_A2_M1001_g N_A2_M1000_g
+ N_A2_c_238_n N_A2_M1022_g N_A2_M1004_g N_A2_c_239_n N_A2_M1024_g N_A2_M1007_g
+ N_A2_c_240_n N_A2_M1025_g N_A2_M1010_g A2 N_A2_c_241_n N_A2_c_242_n
+ PM_SKY130_FD_SC_HD__O22AI_4%A2
x_PM_SKY130_FD_SC_HD__O22AI_4%B1 N_B1_c_319_n N_B1_M1018_g N_B1_M1003_g
+ N_B1_c_320_n N_B1_M1021_g N_B1_M1008_g N_B1_c_321_n N_B1_M1029_g N_B1_M1020_g
+ N_B1_M1030_g N_B1_M1026_g N_B1_c_331_n N_B1_c_322_n N_B1_c_323_n B1
+ N_B1_c_324_n N_B1_c_325_n N_B1_c_326_n PM_SKY130_FD_SC_HD__O22AI_4%B1
x_PM_SKY130_FD_SC_HD__O22AI_4%B2 N_B2_c_436_n N_B2_M1014_g N_B2_M1006_g
+ N_B2_c_437_n N_B2_M1019_g N_B2_M1011_g N_B2_c_438_n N_B2_M1028_g N_B2_M1012_g
+ N_B2_c_439_n N_B2_M1031_g N_B2_M1016_g B2 N_B2_c_440_n
+ PM_SKY130_FD_SC_HD__O22AI_4%B2
x_PM_SKY130_FD_SC_HD__O22AI_4%VPWR N_VPWR_M1002_s N_VPWR_M1005_s N_VPWR_M1015_s
+ N_VPWR_M1008_s N_VPWR_M1026_s N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n
+ N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n
+ N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n VPWR N_VPWR_c_510_n
+ N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_498_n PM_SKY130_FD_SC_HD__O22AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O22AI_4%A_115_297# N_A_115_297#_M1002_d
+ N_A_115_297#_M1009_d N_A_115_297#_M1004_s N_A_115_297#_M1010_s
+ N_A_115_297#_c_614_n N_A_115_297#_c_639_n N_A_115_297#_c_623_n
+ N_A_115_297#_c_630_n N_A_115_297#_c_646_n N_A_115_297#_c_632_n
+ N_A_115_297#_c_650_n N_A_115_297#_c_629_n
+ PM_SKY130_FD_SC_HD__O22AI_4%A_115_297#
x_PM_SKY130_FD_SC_HD__O22AI_4%Y N_Y_M1018_s N_Y_M1029_s N_Y_M1019_d N_Y_M1031_d
+ N_Y_M1000_d N_Y_M1007_d N_Y_M1006_s N_Y_M1012_s N_Y_c_674_n N_Y_c_675_n
+ N_Y_c_695_n N_Y_c_665_n N_Y_c_666_n N_Y_c_710_n N_Y_c_669_n N_Y_c_667_n
+ N_Y_c_680_n N_Y_c_671_n N_Y_c_683_n N_Y_c_724_n N_Y_c_725_n Y Y
+ PM_SKY130_FD_SC_HD__O22AI_4%Y
x_PM_SKY130_FD_SC_HD__O22AI_4%A_797_297# N_A_797_297#_M1003_d
+ N_A_797_297#_M1020_d N_A_797_297#_M1011_d N_A_797_297#_M1016_d
+ N_A_797_297#_c_800_n N_A_797_297#_c_804_n N_A_797_297#_c_809_n
+ N_A_797_297#_c_822_n N_A_797_297#_c_811_n N_A_797_297#_c_807_n
+ N_A_797_297#_c_808_n N_A_797_297#_c_828_n N_A_797_297#_c_830_n
+ PM_SKY130_FD_SC_HD__O22AI_4%A_797_297#
x_PM_SKY130_FD_SC_HD__O22AI_4%A_33_47# N_A_33_47#_M1013_s N_A_33_47#_M1017_s
+ N_A_33_47#_M1001_d N_A_33_47#_M1024_d N_A_33_47#_M1027_s N_A_33_47#_M1021_d
+ N_A_33_47#_M1014_s N_A_33_47#_M1028_s N_A_33_47#_M1030_d N_A_33_47#_c_847_n
+ N_A_33_47#_c_848_n N_A_33_47#_c_849_n N_A_33_47#_c_866_n N_A_33_47#_c_850_n
+ N_A_33_47#_c_872_n N_A_33_47#_c_851_n N_A_33_47#_c_873_n N_A_33_47#_c_852_n
+ N_A_33_47#_c_878_n N_A_33_47#_c_879_n N_A_33_47#_c_853_n N_A_33_47#_c_854_n
+ N_A_33_47#_c_855_n N_A_33_47#_c_856_n PM_SKY130_FD_SC_HD__O22AI_4%A_33_47#
x_PM_SKY130_FD_SC_HD__O22AI_4%VGND N_VGND_M1013_d N_VGND_M1023_d N_VGND_M1022_s
+ N_VGND_M1025_s N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n
+ N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n
+ N_VGND_c_980_n VGND N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n
+ PM_SKY130_FD_SC_HD__O22AI_4%VGND
cc_1 VNB N_A1_c_105_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_2 VNB N_A1_c_106_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=0.995
cc_3 VNB N_A1_c_107_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.995
cc_4 VNB N_A1_c_108_n 0.0166725f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=0.995
cc_5 VNB N_A1_c_109_n 4.94559e-19 $X=-0.19 $Y=-0.24 $X2=3.425 $Y2=1.445
cc_6 VNB N_A1_c_110_n 0.00338786f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.16
cc_7 VNB N_A1_c_111_n 0.0200608f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.16
cc_8 VNB A1 0.0189511f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_9 VNB N_A1_c_113_n 0.0558437f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=1.16
cc_10 VNB N_A2_c_237_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_11 VNB N_A2_c_238_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=0.995
cc_12 VNB N_A2_c_239_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.995
cc_13 VNB N_A2_c_240_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=0.995
cc_14 VNB N_A2_c_241_n 0.00275279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_242_n 0.0613231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_c_319_n 0.016224f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_17 VNB N_B1_c_320_n 0.0159777f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=0.995
cc_18 VNB N_B1_c_321_n 0.0162467f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.995
cc_19 VNB N_B1_c_322_n 6.43834e-19 $X=-0.19 $Y=-0.24 $X2=1.282 $Y2=1.445
cc_20 VNB N_B1_c_323_n 0.0260784f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.16
cc_21 VNB N_B1_c_324_n 0.049609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B1_c_325_n 0.0195375f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_23 VNB N_B1_c_326_n 0.00296821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_B2_c_436_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_25 VNB N_B2_c_437_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=0.995
cc_26 VNB N_B2_c_438_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.995
cc_27 VNB N_B2_c_439_n 0.0162474f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=0.995
cc_28 VNB N_B2_c_440_n 0.0634264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_498_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_665_n 0.00103009f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=1.53
cc_31 VNB N_Y_c_666_n 0.0086211f $X=-0.19 $Y=-0.24 $X2=3.425 $Y2=1.245
cc_32 VNB N_Y_c_667_n 0.0221948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_33_47#_c_847_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=1.53
cc_34 VNB N_A_33_47#_c_848_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=3.425 $Y2=1.445
cc_35 VNB N_A_33_47#_c_849_n 0.0102929f $X=-0.19 $Y=-0.24 $X2=1.282 $Y2=1.445
cc_36 VNB N_A_33_47#_c_850_n 0.00406612f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.245
cc_37 VNB N_A_33_47#_c_851_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_33_47#_c_852_n 0.0104349f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.16
cc_39 VNB N_A_33_47#_c_853_n 0.0103442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_33_47#_c_854_n 0.00222331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_33_47#_c_855_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_33_47#_c_856_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_971_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.34 $Y2=0.56
cc_44 VNB N_VGND_c_972_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_973_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.325
cc_46 VNB N_VGND_c_974_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=3.275 $Y2=1.53
cc_47 VNB N_VGND_c_975_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=3.425 $Y2=1.445
cc_48 VNB N_VGND_c_976_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=1.282 $Y2=1.445
cc_49 VNB N_VGND_c_977_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.16
cc_50 VNB N_VGND_c_978_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.16
cc_51 VNB N_VGND_c_979_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.245
cc_52 VNB N_VGND_c_980_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_53 VNB N_VGND_c_981_n 0.0936731f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.175
cc_54 VNB N_VGND_c_982_n 0.353813f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_983_n 0.0214165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VPB N_A1_M1002_g 0.0249322f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_57 VPB N_A1_M1005_g 0.0184569f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_58 VPB N_A1_M1009_g 0.0178828f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_59 VPB N_A1_M1015_g 0.0177905f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.985
cc_60 VPB N_A1_c_118_n 0.0135476f $X=-0.19 $Y=1.305 $X2=3.275 $Y2=1.53
cc_61 VPB N_A1_c_119_n 3.01294e-19 $X=-0.19 $Y=1.305 $X2=1.415 $Y2=1.53
cc_62 VPB N_A1_c_109_n 0.00244334f $X=-0.19 $Y=1.305 $X2=3.425 $Y2=1.445
cc_63 VPB N_A1_c_121_n 0.00119441f $X=-0.19 $Y=1.305 $X2=1.282 $Y2=1.445
cc_64 VPB N_A1_c_111_n 0.00455127f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.16
cc_65 VPB N_A1_c_113_n 0.00982609f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.16
cc_66 VPB N_A2_M1000_g 0.0183663f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_67 VPB N_A2_M1004_g 0.01812f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_68 VPB N_A2_M1007_g 0.018119f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_69 VPB N_A2_M1010_g 0.0183572f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.985
cc_70 VPB N_A2_c_242_n 0.0100831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_B1_M1003_g 0.0183913f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_72 VPB N_B1_M1008_g 0.0177586f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_73 VPB N_B1_M1020_g 0.0171878f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_74 VPB N_B1_M1026_g 0.0223541f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.985
cc_75 VPB N_B1_c_331_n 0.012802f $X=-0.19 $Y=1.305 $X2=3.275 $Y2=1.53
cc_76 VPB N_B1_c_322_n 0.00231177f $X=-0.19 $Y=1.305 $X2=1.282 $Y2=1.445
cc_77 VPB N_B1_c_323_n 0.00578485f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.16
cc_78 VPB N_B1_c_324_n 0.00972087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_B1_c_326_n 0.00156635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_B2_M1006_g 0.0183545f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_81 VPB N_B2_M1011_g 0.0181185f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_82 VPB N_B2_M1012_g 0.0181194f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.985
cc_83 VPB N_B2_M1016_g 0.0183603f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.985
cc_84 VPB N_B2_c_440_n 0.0100326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_499_n 0.012247f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.56
cc_86 VPB N_VPWR_c_500_n 0.00873736f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.325
cc_87 VPB N_VPWR_c_501_n 0.00454762f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=0.56
cc_88 VPB N_VPWR_c_502_n 0.00435494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_503_n 0.00455163f $X=-0.19 $Y=1.305 $X2=3.425 $Y2=1.445
cc_90 VPB N_VPWR_c_504_n 0.0119702f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.16
cc_91 VPB N_VPWR_c_505_n 0.0190373f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.16
cc_92 VPB N_VPWR_c_506_n 0.05431f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_93 VPB N_VPWR_c_507_n 0.0041991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_508_n 0.0173603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_509_n 0.00459045f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.16
cc_96 VPB N_VPWR_c_510_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_97 VPB N_VPWR_c_511_n 0.0535132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_512_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_498_n 0.045642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_115_297#_c_614_n 0.00281045f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=0.995
cc_101 VPB N_Y_c_665_n 0.00110481f $X=-0.19 $Y=1.305 $X2=1.415 $Y2=1.53
cc_102 VPB N_Y_c_669_n 0.00865182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_Y_c_667_n 0.0195807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_Y_c_671_n 0.00314618f $X=-0.19 $Y=1.305 $X2=1.34 $Y2=1.16
cc_105 N_A1_c_107_n N_A2_c_237_n 0.0239518f $X=1.34 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_106 N_A1_M1009_g N_A2_M1000_g 0.0239518f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A1_c_118_n N_A2_M1000_g 0.0149047f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_108 N_A1_c_118_n N_A2_M1004_g 0.0103677f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_109 N_A1_c_118_n N_A2_M1007_g 0.0103677f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_110 N_A1_c_108_n N_A2_c_240_n 0.0258191f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A1_M1015_g N_A2_M1010_g 0.0434932f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A1_c_118_n N_A2_M1010_g 0.0103235f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_113 N_A1_c_118_n N_A2_c_241_n 0.0998202f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_114 N_A1_c_110_n N_A2_c_241_n 0.0158542f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A1_c_111_n N_A2_c_241_n 2.34957e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_116 A1 N_A2_c_241_n 0.0115402f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A1_c_113_n N_A2_c_241_n 2.49913e-19 $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A1_c_118_n N_A2_c_242_n 0.00642092f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_119 N_A1_c_109_n N_A2_c_242_n 0.0038846f $X=3.425 $Y=1.445 $X2=0 $Y2=0
cc_120 N_A1_c_121_n N_A2_c_242_n 0.00112116f $X=1.282 $Y=1.445 $X2=0 $Y2=0
cc_121 N_A1_c_110_n N_A2_c_242_n 6.53899e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A1_c_111_n N_A2_c_242_n 0.0225674f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_123 A1 N_A2_c_242_n 2.49913e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A1_c_113_n N_A2_c_242_n 0.0239518f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A1_c_108_n N_B1_c_319_n 0.00984352f $X=3.44 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_126 N_A1_M1015_g N_B1_M1003_g 0.0346017f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A1_c_118_n N_B1_M1003_g 5.59915e-19 $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_128 N_A1_c_109_n N_B1_M1003_g 8.92305e-19 $X=3.425 $Y=1.445 $X2=0 $Y2=0
cc_129 N_A1_c_109_n N_B1_c_324_n 3.7227e-19 $X=3.425 $Y=1.445 $X2=0 $Y2=0
cc_130 N_A1_c_110_n N_B1_c_324_n 0.00141733f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A1_c_111_n N_B1_c_324_n 0.0173674f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A1_c_119_n N_VPWR_M1005_s 0.00209238f $X=1.415 $Y=1.53 $X2=0 $Y2=0
cc_133 N_A1_c_118_n N_VPWR_M1015_s 0.00115961f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_134 N_A1_M1002_g N_VPWR_c_500_n 0.00431697f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_135 A1 N_VPWR_c_500_n 0.0210492f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A1_c_113_n N_VPWR_c_500_n 8.41451e-19 $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_M1005_g N_VPWR_c_501_n 0.00157837f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_M1009_g N_VPWR_c_501_n 0.00302074f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_M1015_g N_VPWR_c_502_n 0.00283367f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_M1009_g N_VPWR_c_506_n 0.00585385f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_M1015_g N_VPWR_c_506_n 0.00541359f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A1_M1002_g N_VPWR_c_510_n 0.00585385f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A1_M1005_g N_VPWR_c_510_n 0.00585385f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A1_M1002_g N_VPWR_c_498_n 0.0114186f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1005_g N_VPWR_c_498_n 0.00588483f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1009_g N_VPWR_c_498_n 0.00591203f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_M1015_g N_VPWR_c_498_n 0.00598342f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A1_c_118_n N_A_115_297#_M1009_d 0.00165831f $X=3.275 $Y=1.53 $X2=0
+ $Y2=0
cc_149 N_A1_c_118_n N_A_115_297#_M1004_s 0.00166235f $X=3.275 $Y=1.53 $X2=0
+ $Y2=0
cc_150 N_A1_c_118_n N_A_115_297#_M1010_s 0.00165255f $X=3.275 $Y=1.53 $X2=0
+ $Y2=0
cc_151 N_A1_M1002_g N_A_115_297#_c_614_n 3.09636e-19 $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1005_g N_A_115_297#_c_614_n 4.03862e-19 $X=0.92 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A1_c_119_n N_A_115_297#_c_614_n 0.00592489f $X=1.415 $Y=1.53 $X2=0
+ $Y2=0
cc_154 A1 N_A_115_297#_c_614_n 0.020226f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A1_c_113_n N_A_115_297#_c_614_n 0.00222737f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A1_M1005_g N_A_115_297#_c_623_n 0.0112521f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A1_M1009_g N_A_115_297#_c_623_n 0.0095558f $X=1.34 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A1_c_118_n N_A_115_297#_c_623_n 0.0126919f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_159 N_A1_c_119_n N_A_115_297#_c_623_n 0.0157651f $X=1.415 $Y=1.53 $X2=0 $Y2=0
cc_160 A1 N_A_115_297#_c_623_n 0.00808474f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A1_c_113_n N_A_115_297#_c_623_n 0.00129797f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A1_M1015_g N_A_115_297#_c_629_n 0.00420836f $X=3.44 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A1_c_118_n N_Y_M1000_d 0.00165831f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_164 N_A1_c_118_n N_Y_M1007_d 0.00165831f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A1_c_118_n N_Y_c_674_n 0.0315971f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A1_M1015_g N_Y_c_675_n 0.00331717f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_c_108_n N_Y_c_665_n 4.65391e-19 $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_109_n N_Y_c_665_n 0.00785664f $X=3.425 $Y=1.445 $X2=0 $Y2=0
cc_169 N_A1_c_110_n N_Y_c_665_n 0.00751516f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A1_c_111_n N_Y_c_665_n 8.46851e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A1_c_118_n N_Y_c_680_n 0.0120079f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_172 N_A1_M1015_g N_Y_c_671_n 5.38459e-19 $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A1_c_118_n N_Y_c_671_n 0.0146501f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_174 N_A1_M1015_g N_Y_c_683_n 0.0115507f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A1_c_118_n N_Y_c_683_n 0.0331153f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A1_c_110_n N_Y_c_683_n 9.38486e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A1_c_111_n N_Y_c_683_n 2.9763e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A1_c_118_n Y 0.0120079f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_179 N_A1_c_105_n N_A_33_47#_c_847_n 0.00630972f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_106_n N_A_33_47#_c_847_n 5.22228e-19 $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_105_n N_A_33_47#_c_848_n 0.00870364f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_106_n N_A_33_47#_c_848_n 0.00870364f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_183 A1 N_A_33_47#_c_848_n 0.036111f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A1_c_113_n N_A_33_47#_c_848_n 0.00222133f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A1_c_105_n N_A_33_47#_c_849_n 0.00129539f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_186 A1 N_A_33_47#_c_849_n 0.0276561f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A1_c_113_n N_A_33_47#_c_849_n 0.00115169f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A1_c_105_n N_A_33_47#_c_866_n 5.22228e-19 $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_106_n N_A_33_47#_c_866_n 0.00630972f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A1_c_107_n N_A_33_47#_c_866_n 0.00630972f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A1_c_107_n N_A_33_47#_c_850_n 0.00845282f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_118_n N_A_33_47#_c_850_n 0.00911016f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_193 A1 N_A_33_47#_c_850_n 0.00893273f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_194 N_A1_c_107_n N_A_33_47#_c_872_n 5.22228e-19 $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_108_n N_A_33_47#_c_873_n 5.22228e-19 $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_108_n N_A_33_47#_c_852_n 0.00955706f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_118_n N_A_33_47#_c_852_n 0.0060678f $X=3.275 $Y=1.53 $X2=0 $Y2=0
cc_198 N_A1_c_110_n N_A_33_47#_c_852_n 0.026225f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A1_c_111_n N_A_33_47#_c_852_n 0.00301245f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A1_c_108_n N_A_33_47#_c_878_n 0.00255288f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_108_n N_A_33_47#_c_879_n 0.00393886f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A1_c_106_n N_A_33_47#_c_854_n 0.00113286f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_107_n N_A_33_47#_c_854_n 0.00127865f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_204 A1 N_A_33_47#_c_854_n 0.0273972f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_205 N_A1_c_113_n N_A_33_47#_c_854_n 0.00230291f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A1_c_105_n N_VGND_c_971_n 0.00268723f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_c_106_n N_VGND_c_971_n 0.00146448f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A1_c_107_n N_VGND_c_972_n 0.00146448f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_108_n N_VGND_c_974_n 0.00268723f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_106_n N_VGND_c_975_n 0.00423334f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A1_c_107_n N_VGND_c_975_n 0.00424416f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A1_c_108_n N_VGND_c_981_n 0.00422898f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A1_c_105_n N_VGND_c_982_n 0.00669811f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A1_c_106_n N_VGND_c_982_n 0.0057163f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A1_c_107_n N_VGND_c_982_n 0.00576327f $X=1.34 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A1_c_108_n N_VGND_c_982_n 0.00591777f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A1_c_105_n N_VGND_c_983_n 0.00423334f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A2_M1000_g N_VPWR_c_506_n 0.00357877f $X=1.76 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A2_M1004_g N_VPWR_c_506_n 0.00357877f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A2_M1007_g N_VPWR_c_506_n 0.00357877f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A2_M1010_g N_VPWR_c_506_n 0.00357877f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A2_M1000_g N_VPWR_c_498_n 0.00525237f $X=1.76 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A2_M1004_g N_VPWR_c_498_n 0.00522516f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A2_M1007_g N_VPWR_c_498_n 0.00522516f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A2_M1010_g N_VPWR_c_498_n 0.00525237f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A2_M1000_g N_A_115_297#_c_630_n 0.0121306f $X=1.76 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A2_M1004_g N_A_115_297#_c_630_n 0.00851673f $X=2.18 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A2_M1007_g N_A_115_297#_c_632_n 0.00851673f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A2_M1010_g N_A_115_297#_c_632_n 0.00851673f $X=3.02 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A2_M1004_g N_Y_c_674_n 0.00924026f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A2_M1007_g N_Y_c_674_n 0.00924026f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A2_M1010_g N_Y_c_683_n 0.00924026f $X=3.02 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A2_c_237_n N_A_33_47#_c_866_n 5.22228e-19 $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_237_n N_A_33_47#_c_850_n 0.00845772f $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_241_n N_A_33_47#_c_850_n 0.00820272f $X=2.93 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A2_c_237_n N_A_33_47#_c_872_n 0.00630972f $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A2_c_238_n N_A_33_47#_c_872_n 0.00630972f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A2_c_239_n N_A_33_47#_c_872_n 5.22228e-19 $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A2_c_238_n N_A_33_47#_c_851_n 0.00870364f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_239_n N_A_33_47#_c_851_n 0.00870364f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A2_c_241_n N_A_33_47#_c_851_n 0.036111f $X=2.93 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A2_c_242_n N_A_33_47#_c_851_n 0.00222133f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A2_c_238_n N_A_33_47#_c_873_n 5.22228e-19 $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A2_c_239_n N_A_33_47#_c_873_n 0.00630972f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A2_c_240_n N_A_33_47#_c_873_n 0.00630972f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A2_c_240_n N_A_33_47#_c_852_n 0.00845772f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A2_c_241_n N_A_33_47#_c_852_n 0.00820272f $X=2.93 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A2_c_240_n N_A_33_47#_c_879_n 4.86829e-19 $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A2_c_237_n N_A_33_47#_c_855_n 0.00127992f $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A2_c_238_n N_A_33_47#_c_855_n 0.00113286f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A2_c_241_n N_A_33_47#_c_855_n 0.0265405f $X=2.93 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A2_c_242_n N_A_33_47#_c_855_n 0.00230339f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A2_c_239_n N_A_33_47#_c_856_n 0.00113286f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A2_c_240_n N_A_33_47#_c_856_n 0.00128009f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A2_c_241_n N_A_33_47#_c_856_n 0.0265405f $X=2.93 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A2_c_242_n N_A_33_47#_c_856_n 0.00230339f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A2_c_237_n N_VGND_c_972_n 0.00146448f $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A2_c_238_n N_VGND_c_973_n 0.00146448f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A2_c_239_n N_VGND_c_973_n 0.00146448f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A2_c_240_n N_VGND_c_974_n 0.00146448f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A2_c_237_n N_VGND_c_977_n 0.00424416f $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A2_c_238_n N_VGND_c_977_n 0.00423334f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A2_c_239_n N_VGND_c_979_n 0.00423334f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A2_c_240_n N_VGND_c_979_n 0.00424416f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A2_c_237_n N_VGND_c_982_n 0.00576327f $X=1.76 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A2_c_238_n N_VGND_c_982_n 0.0057163f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A2_c_239_n N_VGND_c_982_n 0.0057163f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A2_c_240_n N_VGND_c_982_n 0.00576327f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B1_c_321_n N_B2_c_436_n 0.0271098f $X=4.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_270 N_B1_M1020_g N_B2_M1006_g 0.0277573f $X=4.75 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B1_c_331_n N_B2_M1006_g 0.0151175f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_272 N_B1_c_331_n N_B2_M1011_g 0.0103677f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_273 N_B1_c_331_n N_B2_M1012_g 0.0103677f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_274 N_B1_c_325_n N_B2_c_439_n 0.0267447f $X=6.865 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B1_M1026_g N_B2_M1016_g 0.0434538f $X=6.85 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B1_c_331_n N_B2_M1016_g 0.0109619f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_277 N_B1_c_322_n N_B2_M1016_g 0.00245342f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_278 N_B1_c_331_n B2 0.0957019f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_279 N_B1_c_322_n B2 0.0110886f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B1_c_323_n B2 6.32117e-19 $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_281 N_B1_c_324_n B2 2.11472e-19 $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_282 N_B1_c_326_n B2 0.0175788f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_283 N_B1_c_331_n N_B2_c_440_n 0.00642092f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_284 N_B1_c_322_n N_B2_c_440_n 0.00184556f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B1_c_323_n N_B2_c_440_n 0.0221893f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B1_c_324_n N_B2_c_440_n 0.0219214f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_287 N_B1_c_326_n N_B2_c_440_n 0.00826833f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_288 N_B1_c_326_n N_VPWR_M1008_s 0.00172977f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_289 N_B1_M1003_g N_VPWR_c_502_n 0.00153693f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_290 N_B1_M1008_g N_VPWR_c_503_n 0.00159538f $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_291 N_B1_M1020_g N_VPWR_c_503_n 0.00300811f $X=4.75 $Y=1.985 $X2=0 $Y2=0
cc_292 N_B1_M1026_g N_VPWR_c_505_n 0.00485906f $X=6.85 $Y=1.985 $X2=0 $Y2=0
cc_293 N_B1_M1003_g N_VPWR_c_508_n 0.00541359f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_294 N_B1_M1008_g N_VPWR_c_508_n 0.00585385f $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_295 N_B1_M1020_g N_VPWR_c_511_n 0.00585385f $X=4.75 $Y=1.985 $X2=0 $Y2=0
cc_296 N_B1_M1026_g N_VPWR_c_511_n 0.00585385f $X=6.85 $Y=1.985 $X2=0 $Y2=0
cc_297 N_B1_M1003_g N_VPWR_c_498_n 0.0072159f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_298 N_B1_M1008_g N_VPWR_c_498_n 0.00590992f $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_299 N_B1_M1020_g N_VPWR_c_498_n 0.00591203f $X=4.75 $Y=1.985 $X2=0 $Y2=0
cc_300 N_B1_M1026_g N_VPWR_c_498_n 0.0069025f $X=6.85 $Y=1.985 $X2=0 $Y2=0
cc_301 N_B1_c_331_n N_Y_M1006_s 0.00165831f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_302 N_B1_c_331_n N_Y_M1012_s 0.00165831f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_303 N_B1_M1003_g N_Y_c_675_n 0.00496693f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_304 N_B1_M1008_g N_Y_c_675_n 9.3226e-19 $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_305 N_B1_c_319_n N_Y_c_695_n 0.00226162f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B1_c_319_n N_Y_c_665_n 0.0032387f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_M1003_g N_Y_c_665_n 0.00273282f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_308 N_B1_c_320_n N_Y_c_665_n 0.00353216f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B1_M1008_g N_Y_c_665_n 7.00148e-19 $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_310 N_B1_c_324_n N_Y_c_665_n 0.0156975f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_311 N_B1_c_326_n N_Y_c_665_n 0.0344578f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_312 N_B1_c_320_n N_Y_c_666_n 0.00971041f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B1_c_321_n N_Y_c_666_n 0.00852218f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B1_c_331_n N_Y_c_666_n 0.0103306f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_315 N_B1_c_322_n N_Y_c_666_n 0.0138956f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_316 N_B1_c_323_n N_Y_c_666_n 0.0024893f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_317 N_B1_c_324_n N_Y_c_666_n 0.00470837f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_318 N_B1_c_325_n N_Y_c_666_n 0.0101218f $X=6.865 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B1_c_326_n N_Y_c_666_n 0.0425389f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_320 N_B1_c_331_n N_Y_c_710_n 0.0315971f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_321 N_B1_M1026_g N_Y_c_669_n 0.0131107f $X=6.85 $Y=1.985 $X2=0 $Y2=0
cc_322 N_B1_c_331_n N_Y_c_669_n 0.0327907f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_323 N_B1_c_323_n N_Y_c_669_n 0.00177598f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_324 N_B1_M1026_g N_Y_c_667_n 0.00776159f $X=6.85 $Y=1.985 $X2=0 $Y2=0
cc_325 N_B1_c_331_n N_Y_c_667_n 0.00807294f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_326 N_B1_c_322_n N_Y_c_667_n 0.0332285f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_327 N_B1_c_323_n N_Y_c_667_n 0.00797697f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_328 N_B1_c_325_n N_Y_c_667_n 0.00589321f $X=6.865 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B1_M1003_g N_Y_c_671_n 0.0129404f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_330 N_B1_M1008_g N_Y_c_671_n 0.00106596f $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_331 N_B1_c_324_n N_Y_c_671_n 2.90548e-19 $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_332 N_B1_c_326_n N_Y_c_671_n 0.0141181f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_333 N_B1_M1003_g N_Y_c_683_n 0.00642799f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_334 N_B1_c_331_n N_Y_c_724_n 0.0120079f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_335 N_B1_c_331_n N_Y_c_725_n 0.0120079f $X=6.715 $Y=1.53 $X2=0 $Y2=0
cc_336 N_B1_c_331_n N_A_797_297#_M1020_d 0.00103113f $X=6.715 $Y=1.53 $X2=0
+ $Y2=0
cc_337 N_B1_c_326_n N_A_797_297#_M1020_d 6.41547e-19 $X=4.94 $Y=1.305 $X2=0
+ $Y2=0
cc_338 N_B1_c_331_n N_A_797_297#_M1011_d 0.00166235f $X=6.715 $Y=1.53 $X2=0
+ $Y2=0
cc_339 N_B1_c_331_n N_A_797_297#_M1016_d 0.00161973f $X=6.715 $Y=1.53 $X2=0
+ $Y2=0
cc_340 N_B1_M1008_g N_A_797_297#_c_800_n 0.0107531f $X=4.33 $Y=1.985 $X2=0 $Y2=0
cc_341 N_B1_M1020_g N_A_797_297#_c_800_n 0.00956194f $X=4.75 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_B1_c_324_n N_A_797_297#_c_800_n 4.63201e-19 $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_343 N_B1_c_326_n N_A_797_297#_c_800_n 0.0451651f $X=4.94 $Y=1.305 $X2=0 $Y2=0
cc_344 N_B1_M1003_g N_A_797_297#_c_804_n 0.00122697f $X=3.91 $Y=1.985 $X2=0
+ $Y2=0
cc_345 N_B1_M1008_g N_A_797_297#_c_804_n 0.00128716f $X=4.33 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_B1_c_324_n N_A_797_297#_c_804_n 0.00131736f $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_347 N_B1_M1003_g N_A_797_297#_c_807_n 0.00453735f $X=3.91 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_B1_M1003_g N_A_797_297#_c_808_n 0.00370075f $X=3.91 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_B1_c_319_n N_A_33_47#_c_853_n 0.0127015f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_350 N_B1_c_320_n N_A_33_47#_c_853_n 0.00892725f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_351 N_B1_c_321_n N_A_33_47#_c_853_n 0.00886996f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_352 N_B1_c_324_n N_A_33_47#_c_853_n 2.31645e-19 $X=4.75 $Y=1.16 $X2=0 $Y2=0
cc_353 N_B1_c_325_n N_A_33_47#_c_853_n 0.00886996f $X=6.865 $Y=0.995 $X2=0 $Y2=0
cc_354 N_B1_c_319_n N_VGND_c_981_n 0.00357877f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_355 N_B1_c_320_n N_VGND_c_981_n 0.00357877f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_356 N_B1_c_321_n N_VGND_c_981_n 0.00357877f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_357 N_B1_c_325_n N_VGND_c_981_n 0.00357877f $X=6.865 $Y=0.995 $X2=0 $Y2=0
cc_358 N_B1_c_319_n N_VGND_c_982_n 0.00537058f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_359 N_B1_c_320_n N_VGND_c_982_n 0.00522516f $X=4.33 $Y=0.995 $X2=0 $Y2=0
cc_360 N_B1_c_321_n N_VGND_c_982_n 0.00525341f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_361 N_B1_c_325_n N_VGND_c_982_n 0.00624388f $X=6.865 $Y=0.995 $X2=0 $Y2=0
cc_362 N_B2_M1006_g N_VPWR_c_511_n 0.00357877f $X=5.17 $Y=1.985 $X2=0 $Y2=0
cc_363 N_B2_M1011_g N_VPWR_c_511_n 0.00357877f $X=5.59 $Y=1.985 $X2=0 $Y2=0
cc_364 N_B2_M1012_g N_VPWR_c_511_n 0.00357877f $X=6.01 $Y=1.985 $X2=0 $Y2=0
cc_365 N_B2_M1016_g N_VPWR_c_511_n 0.00357877f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_366 N_B2_M1006_g N_VPWR_c_498_n 0.00525237f $X=5.17 $Y=1.985 $X2=0 $Y2=0
cc_367 N_B2_M1011_g N_VPWR_c_498_n 0.00522516f $X=5.59 $Y=1.985 $X2=0 $Y2=0
cc_368 N_B2_M1012_g N_VPWR_c_498_n 0.00522516f $X=6.01 $Y=1.985 $X2=0 $Y2=0
cc_369 N_B2_M1016_g N_VPWR_c_498_n 0.00525237f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_370 N_B2_c_436_n N_Y_c_666_n 0.00913856f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_371 N_B2_c_437_n N_Y_c_666_n 0.00898612f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_372 N_B2_c_438_n N_Y_c_666_n 0.00898612f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_373 N_B2_c_439_n N_Y_c_666_n 0.00946523f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_374 B2 N_Y_c_666_n 0.0598376f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_375 N_B2_c_440_n N_Y_c_666_n 0.00628591f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_376 N_B2_M1011_g N_Y_c_710_n 0.00924026f $X=5.59 $Y=1.985 $X2=0 $Y2=0
cc_377 N_B2_M1012_g N_Y_c_710_n 0.00924026f $X=6.01 $Y=1.985 $X2=0 $Y2=0
cc_378 N_B2_M1016_g N_Y_c_669_n 0.00924026f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_379 N_B2_M1006_g N_A_797_297#_c_809_n 0.0121306f $X=5.17 $Y=1.985 $X2=0 $Y2=0
cc_380 N_B2_M1011_g N_A_797_297#_c_809_n 0.00851673f $X=5.59 $Y=1.985 $X2=0
+ $Y2=0
cc_381 N_B2_M1012_g N_A_797_297#_c_811_n 0.00851673f $X=6.01 $Y=1.985 $X2=0
+ $Y2=0
cc_382 N_B2_M1016_g N_A_797_297#_c_811_n 0.00851673f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_383 N_B2_c_436_n N_A_33_47#_c_853_n 0.00886996f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_384 N_B2_c_437_n N_A_33_47#_c_853_n 0.00892725f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_385 N_B2_c_438_n N_A_33_47#_c_853_n 0.00892725f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_386 N_B2_c_439_n N_A_33_47#_c_853_n 0.00886996f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_387 N_B2_c_436_n N_VGND_c_981_n 0.00357877f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_388 N_B2_c_437_n N_VGND_c_981_n 0.00357877f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_389 N_B2_c_438_n N_VGND_c_981_n 0.00357877f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_390 N_B2_c_439_n N_VGND_c_981_n 0.00357877f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_391 N_B2_c_436_n N_VGND_c_982_n 0.00525341f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_392 N_B2_c_437_n N_VGND_c_982_n 0.00522516f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_393 N_B2_c_438_n N_VGND_c_982_n 0.00522516f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_394 N_B2_c_439_n N_VGND_c_982_n 0.00525341f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_395 N_VPWR_c_498_n N_A_115_297#_M1002_d 0.00254126f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_396 N_VPWR_c_498_n N_A_115_297#_M1009_d 0.00220214f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_498_n N_A_115_297#_M1004_s 0.00213597f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_498_n N_A_115_297#_M1010_s 0.00214399f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_500_n N_A_115_297#_c_614_n 0.00311153f $X=0.29 $Y=1.62 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_510_n N_A_115_297#_c_639_n 0.0142343f $X=1.005 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_498_n N_A_115_297#_c_639_n 0.00955092f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_M1005_s N_A_115_297#_c_623_n 0.00378557f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_501_n N_A_115_297#_c_623_n 0.0123301f $X=1.13 $Y=2.3 $X2=0 $Y2=0
cc_404 N_VPWR_c_498_n N_A_115_297#_c_623_n 0.0109281f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_506_n N_A_115_297#_c_630_n 0.0330174f $X=3.565 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_498_n N_A_115_297#_c_630_n 0.0204667f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_506_n N_A_115_297#_c_646_n 0.0143053f $X=3.565 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_498_n N_A_115_297#_c_646_n 0.00962794f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_506_n N_A_115_297#_c_632_n 0.0330174f $X=3.565 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_498_n N_A_115_297#_c_632_n 0.0204707f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_506_n N_A_115_297#_c_650_n 0.0137033f $X=3.565 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_498_n N_A_115_297#_c_650_n 0.00938745f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_506_n N_A_115_297#_c_629_n 0.0159465f $X=3.565 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_498_n N_A_115_297#_c_629_n 0.0106981f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_498_n N_Y_M1000_d 0.0021603f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_498_n N_Y_M1007_d 0.00215227f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_498_n N_Y_M1006_s 0.0021603f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_498_n N_Y_M1012_s 0.00215227f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_419 N_VPWR_c_498_n N_Y_c_674_n 0.00127799f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_M1015_s N_Y_c_675_n 0.00214305f $X=3.515 $Y=1.485 $X2=0 $Y2=0
cc_421 N_VPWR_c_498_n N_Y_c_710_n 0.00127799f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_M1026_s N_Y_c_669_n 0.00676748f $X=6.925 $Y=1.485 $X2=0 $Y2=0
cc_423 N_VPWR_c_504_n N_Y_c_669_n 9.43314e-19 $X=7.075 $Y=2.635 $X2=0 $Y2=0
cc_424 N_VPWR_c_505_n N_Y_c_669_n 0.0192638f $X=7.06 $Y=2.3 $X2=0 $Y2=0
cc_425 N_VPWR_c_498_n N_Y_c_669_n 0.00867427f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_M1026_s N_Y_c_667_n 0.00435292f $X=6.925 $Y=1.485 $X2=0 $Y2=0
cc_427 N_VPWR_M1015_s N_Y_c_671_n 0.00122049f $X=3.515 $Y=1.485 $X2=0 $Y2=0
cc_428 N_VPWR_M1015_s N_Y_c_683_n 0.00798796f $X=3.515 $Y=1.485 $X2=0 $Y2=0
cc_429 N_VPWR_c_502_n N_Y_c_683_n 0.0163894f $X=3.69 $Y=2.3 $X2=0 $Y2=0
cc_430 N_VPWR_c_498_n N_Y_c_683_n 0.0114731f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_c_498_n N_A_797_297#_M1003_d 0.00215201f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_432 N_VPWR_c_498_n N_A_797_297#_M1020_d 0.00220214f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_498_n N_A_797_297#_M1011_d 0.00213597f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_498_n N_A_797_297#_M1016_d 0.00219968f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_435 N_VPWR_M1008_s N_A_797_297#_c_800_n 0.00317012f $X=4.405 $Y=1.485 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_503_n N_A_797_297#_c_800_n 0.0123301f $X=4.54 $Y=2.3 $X2=0 $Y2=0
cc_437 N_VPWR_c_498_n N_A_797_297#_c_800_n 0.0109456f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_511_n N_A_797_297#_c_809_n 0.0330174f $X=6.935 $Y=2.72 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_498_n N_A_797_297#_c_809_n 0.0204667f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_511_n N_A_797_297#_c_822_n 0.0143053f $X=6.935 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_498_n N_A_797_297#_c_822_n 0.00962794f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_511_n N_A_797_297#_c_811_n 0.0330174f $X=6.935 $Y=2.72 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_498_n N_A_797_297#_c_811_n 0.0204707f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_508_n N_A_797_297#_c_807_n 0.0166859f $X=4.425 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_498_n N_A_797_297#_c_807_n 0.011188f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_c_511_n N_A_797_297#_c_828_n 0.0137033f $X=6.935 $Y=2.72 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_498_n N_A_797_297#_c_828_n 0.00938745f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_511_n N_A_797_297#_c_830_n 0.0136817f $X=6.935 $Y=2.72 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_498_n N_A_797_297#_c_830_n 0.00938089f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_450 N_A_115_297#_c_630_n N_Y_M1000_d 0.00312348f $X=2.265 $Y=2.38 $X2=0 $Y2=0
cc_451 N_A_115_297#_c_632_n N_Y_M1007_d 0.00312348f $X=3.105 $Y=2.38 $X2=0 $Y2=0
cc_452 N_A_115_297#_M1004_s N_Y_c_674_n 0.00317012f $X=2.255 $Y=1.485 $X2=0
+ $Y2=0
cc_453 N_A_115_297#_c_630_n N_Y_c_674_n 0.00506389f $X=2.265 $Y=2.38 $X2=0 $Y2=0
cc_454 N_A_115_297#_c_632_n N_Y_c_674_n 0.00506389f $X=3.105 $Y=2.38 $X2=0 $Y2=0
cc_455 N_A_115_297#_c_650_n N_Y_c_674_n 0.0116461f $X=2.39 $Y=2.3 $X2=0 $Y2=0
cc_456 N_A_115_297#_c_630_n N_Y_c_680_n 0.0112811f $X=2.265 $Y=2.38 $X2=0 $Y2=0
cc_457 N_A_115_297#_M1010_s N_Y_c_683_n 0.00325521f $X=3.095 $Y=1.485 $X2=0
+ $Y2=0
cc_458 N_A_115_297#_c_632_n N_Y_c_683_n 0.00506389f $X=3.105 $Y=2.38 $X2=0 $Y2=0
cc_459 N_A_115_297#_c_629_n N_Y_c_683_n 0.0136322f $X=3.23 $Y=2.3 $X2=0 $Y2=0
cc_460 N_A_115_297#_c_632_n Y 0.0112811f $X=3.105 $Y=2.38 $X2=0 $Y2=0
cc_461 N_Y_c_671_n N_A_797_297#_M1003_d 0.00229744f $X=4.04 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_462 N_Y_c_710_n N_A_797_297#_M1011_d 0.00317012f $X=6.095 $Y=1.87 $X2=0 $Y2=0
cc_463 N_Y_c_669_n N_A_797_297#_M1016_d 0.00329438f $X=7.105 $Y=1.87 $X2=0 $Y2=0
cc_464 N_Y_c_671_n N_A_797_297#_c_804_n 0.00325434f $X=4.04 $Y=1.53 $X2=0 $Y2=0
cc_465 N_Y_c_683_n N_A_797_297#_c_804_n 0.0148586f $X=3.745 $Y=1.87 $X2=0 $Y2=0
cc_466 N_Y_M1006_s N_A_797_297#_c_809_n 0.00312348f $X=5.245 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_Y_c_710_n N_A_797_297#_c_809_n 0.00506389f $X=6.095 $Y=1.87 $X2=0 $Y2=0
cc_468 N_Y_c_724_n N_A_797_297#_c_809_n 0.0112811f $X=5.38 $Y=1.87 $X2=0 $Y2=0
cc_469 N_Y_M1012_s N_A_797_297#_c_811_n 0.00312348f $X=6.085 $Y=1.485 $X2=0
+ $Y2=0
cc_470 N_Y_c_710_n N_A_797_297#_c_811_n 0.00506389f $X=6.095 $Y=1.87 $X2=0 $Y2=0
cc_471 N_Y_c_669_n N_A_797_297#_c_811_n 0.00506389f $X=7.105 $Y=1.87 $X2=0 $Y2=0
cc_472 N_Y_c_725_n N_A_797_297#_c_811_n 0.0112811f $X=6.22 $Y=1.87 $X2=0 $Y2=0
cc_473 N_Y_c_671_n N_A_797_297#_c_807_n 0.00229493f $X=4.04 $Y=1.53 $X2=0 $Y2=0
cc_474 N_Y_c_710_n N_A_797_297#_c_828_n 0.0116461f $X=6.095 $Y=1.87 $X2=0 $Y2=0
cc_475 N_Y_c_669_n N_A_797_297#_c_830_n 0.0110749f $X=7.105 $Y=1.87 $X2=0 $Y2=0
cc_476 N_Y_c_666_n N_A_33_47#_M1021_d 0.00307941f $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_477 N_Y_c_666_n N_A_33_47#_M1014_s 0.00333526f $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_478 N_Y_c_666_n N_A_33_47#_M1028_s 0.00333526f $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_479 N_Y_c_666_n N_A_33_47#_M1030_d 0.00667482f $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_480 N_Y_c_667_n N_A_33_47#_M1030_d 9.98841e-19 $X=7.19 $Y=1.785 $X2=0 $Y2=0
cc_481 N_Y_c_665_n N_A_33_47#_c_852_n 0.00374607f $X=4.04 $Y=1.445 $X2=0 $Y2=0
cc_482 N_Y_c_671_n N_A_33_47#_c_852_n 0.00150667f $X=4.04 $Y=1.53 $X2=0 $Y2=0
cc_483 N_Y_M1018_s N_A_33_47#_c_853_n 0.00303872f $X=3.985 $Y=0.235 $X2=0 $Y2=0
cc_484 N_Y_M1029_s N_A_33_47#_c_853_n 0.00312026f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_485 N_Y_M1019_d N_A_33_47#_c_853_n 0.00305026f $X=5.665 $Y=0.235 $X2=0 $Y2=0
cc_486 N_Y_M1031_d N_A_33_47#_c_853_n 0.00313101f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_487 N_Y_c_695_n N_A_33_47#_c_853_n 0.00867341f $X=4.04 $Y=0.82 $X2=0 $Y2=0
cc_488 N_Y_c_666_n N_A_33_47#_c_853_n 0.159818f $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_489 N_Y_c_666_n N_VGND_c_981_n 5.96728e-19 $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_490 N_Y_M1018_s N_VGND_c_982_n 0.00216833f $X=3.985 $Y=0.235 $X2=0 $Y2=0
cc_491 N_Y_M1029_s N_VGND_c_982_n 0.00216833f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_492 N_Y_M1019_d N_VGND_c_982_n 0.00216833f $X=5.665 $Y=0.235 $X2=0 $Y2=0
cc_493 N_Y_M1031_d N_VGND_c_982_n 0.00216833f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_494 N_Y_c_666_n N_VGND_c_982_n 0.00124674f $X=7.105 $Y=0.732 $X2=0 $Y2=0
cc_495 N_A_33_47#_c_848_n N_VGND_M1013_d 0.00162089f $X=0.965 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_496 N_A_33_47#_c_850_n N_VGND_M1023_d 0.00165819f $X=1.805 $Y=0.82 $X2=0
+ $Y2=0
cc_497 N_A_33_47#_c_851_n N_VGND_M1022_s 0.00162089f $X=2.645 $Y=0.815 $X2=0
+ $Y2=0
cc_498 N_A_33_47#_c_852_n N_VGND_M1025_s 0.00165819f $X=3.485 $Y=0.82 $X2=0
+ $Y2=0
cc_499 N_A_33_47#_c_848_n N_VGND_c_971_n 0.0122559f $X=0.965 $Y=0.815 $X2=0
+ $Y2=0
cc_500 N_A_33_47#_c_850_n N_VGND_c_972_n 0.0116529f $X=1.805 $Y=0.82 $X2=0 $Y2=0
cc_501 N_A_33_47#_c_851_n N_VGND_c_973_n 0.0122559f $X=2.645 $Y=0.815 $X2=0
+ $Y2=0
cc_502 N_A_33_47#_c_852_n N_VGND_c_974_n 0.0116528f $X=3.485 $Y=0.82 $X2=0 $Y2=0
cc_503 N_A_33_47#_c_848_n N_VGND_c_975_n 0.00198695f $X=0.965 $Y=0.815 $X2=0
+ $Y2=0
cc_504 N_A_33_47#_c_866_n N_VGND_c_975_n 0.0188551f $X=1.13 $Y=0.39 $X2=0 $Y2=0
cc_505 N_A_33_47#_c_850_n N_VGND_c_975_n 0.00193763f $X=1.805 $Y=0.82 $X2=0
+ $Y2=0
cc_506 N_A_33_47#_c_850_n N_VGND_c_977_n 0.00193763f $X=1.805 $Y=0.82 $X2=0
+ $Y2=0
cc_507 N_A_33_47#_c_872_n N_VGND_c_977_n 0.0188551f $X=1.97 $Y=0.39 $X2=0 $Y2=0
cc_508 N_A_33_47#_c_851_n N_VGND_c_977_n 0.00198695f $X=2.645 $Y=0.815 $X2=0
+ $Y2=0
cc_509 N_A_33_47#_c_851_n N_VGND_c_979_n 0.00198695f $X=2.645 $Y=0.815 $X2=0
+ $Y2=0
cc_510 N_A_33_47#_c_873_n N_VGND_c_979_n 0.0188551f $X=2.81 $Y=0.39 $X2=0 $Y2=0
cc_511 N_A_33_47#_c_852_n N_VGND_c_979_n 0.00193763f $X=3.485 $Y=0.82 $X2=0
+ $Y2=0
cc_512 N_A_33_47#_c_852_n N_VGND_c_981_n 0.00193763f $X=3.485 $Y=0.82 $X2=0
+ $Y2=0
cc_513 N_A_33_47#_c_878_n N_VGND_c_981_n 0.0187152f $X=3.635 $Y=0.475 $X2=0
+ $Y2=0
cc_514 N_A_33_47#_c_853_n N_VGND_c_981_n 0.194257f $X=7.06 $Y=0.39 $X2=0 $Y2=0
cc_515 N_A_33_47#_M1013_s N_VGND_c_982_n 0.00209319f $X=0.165 $Y=0.235 $X2=0
+ $Y2=0
cc_516 N_A_33_47#_M1017_s N_VGND_c_982_n 0.00215201f $X=0.995 $Y=0.235 $X2=0
+ $Y2=0
cc_517 N_A_33_47#_M1001_d N_VGND_c_982_n 0.00215201f $X=1.835 $Y=0.235 $X2=0
+ $Y2=0
cc_518 N_A_33_47#_M1024_d N_VGND_c_982_n 0.00215201f $X=2.675 $Y=0.235 $X2=0
+ $Y2=0
cc_519 N_A_33_47#_M1027_s N_VGND_c_982_n 0.00255355f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_520 N_A_33_47#_M1021_d N_VGND_c_982_n 0.00215227f $X=4.405 $Y=0.235 $X2=0
+ $Y2=0
cc_521 N_A_33_47#_M1014_s N_VGND_c_982_n 0.00215227f $X=5.245 $Y=0.235 $X2=0
+ $Y2=0
cc_522 N_A_33_47#_M1028_s N_VGND_c_982_n 0.00215227f $X=6.085 $Y=0.235 $X2=0
+ $Y2=0
cc_523 N_A_33_47#_M1030_d N_VGND_c_982_n 0.00209344f $X=6.925 $Y=0.235 $X2=0
+ $Y2=0
cc_524 N_A_33_47#_c_847_n N_VGND_c_982_n 0.0124119f $X=0.29 $Y=0.39 $X2=0 $Y2=0
cc_525 N_A_33_47#_c_848_n N_VGND_c_982_n 0.00835832f $X=0.965 $Y=0.815 $X2=0
+ $Y2=0
cc_526 N_A_33_47#_c_866_n N_VGND_c_982_n 0.0122069f $X=1.13 $Y=0.39 $X2=0 $Y2=0
cc_527 N_A_33_47#_c_850_n N_VGND_c_982_n 0.00827287f $X=1.805 $Y=0.82 $X2=0
+ $Y2=0
cc_528 N_A_33_47#_c_872_n N_VGND_c_982_n 0.0122069f $X=1.97 $Y=0.39 $X2=0 $Y2=0
cc_529 N_A_33_47#_c_851_n N_VGND_c_982_n 0.00835832f $X=2.645 $Y=0.815 $X2=0
+ $Y2=0
cc_530 N_A_33_47#_c_873_n N_VGND_c_982_n 0.0122069f $X=2.81 $Y=0.39 $X2=0 $Y2=0
cc_531 N_A_33_47#_c_852_n N_VGND_c_982_n 0.00827287f $X=3.485 $Y=0.82 $X2=0
+ $Y2=0
cc_532 N_A_33_47#_c_878_n N_VGND_c_982_n 0.0113303f $X=3.635 $Y=0.475 $X2=0
+ $Y2=0
cc_533 N_A_33_47#_c_853_n N_VGND_c_982_n 0.123555f $X=7.06 $Y=0.39 $X2=0 $Y2=0
cc_534 N_A_33_47#_c_847_n N_VGND_c_983_n 0.0209752f $X=0.29 $Y=0.39 $X2=0 $Y2=0
cc_535 N_A_33_47#_c_848_n N_VGND_c_983_n 0.00198695f $X=0.965 $Y=0.815 $X2=0
+ $Y2=0

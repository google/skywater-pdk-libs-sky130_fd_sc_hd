* File: sky130_fd_sc_hd__and2_0.spice.SKY130_FD_SC_HD__AND2_0.pxi
* Created: Thu Aug 27 14:06:42 2020
* 
x_PM_SKY130_FD_SC_HD__AND2_0%A N_A_c_45_n N_A_M1001_g N_A_M1005_g N_A_c_47_n A
+ N_A_c_43_n N_A_c_44_n PM_SKY130_FD_SC_HD__AND2_0%A
x_PM_SKY130_FD_SC_HD__AND2_0%B N_B_M1004_g N_B_M1000_g B B N_B_c_77_n
+ PM_SKY130_FD_SC_HD__AND2_0%B
x_PM_SKY130_FD_SC_HD__AND2_0%A_40_47# N_A_40_47#_M1001_s N_A_40_47#_M1005_d
+ N_A_40_47#_M1003_g N_A_40_47#_M1002_g N_A_40_47#_c_111_n N_A_40_47#_c_112_n
+ N_A_40_47#_c_113_n N_A_40_47#_c_114_n N_A_40_47#_c_115_n N_A_40_47#_c_116_n
+ N_A_40_47#_c_117_n N_A_40_47#_c_118_n N_A_40_47#_c_128_n N_A_40_47#_c_119_n
+ PM_SKY130_FD_SC_HD__AND2_0%A_40_47#
x_PM_SKY130_FD_SC_HD__AND2_0%VPWR N_VPWR_M1005_s N_VPWR_M1000_d N_VPWR_c_184_n
+ N_VPWR_c_185_n N_VPWR_c_186_n N_VPWR_c_187_n VPWR N_VPWR_c_188_n
+ N_VPWR_c_183_n N_VPWR_c_190_n PM_SKY130_FD_SC_HD__AND2_0%VPWR
x_PM_SKY130_FD_SC_HD__AND2_0%X N_X_M1003_d N_X_M1002_d N_X_c_217_n X N_X_c_219_n
+ N_X_c_218_n PM_SKY130_FD_SC_HD__AND2_0%X
x_PM_SKY130_FD_SC_HD__AND2_0%VGND N_VGND_M1004_d VGND N_VGND_c_237_n
+ N_VGND_c_238_n N_VGND_c_239_n N_VGND_c_240_n PM_SKY130_FD_SC_HD__AND2_0%VGND
cc_1 VNB N_A_M1001_g 0.0476667f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.445
cc_2 VNB N_A_c_43_n 0.0161364f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.375
cc_3 VNB N_A_c_44_n 0.0112439f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.375
cc_4 VNB N_B_M1004_g 0.0307298f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.21
cc_5 VNB N_B_c_77_n 0.0284945f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.375
cc_6 VNB N_A_40_47#_c_111_n 0.0212309f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.375
cc_7 VNB N_A_40_47#_c_112_n 0.0212168f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.375
cc_8 VNB N_A_40_47#_c_113_n 0.00296141f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.375
cc_9 VNB N_A_40_47#_c_114_n 0.0164073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_40_47#_c_115_n 0.0174546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_40_47#_c_116_n 0.00353309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_40_47#_c_117_n 0.0257029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_40_47#_c_118_n 0.0170757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_40_47#_c_119_n 0.00292267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_183_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_217_n 0.0207333f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.88
cc_17 VNB N_X_c_218_n 0.0413069f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.21
cc_18 VNB N_VGND_c_237_n 0.0268085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_238_n 0.0241965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_239_n 0.14877f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.375
cc_21 VNB N_VGND_c_240_n 0.0106641f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.375
cc_22 VPB N_A_c_45_n 0.0198675f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.663
cc_23 VPB N_A_M1005_g 0.0256089f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=2.275
cc_24 VPB N_A_c_47_n 0.0276554f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.88
cc_25 VPB N_A_c_43_n 0.0103583f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.375
cc_26 VPB N_A_c_44_n 0.0284996f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.375
cc_27 VPB N_B_M1000_g 0.0346612f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.88
cc_28 VPB N_B_c_77_n 0.0453285f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.375
cc_29 VPB N_A_40_47#_M1002_g 0.0405232f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.785
cc_30 VPB N_A_40_47#_c_113_n 0.0147318f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.375
cc_31 VPB N_A_40_47#_c_116_n 0.00533071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_40_47#_c_119_n 0.0055554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_184_n 0.0122121f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.88
cc_34 VPB N_VPWR_c_185_n 0.0171887f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=2.275
cc_35 VPB N_VPWR_c_186_n 0.0189803f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.88
cc_36 VPB N_VPWR_c_187_n 0.0192412f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.375
cc_37 VPB N_VPWR_c_188_n 0.0196753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_183_n 0.0443452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_190_n 0.0097805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_X_c_219_n 0.0330851f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.375
cc_41 VPB N_X_c_218_n 0.0285967f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.21
cc_42 N_A_M1001_g N_B_M1004_g 0.0498104f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_43 N_A_c_47_n N_B_M1000_g 0.0215005f $X=0.397 $Y=1.88 $X2=0 $Y2=0
cc_44 N_A_M1001_g B 4.18345e-19 $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_45 N_A_c_45_n N_B_c_77_n 0.0498104f $X=0.397 $Y=1.663 $X2=0 $Y2=0
cc_46 N_A_M1001_g N_A_40_47#_c_114_n 0.00820836f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_47 N_A_M1001_g N_A_40_47#_c_118_n 0.0203126f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_48 N_A_c_43_n N_A_40_47#_c_118_n 0.00295742f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_49 N_A_c_44_n N_A_40_47#_c_118_n 0.0168822f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_50 N_A_M1005_g N_A_40_47#_c_128_n 0.00466007f $X=0.54 $Y=2.275 $X2=0 $Y2=0
cc_51 N_A_c_45_n N_A_40_47#_c_119_n 0.00485784f $X=0.397 $Y=1.663 $X2=0 $Y2=0
cc_52 N_A_M1001_g N_A_40_47#_c_119_n 0.0110686f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_A_40_47#_c_119_n 0.00955613f $X=0.54 $Y=2.275 $X2=0 $Y2=0
cc_54 N_A_c_47_n N_A_40_47#_c_119_n 0.00484444f $X=0.397 $Y=1.88 $X2=0 $Y2=0
cc_55 N_A_c_43_n N_A_40_47#_c_119_n 0.00450492f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_56 N_A_c_44_n N_A_40_47#_c_119_n 0.0553845f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_57 N_A_c_44_n N_VPWR_c_184_n 0.0011743f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_58 N_A_M1005_g N_VPWR_c_185_n 0.00463875f $X=0.54 $Y=2.275 $X2=0 $Y2=0
cc_59 N_A_c_47_n N_VPWR_c_185_n 0.00151118f $X=0.397 $Y=1.88 $X2=0 $Y2=0
cc_60 N_A_c_44_n N_VPWR_c_185_n 0.0183807f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_61 N_A_M1005_g N_VPWR_c_186_n 0.00564131f $X=0.54 $Y=2.275 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_VPWR_c_183_n 0.0111094f $X=0.54 $Y=2.275 $X2=0 $Y2=0
cc_63 N_A_c_47_n N_VPWR_c_183_n 8.69229e-19 $X=0.397 $Y=1.88 $X2=0 $Y2=0
cc_64 N_A_c_44_n N_VPWR_c_183_n 0.0033011f $X=0.345 $Y=1.375 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_VGND_c_237_n 0.00422379f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_M1001_g N_VGND_c_239_n 0.00682282f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_VGND_c_240_n 0.00203008f $X=0.54 $Y=0.445 $X2=0 $Y2=0
cc_68 N_B_M1000_g N_A_40_47#_M1002_g 0.00701651f $X=0.98 $Y=2.275 $X2=0 $Y2=0
cc_69 B N_A_40_47#_M1002_g 0.00102708f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_70 N_B_c_77_n N_A_40_47#_M1002_g 0.00847043f $X=1.105 $Y=1.18 $X2=0 $Y2=0
cc_71 N_B_M1004_g N_A_40_47#_c_111_n 0.0193076f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_72 N_B_M1004_g N_A_40_47#_c_114_n 0.00152097f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_73 N_B_M1004_g N_A_40_47#_c_115_n 0.0176202f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_74 B N_A_40_47#_c_115_n 0.0260352f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_75 N_B_c_77_n N_A_40_47#_c_115_n 0.00805337f $X=1.105 $Y=1.18 $X2=0 $Y2=0
cc_76 N_B_M1004_g N_A_40_47#_c_116_n 0.00234703f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_77 B N_A_40_47#_c_116_n 0.0269139f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_78 N_B_c_77_n N_A_40_47#_c_116_n 0.00289746f $X=1.105 $Y=1.18 $X2=0 $Y2=0
cc_79 N_B_M1004_g N_A_40_47#_c_117_n 0.00240602f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_80 B N_A_40_47#_c_117_n 4.1872e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_81 N_B_c_77_n N_A_40_47#_c_117_n 0.0249349f $X=1.105 $Y=1.18 $X2=0 $Y2=0
cc_82 N_B_M1004_g N_A_40_47#_c_118_n 0.00114724f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_83 N_B_c_77_n N_A_40_47#_c_128_n 0.00107645f $X=1.105 $Y=1.18 $X2=0 $Y2=0
cc_84 N_B_M1004_g N_A_40_47#_c_119_n 0.00898667f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_85 N_B_M1000_g N_A_40_47#_c_119_n 0.0050147f $X=0.98 $Y=2.275 $X2=0 $Y2=0
cc_86 B N_A_40_47#_c_119_n 0.0402034f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B_M1000_g N_VPWR_c_186_n 0.00585385f $X=0.98 $Y=2.275 $X2=0 $Y2=0
cc_88 N_B_M1000_g N_VPWR_c_187_n 0.00745696f $X=0.98 $Y=2.275 $X2=0 $Y2=0
cc_89 B N_VPWR_c_187_n 0.0113969f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B_c_77_n N_VPWR_c_187_n 0.004657f $X=1.105 $Y=1.18 $X2=0 $Y2=0
cc_91 N_B_M1000_g N_VPWR_c_183_n 0.011293f $X=0.98 $Y=2.275 $X2=0 $Y2=0
cc_92 N_B_M1004_g N_VGND_c_237_n 0.00361431f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_93 N_B_M1004_g N_VGND_c_239_n 0.00411857f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_94 N_B_M1004_g N_VGND_c_240_n 0.0148196f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_40_47#_c_128_n N_VPWR_c_186_n 0.0156121f $X=0.765 $Y=2.3 $X2=0 $Y2=0
cc_96 N_A_40_47#_M1002_g N_VPWR_c_187_n 0.00354558f $X=1.75 $Y=2.165 $X2=0 $Y2=0
cc_97 N_A_40_47#_c_113_n N_VPWR_c_187_n 9.72181e-19 $X=1.652 $Y=1.435 $X2=0
+ $Y2=0
cc_98 N_A_40_47#_c_116_n N_VPWR_c_187_n 0.00801912f $X=1.615 $Y=0.93 $X2=0 $Y2=0
cc_99 N_A_40_47#_c_119_n N_VPWR_c_187_n 0.0131293f $X=0.732 $Y=2.135 $X2=0 $Y2=0
cc_100 N_A_40_47#_M1002_g N_VPWR_c_188_n 0.00533769f $X=1.75 $Y=2.165 $X2=0
+ $Y2=0
cc_101 N_A_40_47#_M1005_d N_VPWR_c_183_n 0.00370124f $X=0.615 $Y=2.065 $X2=0
+ $Y2=0
cc_102 N_A_40_47#_M1002_g N_VPWR_c_183_n 0.0110193f $X=1.75 $Y=2.165 $X2=0 $Y2=0
cc_103 N_A_40_47#_c_128_n N_VPWR_c_183_n 0.00992767f $X=0.765 $Y=2.3 $X2=0 $Y2=0
cc_104 N_A_40_47#_c_111_n N_X_c_217_n 0.0033293f $X=1.63 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A_40_47#_c_112_n N_X_c_217_n 0.00286013f $X=1.63 $Y=0.915 $X2=0 $Y2=0
cc_106 N_A_40_47#_c_115_n N_X_c_217_n 0.0155883f $X=1.45 $Y=0.802 $X2=0 $Y2=0
cc_107 N_A_40_47#_M1002_g N_X_c_219_n 0.00936712f $X=1.75 $Y=2.165 $X2=0 $Y2=0
cc_108 N_A_40_47#_c_111_n N_X_c_218_n 0.00461079f $X=1.63 $Y=0.765 $X2=0 $Y2=0
cc_109 N_A_40_47#_c_112_n N_X_c_218_n 0.0313294f $X=1.63 $Y=0.915 $X2=0 $Y2=0
cc_110 N_A_40_47#_c_115_n N_X_c_218_n 0.0180656f $X=1.45 $Y=0.802 $X2=0 $Y2=0
cc_111 N_A_40_47#_c_116_n N_X_c_218_n 0.0407195f $X=1.615 $Y=0.93 $X2=0 $Y2=0
cc_112 N_A_40_47#_c_114_n N_VGND_c_237_n 0.0160954f $X=0.325 $Y=0.445 $X2=0
+ $Y2=0
cc_113 N_A_40_47#_c_118_n N_VGND_c_237_n 0.00715612f $X=0.77 $Y=0.822 $X2=0
+ $Y2=0
cc_114 N_A_40_47#_c_111_n N_VGND_c_238_n 0.00420974f $X=1.63 $Y=0.765 $X2=0
+ $Y2=0
cc_115 N_A_40_47#_c_115_n N_VGND_c_238_n 0.00268125f $X=1.45 $Y=0.802 $X2=0
+ $Y2=0
cc_116 N_A_40_47#_M1001_s N_VGND_c_239_n 0.00215353f $X=0.2 $Y=0.235 $X2=0 $Y2=0
cc_117 N_A_40_47#_c_111_n N_VGND_c_239_n 0.00731308f $X=1.63 $Y=0.765 $X2=0
+ $Y2=0
cc_118 N_A_40_47#_c_114_n N_VGND_c_239_n 0.011251f $X=0.325 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_40_47#_c_115_n N_VGND_c_239_n 0.00643196f $X=1.45 $Y=0.802 $X2=0
+ $Y2=0
cc_120 N_A_40_47#_c_118_n N_VGND_c_239_n 0.0114393f $X=0.77 $Y=0.822 $X2=0 $Y2=0
cc_121 N_A_40_47#_c_111_n N_VGND_c_240_n 0.00515447f $X=1.63 $Y=0.765 $X2=0
+ $Y2=0
cc_122 N_A_40_47#_c_114_n N_VGND_c_240_n 0.0083323f $X=0.325 $Y=0.445 $X2=0
+ $Y2=0
cc_123 N_A_40_47#_c_115_n N_VGND_c_240_n 0.0319459f $X=1.45 $Y=0.802 $X2=0 $Y2=0
cc_124 N_VPWR_c_183_n N_X_M1002_d 0.00213418f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_125 N_VPWR_c_187_n N_X_c_219_n 0.0249719f $X=1.525 $Y=2 $X2=0 $Y2=0
cc_126 N_VPWR_c_188_n N_X_c_219_n 0.0277856f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_127 N_VPWR_c_183_n N_X_c_219_n 0.0160505f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_128 N_X_c_217_n N_VGND_c_238_n 0.0427963f $X=1.95 $Y=0.39 $X2=0 $Y2=0
cc_129 N_X_M1003_d N_VGND_c_239_n 0.00213443f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_130 N_X_c_217_n N_VGND_c_239_n 0.0246904f $X=1.95 $Y=0.39 $X2=0 $Y2=0
cc_131 A_123_47# N_VGND_c_239_n 0.00263669f $X=0.615 $Y=0.235 $X2=2.07 $Y2=0

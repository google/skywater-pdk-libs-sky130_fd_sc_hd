* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_16.pex.spice
* Created: Thu Aug 27 14:23:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%A 3 5 7 10 12 14 17 19 21 24
+ 26 28 29 30 40
r68 39 40 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=1.335 $Y=1.155
+ $X2=1.765 $Y2=1.155
r69 38 39 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=1.155
+ $X2=1.335 $Y2=1.155
r70 37 38 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.155
+ $X2=0.905 $Y2=1.155
r71 34 37 21.5061 $w=5.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.155
+ $X2=0.475 $Y2=1.155
r72 30 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r73 29 30 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r74 26 40 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.765 $Y=1.41
+ $X2=1.765 $Y2=1.155
r75 26 28 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.765 $Y=1.41
+ $X2=1.765 $Y2=1.985
r76 22 40 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.765 $Y=0.9
+ $X2=1.765 $Y2=1.155
r77 22 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.765 $Y=0.9
+ $X2=1.765 $Y2=0.445
r78 19 39 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.335 $Y=1.41
+ $X2=1.335 $Y2=1.155
r79 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.335 $Y=1.41
+ $X2=1.335 $Y2=1.985
r80 15 39 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.335 $Y=0.9
+ $X2=1.335 $Y2=1.155
r81 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=0.9
+ $X2=1.335 $Y2=0.445
r82 12 38 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.155
r83 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
r84 8 38 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=1.155
r85 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=0.445
r86 5 37 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.155
r87 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.985
r88 1 37 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=1.155
r89 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%A_110_47# 1 2 3 4 15 19 23 27
+ 31 35 39 43 47 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123
+ 127 131 133 135 139 143 147 151 155 159 168 171 172
r335 168 169 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=7.505
+ $Y=1.16 $X2=7.505 $Y2=1.16
r336 165 168 235.098 $w=2.48e-07 $l=5.1e-06 $layer=LI1_cond $X=2.405 $Y=1.2
+ $X2=7.505 $Y2=1.2
r337 165 166 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=2.405
+ $Y=1.16 $X2=2.405 $Y2=1.16
r338 163 172 2.66945 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=1.2
+ $X2=1.555 $Y2=1.2
r339 163 165 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=1.68 $Y=1.2
+ $X2=2.405 $Y2=1.2
r340 159 161 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=1.55 $Y=1.615
+ $X2=1.55 $Y2=2.295
r341 157 172 3.44865 $w=1.9e-07 $l=1.27475e-07 $layer=LI1_cond $X=1.55 $Y=1.325
+ $X2=1.555 $Y2=1.2
r342 157 159 16.9282 $w=1.88e-07 $l=2.9e-07 $layer=LI1_cond $X=1.55 $Y=1.325
+ $X2=1.55 $Y2=1.615
r343 153 172 3.44865 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.075
+ $X2=1.555 $Y2=1.2
r344 153 155 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=1.555 $Y=1.075
+ $X2=1.555 $Y2=0.445
r345 152 171 0.681005 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=0.82 $Y=1.2
+ $X2=0.707 $Y2=1.2
r346 151 172 2.66945 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.43 $Y=1.2
+ $X2=1.555 $Y2=1.2
r347 151 152 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=1.43 $Y=1.2
+ $X2=0.82 $Y2=1.2
r348 147 149 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.615
+ $X2=0.69 $Y2=2.295
r349 145 171 6.01496 $w=2.07e-07 $l=1.33229e-07 $layer=LI1_cond $X=0.69 $Y=1.325
+ $X2=0.707 $Y2=1.2
r350 145 147 16.9282 $w=1.88e-07 $l=2.9e-07 $layer=LI1_cond $X=0.69 $Y=1.325
+ $X2=0.69 $Y2=1.615
r351 141 171 6.01496 $w=2.07e-07 $l=1.25e-07 $layer=LI1_cond $X=0.707 $Y=1.075
+ $X2=0.707 $Y2=1.2
r352 141 143 32.2684 $w=2.23e-07 $l=6.3e-07 $layer=LI1_cond $X=0.707 $Y=1.075
+ $X2=0.707 $Y2=0.445
r353 137 139 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.64 $Y=1.325
+ $X2=8.64 $Y2=1.985
r354 133 137 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.64 $Y=1.137
+ $X2=8.64 $Y2=1.325
r355 133 135 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.64 $Y=0.95
+ $X2=8.64 $Y2=0.445
r356 129 131 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.21 $Y=1.325
+ $X2=8.21 $Y2=1.985
r357 125 133 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=8.21 $Y=1.137
+ $X2=8.64 $Y2=1.137
r358 125 129 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.21 $Y=1.137
+ $X2=8.21 $Y2=1.325
r359 125 127 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.21 $Y=0.95
+ $X2=8.21 $Y2=0.445
r360 121 123 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.78 $Y=1.325
+ $X2=7.78 $Y2=1.985
r361 117 125 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=7.78 $Y=1.137
+ $X2=8.21 $Y2=1.137
r362 117 121 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=7.78 $Y=1.137
+ $X2=7.78 $Y2=1.325
r363 117 169 40.7846 $w=3.75e-07 $l=2.75e-07 $layer=POLY_cond $X=7.78 $Y=1.137
+ $X2=7.505 $Y2=1.137
r364 117 119 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.78 $Y=0.95
+ $X2=7.78 $Y2=0.445
r365 113 115 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.35 $Y=1.325
+ $X2=7.35 $Y2=1.985
r366 109 169 22.9877 $w=3.75e-07 $l=1.55e-07 $layer=POLY_cond $X=7.35 $Y=1.137
+ $X2=7.505 $Y2=1.137
r367 109 113 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=7.35 $Y=1.137
+ $X2=7.35 $Y2=1.325
r368 109 111 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.35 $Y=0.95
+ $X2=7.35 $Y2=0.445
r369 105 107 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.92 $Y=1.325
+ $X2=6.92 $Y2=1.985
r370 101 109 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=6.92 $Y=1.137
+ $X2=7.35 $Y2=1.137
r371 101 105 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.92 $Y=1.137
+ $X2=6.92 $Y2=1.325
r372 101 103 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.92 $Y=0.95
+ $X2=6.92 $Y2=0.445
r373 97 99 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.49 $Y=1.325
+ $X2=6.49 $Y2=1.985
r374 93 101 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=6.49 $Y=1.137
+ $X2=6.92 $Y2=1.137
r375 93 97 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.49 $Y=1.137
+ $X2=6.49 $Y2=1.325
r376 93 95 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.49 $Y=0.95
+ $X2=6.49 $Y2=0.445
r377 89 91 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.06 $Y=1.325
+ $X2=6.06 $Y2=1.985
r378 85 93 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=6.06 $Y=1.137
+ $X2=6.49 $Y2=1.137
r379 85 89 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.06 $Y=1.137
+ $X2=6.06 $Y2=1.325
r380 85 87 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.06 $Y=0.95
+ $X2=6.06 $Y2=0.445
r381 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.985
r382 77 85 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=5.63 $Y=1.137
+ $X2=6.06 $Y2=1.137
r383 77 81 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=5.63 $Y=1.137
+ $X2=5.63 $Y2=1.325
r384 77 79 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.63 $Y=0.95
+ $X2=5.63 $Y2=0.445
r385 73 75 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.205 $Y=1.325
+ $X2=5.205 $Y2=1.985
r386 69 77 63.0308 $w=3.75e-07 $l=4.25e-07 $layer=POLY_cond $X=5.205 $Y=1.137
+ $X2=5.63 $Y2=1.137
r387 69 73 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=5.205 $Y=1.137
+ $X2=5.205 $Y2=1.325
r388 69 71 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.205 $Y=0.95
+ $X2=5.205 $Y2=0.445
r389 65 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.775 $Y=1.325
+ $X2=4.775 $Y2=1.985
r390 61 69 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=4.775 $Y=1.137
+ $X2=5.205 $Y2=1.137
r391 61 65 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=4.775 $Y=1.137
+ $X2=4.775 $Y2=1.325
r392 61 63 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.775 $Y=0.95
+ $X2=4.775 $Y2=0.445
r393 57 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.345 $Y=1.325
+ $X2=4.345 $Y2=1.985
r394 53 61 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=4.345 $Y=1.137
+ $X2=4.775 $Y2=1.137
r395 53 57 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=4.345 $Y=1.137
+ $X2=4.345 $Y2=1.325
r396 53 55 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.345 $Y=0.95
+ $X2=4.345 $Y2=0.445
r397 49 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.915 $Y=1.325
+ $X2=3.915 $Y2=1.985
r398 45 53 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=4.345 $Y2=1.137
r399 45 49 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=3.915 $Y2=1.325
r400 45 47 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.915 $Y=0.95
+ $X2=3.915 $Y2=0.445
r401 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=1.985
r402 37 45 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.915 $Y2=1.137
r403 37 41 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.485 $Y2=1.325
r404 37 39 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.485 $Y=0.95
+ $X2=3.485 $Y2=0.445
r405 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.325
+ $X2=3.055 $Y2=1.985
r406 29 37 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.485 $Y2=1.137
r407 29 33 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.055 $Y2=1.325
r408 29 31 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.055 $Y=0.95
+ $X2=3.055 $Y2=0.445
r409 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.625 $Y=1.325
+ $X2=2.625 $Y2=1.985
r410 21 29 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=3.055 $Y2=1.137
r411 21 25 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=2.625 $Y2=1.325
r412 21 166 32.6277 $w=3.75e-07 $l=2.2e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=2.405 $Y2=1.137
r413 21 23 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.625 $Y=0.95
+ $X2=2.625 $Y2=0.445
r414 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.195 $Y=1.325
+ $X2=2.195 $Y2=1.985
r415 13 166 31.1446 $w=3.75e-07 $l=2.1e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.405 $Y2=1.137
r416 13 17 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.195 $Y2=1.325
r417 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.195 $Y=0.95
+ $X2=2.195 $Y2=0.445
r418 4 161 400 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=2.295
r419 4 159 400 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=1.615
r420 3 149 400 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2.295
r421 3 147 400 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.615
r422 2 155 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.445
r423 1 143 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%KAPWR 1 2 3 4 5 6 7 8 9 10 11
+ 35 52 57 58 62 63 66 67 68 71 72 73 76 77 78 81 82 83 86 87 88 91 92 93 96 97
+ 98 101 102 105 113 119 158
c198 68 0 1.77237e-19 $X=2.97 $Y=2.21
c199 52 0 1.27506e-19 $X=8.72 $Y=2.24
c200 11 0 4.2343e-20 $X=8.715 $Y=1.485
r201 105 108 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.21
r202 102 158 0.00249004 $w=2.51e-07 $l=5e-09 $layer=MET1_cond $X=0.26 $Y=2.21
+ $X2=0.265 $Y2=2.21
r203 102 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.21
+ $X2=0.26 $Y2=2.21
r204 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.865 $Y=2.21
+ $X2=8.865 $Y2=2.21
r205 95 98 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.985 $Y=2.21
+ $X2=8.13 $Y2=2.21
r206 95 97 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.985 $Y=2.21
+ $X2=7.84 $Y2=2.21
r207 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.985 $Y=2.21
+ $X2=7.985 $Y2=2.21
r208 93 97 0.429825 $w=2e-07 $l=5.6e-07 $layer=MET1_cond $X=7.28 $Y=2.24
+ $X2=7.84 $Y2=2.24
r209 90 93 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.135 $Y=2.21
+ $X2=7.28 $Y2=2.21
r210 90 92 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.135 $Y=2.21
+ $X2=6.99 $Y2=2.21
r211 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.135 $Y=2.21
+ $X2=7.135 $Y2=2.21
r212 88 92 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=6.425 $Y=2.24
+ $X2=6.99 $Y2=2.24
r213 85 88 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=6.28 $Y=2.21
+ $X2=6.425 $Y2=2.21
r214 85 87 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=6.28 $Y=2.21
+ $X2=6.135 $Y2=2.21
r215 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.28 $Y=2.21
+ $X2=6.28 $Y2=2.21
r216 83 87 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=5.565 $Y=2.24
+ $X2=6.135 $Y2=2.24
r217 80 83 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.42 $Y=2.21
+ $X2=5.565 $Y2=2.21
r218 80 82 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.42 $Y=2.21
+ $X2=5.275 $Y2=2.21
r219 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.42 $Y=2.21
+ $X2=5.42 $Y2=2.21
r220 78 82 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=4.71 $Y=2.24
+ $X2=5.275 $Y2=2.24
r221 75 78 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.565 $Y=2.21
+ $X2=4.71 $Y2=2.21
r222 75 77 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.565 $Y=2.21
+ $X2=4.42 $Y2=2.21
r223 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.565 $Y=2.21
+ $X2=4.565 $Y2=2.21
r224 73 77 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=3.85 $Y=2.24
+ $X2=4.42 $Y2=2.24
r225 70 73 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.705 $Y=2.21
+ $X2=3.85 $Y2=2.21
r226 70 72 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.705 $Y=2.21
+ $X2=3.56 $Y2=2.21
r227 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.705 $Y=2.21
+ $X2=3.705 $Y2=2.21
r228 68 72 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=2.97 $Y=2.24
+ $X2=3.56 $Y2=2.24
r229 65 68 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.825 $Y=2.21
+ $X2=2.97 $Y2=2.21
r230 65 67 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.825 $Y=2.21
+ $X2=2.68 $Y2=2.21
r231 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.825 $Y=2.21
+ $X2=2.825 $Y2=2.21
r232 63 67 0.429825 $w=2e-07 $l=5.6e-07 $layer=MET1_cond $X=2.12 $Y=2.24
+ $X2=2.68 $Y2=2.24
r233 61 119 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.98 $Y=2.21
+ $X2=1.98 $Y2=1.66
r234 60 63 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=2.12 $Y2=2.21
r235 60 62 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=1.83 $Y2=2.21
r236 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.975 $Y=2.21
+ $X2=1.975 $Y2=2.21
r237 58 62 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=1.265 $Y=2.24
+ $X2=1.83 $Y2=2.24
r238 56 113 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.12 $Y=2.21
+ $X2=1.12 $Y2=1.66
r239 55 58 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.12 $Y=2.21
+ $X2=1.265 $Y2=2.21
r240 55 57 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.12 $Y=2.21
+ $X2=0.975 $Y2=2.21
r241 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.21
+ $X2=1.12 $Y2=2.21
r242 52 100 0.0790316 $w=2.42e-07 $l=1.59295e-07 $layer=MET1_cond $X=8.72
+ $Y=2.24 $X2=8.865 $Y2=2.21
r243 52 98 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=8.72 $Y=2.24
+ $X2=8.13 $Y2=2.24
r244 35 158 0.0752387 $w=2.51e-07 $l=1.54272e-07 $layer=MET1_cond $X=0.405
+ $Y=2.24 $X2=0.265 $Y2=2.21
r245 35 57 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=0.405 $Y=2.24
+ $X2=0.975 $Y2=2.24
r246 11 101 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.485 $X2=8.855 $Y2=2.22
r247 10 96 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.485 $X2=7.995 $Y2=2.22
r248 9 91 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=6.995
+ $Y=1.485 $X2=7.135 $Y2=2.22
r249 8 86 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=6.135
+ $Y=1.485 $X2=6.275 $Y2=2.22
r250 7 81 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.485 $X2=5.42 $Y2=2.22
r251 6 76 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.485 $X2=4.56 $Y2=2.22
r252 5 71 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.7 $Y2=2.22
r253 4 66 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.84 $Y2=2.22
r254 3 61 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.485 $X2=1.98 $Y2=2.34
r255 3 119 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.485 $X2=1.98 $Y2=1.66
r256 2 56 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=2.34
r257 2 113 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=1.66
r258 1 108 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r259 1 105 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%X 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 51 55 56 57 61 65 67 71 75 77 81 85 87 91 95 97 101 105 107 111
+ 115 119 124 125 127 128 130 131 133 134 136 137 139 140 141 142 143 168 173
c300 141 0 1.18325e-19 $X=8.51 $Y=0.85
c301 16 0 1.27506e-19 $X=8.285 $Y=1.485
r302 171 173 0.362137 $w=1.516e-06 $l=4.5e-08 $layer=LI1_cond $X=8.225 $Y=1.615
+ $X2=8.225 $Y2=1.66
r303 158 168 0.966712 $w=1.516e-06 $l=2.33846e-07 $layer=LI1_cond $X=8.442
+ $Y=1.495 $X2=8.225 $Y2=1.53
r304 143 171 0.48285 $w=1.516e-06 $l=6e-08 $layer=LI1_cond $X=8.225 $Y=1.555
+ $X2=8.225 $Y2=1.615
r305 143 168 0.201187 $w=1.516e-06 $l=2.5e-08 $layer=LI1_cond $X=8.225 $Y=1.555
+ $X2=8.225 $Y2=1.53
r306 143 158 0.261803 $w=1.163e-06 $l=2.5e-08 $layer=LI1_cond $X=8.442 $Y=1.47
+ $X2=8.442 $Y2=1.495
r307 142 143 2.93219 $w=1.163e-06 $l=2.8e-07 $layer=LI1_cond $X=8.442 $Y=1.19
+ $X2=8.442 $Y2=1.47
r308 141 157 1.4003 $w=7.12e-07 $l=8.5e-08 $layer=LI1_cond $X=8.442 $Y=0.82
+ $X2=8.442 $Y2=0.905
r309 141 142 2.82747 $w=1.163e-06 $l=2.7e-07 $layer=LI1_cond $X=8.442 $Y=0.92
+ $X2=8.442 $Y2=1.19
r310 141 157 0.157082 $w=1.163e-06 $l=1.5e-08 $layer=LI1_cond $X=8.442 $Y=0.92
+ $X2=8.442 $Y2=0.905
r311 117 141 1.4003 $w=7.12e-07 $l=9.31128e-08 $layer=LI1_cond $X=8.425 $Y=0.735
+ $X2=8.442 $Y2=0.82
r312 117 119 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=8.425 $Y=0.735
+ $X2=8.425 $Y2=0.445
r313 116 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.685 $Y=0.82
+ $X2=7.555 $Y2=0.82
r314 115 141 6.76561 $w=1.7e-07 $l=5.82e-07 $layer=LI1_cond $X=7.86 $Y=0.82
+ $X2=8.442 $Y2=0.82
r315 115 116 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.86 $Y=0.82
+ $X2=7.685 $Y2=0.82
r316 109 140 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.735
+ $X2=7.555 $Y2=0.82
r317 109 111 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=7.555 $Y=0.735
+ $X2=7.555 $Y2=0.445
r318 108 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=6.825 $Y=1.615
+ $X2=6.695 $Y2=1.615
r319 107 171 12.2163 $w=2.4e-07 $l=8e-07 $layer=LI1_cond $X=7.425 $Y=1.615
+ $X2=8.225 $Y2=1.615
r320 107 108 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=7.425 $Y=1.615
+ $X2=6.825 $Y2=1.615
r321 106 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.825 $Y=0.82
+ $X2=6.695 $Y2=0.82
r322 105 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.425 $Y=0.82
+ $X2=7.555 $Y2=0.82
r323 105 106 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.425 $Y=0.82
+ $X2=6.825 $Y2=0.82
r324 99 137 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=0.735
+ $X2=6.695 $Y2=0.82
r325 99 101 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=6.695 $Y=0.735
+ $X2=6.695 $Y2=0.445
r326 98 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.965 $Y=1.615
+ $X2=5.835 $Y2=1.615
r327 97 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=6.565 $Y=1.615
+ $X2=6.695 $Y2=1.615
r328 97 98 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=6.565 $Y=1.615
+ $X2=5.965 $Y2=1.615
r329 96 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.965 $Y=0.82
+ $X2=5.835 $Y2=0.82
r330 95 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.565 $Y=0.82
+ $X2=6.695 $Y2=0.82
r331 95 96 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.565 $Y=0.82
+ $X2=5.965 $Y2=0.82
r332 89 134 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0.735
+ $X2=5.835 $Y2=0.82
r333 89 91 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=5.835 $Y=0.735
+ $X2=5.835 $Y2=0.445
r334 88 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.12 $Y=1.615
+ $X2=4.99 $Y2=1.615
r335 87 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.705 $Y=1.615
+ $X2=5.835 $Y2=1.615
r336 87 88 28.0908 $w=2.38e-07 $l=5.85e-07 $layer=LI1_cond $X=5.705 $Y=1.615
+ $X2=5.12 $Y2=1.615
r337 86 131 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.12 $Y=0.82
+ $X2=4.982 $Y2=0.82
r338 85 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.705 $Y=0.82
+ $X2=5.835 $Y2=0.82
r339 85 86 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.705 $Y=0.82
+ $X2=5.12 $Y2=0.82
r340 79 131 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.982 $Y=0.735
+ $X2=4.982 $Y2=0.82
r341 79 81 12.153 $w=2.73e-07 $l=2.9e-07 $layer=LI1_cond $X=4.982 $Y=0.735
+ $X2=4.982 $Y2=0.445
r342 78 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=1.615
+ $X2=4.13 $Y2=1.615
r343 77 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4.86 $Y=1.615
+ $X2=4.99 $Y2=1.615
r344 77 78 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=4.86 $Y=1.615
+ $X2=4.26 $Y2=1.615
r345 76 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=0.82
+ $X2=4.13 $Y2=0.82
r346 75 131 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.845 $Y=0.82
+ $X2=4.982 $Y2=0.82
r347 75 76 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.845 $Y=0.82
+ $X2=4.26 $Y2=0.82
r348 69 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.82
r349 69 71 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.445
r350 68 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=1.615
+ $X2=3.27 $Y2=1.615
r351 67 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=1.615 $X2=4.13
+ $Y2=1.615
r352 67 68 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=4 $Y=1.615 $X2=3.4
+ $Y2=1.615
r353 66 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=0.82
+ $X2=3.27 $Y2=0.82
r354 65 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=0.82 $X2=4.13
+ $Y2=0.82
r355 65 66 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4 $Y=0.82 $X2=3.4
+ $Y2=0.82
r356 59 125 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.82
r357 59 61 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.445
r358 58 124 3.31033 $w=2.4e-07 $l=1.13e-07 $layer=LI1_cond $X=2.54 $Y=1.615
+ $X2=2.427 $Y2=1.615
r359 57 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=3.27 $Y2=1.615
r360 57 58 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=2.54 $Y2=1.615
r361 55 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=0.82
+ $X2=3.27 $Y2=0.82
r362 55 56 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.82 $X2=2.54
+ $Y2=0.82
r363 49 56 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.54 $Y2=0.82
r364 49 51 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.445
r365 16 173 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=8.285
+ $Y=1.485 $X2=8.425 $Y2=1.66
r366 15 173 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=7.425
+ $Y=1.485 $X2=7.565 $Y2=1.66
r367 14 139 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=6.565
+ $Y=1.485 $X2=6.705 $Y2=1.66
r368 13 136 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=5.705
+ $Y=1.485 $X2=5.845 $Y2=1.66
r369 12 133 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=4.85
+ $Y=1.485 $X2=4.99 $Y2=1.66
r370 11 130 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.485 $X2=4.13 $Y2=1.66
r371 10 127 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.485 $X2=3.27 $Y2=1.66
r372 9 124 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.485 $X2=2.41 $Y2=1.66
r373 8 119 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.285
+ $Y=0.235 $X2=8.425 $Y2=0.445
r374 7 111 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.565 $Y2=0.445
r375 6 101 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.705 $Y2=0.445
r376 5 91 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.845 $Y2=0.445
r377 4 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.85
+ $Y=0.235 $X2=4.99 $Y2=0.445
r378 3 71 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.445
r379 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.445
r380 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%VGND 1 2 3 4 5 6 7 8 9 10 11
+ 34 36 40 44 48 52 56 58 62 64 68 72 76 78 80 83 84 86 87 89 90 91 92 94 95 96
+ 98 116 125 133 136 139 142 146
c160 94 0 7.59816e-20 $X=7.865 $Y=0
r161 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r162 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r163 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r164 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r165 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r166 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r167 128 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r168 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r169 125 145 4.35621 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=8.725 $Y=0
+ $X2=8.962 $Y2=0
r170 125 127 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.725 $Y=0
+ $X2=8.51 $Y2=0
r171 124 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r172 124 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r173 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r174 121 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=0
+ $X2=7.13 $Y2=0
r175 121 123 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.255 $Y=0
+ $X2=7.59 $Y2=0
r176 120 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r177 120 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r178 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r179 117 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.395 $Y=0
+ $X2=6.27 $Y2=0
r180 117 119 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.395 $Y=0
+ $X2=6.67 $Y2=0
r181 116 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.13 $Y2=0
r182 116 119 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=6.67 $Y2=0
r183 115 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r184 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r185 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r186 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r187 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r188 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r189 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r190 106 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r191 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r192 103 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r193 103 105 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=0
+ $X2=1.61 $Y2=0
r194 102 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r195 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r196 99 130 4.57719 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0
+ $X2=0.195 $Y2=0
r197 99 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r198 98 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r199 98 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.69
+ $Y2=0
r200 96 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r201 96 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r202 94 123 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.865 $Y=0
+ $X2=7.59 $Y2=0
r203 94 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.865 $Y=0 $X2=7.995
+ $Y2=0
r204 93 127 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.125 $Y=0
+ $X2=8.51 $Y2=0
r205 93 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.125 $Y=0 $X2=7.995
+ $Y2=0
r206 91 114 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.37
+ $Y2=0
r207 91 92 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.552
+ $Y2=0
r208 89 111 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r209 89 90 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.7
+ $Y2=0
r210 88 114 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.37
+ $Y2=0
r211 88 90 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.7
+ $Y2=0
r212 86 108 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r213 86 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.84
+ $Y2=0
r214 85 111 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.45
+ $Y2=0
r215 85 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.84
+ $Y2=0
r216 83 105 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.61
+ $Y2=0
r217 83 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.98
+ $Y2=0
r218 82 108 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.53
+ $Y2=0
r219 82 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.98
+ $Y2=0
r220 78 145 3.16147 $w=3e-07 $l=1.22327e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.962 $Y2=0
r221 78 80 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0.4
r222 74 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.995 $Y=0.085
+ $X2=7.995 $Y2=0
r223 74 76 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=7.995 $Y=0.085
+ $X2=7.995 $Y2=0.4
r224 70 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.13 $Y=0.085
+ $X2=7.13 $Y2=0
r225 70 72 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=7.13 $Y=0.085
+ $X2=7.13 $Y2=0.4
r226 66 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0
r227 66 68 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0.4
r228 65 136 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=5.535 $Y=0
+ $X2=5.412 $Y2=0
r229 64 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=6.27 $Y2=0
r230 64 65 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=5.535 $Y2=0
r231 60 136 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.412 $Y=0.085
+ $X2=5.412 $Y2=0
r232 60 62 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=5.412 $Y=0.085
+ $X2=5.412 $Y2=0.4
r233 59 92 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4.675 $Y=0
+ $X2=4.552 $Y2=0
r234 58 136 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.412 $Y2=0
r235 58 59 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=4.675
+ $Y2=0
r236 54 92 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.552 $Y=0.085
+ $X2=4.552 $Y2=0
r237 54 56 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=4.552 $Y=0.085
+ $X2=4.552 $Y2=0.4
r238 50 90 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r239 50 52 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.4
r240 46 87 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r241 46 48 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.4
r242 42 84 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r243 42 44 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.445
r244 38 133 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r245 38 40 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.445
r246 34 130 2.98104 $w=3.05e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.195 $Y2=0
r247 34 36 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.38
r248 11 80 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.715
+ $Y=0.235 $X2=8.855 $Y2=0.4
r249 10 76 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.855
+ $Y=0.235 $X2=7.995 $Y2=0.4
r250 9 72 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.995
+ $Y=0.235 $X2=7.135 $Y2=0.4
r251 8 68 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.135
+ $Y=0.235 $X2=6.275 $Y2=0.4
r252 7 62 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.28
+ $Y=0.235 $X2=5.42 $Y2=0.4
r253 6 56 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.235 $X2=4.56 $Y2=0.4
r254 5 52 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.4
r255 4 48 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.4
r256 3 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.445
r257 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
r258 1 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%VPWR 1 8 9
c122 8 0 1.77237e-19 $X=8.97 $Y=2.72
r123 8 9 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r124 4 8 570.203 $w=1.68e-07 $l=8.74e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=8.97 $Y2=2.72
r125 1 9 2.48689 $w=4.8e-07 $l=8.74e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=8.97 $Y2=2.72
r126 1 4 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__and3b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__and3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715000 0.615000 3.995000 1.705000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.725000 1.235000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.715000 1.340000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.535000 3.535000 1.705000 ;
        RECT 2.285000 0.515000 2.475000 0.615000 ;
        RECT 2.285000 0.615000 3.535000 0.845000 ;
        RECT 3.145000 0.255000 3.335000 0.615000 ;
        RECT 3.270000 0.845000 3.535000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.150000  0.255000 0.635000 0.355000 ;
      RECT 0.150000  0.355000 1.600000 0.545000 ;
      RECT 0.150000  0.545000 0.635000 0.805000 ;
      RECT 0.150000  0.805000 0.370000 1.495000 ;
      RECT 0.150000  1.495000 0.510000 2.165000 ;
      RECT 0.540000  0.995000 0.850000 1.325000 ;
      RECT 0.680000  1.325000 0.850000 1.875000 ;
      RECT 0.680000  1.875000 4.445000 2.105000 ;
      RECT 0.730000  2.275000 1.180000 2.635000 ;
      RECT 1.280000  1.525000 2.055000 1.695000 ;
      RECT 1.420000  0.545000 1.600000 0.615000 ;
      RECT 1.420000  0.615000 2.115000 0.805000 ;
      RECT 1.745000  2.275000 2.075000 2.635000 ;
      RECT 1.780000  0.085000 2.110000 0.445000 ;
      RECT 1.885000  0.805000 2.115000 1.020000 ;
      RECT 1.885000  1.020000 3.100000 1.355000 ;
      RECT 1.885000  1.355000 2.055000 1.525000 ;
      RECT 2.645000  0.085000 2.975000 0.445000 ;
      RECT 2.645000  2.275000 2.980000 2.635000 ;
      RECT 3.505000  0.085000 3.835000 0.445000 ;
      RECT 3.505000  2.275000 3.835000 2.635000 ;
      RECT 4.165000  0.425000 4.445000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_4
END LIBRARY

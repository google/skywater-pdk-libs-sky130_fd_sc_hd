# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.075000 4.455000 1.245000 ;
        RECT 3.560000 1.245000 4.455000 1.295000 ;
        RECT 4.115000 0.765000 4.455000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.075000 3.335000 1.355000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.905000 1.365000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.375000 1.970000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.022000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.670000 0.875000 1.540000 ;
        RECT 0.545000 1.540000 3.155000 1.710000 ;
        RECT 0.545000 1.710000 0.805000 2.465000 ;
        RECT 1.475000 1.710000 1.665000 2.465000 ;
        RECT 2.825000 1.710000 3.155000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.255000 2.165000 0.445000 ;
      RECT 0.115000  2.175000 0.375000 2.635000 ;
      RECT 0.975000  1.915000 1.305000 2.635000 ;
      RECT 1.045000  0.445000 2.165000 0.465000 ;
      RECT 1.045000  0.465000 1.235000 0.890000 ;
      RECT 1.405000  0.635000 3.945000 0.845000 ;
      RECT 1.835000  1.915000 2.165000 2.635000 ;
      RECT 2.395000  0.085000 2.725000 0.445000 ;
      RECT 2.395000  2.100000 2.655000 2.295000 ;
      RECT 2.395000  2.295000 3.515000 2.465000 ;
      RECT 3.255000  0.085000 3.585000 0.445000 ;
      RECT 3.325000  1.525000 4.445000 1.695000 ;
      RECT 3.325000  1.695000 3.515000 2.295000 ;
      RECT 3.685000  1.865000 4.015000 2.635000 ;
      RECT 3.755000  0.515000 3.945000 0.635000 ;
      RECT 4.115000  0.085000 4.445000 0.445000 ;
      RECT 4.185000  1.695000 4.445000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o211ai_2
END LIBRARY

* File: sky130_fd_sc_hd__dfrtp_1.spice
* Created: Thu Aug 27 14:14:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dfrtp_1.pex.spice"
.subckt sky130_fd_sc_hd__dfrtp_1  VNB VPB CLK D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_27_47#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_193_47#_M1012_d N_A_27_47#_M1012_g N_VGND_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_448_47#_M1025_d N_D_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.2205 PD=0.802308 PS=1.89 NRD=0 NRS=68.568 M=1 R=2.8
+ SA=75000.4 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_543_47#_M1008_d N_A_27_47#_M1008_g N_A_448_47#_M1025_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0594 AS=0.0609231 PD=0.69 PS=0.687692 NRD=18.324 NRS=16.656
+ M=1 R=2.4 SA=75000.9 SB=75005.2 A=0.054 P=1.02 MULT=1
MM1017 A_639_47# N_A_193_47#_M1017_g N_A_543_47#_M1008_d VNB NSHORT L=0.15
+ W=0.36 AD=0.129323 AS=0.0594 PD=1.01538 PS=0.69 NRD=101.4 NRS=0 M=1 R=2.4
+ SA=75001.4 SB=75004.8 A=0.054 P=1.02 MULT=1
MM1002 A_805_47# N_A_761_289#_M1002_g A_639_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.150877 PD=0.63 PS=1.18462 NRD=14.28 NRS=86.916 M=1 R=2.8
+ SA=75002 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_805_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.106664 AS=0.0441 PD=0.911321 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75002.3 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_761_289#_M1019_d N_A_543_47#_M1019_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.64 AD=0.127872 AS=0.162536 PD=1.2608 PS=1.38868 NRD=2.808 NRS=21.552 M=1
+ R=4.26667 SA=75002 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_1108_47#_M1020_d N_A_193_47#_M1020_g N_A_761_289#_M1019_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0711 AS=0.071928 PD=0.755 PS=0.7092 NRD=23.328 NRS=16.656
+ M=1 R=2.4 SA=75003.7 SB=75002.4 A=0.054 P=1.02 MULT=1
MM1018 A_1217_47# N_A_27_47#_M1018_g N_A_1108_47#_M1020_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0617538 AS=0.0711 PD=0.692308 PS=0.755 NRD=38.844 NRS=14.988 M=1
+ R=2.4 SA=75004.3 SB=75001.9 A=0.054 P=1.02 MULT=1
MM1022 N_VGND_M1022_d N_A_1283_21#_M1022_g A_1217_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.12495 AS=0.0720462 PD=1.015 PS=0.807692 NRD=30 NRS=33.288 M=1 R=2.8
+ SA=75004.1 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 A_1462_47# N_RESET_B_M1004_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06405 AS=0.12495 PD=0.725 PS=1.015 NRD=27.852 NRS=59.988 M=1 R=2.8
+ SA=75004.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_1283_21#_M1001_d N_A_1108_47#_M1001_g A_1462_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.06405 PD=1.36 PS=0.725 NRD=0 NRS=27.852 M=1 R=2.8
+ SA=75005.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_Q_M1005_d N_A_1283_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.2087 PD=1.82 PS=2.02 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_CLK_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_A_448_47#_M1024_d N_D_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0651 AS=0.1092 PD=0.73 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1026 N_A_543_47#_M1026_d N_A_193_47#_M1026_g N_A_448_47#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.07245 AS=0.0651 PD=0.765 PS=0.73 NRD=0 NRS=16.4101 M=1
+ R=2.8 SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_651_413#_M1006_d N_A_27_47#_M1006_g N_A_543_47#_M1026_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1155 AS=0.07245 PD=0.97 PS=0.765 NRD=128.976 NRS=30.4759
+ M=1 R=2.8 SA=75001.1 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_761_289#_M1009_g N_A_651_413#_M1006_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.07035 AS=0.1155 PD=0.755 PS=0.97 NRD=28.1316 NRS=0 M=1
+ R=2.8 SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_A_651_413#_M1027_d N_RESET_B_M1027_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.07035 PD=1.36 PS=0.755 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_761_289#_M1014_d N_A_543_47#_M1014_g N_VPWR_M1014_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1722 AS=0.2184 PD=1.58 PS=2.2 NRD=3.5066 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1021 N_A_1108_47#_M1021_d N_A_27_47#_M1021_g N_A_761_289#_M1014_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0861 PD=0.7 PS=0.79 NRD=2.3443 NRS=23.443 M=1
+ R=2.8 SA=75000.7 SB=75002 A=0.063 P=1.14 MULT=1
MM1010 A_1270_413# N_A_193_47#_M1010_g N_A_1108_47#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0588 PD=0.69 PS=0.7 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_1283_21#_M1007_g A_1270_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0567 PD=0.81 PS=0.69 NRD=53.9386 NRS=37.5088 M=1 R=2.8
+ SA=75001.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_1283_21#_M1016_d N_RESET_B_M1016_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0819 PD=0.69 PS=0.81 NRD=0 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_1108_47#_M1013_g N_A_1283_21#_M1016_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1134 AS=0.0567 PD=1.38 PS=0.69 NRD=2.3443 NRS=0 M=1 R=2.8
+ SA=75002.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_Q_M1015_d N_A_1283_21#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.3012 PD=2.52 PS=2.66 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.3759 P=22.37
c_93 VNB 0 1.85993e-19 $X=0.145 $Y=-0.085
c_192 VPB 0 1.60161e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dfrtp_1.pxi.spice"
*
.ends
*
*

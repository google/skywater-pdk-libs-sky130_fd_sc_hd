* File: sky130_fd_sc_hd__mux2i_1.spice
* Created: Thu Aug 27 14:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2i_1.pex.spice"
.subckt sky130_fd_sc_hd__mux2i_1  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_A0_M1007_g N_A_27_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1005 N_A_193_47#_M1005_d N_A1_M1005_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_283_205#_M1009_g N_A_27_47#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_193_47#_M1002_d N_S_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_S_M1006_g N_A_283_205#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_A0_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.28 PD=1.305 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1001 A_204_297# N_A1_M1001_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.1975
+ AS=0.1525 PD=1.395 PS=1.305 NRD=28.0528 NRS=5.8903 M=1 R=6.66667 SA=75000.7
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_283_205#_M1004_g A_204_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.3 AS=0.1975 PD=1.6 PS=1.395 NRD=24.6053 NRS=28.0528 M=1 R=6.66667
+ SA=75001.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_297#_M1008_d N_S_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.3 PD=2.52 PS=1.6 NRD=0 NRS=38.3953 M=1 R=6.66667 SA=75002
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_S_M1000_g N_A_283_205#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.29 PD=2.52 PS=2.58 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_64 VPB 0 1.55727e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__mux2i_1.pxi.spice"
*
.ends
*
*

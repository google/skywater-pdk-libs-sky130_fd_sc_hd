* File: sky130_fd_sc_hd__a31o_2.spice
* Created: Thu Aug 27 14:04:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a31o_2.pex.spice"
.subckt sky130_fd_sc_hd__a31o_2  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_79_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_79_21#_M1011_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1008 A_277_47# N_A3_M1008_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1007 A_361_47# N_A2_M1007_g A_277_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=14.76 M=1 R=4.33333 SA=75001.4
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_79_21#_M1000_d N_A1_M1000_g A_361_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.10725 PD=1.04 PS=0.98 NRD=21.228 NRS=20.304 M=1 R=4.33333
+ SA=75001.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_A_79_21#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12675 PD=1.82 PS=1.04 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_79_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_79_21#_M1009_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_A_277_297#_M1001_d N_A3_M1001_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A2_M1010_g N_A_277_297#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_277_297#_M1006_d N_A1_M1006_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.165 PD=1.33 PS=1.33 NRD=10.8153 NRS=2.9353 M=1 R=6.66667
+ SA=75001.9 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1002 N_A_79_21#_M1002_d N_B1_M1002_g N_A_277_297#_M1006_d VPB PHIGHVT L=0.15
+ W=1 AD=0.32 AS=0.165 PD=2.64 PS=1.33 NRD=10.8153 NRS=0 M=1 R=6.66667
+ SA=75002.4 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a31o_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__or2b_4.spice
* Created: Tue Sep  1 19:27:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or2b_4.pex.spice"
.subckt sky130_fd_sc_hd__or2b_4  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B_N_M1002_g N_A_27_53#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.158403 AS=0.1092 PD=1.09907 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1012 N_A_219_297#_M1012_d N_A_27_53#_M1012_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.245147 PD=0.92 PS=1.70093 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.8 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_219_297#_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1105 AS=0.08775 PD=0.99 PS=0.92 NRD=11.988 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_219_297#_M1003_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1105 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1003_d N_A_219_297#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_219_297#_M1006_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1006_d N_A_219_297#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2145 PD=0.92 PS=1.96 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_53#_M1005_d N_B_N_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1176 AS=0.1092 PD=1.4 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 A_301_297# N_A_27_53#_M1007_g N_A_219_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.26 PD=1.21 PS=2.52 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_301_297# VPB PHIGHVT L=0.15 W=1 AD=0.17
+ AS=0.105 PD=1.34 PS=1.21 NRD=11.8003 NRS=9.8303 M=1 R=6.66667 SA=75000.5
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_219_297#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.17 PD=1.27 PS=1.34 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1001 N_X_M1000_d N_A_219_297#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1011_d N_A_219_297#_M1011_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1011_d N_A_219_297#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__or2b_4.pxi.spice"
*
.ends
*
*

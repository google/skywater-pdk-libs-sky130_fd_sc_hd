* File: sky130_fd_sc_hd__o311a_1.spice.SKY130_FD_SC_HD__O311A_1.pxi
* Created: Thu Aug 27 14:38:56 2020
* 
x_PM_SKY130_FD_SC_HD__O311A_1%A_81_21# N_A_81_21#_M1010_d N_A_81_21#_M1011_d
+ N_A_81_21#_M1000_d N_A_81_21#_c_64_n N_A_81_21#_M1001_g N_A_81_21#_M1005_g
+ N_A_81_21#_c_65_n N_A_81_21#_c_66_n N_A_81_21#_c_77_p N_A_81_21#_c_124_p
+ N_A_81_21#_c_78_p N_A_81_21#_c_87_p N_A_81_21#_c_79_p N_A_81_21#_c_91_p
+ N_A_81_21#_c_88_p N_A_81_21#_c_97_p N_A_81_21#_c_93_p N_A_81_21#_c_67_n
+ N_A_81_21#_c_73_n N_A_81_21#_c_74_n N_A_81_21#_c_68_n
+ PM_SKY130_FD_SC_HD__O311A_1%A_81_21#
x_PM_SKY130_FD_SC_HD__O311A_1%A1 N_A1_M1003_g N_A1_M1002_g A1 N_A1_c_164_n
+ N_A1_c_165_n PM_SKY130_FD_SC_HD__O311A_1%A1
x_PM_SKY130_FD_SC_HD__O311A_1%A2 N_A2_M1006_g N_A2_M1004_g A2 A2 A2 N_A2_c_196_n
+ N_A2_c_197_n N_A2_c_198_n PM_SKY130_FD_SC_HD__O311A_1%A2
x_PM_SKY130_FD_SC_HD__O311A_1%A3 N_A3_M1008_g N_A3_M1011_g A3 A3 A3 N_A3_c_232_n
+ N_A3_c_233_n N_A3_c_234_n PM_SKY130_FD_SC_HD__O311A_1%A3
x_PM_SKY130_FD_SC_HD__O311A_1%B1 N_B1_M1007_g N_B1_M1009_g B1 N_B1_c_267_n
+ N_B1_c_268_n N_B1_c_269_n PM_SKY130_FD_SC_HD__O311A_1%B1
x_PM_SKY130_FD_SC_HD__O311A_1%C1 N_C1_c_302_n N_C1_M1010_g N_C1_M1000_g C1
+ N_C1_c_304_n PM_SKY130_FD_SC_HD__O311A_1%C1
x_PM_SKY130_FD_SC_HD__O311A_1%X N_X_M1001_s N_X_M1005_s X X X X X X X
+ PM_SKY130_FD_SC_HD__O311A_1%X
x_PM_SKY130_FD_SC_HD__O311A_1%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_c_343_n
+ N_VPWR_c_344_n VPWR N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n
+ N_VPWR_c_342_n N_VPWR_c_349_n N_VPWR_c_350_n VPWR
+ PM_SKY130_FD_SC_HD__O311A_1%VPWR
x_PM_SKY130_FD_SC_HD__O311A_1%VGND N_VGND_M1001_d N_VGND_M1006_d N_VGND_c_401_n
+ N_VGND_c_402_n VGND N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n
+ N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n VGND
+ PM_SKY130_FD_SC_HD__O311A_1%VGND
x_PM_SKY130_FD_SC_HD__O311A_1%A_266_47# N_A_266_47#_M1003_d N_A_266_47#_M1008_d
+ N_A_266_47#_c_461_n N_A_266_47#_c_449_n N_A_266_47#_c_452_n
+ N_A_266_47#_c_457_n N_A_266_47#_c_468_n PM_SKY130_FD_SC_HD__O311A_1%A_266_47#
cc_1 VNB N_A_81_21#_c_64_n 0.0215929f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_A_81_21#_c_65_n 0.00157408f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_3 VNB N_A_81_21#_c_66_n 0.0350059f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_4 VNB N_A_81_21#_c_67_n 0.00281491f $X=-0.19 $Y=-0.24 $X2=3.095 $Y2=1.495
cc_5 VNB N_A_81_21#_c_68_n 0.0245152f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.4
cc_6 VNB A1 0.00290387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A1_c_164_n 0.0207716f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_8 VNB N_A1_c_165_n 0.0195561f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_9 VNB N_A2_c_196_n 0.020988f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.985
cc_10 VNB N_A2_c_197_n 0.00407077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_198_n 0.0185336f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.495
cc_12 VNB N_A3_c_232_n 0.0261176f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.985
cc_13 VNB N_A3_c_233_n 0.00452535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A3_c_234_n 0.0185884f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.495
cc_15 VNB N_B1_c_267_n 0.0226542f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_16 VNB N_B1_c_268_n 0.00347516f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_17 VNB N_B1_c_269_n 0.0167081f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_18 VNB N_C1_c_302_n 0.0209378f $X=-0.19 $Y=-0.24 $X2=3.285 $Y2=0.235
cc_19 VNB C1 0.0133884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_C1_c_304_n 0.0344721f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_21 VNB X 0.0339008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB X 0.0120233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_342_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.715 $Y2=1.58
cc_24 VNB N_VGND_c_401_n 0.00187948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_402_n 0.00530857f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_26 VNB N_VGND_c_403_n 0.0152818f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.495
cc_27 VNB N_VGND_c_404_n 0.0161623f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.58
cc_28 VNB N_VGND_c_405_n 0.0394108f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.58
cc_29 VNB N_VGND_c_406_n 0.199543f $X=-0.19 $Y=-0.24 $X2=2.715 $Y2=1.58
cc_30 VNB N_VGND_c_407_n 0.0104906f $X=-0.19 $Y=-0.24 $X2=3.45 $Y2=1.665
cc_31 VNB N_VGND_c_408_n 0.00718038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_81_21#_M1005_g 0.0261763f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_33 VPB N_A_81_21#_c_65_n 0.00280012f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_34 VPB N_A_81_21#_c_66_n 0.0104131f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_35 VPB N_A_81_21#_c_67_n 0.00165139f $X=-0.19 $Y=1.305 $X2=3.095 $Y2=1.495
cc_36 VPB N_A_81_21#_c_73_n 0.00763029f $X=-0.19 $Y=1.305 $X2=3.45 $Y2=1.665
cc_37 VPB N_A_81_21#_c_74_n 0.0312708f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=1.815
cc_38 VPB N_A1_M1002_g 0.0230681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB A1 0.0011816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A1_c_164_n 0.00404249f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_41 VPB N_A2_M1004_g 0.0206081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB A2 0.00163815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A2_c_196_n 0.00453712f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_44 VPB N_A2_c_197_n 0.00268647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A3_M1011_g 0.0206248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB A3 0.00247089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A3_c_232_n 0.00728583f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_48 VPB N_A3_c_233_n 0.0018022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_B1_M1007_g 0.0195048f $X=-0.19 $Y=1.305 $X2=3.285 $Y2=1.485
cc_50 VPB N_B1_c_267_n 0.00509613f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_51 VPB N_B1_c_268_n 0.00178038f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_52 VPB N_C1_M1000_g 0.0257003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB C1 0.00297249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_C1_c_304_n 0.0096974f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.325
cc_55 VPB X 0.0470377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_343_n 0.00595658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_344_n 0.00509471f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.325
cc_58 VPB N_VPWR_c_345_n 0.0179959f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.495
cc_59 VPB N_VPWR_c_346_n 0.0450745f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.58
cc_60 VPB N_VPWR_c_347_n 0.0167769f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.58
cc_61 VPB N_VPWR_c_342_n 0.0437521f $X=-0.19 $Y=1.305 $X2=2.715 $Y2=1.58
cc_62 VPB N_VPWR_c_349_n 0.00775716f $X=-0.19 $Y=1.305 $X2=3.45 $Y2=1.665
cc_63 VPB N_VPWR_c_350_n 0.00449427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 N_A_81_21#_M1005_g N_A1_M1002_g 0.0161896f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A_81_21#_c_65_n N_A1_M1002_g 0.00301901f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_81_21#_c_77_p N_A1_M1002_g 0.0105598f $X=1.18 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A_81_21#_c_78_p N_A1_M1002_g 0.0171212f $X=1.265 $Y=2.295 $X2=0 $Y2=0
cc_68 N_A_81_21#_c_79_p N_A1_M1002_g 0.00610252f $X=1.35 $Y=2.38 $X2=0 $Y2=0
cc_69 N_A_81_21#_c_65_n A1 0.024918f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_81_21#_c_66_n A1 0.00223817f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_81_21#_c_77_p A1 0.0237374f $X=1.18 $Y=1.58 $X2=0 $Y2=0
cc_72 N_A_81_21#_c_65_n N_A1_c_164_n 3.10952e-19 $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_81_21#_c_66_n N_A1_c_164_n 0.0180431f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_81_21#_c_77_p N_A1_c_164_n 0.00256542f $X=1.18 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A_81_21#_c_64_n N_A1_c_165_n 0.00425898f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_81_21#_c_87_p N_A2_M1004_g 0.0125311f $X=2.385 $Y=2.38 $X2=0 $Y2=0
cc_77 N_A_81_21#_c_88_p N_A2_M1004_g 0.00110498f $X=2.55 $Y=1.68 $X2=0 $Y2=0
cc_78 N_A_81_21#_c_87_p A2 0.0121614f $X=2.385 $Y=2.38 $X2=0 $Y2=0
cc_79 N_A_81_21#_c_87_p N_A3_M1011_g 0.011169f $X=2.385 $Y=2.38 $X2=0 $Y2=0
cc_80 N_A_81_21#_c_91_p N_A3_M1011_g 5.89792e-19 $X=2.55 $Y=2.295 $X2=0 $Y2=0
cc_81 N_A_81_21#_c_88_p N_A3_M1011_g 0.00872665f $X=2.55 $Y=1.68 $X2=0 $Y2=0
cc_82 N_A_81_21#_c_93_p N_A3_M1011_g 0.00249995f $X=2.715 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_81_21#_c_87_p A3 0.0132929f $X=2.385 $Y=2.38 $X2=0 $Y2=0
cc_84 N_A_81_21#_c_91_p N_B1_M1007_g 0.00209677f $X=2.55 $Y=2.295 $X2=0 $Y2=0
cc_85 N_A_81_21#_c_88_p N_B1_M1007_g 0.00815505f $X=2.55 $Y=1.68 $X2=0 $Y2=0
cc_86 N_A_81_21#_c_97_p N_B1_M1007_g 0.0108502f $X=3.01 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_81_21#_c_93_p N_B1_M1007_g 8.84614e-19 $X=2.715 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_81_21#_c_67_n N_B1_M1007_g 0.00352622f $X=3.095 $Y=1.495 $X2=0 $Y2=0
cc_89 N_A_81_21#_c_97_p N_B1_c_267_n 0.0027472f $X=3.01 $Y=1.58 $X2=0 $Y2=0
cc_90 N_A_81_21#_c_93_p N_B1_c_267_n 0.00134053f $X=2.715 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_81_21#_c_67_n N_B1_c_267_n 0.00573092f $X=3.095 $Y=1.495 $X2=0 $Y2=0
cc_92 N_A_81_21#_c_97_p N_B1_c_268_n 0.00872323f $X=3.01 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A_81_21#_c_93_p N_B1_c_268_n 0.0195547f $X=2.715 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_81_21#_c_67_n N_B1_c_268_n 0.0251379f $X=3.095 $Y=1.495 $X2=0 $Y2=0
cc_95 N_A_81_21#_c_68_n N_B1_c_269_n 0.00573092f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_96 N_A_81_21#_c_67_n N_C1_c_302_n 0.00789512f $X=3.095 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_81_21#_c_68_n N_C1_c_302_n 0.0150777f $X=3.42 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_81_21#_c_88_p N_C1_M1000_g 5.87886e-19 $X=2.55 $Y=1.68 $X2=0 $Y2=0
cc_99 N_A_81_21#_c_67_n N_C1_M1000_g 0.0084555f $X=3.095 $Y=1.495 $X2=0 $Y2=0
cc_100 N_A_81_21#_c_73_n N_C1_M1000_g 0.0166705f $X=3.45 $Y=1.665 $X2=0 $Y2=0
cc_101 N_A_81_21#_c_67_n C1 0.0230137f $X=3.095 $Y=1.495 $X2=0 $Y2=0
cc_102 N_A_81_21#_c_73_n C1 0.0181761f $X=3.45 $Y=1.665 $X2=0 $Y2=0
cc_103 N_A_81_21#_c_68_n C1 0.0200459f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_104 N_A_81_21#_c_67_n N_C1_c_304_n 0.00752413f $X=3.095 $Y=1.495 $X2=0 $Y2=0
cc_105 N_A_81_21#_c_73_n N_C1_c_304_n 0.00297804f $X=3.45 $Y=1.665 $X2=0 $Y2=0
cc_106 N_A_81_21#_c_68_n N_C1_c_304_n 0.00315879f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_107 N_A_81_21#_c_64_n X 0.0112728f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_81_21#_c_65_n X 0.00414841f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_81_21#_M1005_g X 0.0216151f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_81_21#_c_65_n X 0.0306398f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_81_21#_c_66_n X 0.0108521f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_81_21#_c_77_p N_VPWR_M1005_d 0.0138071f $X=1.18 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_81_21#_c_124_p N_VPWR_M1005_d 0.00321774f $X=0.775 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_81_21#_c_97_p N_VPWR_M1007_d 0.00507927f $X=3.01 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A_81_21#_c_67_n N_VPWR_M1007_d 3.14485e-19 $X=3.095 $Y=1.495 $X2=0
+ $Y2=0
cc_116 N_A_81_21#_c_73_n N_VPWR_M1007_d 9.10335e-19 $X=3.45 $Y=1.665 $X2=0 $Y2=0
cc_117 N_A_81_21#_M1005_g N_VPWR_c_343_n 0.00874064f $X=0.48 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_81_21#_c_66_n N_VPWR_c_343_n 7.36359e-19 $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_81_21#_c_77_p N_VPWR_c_343_n 0.0190014f $X=1.18 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A_81_21#_c_124_p N_VPWR_c_343_n 0.0146353f $X=0.775 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A_81_21#_c_78_p N_VPWR_c_343_n 0.0345753f $X=1.265 $Y=2.295 $X2=0 $Y2=0
cc_122 N_A_81_21#_c_79_p N_VPWR_c_343_n 0.0142211f $X=1.35 $Y=2.38 $X2=0 $Y2=0
cc_123 N_A_81_21#_c_91_p N_VPWR_c_344_n 0.0127992f $X=2.55 $Y=2.295 $X2=0 $Y2=0
cc_124 N_A_81_21#_c_88_p N_VPWR_c_344_n 0.032561f $X=2.55 $Y=1.68 $X2=0 $Y2=0
cc_125 N_A_81_21#_c_97_p N_VPWR_c_344_n 0.0143275f $X=3.01 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A_81_21#_M1005_g N_VPWR_c_345_n 0.00541359f $X=0.48 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_81_21#_c_87_p N_VPWR_c_346_n 0.0592194f $X=2.385 $Y=2.38 $X2=0 $Y2=0
cc_128 N_A_81_21#_c_79_p N_VPWR_c_346_n 0.0109366f $X=1.35 $Y=2.38 $X2=0 $Y2=0
cc_129 N_A_81_21#_c_91_p N_VPWR_c_346_n 0.019051f $X=2.55 $Y=2.295 $X2=0 $Y2=0
cc_130 N_A_81_21#_c_74_n N_VPWR_c_347_n 0.0190655f $X=3.42 $Y=1.815 $X2=0 $Y2=0
cc_131 N_A_81_21#_M1011_d N_VPWR_c_342_n 0.00219216f $X=2.41 $Y=1.485 $X2=0
+ $Y2=0
cc_132 N_A_81_21#_M1000_d N_VPWR_c_342_n 0.00283025f $X=3.285 $Y=1.485 $X2=0
+ $Y2=0
cc_133 N_A_81_21#_M1005_g N_VPWR_c_342_n 0.0112409f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_81_21#_c_87_p N_VPWR_c_342_n 0.0372911f $X=2.385 $Y=2.38 $X2=0 $Y2=0
cc_135 N_A_81_21#_c_79_p N_VPWR_c_342_n 0.00586103f $X=1.35 $Y=2.38 $X2=0 $Y2=0
cc_136 N_A_81_21#_c_91_p N_VPWR_c_342_n 0.0123125f $X=2.55 $Y=2.295 $X2=0 $Y2=0
cc_137 N_A_81_21#_c_74_n N_VPWR_c_342_n 0.0110914f $X=3.42 $Y=1.815 $X2=0 $Y2=0
cc_138 N_A_81_21#_c_87_p A_266_297# 0.00876975f $X=2.385 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_139 N_A_81_21#_c_87_p A_368_297# 0.00930583f $X=2.385 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_81_21#_c_64_n N_VGND_c_401_n 0.0144594f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_81_21#_c_65_n N_VGND_c_401_n 0.0143975f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_81_21#_c_66_n N_VGND_c_401_n 0.00286475f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_81_21#_c_77_p N_VGND_c_401_n 0.00488088f $X=1.18 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A_81_21#_c_64_n N_VGND_c_403_n 0.0046653f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_81_21#_c_68_n N_VGND_c_405_n 0.0364195f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_146 N_A_81_21#_M1010_d N_VGND_c_406_n 0.00209319f $X=3.285 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_81_21#_c_64_n N_VGND_c_406_n 0.00896841f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_81_21#_c_68_n N_VGND_c_406_n 0.0216215f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_149 N_A_81_21#_c_93_p N_A_266_47#_c_449_n 5.79016e-19 $X=2.715 $Y=1.58 $X2=0
+ $Y2=0
cc_150 N_A_81_21#_c_67_n A_585_47# 6.54266e-19 $X=3.095 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_81_21#_c_68_n A_585_47# 0.00644001f $X=3.42 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A1_M1002_g N_A2_M1004_g 0.0412933f $X=1.255 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A1_M1002_g A2 0.00586542f $X=1.255 $Y=1.985 $X2=0 $Y2=0
cc_154 A1 N_A2_c_196_n 3.08149e-19 $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A1_c_164_n N_A2_c_196_n 0.0169926f $X=1.195 $Y=1.16 $X2=0 $Y2=0
cc_156 A1 N_A2_c_197_n 0.0261733f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A1_c_164_n N_A2_c_197_n 0.0021587f $X=1.195 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A1_c_165_n N_A2_c_198_n 0.0173814f $X=1.195 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A1_M1002_g N_VPWR_c_343_n 0.00820357f $X=1.255 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A1_M1002_g N_VPWR_c_346_n 0.00357668f $X=1.255 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A1_M1002_g N_VPWR_c_342_n 0.00620538f $X=1.255 $Y=1.985 $X2=0 $Y2=0
cc_162 A1 N_VGND_c_401_n 0.0183964f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A1_c_164_n N_VGND_c_401_n 0.00262179f $X=1.195 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A1_c_165_n N_VGND_c_401_n 0.011102f $X=1.195 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_165_n N_VGND_c_404_n 0.00525069f $X=1.195 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_165_n N_VGND_c_406_n 0.00913058f $X=1.195 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_M1004_g N_A3_M1011_g 0.0302643f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A2_M1004_g A3 0.00390408f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_169 A2 A3 0.0374687f $X=1.52 $Y=1.445 $X2=0 $Y2=0
cc_170 N_A2_c_196_n N_A3_c_232_n 0.0202578f $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A2_c_197_n N_A3_c_232_n 3.33292e-19 $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_c_196_n N_A3_c_233_n 0.00390408f $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A2_c_197_n N_A3_c_233_n 0.0374687f $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A2_c_198_n N_A3_c_234_n 0.0235995f $X=1.705 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_VPWR_c_346_n 0.00357877f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A2_M1004_g N_VPWR_c_342_n 0.00587103f $X=1.765 $Y=1.985 $X2=0 $Y2=0
cc_177 A2 A_266_297# 0.00638515f $X=1.52 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_178 N_A2_c_198_n N_VGND_c_401_n 8.01811e-19 $X=1.705 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A2_c_198_n N_VGND_c_402_n 0.00365716f $X=1.705 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_198_n N_VGND_c_404_n 0.00427293f $X=1.705 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A2_c_198_n N_VGND_c_406_n 0.00628404f $X=1.705 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_197_n N_A_266_47#_c_449_n 0.00880508f $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A2_c_198_n N_A_266_47#_c_449_n 0.0129853f $X=1.705 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_196_n N_A_266_47#_c_452_n 6.16454e-19 $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A2_c_197_n N_A_266_47#_c_452_n 0.0169246f $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A3_M1011_g N_B1_M1007_g 0.0136218f $X=2.335 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A3_c_232_n N_B1_c_267_n 0.0204866f $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A3_c_233_n N_B1_c_267_n 2.38775e-19 $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A3_c_232_n N_B1_c_268_n 0.0025442f $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A3_c_233_n N_B1_c_268_n 0.0262419f $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A3_c_234_n N_B1_c_269_n 0.0087356f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A3_M1011_g N_VPWR_c_346_n 0.00357842f $X=2.335 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A3_M1011_g N_VPWR_c_342_n 0.00563013f $X=2.335 $Y=1.985 $X2=0 $Y2=0
cc_194 A3 A_368_297# 0.014726f $X=1.98 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_195 N_A3_c_234_n N_VGND_c_402_n 0.00467408f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A3_c_234_n N_VGND_c_405_n 0.00428022f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A3_c_234_n N_VGND_c_406_n 0.00635517f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A3_c_232_n N_A_266_47#_c_449_n 0.00135602f $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A3_c_233_n N_A_266_47#_c_449_n 0.0206113f $X=2.185 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A3_c_234_n N_A_266_47#_c_449_n 0.0144537f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B1_c_269_n N_C1_c_302_n 0.0368767f $X=2.772 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_202 N_B1_M1007_g N_C1_M1000_g 0.0246074f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_c_267_n N_C1_c_304_n 0.0368767f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B1_c_268_n N_C1_c_304_n 2.80449e-19 $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B1_M1007_g N_VPWR_c_344_n 0.00510038f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B1_M1007_g N_VPWR_c_346_n 0.00539841f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1007_g N_VPWR_c_342_n 0.00964112f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_c_269_n N_VGND_c_405_n 0.00585385f $X=2.772 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B1_c_269_n N_VGND_c_406_n 0.0108442f $X=2.772 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B1_c_267_n N_A_266_47#_c_457_n 0.00340725f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B1_c_268_n N_A_266_47#_c_457_n 0.0236139f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_212 N_C1_M1000_g N_VPWR_c_344_n 0.00307308f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_213 N_C1_M1000_g N_VPWR_c_347_n 0.00583607f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_214 N_C1_M1000_g N_VPWR_c_342_n 0.0115712f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_215 N_C1_c_302_n N_VGND_c_405_n 0.00357668f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_216 N_C1_c_302_n N_VGND_c_406_n 0.00604465f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_217 X N_VPWR_c_345_n 0.0224721f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_218 N_X_M1005_s N_VPWR_c_342_n 0.00209319f $X=0.145 $Y=1.485 $X2=0 $Y2=0
cc_219 X N_VPWR_c_342_n 0.013197f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_220 X N_VGND_c_403_n 0.018718f $X=0.14 $Y=0.425 $X2=0 $Y2=0
cc_221 N_X_M1001_s N_VGND_c_406_n 0.00387172f $X=0.145 $Y=0.235 $X2=0 $Y2=0
cc_222 X N_VGND_c_406_n 0.0103212f $X=0.14 $Y=0.425 $X2=0 $Y2=0
cc_223 N_VPWR_c_342_n A_266_297# 0.00289109f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_224 N_VPWR_c_342_n A_368_297# 0.00338304f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_225 N_VGND_c_406_n N_A_266_47#_M1003_d 0.00429284f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_226 N_VGND_c_406_n N_A_266_47#_M1008_d 0.00354962f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_404_n N_A_266_47#_c_461_n 0.0137779f $X=1.84 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_406_n N_A_266_47#_c_461_n 0.0108787f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_M1006_d N_A_266_47#_c_449_n 0.00888498f $X=1.84 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_VGND_c_402_n N_A_266_47#_c_449_n 0.0234908f $X=2.05 $Y=0.36 $X2=0 $Y2=0
cc_231 N_VGND_c_404_n N_A_266_47#_c_449_n 0.00260706f $X=1.84 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_405_n N_A_266_47#_c_449_n 0.00293207f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_406_n N_A_266_47#_c_449_n 0.0110612f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_405_n N_A_266_47#_c_468_n 0.0148394f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_406_n N_A_266_47#_c_468_n 0.0121783f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_406_n A_585_47# 0.00467183f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 1.005000 2.170000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.115000 0.255000 12.345000 0.825000 ;
        RECT 12.115000 1.445000 12.345000 2.465000 ;
        RECT 12.160000 0.825000 12.345000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.240000 0.255000 10.500000 0.715000 ;
        RECT 10.240000 1.630000 10.500000 2.465000 ;
        RECT 10.320000 0.715000 10.500000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.250000 1.095000 9.730000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.600000 0.735000 4.010000 0.965000 ;
        RECT 3.600000 0.965000 3.930000 1.065000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.470000 0.735000 7.845000 1.065000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.780000 0.735000 4.070000 0.780000 ;
        RECT 3.780000 0.780000 7.750000 0.920000 ;
        RECT 3.780000 0.920000 4.070000 0.965000 ;
        RECT 7.460000 0.735000 7.750000 0.780000 ;
        RECT 7.460000 0.920000 7.750000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.440000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.880000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  1.445000  0.085000  1.785000 0.465000 ;
        RECT  3.580000  0.085000  3.750000 0.525000 ;
        RECT  5.360000  0.085000  5.690000 0.465000 ;
        RECT  7.275000  0.085000  7.535000 0.525000 ;
        RECT  9.740000  0.085000 10.070000 0.805000 ;
        RECT 10.680000  0.085000 10.910000 0.885000 ;
        RECT 11.650000  0.085000 11.945000 0.545000 ;
        RECT 12.515000  0.085000 12.795000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 12.880000 2.805000 ;
        RECT  0.515000 2.135000  0.845000 2.635000 ;
        RECT  1.445000 2.135000  1.785000 2.635000 ;
        RECT  3.420000 2.205000  3.800000 2.635000 ;
        RECT  4.890000 1.915000  5.220000 2.635000 ;
        RECT  7.335000 2.255000  7.715000 2.635000 ;
        RECT  8.655000 2.255000 10.070000 2.635000 ;
        RECT 10.680000 1.465000 10.910000 2.635000 ;
        RECT 11.650000 1.765000 11.945000 2.635000 ;
        RECT 12.515000 1.465000 12.795000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.345000  0.345000 0.635000 ;
      RECT  0.085000 0.635000  0.840000 0.805000 ;
      RECT  0.085000 1.795000  0.840000 1.965000 ;
      RECT  0.085000 1.965000  0.345000 2.465000 ;
      RECT  0.610000 0.805000  0.840000 1.795000 ;
      RECT  1.015000 0.345000  1.240000 2.465000 ;
      RECT  1.420000 0.635000  2.125000 0.825000 ;
      RECT  1.420000 0.825000  1.590000 1.795000 ;
      RECT  1.420000 1.795000  2.125000 1.965000 ;
      RECT  1.955000 0.305000  2.125000 0.635000 ;
      RECT  1.955000 1.965000  2.125000 2.465000 ;
      RECT  2.340000 0.705000  2.560000 1.575000 ;
      RECT  2.340000 1.575000  2.840000 1.955000 ;
      RECT  2.350000 2.250000  3.180000 2.420000 ;
      RECT  2.415000 0.265000  3.410000 0.465000 ;
      RECT  2.740000 0.645000  3.070000 1.015000 ;
      RECT  3.010000 1.195000  3.410000 1.235000 ;
      RECT  3.010000 1.235000  4.360000 1.405000 ;
      RECT  3.010000 1.405000  3.180000 2.250000 ;
      RECT  3.240000 0.465000  3.410000 1.195000 ;
      RECT  3.350000 1.575000  3.600000 1.785000 ;
      RECT  3.350000 1.785000  4.700000 2.035000 ;
      RECT  3.920000 0.255000  5.170000 0.425000 ;
      RECT  3.920000 0.425000  4.250000 0.545000 ;
      RECT  4.100000 2.035000  4.270000 2.375000 ;
      RECT  4.110000 1.405000  4.360000 1.485000 ;
      RECT  4.140000 1.155000  4.360000 1.235000 ;
      RECT  4.420000 0.595000  4.750000 0.765000 ;
      RECT  4.530000 0.765000  4.750000 0.895000 ;
      RECT  4.530000 0.895000  5.840000 1.065000 ;
      RECT  4.530000 1.065000  4.700000 1.785000 ;
      RECT  4.870000 1.235000  5.200000 1.415000 ;
      RECT  4.870000 1.415000  5.875000 1.655000 ;
      RECT  4.920000 0.425000  5.170000 0.715000 ;
      RECT  5.510000 1.065000  5.840000 1.235000 ;
      RECT  6.075000 1.575000  6.310000 1.985000 ;
      RECT  6.135000 0.705000  6.420000 1.125000 ;
      RECT  6.135000 1.125000  6.755000 1.305000 ;
      RECT  6.265000 2.250000  7.095000 2.420000 ;
      RECT  6.330000 0.265000  7.095000 0.465000 ;
      RECT  6.550000 1.305000  6.755000 1.905000 ;
      RECT  6.925000 0.465000  7.095000 1.235000 ;
      RECT  6.925000 1.235000  8.275000 1.405000 ;
      RECT  6.925000 1.405000  7.095000 2.250000 ;
      RECT  7.265000 1.575000  7.515000 1.915000 ;
      RECT  7.265000 1.915000 10.070000 2.085000 ;
      RECT  7.795000 0.255000  8.965000 0.425000 ;
      RECT  7.795000 0.425000  8.125000 0.545000 ;
      RECT  7.955000 2.085000  8.125000 2.375000 ;
      RECT  8.055000 1.075000  8.275000 1.235000 ;
      RECT  8.295000 0.595000  8.625000 0.780000 ;
      RECT  8.445000 0.780000  8.625000 1.915000 ;
      RECT  8.795000 0.425000  8.965000 0.585000 ;
      RECT  8.795000 0.755000  9.500000 0.925000 ;
      RECT  8.795000 0.925000  9.070000 1.575000 ;
      RECT  8.795000 1.575000  9.570000 1.745000 ;
      RECT  9.280000 0.265000  9.500000 0.755000 ;
      RECT  9.900000 0.995000 10.140000 1.325000 ;
      RECT  9.900000 1.325000 10.070000 1.915000 ;
      RECT 11.215000 0.255000 11.470000 0.995000 ;
      RECT 11.215000 0.995000 11.990000 1.325000 ;
      RECT 11.215000 1.325000 11.470000 2.415000 ;
    LAYER mcon ;
      RECT 0.610000 0.765000 0.780000 0.935000 ;
      RECT 1.070000 1.785000 1.240000 1.955000 ;
      RECT 2.460000 1.785000 2.630000 1.955000 ;
      RECT 2.900000 0.765000 3.070000 0.935000 ;
      RECT 5.680000 1.445000 5.850000 1.615000 ;
      RECT 6.140000 1.105000 6.310000 1.275000 ;
      RECT 6.140000 1.785000 6.310000 1.955000 ;
      RECT 8.900000 1.445000 9.070000 1.615000 ;
    LAYER met1 ;
      RECT 0.550000 0.735000 0.840000 0.780000 ;
      RECT 0.550000 0.780000 3.130000 0.920000 ;
      RECT 0.550000 0.920000 0.840000 0.965000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 6.370000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.400000 1.755000 2.690000 1.800000 ;
      RECT 2.400000 1.940000 2.690000 1.985000 ;
      RECT 2.840000 0.735000 3.130000 0.780000 ;
      RECT 2.840000 0.920000 3.130000 0.965000 ;
      RECT 2.935000 0.965000 3.130000 1.120000 ;
      RECT 2.935000 1.120000 6.370000 1.260000 ;
      RECT 5.620000 1.415000 5.910000 1.460000 ;
      RECT 5.620000 1.460000 9.130000 1.600000 ;
      RECT 5.620000 1.600000 5.910000 1.645000 ;
      RECT 6.080000 1.075000 6.370000 1.120000 ;
      RECT 6.080000 1.260000 6.370000 1.305000 ;
      RECT 6.080000 1.755000 6.370000 1.800000 ;
      RECT 6.080000 1.940000 6.370000 1.985000 ;
      RECT 8.840000 1.415000 9.130000 1.460000 ;
      RECT 8.840000 1.600000 9.130000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbn_2

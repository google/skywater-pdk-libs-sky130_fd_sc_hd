* NGSPICE file created from sky130_fd_sc_hd__dfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.5449e+12p ps=1.575e+07u
M1001 VPWR SET_B a_1028_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.73e+11p ps=2.98e+06u
M1002 VGND SET_B a_1300_47# VNB nshort w=420000u l=150000u
+  ad=1.1373e+12p pd=1.19e+07u as=8.82e+10p ps=1.26e+06u
M1003 VGND a_1602_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1004 a_796_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 a_1028_413# a_27_47# a_956_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VPWR a_1028_413# a_1602_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1007 a_652_21# a_476_47# a_796_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1008 Q a_1602_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_652_21# a_562_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.89e+11p ps=1.74e+06u
M1010 a_381_47# D VGND VNB nshort w=640000u l=150000u
+  ad=1.87e+11p pd=1.93e+06u as=0p ps=0u
M1011 a_476_47# a_193_47# a_381_47# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=2.499e+11p ps=2.35e+06u
M1012 a_1228_47# a_27_47# a_1028_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.47e+11p ps=1.54e+06u
M1013 a_1178_261# a_1028_413# VGND VNB nshort w=540000u l=150000u
+  ad=1.404e+11p pd=1.6e+06u as=0p ps=0u
M1014 a_1028_413# a_193_47# a_1056_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1015 VPWR a_1178_261# a_1136_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1016 a_956_413# a_476_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR CLK a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1018 a_586_47# a_193_47# a_476_47# VNB nshort w=360000u l=150000u
+  ad=1.341e+11p pd=1.5e+06u as=1.44e+11p ps=1.52e+06u
M1019 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1020 VPWR a_476_47# a_652_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1021 a_1056_47# a_476_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_652_21# a_586_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_381_47# D VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1136_413# a_193_47# a_1028_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1602_47# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1026 a_652_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1178_261# a_1028_413# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1028 a_476_47# a_27_47# a_381_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1030 VGND a_1028_413# a_1602_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1031 a_562_413# a_27_47# a_476_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_1602_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1300_47# a_1178_261# a_1228_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


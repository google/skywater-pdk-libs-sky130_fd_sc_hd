* File: sky130_fd_sc_hd__sdfrtp_4.pxi.spice
* Created: Tue Sep  1 19:30:24 2020
* 
x_PM_SKY130_FD_SC_HD__SDFRTP_4%CLK N_CLK_c_273_n N_CLK_M1036_g N_CLK_M1029_g CLK
+ CLK N_CLK_c_275_n PM_SKY130_FD_SC_HD__SDFRTP_4%CLK
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_27_47# N_A_27_47#_M1036_s N_A_27_47#_M1029_s
+ N_A_27_47#_c_304_n N_A_27_47#_M1022_g N_A_27_47#_M1041_g N_A_27_47#_c_305_n
+ N_A_27_47#_c_306_n N_A_27_47#_M1023_g N_A_27_47#_M1005_g N_A_27_47#_c_307_n
+ N_A_27_47#_M1001_g N_A_27_47#_M1011_g N_A_27_47#_c_309_n N_A_27_47#_c_310_n
+ N_A_27_47#_c_339_n N_A_27_47#_c_311_n N_A_27_47#_c_343_n N_A_27_47#_c_328_n
+ N_A_27_47#_c_329_n N_A_27_47#_c_312_n N_A_27_47#_c_313_n N_A_27_47#_c_314_n
+ N_A_27_47#_c_424_p N_A_27_47#_c_315_n N_A_27_47#_c_316_n N_A_27_47#_c_317_n
+ N_A_27_47#_c_318_n N_A_27_47#_c_319_n N_A_27_47#_c_320_n N_A_27_47#_c_321_n
+ N_A_27_47#_c_322_n PM_SKY130_FD_SC_HD__SDFRTP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_299_66# N_A_299_66#_M1025_s N_A_299_66#_M1006_s
+ N_A_299_66#_c_567_n N_A_299_66#_M1009_g N_A_299_66#_c_568_n
+ N_A_299_66#_M1004_g N_A_299_66#_c_646_p N_A_299_66#_c_569_n
+ N_A_299_66#_c_570_n N_A_299_66#_c_571_n N_A_299_66#_c_572_n
+ N_A_299_66#_c_573_n N_A_299_66#_c_574_n N_A_299_66#_c_575_n
+ N_A_299_66#_c_576_n N_A_299_66#_c_615_p N_A_299_66#_c_582_n
+ N_A_299_66#_c_577_n PM_SKY130_FD_SC_HD__SDFRTP_4%A_299_66#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%D N_D_M1026_g N_D_M1018_g D D N_D_c_710_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%D
x_PM_SKY130_FD_SC_HD__SDFRTP_4%SCE N_SCE_M1025_g N_SCE_c_751_n N_SCE_c_752_n
+ N_SCE_c_756_n N_SCE_M1006_g N_SCE_c_758_n N_SCE_M1003_g N_SCE_c_753_n
+ N_SCE_M1017_g N_SCE_c_760_n N_SCE_c_761_n SCE SCE N_SCE_c_754_n N_SCE_c_755_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%SCE
x_PM_SKY130_FD_SC_HD__SDFRTP_4%SCD N_SCD_M1035_g N_SCD_M1030_g SCD N_SCD_c_851_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%SCD
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_193_47# N_A_193_47#_M1022_d N_A_193_47#_M1041_d
+ N_A_193_47#_M1007_g N_A_193_47#_M1020_g N_A_193_47#_c_893_n
+ N_A_193_47#_M1014_g N_A_193_47#_M1031_g N_A_193_47#_c_924_n
+ N_A_193_47#_c_894_n N_A_193_47#_c_895_n N_A_193_47#_c_896_n
+ N_A_193_47#_c_897_n N_A_193_47#_c_898_n N_A_193_47#_c_899_n
+ N_A_193_47#_c_907_n N_A_193_47#_c_908_n N_A_193_47#_c_900_n
+ N_A_193_47#_c_909_n N_A_193_47#_c_910_n N_A_193_47#_c_911_n
+ N_A_193_47#_c_912_n N_A_193_47#_c_913_n N_A_193_47#_c_914_n
+ N_A_193_47#_c_915_n N_A_193_47#_c_916_n N_A_193_47#_c_917_n
+ N_A_193_47#_c_918_n N_A_193_47#_c_901_n N_A_193_47#_c_919_n
+ N_A_193_47#_c_902_n PM_SKY130_FD_SC_HD__SDFRTP_4%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_1245_303# N_A_1245_303#_M1039_d
+ N_A_1245_303#_M1021_d N_A_1245_303#_M1038_g N_A_1245_303#_M1010_g
+ N_A_1245_303#_c_1167_n N_A_1245_303#_c_1168_n N_A_1245_303#_c_1193_n
+ N_A_1245_303#_c_1169_n N_A_1245_303#_c_1170_n N_A_1245_303#_c_1214_p
+ N_A_1245_303#_c_1181_n N_A_1245_303#_c_1171_n N_A_1245_303#_c_1164_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%A_1245_303#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%RESET_B N_RESET_B_M1013_g N_RESET_B_M1033_g
+ N_RESET_B_c_1276_n N_RESET_B_c_1290_n N_RESET_B_M1000_g N_RESET_B_c_1291_n
+ N_RESET_B_M1012_g N_RESET_B_c_1292_n RESET_B RESET_B N_RESET_B_c_1280_n
+ N_RESET_B_c_1281_n N_RESET_B_c_1282_n N_RESET_B_c_1283_n N_RESET_B_c_1284_n
+ N_RESET_B_c_1285_n N_RESET_B_c_1286_n N_RESET_B_c_1287_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%RESET_B
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_1079_413# N_A_1079_413#_M1023_d
+ N_A_1079_413#_M1007_d N_A_1079_413#_M1039_g N_A_1079_413#_c_1451_n
+ N_A_1079_413#_c_1452_n N_A_1079_413#_M1021_g N_A_1079_413#_c_1479_n
+ N_A_1079_413#_c_1445_n N_A_1079_413#_c_1446_n N_A_1079_413#_c_1447_n
+ N_A_1079_413#_c_1448_n N_A_1079_413#_c_1467_n N_A_1079_413#_c_1455_n
+ N_A_1079_413#_c_1456_n N_A_1079_413#_c_1449_n N_A_1079_413#_c_1450_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%A_1079_413#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_1767_21# N_A_1767_21#_M1015_d
+ N_A_1767_21#_M1012_d N_A_1767_21#_M1027_g N_A_1767_21#_M1028_g
+ N_A_1767_21#_c_1585_n N_A_1767_21#_M1016_g N_A_1767_21#_M1002_g
+ N_A_1767_21#_c_1586_n N_A_1767_21#_M1019_g N_A_1767_21#_M1008_g
+ N_A_1767_21#_c_1587_n N_A_1767_21#_M1037_g N_A_1767_21#_M1024_g
+ N_A_1767_21#_c_1588_n N_A_1767_21#_M1040_g N_A_1767_21#_M1034_g
+ N_A_1767_21#_c_1589_n N_A_1767_21#_c_1590_n N_A_1767_21#_c_1591_n
+ N_A_1767_21#_c_1592_n N_A_1767_21#_c_1593_n N_A_1767_21#_c_1643_n
+ N_A_1767_21#_c_1702_p N_A_1767_21#_c_1604_n N_A_1767_21#_c_1605_n
+ N_A_1767_21#_c_1594_n N_A_1767_21#_c_1606_n N_A_1767_21#_c_1595_n
+ N_A_1767_21#_c_1596_n N_A_1767_21#_c_1597_n N_A_1767_21#_c_1598_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%A_1767_21#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_1592_47# N_A_1592_47#_M1014_d
+ N_A_1592_47#_M1001_d N_A_1592_47#_c_1773_n N_A_1592_47#_M1015_g
+ N_A_1592_47#_c_1776_n N_A_1592_47#_M1032_g N_A_1592_47#_c_1774_n
+ N_A_1592_47#_c_1783_n N_A_1592_47#_c_1779_n N_A_1592_47#_c_1775_n
+ N_A_1592_47#_c_1780_n N_A_1592_47#_c_1781_n N_A_1592_47#_c_1782_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%A_1592_47#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%VPWR N_VPWR_M1029_d N_VPWR_M1006_d N_VPWR_M1035_d
+ N_VPWR_M1038_d N_VPWR_M1021_s N_VPWR_M1028_d N_VPWR_M1032_d N_VPWR_M1002_d
+ N_VPWR_M1008_d N_VPWR_M1034_d N_VPWR_c_1892_n N_VPWR_c_1893_n N_VPWR_c_1894_n
+ N_VPWR_c_1895_n N_VPWR_c_1896_n N_VPWR_c_1897_n N_VPWR_c_1898_n
+ N_VPWR_c_1899_n N_VPWR_c_1900_n N_VPWR_c_1901_n N_VPWR_c_1902_n
+ N_VPWR_c_1903_n N_VPWR_c_1904_n N_VPWR_c_1905_n N_VPWR_c_1906_n VPWR
+ N_VPWR_c_1907_n N_VPWR_c_1908_n N_VPWR_c_1909_n N_VPWR_c_1910_n
+ N_VPWR_c_1911_n N_VPWR_c_1912_n N_VPWR_c_1913_n N_VPWR_c_1914_n
+ N_VPWR_c_1915_n N_VPWR_c_1916_n N_VPWR_c_1917_n N_VPWR_c_1918_n
+ N_VPWR_c_1919_n N_VPWR_c_1920_n N_VPWR_c_1891_n VPWR
+ PM_SKY130_FD_SC_HD__SDFRTP_4%VPWR
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_620_389# N_A_620_389#_M1018_d
+ N_A_620_389#_M1023_s N_A_620_389#_M1026_d N_A_620_389#_M1007_s
+ N_A_620_389#_c_2129_n N_A_620_389#_c_2098_n N_A_620_389#_c_2133_n
+ N_A_620_389#_c_2106_n N_A_620_389#_c_2107_n N_A_620_389#_c_2099_n
+ N_A_620_389#_c_2100_n N_A_620_389#_c_2101_n N_A_620_389#_c_2102_n
+ N_A_620_389#_c_2103_n N_A_620_389#_c_2104_n
+ PM_SKY130_FD_SC_HD__SDFRTP_4%A_620_389#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%A_1191_413# N_A_1191_413#_M1005_d
+ N_A_1191_413#_M1033_d N_A_1191_413#_c_2203_n N_A_1191_413#_c_2204_n
+ N_A_1191_413#_c_2205_n PM_SKY130_FD_SC_HD__SDFRTP_4%A_1191_413#
x_PM_SKY130_FD_SC_HD__SDFRTP_4%Q N_Q_M1016_s N_Q_M1037_s N_Q_M1002_s N_Q_M1024_s
+ N_Q_c_2236_n N_Q_c_2243_n N_Q_c_2237_n N_Q_c_2238_n N_Q_c_2248_n N_Q_c_2250_n
+ Q Q Q Q N_Q_c_2239_n Q PM_SKY130_FD_SC_HD__SDFRTP_4%Q
x_PM_SKY130_FD_SC_HD__SDFRTP_4%VGND N_VGND_M1036_d N_VGND_M1025_d N_VGND_M1009_s
+ N_VGND_M1030_d N_VGND_M1013_d N_VGND_M1027_d N_VGND_M1016_d N_VGND_M1019_d
+ N_VGND_M1040_d N_VGND_c_2277_n N_VGND_c_2278_n N_VGND_c_2279_n N_VGND_c_2280_n
+ N_VGND_c_2281_n N_VGND_c_2282_n N_VGND_c_2283_n N_VGND_c_2284_n
+ N_VGND_c_2285_n N_VGND_c_2286_n N_VGND_c_2287_n N_VGND_c_2288_n
+ N_VGND_c_2289_n N_VGND_c_2290_n N_VGND_c_2291_n N_VGND_c_2292_n
+ N_VGND_c_2293_n N_VGND_c_2294_n N_VGND_c_2295_n N_VGND_c_2296_n VGND
+ N_VGND_c_2297_n N_VGND_c_2298_n N_VGND_c_2299_n N_VGND_c_2300_n
+ N_VGND_c_2301_n N_VGND_c_2302_n N_VGND_c_2303_n N_VGND_c_2304_n
+ N_VGND_c_2305_n VGND PM_SKY130_FD_SC_HD__SDFRTP_4%VGND
cc_1 VNB N_CLK_c_273_n 0.0205109f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.98
cc_2 VNB CLK 0.00313032f $X=-0.19 $Y=-0.24 $X2=0.2 $Y2=1.105
cc_3 VNB N_CLK_c_275_n 0.0452947f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.162
cc_4 VNB N_A_27_47#_c_304_n 0.0186136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_c_305_n 0.0222058f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_6 VNB N_A_27_47#_c_306_n 0.0181117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_307_n 0.039334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1011_g 0.0291916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_309_n 0.0255512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_310_n 0.011157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_311_n 0.00784715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_312_n 0.0342871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_313_n 7.22032e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_314_n 0.0190351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_315_n 8.25118e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_316_n 0.00212824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_317_n 0.0233797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_318_n 0.00217752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_319_n 0.0194531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_320_n 0.0137739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_321_n 7.19339e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_322_n 9.50937e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_66#_c_567_n 0.0142002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_299_66#_c_568_n 0.0121103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_299_66#_c_569_n 0.00168045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_299_66#_c_570_n 0.00234188f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_27 VNB N_A_299_66#_c_571_n 0.0162157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_299_66#_c_572_n 7.10207e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_299_66#_c_573_n 0.00155275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_299_66#_c_574_n 0.00618254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_299_66#_c_575_n 0.00184774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_299_66#_c_576_n 0.0064465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_299_66#_c_577_n 0.049101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_D_M1018_g 0.0325237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB D 0.00255827f $X=-0.19 $Y=-0.24 $X2=0.2 $Y2=1.445
cc_36 VNB N_SCE_M1025_g 0.0316479f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.345
cc_37 VNB N_SCE_c_751_n 0.150126f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_38 VNB N_SCE_c_752_n 0.0127193f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_39 VNB N_SCE_c_753_n 0.0323957f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_40 VNB N_SCE_c_754_n 0.0250033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_SCE_c_755_n 0.00473389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_SCD_M1030_g 0.0529849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB SCD 0.00594926f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_44 VNB N_SCD_c_851_n 0.00548947f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_45 VNB N_A_193_47#_c_893_n 0.0180202f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_46 VNB N_A_193_47#_c_894_n 0.0103282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_895_n 0.00319457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_896_n 0.00491988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_193_47#_c_897_n 0.0289642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_193_47#_c_898_n 0.00511336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_193_47#_c_899_n 0.0368515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_193_47#_c_900_n 0.00474915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_193_47#_c_901_n 0.0181157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_193_47#_c_902_n 0.00375532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1245_303#_M1010_g 0.0437454f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_56 VNB N_A_1245_303#_c_1164_n 0.00620267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_M1033_g 0.00749317f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_58 VNB N_RESET_B_c_1276_n 0.0241938f $X=-0.19 $Y=-0.24 $X2=0.2 $Y2=1.105
cc_59 VNB N_RESET_B_M1000_g 0.0279211f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.162
cc_60 VNB RESET_B 0.00195157f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_61 VNB RESET_B 0.00264667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_RESET_B_c_1280_n 0.00409977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_RESET_B_c_1281_n 0.00761703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_c_1282_n 0.0164959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_RESET_B_c_1283_n 0.00128772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_1284_n 8.96978e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_RESET_B_c_1285_n 0.0290107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_RESET_B_c_1286_n 0.0169629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_RESET_B_c_1287_n 0.0013981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1079_413#_M1039_g 0.0191314f $X=-0.19 $Y=-0.24 $X2=0.2 $Y2=1.445
cc_71 VNB N_A_1079_413#_c_1445_n 0.00291989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1079_413#_c_1446_n 7.14483e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1079_413#_c_1447_n 0.00491059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1079_413#_c_1448_n 0.00293419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1079_413#_c_1449_n 0.00142696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1079_413#_c_1450_n 0.0279451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1767_21#_M1027_g 0.0214619f $X=-0.19 $Y=-0.24 $X2=0.2 $Y2=1.445
cc_78 VNB N_A_1767_21#_M1028_g 0.00966172f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_79 VNB N_A_1767_21#_c_1585_n 0.0197342f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.162
cc_80 VNB N_A_1767_21#_c_1586_n 0.0156266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1767_21#_c_1587_n 0.0160644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1767_21#_c_1588_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1767_21#_c_1589_n 0.00124594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1767_21#_c_1590_n 0.0051153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1767_21#_c_1591_n 0.00233676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1767_21#_c_1592_n 4.41081e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1767_21#_c_1593_n 0.00282287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1767_21#_c_1594_n 0.010488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1767_21#_c_1595_n 0.00846913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1767_21#_c_1596_n 0.00576234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1767_21#_c_1597_n 0.0463941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_1767_21#_c_1598_n 0.0886768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1592_47#_c_1773_n 0.0267637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1592_47#_c_1774_n 0.0244895f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.162
cc_95 VNB N_A_1592_47#_c_1775_n 0.00787141f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VPWR_c_1891_n 0.535415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_620_389#_c_2098_n 0.0053174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_620_389#_c_2099_n 0.00697414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_620_389#_c_2100_n 0.00522158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_620_389#_c_2101_n 0.00172242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_620_389#_c_2102_n 0.00327401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_A_620_389#_c_2103_n 0.00380619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_620_389#_c_2104_n 0.00207284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_Q_c_2236_n 0.00105631f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_105 VNB N_Q_c_2237_n 8.70049e-19 $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_106 VNB N_VGND_c_2277_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2278_n 0.00281411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2279_n 0.00480695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2280_n 0.00839765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2281_n 0.00774496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2282_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2283_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2284_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2285_n 0.00416502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2286_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2287_n 0.0415149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2288_n 0.00581387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2289_n 0.0462287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2290_n 0.00323844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2291_n 0.036703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2292_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2293_n 0.0191951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2294_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2295_n 0.0189691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2296_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2297_n 0.0147647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2298_n 0.0264169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2299_n 0.0566868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2300_n 0.0116899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2301_n 0.611668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2302_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2303_n 0.0043669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2304_n 0.00439458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2305_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VPB N_CLK_M1029_g 0.0220032f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_136 VPB CLK 0.00600609f $X=-0.19 $Y=1.305 $X2=0.2 $Y2=1.105
cc_137 VPB N_CLK_c_275_n 0.0122863f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.162
cc_138 VPB N_A_27_47#_M1041_g 0.0215501f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.162
cc_139 VPB N_A_27_47#_c_305_n 0.0240915f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_140 VPB N_A_27_47#_M1005_g 0.0473324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_307_n 0.0106083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_M1001_g 0.0448228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_328_n 9.37717e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_329_n 0.0273694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_315_n 0.00218623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_316_n 3.61249e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_317_n 0.00506712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_27_47#_c_319_n 0.0150989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_321_n 8.40813e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_299_66#_c_568_n 0.0218976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_299_66#_M1004_g 0.0269778f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.162
cc_152 VPB N_A_299_66#_c_571_n 0.00245276f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_299_66#_c_576_n 5.82055e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_299_66#_c_582_n 0.00522461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_299_66#_c_577_n 0.00388256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_D_M1026_g 0.020144f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_157 VPB N_D_M1018_g 0.00197249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB D 0.00603351f $X=-0.19 $Y=1.305 $X2=0.2 $Y2=1.445
cc_159 VPB D 0.00255959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_D_c_710_n 0.0353039f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_161 VPB N_SCE_c_756_n 0.0156381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_SCE_M1006_g 0.0224518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_SCE_c_758_n 0.0193512f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_164 VPB N_SCE_M1003_g 0.017331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_SCE_c_760_n 0.00590469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_SCE_c_761_n 0.00342234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB SCE 0.0107872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_SCE_c_754_n 0.0539173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_SCE_c_755_n 0.0044346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_SCD_M1035_g 0.027313f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_171 VPB N_SCD_M1030_g 0.00185092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB SCD 0.00352162f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_173 VPB N_SCD_c_851_n 0.025183f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_174 VPB N_A_193_47#_M1007_g 0.0257475f $X=-0.19 $Y=1.305 $X2=0.2 $Y2=1.445
cc_175 VPB N_A_193_47#_M1031_g 0.0184116f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.53
cc_176 VPB N_A_193_47#_c_894_n 0.00555562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_193_47#_c_898_n 0.00395561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_193_47#_c_907_n 0.00175719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_193_47#_c_908_n 7.52751e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_193_47#_c_909_n 0.00316594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_193_47#_c_910_n 0.00372313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_193_47#_c_911_n 0.030488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_193_47#_c_912_n 0.0328457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_193_47#_c_913_n 6.49743e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_193_47#_c_914_n 0.0124185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_193_47#_c_915_n 0.00250224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_193_47#_c_916_n 0.00151832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_193_47#_c_917_n 0.0321438f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_193_47#_c_918_n 0.00229435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_193_47#_c_919_n 0.0023012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_193_47#_c_902_n 0.00397602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1245_303#_M1038_g 0.0212174f $X=-0.19 $Y=1.305 $X2=0.2 $Y2=1.445
cc_193 VPB N_A_1245_303#_M1010_g 0.0114089f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_194 VPB N_A_1245_303#_c_1167_n 0.0127484f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.162
cc_195 VPB N_A_1245_303#_c_1168_n 0.0357454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1245_303#_c_1169_n 7.24024e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1245_303#_c_1170_n 5.38139e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1245_303#_c_1171_n 0.00414915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1245_303#_c_1164_n 0.00207203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_M1033_g 0.0583973f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_201 VPB N_RESET_B_c_1276_n 0.0172676f $X=-0.19 $Y=1.305 $X2=0.2 $Y2=1.105
cc_202 VPB N_RESET_B_c_1290_n 0.019935f $X=-0.19 $Y=1.305 $X2=0.2 $Y2=1.445
cc_203 VPB N_RESET_B_c_1291_n 0.0151236f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_204 VPB N_RESET_B_c_1292_n 0.0185949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_1284_n 9.23966e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1079_413#_c_1451_n 0.0275308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_1079_413#_c_1452_n 0.0165899f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_208 VPB N_A_1079_413#_c_1445_n 0.00279025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_1079_413#_c_1448_n 0.00495216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_1079_413#_c_1455_n 0.00460975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_A_1079_413#_c_1456_n 0.00144164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1079_413#_c_1449_n 0.00126247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_1079_413#_c_1450_n 0.0216746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_1767_21#_M1028_g 0.0431751f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_215 VPB N_A_1767_21#_M1002_g 0.0217167f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1767_21#_M1008_g 0.0179369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_1767_21#_M1024_g 0.0183405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1767_21#_M1034_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_1767_21#_c_1604_n 0.0099556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1767_21#_c_1605_n 0.00285193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1767_21#_c_1606_n 0.0134808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_1767_21#_c_1595_n 0.00730666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1767_21#_c_1596_n 3.43438e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1767_21#_c_1598_n 0.0157353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1592_47#_c_1776_n 0.0311824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1592_47#_M1032_g 0.0262666f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.162
cc_227 VPB N_A_1592_47#_c_1774_n 0.011759f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.162
cc_228 VPB N_A_1592_47#_c_1779_n 9.33226e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_1592_47#_c_1780_n 0.00458975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_1592_47#_c_1781_n 0.0117011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_1592_47#_c_1782_n 0.0188067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1892_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1893_n 0.00468754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1894_n 0.00531826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1895_n 0.00712128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1896_n 0.00222993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1897_n 0.00372502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1898_n 0.00810983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1899_n 0.00111115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1900_n 0.00167829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1901_n 0.0140014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1902_n 0.0431198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1903_n 0.0391891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1904_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1905_n 0.0104664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1906_n 0.0460908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1907_n 0.0149258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1908_n 0.0484444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1909_n 0.0176581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1910_n 0.0391861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1911_n 0.011983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1912_n 0.0161376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1913_n 0.0158909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1914_n 0.00436818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1915_n 0.00507043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1916_n 0.00596369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1917_n 0.00353358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1918_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1919_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1920_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1891_n 0.0667128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_A_620_389#_c_2098_n 0.0102954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_A_620_389#_c_2106_n 0.00572038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_A_620_389#_c_2107_n 0.0023107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_A_620_389#_c_2099_n 0.0261275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_A_1191_413#_c_2203_n 0.00288813f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_A_1191_413#_c_2204_n 0.00250365f $X=-0.19 $Y=1.305 $X2=0.2
+ $Y2=1.445
cc_268 VPB N_A_1191_413#_c_2205_n 0.00240785f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.16
cc_269 VPB N_Q_c_2238_n 0.00127173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_Q_c_2239_n 0.00216937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 CLK N_A_27_47#_M1029_s 0.00841523f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_272 N_CLK_c_273_n N_A_27_47#_c_304_n 0.0247689f $X=0.47 $Y=0.98 $X2=0 $Y2=0
cc_273 CLK N_A_27_47#_M1041_g 2.66895e-19 $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_274 N_CLK_c_275_n N_A_27_47#_M1041_g 0.0372159f $X=0.47 $Y=1.162 $X2=0 $Y2=0
cc_275 N_CLK_c_273_n N_A_27_47#_c_339_n 0.0131216f $X=0.47 $Y=0.98 $X2=0 $Y2=0
cc_276 CLK N_A_27_47#_c_339_n 0.00945024f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_277 CLK N_A_27_47#_c_311_n 0.017873f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_278 N_CLK_c_275_n N_A_27_47#_c_311_n 0.00296723f $X=0.47 $Y=1.162 $X2=0 $Y2=0
cc_279 N_CLK_M1029_g N_A_27_47#_c_343_n 0.0117673f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_280 CLK N_A_27_47#_c_343_n 0.00709933f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_281 N_CLK_M1029_g N_A_27_47#_c_328_n 0.00393855f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_282 CLK N_A_27_47#_c_329_n 0.0176831f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_283 N_CLK_c_275_n N_A_27_47#_c_329_n 0.0020001f $X=0.47 $Y=1.162 $X2=0 $Y2=0
cc_284 CLK N_A_27_47#_c_313_n 0.00134476f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_285 CLK N_A_27_47#_c_317_n 3.1348e-19 $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_286 N_CLK_c_275_n N_A_27_47#_c_317_n 0.0208917f $X=0.47 $Y=1.162 $X2=0 $Y2=0
cc_287 N_CLK_c_275_n N_A_27_47#_c_318_n 0.00393855f $X=0.47 $Y=1.162 $X2=0 $Y2=0
cc_288 N_CLK_c_273_n N_A_27_47#_c_322_n 0.00393855f $X=0.47 $Y=0.98 $X2=0 $Y2=0
cc_289 CLK N_A_27_47#_c_322_n 0.0489186f $X=0.2 $Y=1.105 $X2=0 $Y2=0
cc_290 N_CLK_M1029_g N_VPWR_c_1892_n 0.00967619f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_291 N_CLK_M1029_g N_VPWR_c_1907_n 0.00396867f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_292 N_CLK_M1029_g N_VPWR_c_1891_n 0.00559284f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_293 N_CLK_c_273_n N_VGND_c_2277_n 0.0112612f $X=0.47 $Y=0.98 $X2=0 $Y2=0
cc_294 N_CLK_c_273_n N_VGND_c_2297_n 0.00339367f $X=0.47 $Y=0.98 $X2=0 $Y2=0
cc_295 N_CLK_c_273_n N_VGND_c_2301_n 0.00497794f $X=0.47 $Y=0.98 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_312_n N_A_299_66#_c_568_n 9.69822e-19 $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_312_n N_A_299_66#_c_569_n 0.011877f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_312_n N_A_299_66#_c_570_n 0.0012622f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_312_n N_A_299_66#_c_571_n 0.0341518f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_312_n N_A_299_66#_c_572_n 0.0309775f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_312_n N_A_299_66#_c_576_n 0.0145537f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_312_n N_A_299_66#_c_577_n 0.00271841f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_312_n N_D_M1018_g 0.00938366f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_312_n D 0.00575784f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_312_n N_SCE_M1025_g 0.00205342f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_312_n N_SCE_c_756_n 9.34876e-19 $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_312_n N_SCE_c_758_n 0.00110755f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_312_n N_SCE_c_753_n 0.00595181f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_309 N_A_27_47#_M1041_g N_SCE_c_754_n 0.00755797f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_312_n N_SCE_c_754_n 0.00648239f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_317_n N_SCE_c_754_n 0.00624852f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_27_47#_M1041_g N_SCE_c_755_n 6.40276e-19 $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_312_n N_SCE_c_755_n 0.0185491f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_314 N_A_27_47#_c_309_n N_SCD_M1030_g 0.00617832f $X=5.36 $Y=0.745 $X2=0 $Y2=0
cc_315 N_A_27_47#_c_312_n N_SCD_M1030_g 0.00469801f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_319_n N_SCD_M1030_g 0.0108611f $X=4.99 $Y=1.23 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_312_n SCD 0.0360755f $X=4.845 $Y=1.19 $X2=0 $Y2=0
cc_318 N_A_27_47#_M1005_g N_A_193_47#_M1007_g 0.0144886f $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_M1011_g N_A_193_47#_c_893_n 0.0127282f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_M1001_g N_A_193_47#_M1031_g 0.0169629f $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_343_n N_A_193_47#_c_924_n 0.00331898f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_304_n N_A_193_47#_c_894_n 0.00601364f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1041_g N_A_193_47#_c_894_n 0.0036639f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_339_n N_A_193_47#_c_894_n 0.00642066f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_328_n N_A_193_47#_c_894_n 0.0198723f $X=0.762 $Y=1.795 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_312_n N_A_193_47#_c_894_n 0.0123974f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_313_n N_A_193_47#_c_894_n 0.00275409f $X=1.035 $Y=1.19 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_317_n N_A_193_47#_c_894_n 0.00425791f $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_318_n N_A_193_47#_c_894_n 0.0226057f $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_322_n N_A_193_47#_c_894_n 0.008551f $X=0.817 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_309_n N_A_193_47#_c_895_n 0.0085464f $X=5.36 $Y=0.745 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_320_n N_A_193_47#_c_895_n 0.00177637f $X=4.987 $Y=1.065
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_305_n N_A_193_47#_c_896_n 0.00585634f $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_314_n N_A_193_47#_c_896_n 0.0176558f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_305_n N_A_193_47#_c_897_n 0.017436f $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_309_n N_A_193_47#_c_897_n 0.00667405f $X=5.36 $Y=0.745 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_314_n N_A_193_47#_c_897_n 0.00371207f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_320_n N_A_193_47#_c_897_n 0.00201772f $X=4.987 $Y=1.065
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_307_n N_A_193_47#_c_898_n 0.00910115f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_M1011_g N_A_193_47#_c_898_n 0.00127125f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_314_n N_A_193_47#_c_898_n 0.015245f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_316_n N_A_193_47#_c_898_n 0.00237014f $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_321_n N_A_193_47#_c_898_n 0.0156117f $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_M1011_g N_A_193_47#_c_899_n 0.0214166f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_314_n N_A_193_47#_c_899_n 0.00135733f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_321_n N_A_193_47#_c_899_n 3.86059e-19 $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_M1001_g N_A_193_47#_c_907_n 0.00731313f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_314_n N_A_193_47#_c_907_n 0.00562532f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_312_n N_A_193_47#_c_900_n 0.00454244f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_313_n N_A_193_47#_c_900_n 7.77055e-19 $X=1.035 $Y=1.19 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_317_n N_A_193_47#_c_900_n 2.24002e-19 $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_307_n N_A_193_47#_c_909_n 0.00514409f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_M1001_g N_A_193_47#_c_909_n 0.0107407f $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_314_n N_A_193_47#_c_909_n 9.49173e-19 $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_316_n N_A_193_47#_c_909_n 0.0025355f $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_321_n N_A_193_47#_c_909_n 0.00818233f $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_307_n N_A_193_47#_c_910_n 5.3506e-19 $X=8.285 $Y=1.395 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1001_g N_A_193_47#_c_910_n 2.52071e-19 $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_316_n N_A_193_47#_c_910_n 0.00168571f $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_321_n N_A_193_47#_c_910_n 0.00197607f $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_307_n N_A_193_47#_c_911_n 0.00262948f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_M1001_g N_A_193_47#_c_911_n 0.0209818f $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_316_n N_A_193_47#_c_911_n 4.59576e-19 $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_312_n N_A_193_47#_c_912_n 0.157967f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_314_n N_A_193_47#_c_912_n 0.00587882f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_424_p N_A_193_47#_c_912_n 0.014344f $X=5.135 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_315_n N_A_193_47#_c_912_n 0.0016551f $X=4.99 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_319_n N_A_193_47#_c_912_n 0.0025783f $X=4.99 $Y=1.23 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_M1041_g N_A_193_47#_c_913_n 0.00240409f $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_343_n N_A_193_47#_c_913_n 0.0053366f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_328_n N_A_193_47#_c_913_n 0.00106255f $X=0.762 $Y=1.795
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_312_n N_A_193_47#_c_913_n 0.0104885f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_313_n N_A_193_47#_c_913_n 0.00362442f $X=1.035 $Y=1.19 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_317_n N_A_193_47#_c_913_n 6.43629e-19 $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_305_n N_A_193_47#_c_914_n 0.00132845f $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_M1005_g N_A_193_47#_c_914_n 0.00420966f $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_M1001_g N_A_193_47#_c_914_n 0.00356005f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_314_n N_A_193_47#_c_914_n 0.118928f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_316_n N_A_193_47#_c_914_n 0.00182236f $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_305_n N_A_193_47#_c_915_n 7.57971e-19 $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_314_n N_A_193_47#_c_915_n 0.0130648f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_M1001_g N_A_193_47#_c_916_n 5.0827e-19 $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_316_n N_A_193_47#_c_916_n 0.0121474f $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_321_n N_A_193_47#_c_916_n 5.23442e-19 $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_305_n N_A_193_47#_c_917_n 0.0211058f $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_M1005_g N_A_193_47#_c_917_n 0.0107367f $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_314_n N_A_193_47#_c_917_n 2.03081e-19 $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_305_n N_A_193_47#_c_918_n 0.00183386f $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1005_g N_A_193_47#_c_918_n 4.97407e-19 $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_314_n N_A_193_47#_c_918_n 0.00222352f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_306_n N_A_193_47#_c_901_n 0.0155794f $X=5.36 $Y=0.67 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_M1041_g N_A_193_47#_c_919_n 4.23008e-19 $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_343_n N_A_193_47#_c_919_n 0.00537623f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_328_n N_A_193_47#_c_919_n 0.00264365f $X=0.762 $Y=1.795
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_312_n N_A_193_47#_c_919_n 0.0024738f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_305_n N_A_193_47#_c_902_n 0.011349f $X=5.805 $Y=1.32 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_M1005_g N_A_193_47#_c_902_n 0.00106158f $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_314_n N_A_193_47#_c_902_n 0.0173608f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_424_p N_A_193_47#_c_902_n 0.00224837f $X=5.135 $Y=1.19 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_315_n N_A_193_47#_c_902_n 0.0148592f $X=4.99 $Y=1.19 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_320_n N_A_193_47#_c_902_n 0.00251608f $X=4.987 $Y=1.065
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_305_n N_A_1245_303#_M1010_g 0.00915737f $X=5.805 $Y=1.32
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_314_n N_A_1245_303#_M1010_g 0.00542236f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_M1005_g N_A_1245_303#_c_1167_n 5.40696e-19 $X=5.88 $Y=2.275
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_314_n N_A_1245_303#_c_1167_n 0.00564111f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_M1005_g N_A_1245_303#_c_1168_n 0.0362882f $X=5.88 $Y=2.275
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_M1001_g N_A_1245_303#_c_1169_n 0.00223454f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_314_n N_A_1245_303#_c_1169_n 0.00195818f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_M1001_g N_A_1245_303#_c_1170_n 0.00375824f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_314_n N_A_1245_303#_c_1181_n 7.74909e-19 $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_314_n N_A_1245_303#_c_1171_n 0.00256862f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_M1011_g N_A_1245_303#_c_1164_n 3.73683e-19 $X=8.43 $Y=0.415
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_314_n N_A_1245_303#_c_1164_n 0.0127435f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_314_n N_RESET_B_M1033_g 0.00108426f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_314_n N_RESET_B_c_1280_n 0.0592788f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_314_n N_RESET_B_c_1281_n 0.00341238f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_307_n N_RESET_B_c_1282_n 0.00154439f $X=8.285 $Y=1.395 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_M1011_g N_RESET_B_c_1282_n 0.00447717f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_314_n N_RESET_B_c_1282_n 0.0993427f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_316_n N_RESET_B_c_1282_n 0.0260309f $X=8.49 $Y=1.19 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_321_n N_RESET_B_c_1282_n 0.0021678f $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_314_n N_RESET_B_c_1285_n 0.00270235f $X=8.345 $Y=1.19 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_M1001_g N_A_1079_413#_c_1451_n 0.0294293f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_314_n N_A_1079_413#_c_1451_n 0.00337185f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_305_n N_A_1079_413#_c_1445_n 0.00649941f $X=5.805 $Y=1.32
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_314_n N_A_1079_413#_c_1445_n 0.0131951f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_305_n N_A_1079_413#_c_1446_n 0.00451192f $X=5.805 $Y=1.32
+ $X2=0 $Y2=0
cc_428 N_A_27_47#_c_314_n N_A_1079_413#_c_1446_n 0.00696389f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_314_n N_A_1079_413#_c_1447_n 0.0156737f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_314_n N_A_1079_413#_c_1448_n 0.0268857f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_M1005_g N_A_1079_413#_c_1467_n 0.00440345f $X=5.88 $Y=2.275
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_305_n N_A_1079_413#_c_1455_n 0.00373226f $X=5.805 $Y=1.32
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_M1005_g N_A_1079_413#_c_1455_n 0.0202605f $X=5.88 $Y=2.275
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_314_n N_A_1079_413#_c_1456_n 0.00403101f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_314_n N_A_1079_413#_c_1449_n 0.0110043f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_314_n N_A_1079_413#_c_1450_n 0.00486738f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_M1011_g N_A_1767_21#_M1027_g 0.0308892f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_307_n N_A_1767_21#_M1028_g 0.00168082f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_M1001_g N_A_1767_21#_M1028_g 0.00181718f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_307_n N_A_1767_21#_c_1597_n 0.00868768f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_307_n N_A_1592_47#_c_1783_n 0.00225842f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_M1011_g N_A_1592_47#_c_1783_n 0.0118273f $X=8.43 $Y=0.415
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_321_n N_A_1592_47#_c_1783_n 0.00348965f $X=8.49 $Y=1.11
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_M1001_g N_A_1592_47#_c_1779_n 0.0049222f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_307_n N_A_1592_47#_c_1775_n 0.00260839f $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_M1011_g N_A_1592_47#_c_1775_n 0.00507754f $X=8.43 $Y=0.415
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_c_316_n N_A_1592_47#_c_1775_n 0.00772758f $X=8.49 $Y=1.19
+ $X2=0 $Y2=0
cc_448 N_A_27_47#_c_321_n N_A_1592_47#_c_1775_n 0.0262865f $X=8.49 $Y=1.11 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_307_n N_A_1592_47#_c_1781_n 9.24049e-19 $X=8.285 $Y=1.395
+ $X2=0 $Y2=0
cc_450 N_A_27_47#_M1001_g N_A_1592_47#_c_1781_n 0.00136255f $X=8.285 $Y=2.275
+ $X2=0 $Y2=0
cc_451 N_A_27_47#_c_321_n N_A_1592_47#_c_1781_n 8.18571e-19 $X=8.49 $Y=1.11
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_343_n N_VPWR_M1029_d 0.0039818f $X=0.66 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_453 N_A_27_47#_c_328_n N_VPWR_M1029_d 0.0031014f $X=0.762 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_454 N_A_27_47#_M1041_g N_VPWR_c_1892_n 0.0105939f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_343_n N_VPWR_c_1892_n 0.017664f $X=0.66 $Y=1.88 $X2=0 $Y2=0
cc_456 N_A_27_47#_M1001_g N_VPWR_c_1895_n 0.00108063f $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_M1041_g N_VPWR_c_1903_n 0.004627f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_M1005_g N_VPWR_c_1906_n 0.00541359f $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_343_n N_VPWR_c_1907_n 0.00204297f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_329_n N_VPWR_c_1907_n 0.0176235f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_461 N_A_27_47#_M1001_g N_VPWR_c_1910_n 0.00524716f $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_M1029_s N_VPWR_c_1891_n 0.00235071f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_M1041_g N_VPWR_c_1891_n 0.00876257f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_M1005_g N_VPWR_c_1891_n 0.00652322f $X=5.88 $Y=2.275 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_M1001_g N_VPWR_c_1891_n 0.00619371f $X=8.285 $Y=2.275 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_343_n N_VPWR_c_1891_n 0.00549713f $X=0.66 $Y=1.88 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_329_n N_VPWR_c_1891_n 0.00973967f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_312_n N_A_620_389#_c_2098_n 0.00959282f $X=4.845 $Y=1.19
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_312_n N_A_620_389#_c_2099_n 0.0134468f $X=4.845 $Y=1.19
+ $X2=0 $Y2=0
cc_470 N_A_27_47#_c_424_p N_A_620_389#_c_2099_n 0.00240264f $X=5.135 $Y=1.19
+ $X2=0 $Y2=0
cc_471 N_A_27_47#_c_315_n N_A_620_389#_c_2099_n 0.0252651f $X=4.99 $Y=1.19 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_319_n N_A_620_389#_c_2099_n 0.00498508f $X=4.99 $Y=1.23
+ $X2=0 $Y2=0
cc_473 N_A_27_47#_c_320_n N_A_620_389#_c_2099_n 0.00176883f $X=4.987 $Y=1.065
+ $X2=0 $Y2=0
cc_474 N_A_27_47#_c_309_n N_A_620_389#_c_2100_n 0.00470436f $X=5.36 $Y=0.745
+ $X2=0 $Y2=0
cc_475 N_A_27_47#_c_312_n N_A_620_389#_c_2100_n 0.00466124f $X=4.845 $Y=1.19
+ $X2=0 $Y2=0
cc_476 N_A_27_47#_c_314_n N_A_620_389#_c_2100_n 3.78682e-19 $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_477 N_A_27_47#_c_424_p N_A_620_389#_c_2100_n 0.00657764f $X=5.135 $Y=1.19
+ $X2=0 $Y2=0
cc_478 N_A_27_47#_c_315_n N_A_620_389#_c_2100_n 0.0116936f $X=4.99 $Y=1.19 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_319_n N_A_620_389#_c_2100_n 0.00350952f $X=4.99 $Y=1.23
+ $X2=0 $Y2=0
cc_480 N_A_27_47#_c_320_n N_A_620_389#_c_2100_n 0.00553901f $X=4.987 $Y=1.065
+ $X2=0 $Y2=0
cc_481 N_A_27_47#_c_306_n N_A_620_389#_c_2102_n 0.00424722f $X=5.36 $Y=0.67
+ $X2=0 $Y2=0
cc_482 N_A_27_47#_c_309_n N_A_620_389#_c_2102_n 0.00434493f $X=5.36 $Y=0.745
+ $X2=0 $Y2=0
cc_483 N_A_27_47#_c_312_n N_A_620_389#_c_2103_n 0.0133431f $X=4.845 $Y=1.19
+ $X2=0 $Y2=0
cc_484 N_A_27_47#_c_306_n N_A_620_389#_c_2104_n 0.00305101f $X=5.36 $Y=0.67
+ $X2=0 $Y2=0
cc_485 N_A_27_47#_c_309_n N_A_620_389#_c_2104_n 0.00459285f $X=5.36 $Y=0.745
+ $X2=0 $Y2=0
cc_486 N_A_27_47#_c_314_n N_A_620_389#_c_2104_n 0.00497164f $X=8.345 $Y=1.19
+ $X2=0 $Y2=0
cc_487 N_A_27_47#_M1005_g N_A_1191_413#_c_2204_n 8.92742e-19 $X=5.88 $Y=2.275
+ $X2=0 $Y2=0
cc_488 N_A_27_47#_c_339_n N_VGND_M1036_d 0.00380105f $X=0.66 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_489 N_A_27_47#_c_322_n N_VGND_M1036_d 8.90628e-19 $X=0.817 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_490 N_A_27_47#_c_304_n N_VGND_c_2277_n 0.011399f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_491 N_A_27_47#_c_339_n N_VGND_c_2277_n 0.0161609f $X=0.66 $Y=0.72 $X2=0 $Y2=0
cc_492 N_A_27_47#_c_313_n N_VGND_c_2277_n 3.6463e-19 $X=1.035 $Y=1.19 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_c_318_n N_VGND_c_2277_n 2.40105e-19 $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_312_n N_VGND_c_2278_n 5.94768e-19 $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_312_n N_VGND_c_2280_n 0.00208311f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_c_306_n N_VGND_c_2281_n 0.00341757f $X=5.36 $Y=0.67 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_312_n N_VGND_c_2281_n 0.0047368f $X=4.845 $Y=1.19 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_M1011_g N_VGND_c_2289_n 0.00357877f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_310_n N_VGND_c_2297_n 0.0106361f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_500 N_A_27_47#_c_339_n N_VGND_c_2297_n 0.00243651f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_c_304_n N_VGND_c_2298_n 0.0046653f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_c_306_n N_VGND_c_2299_n 0.0043254f $X=5.36 $Y=0.67 $X2=0 $Y2=0
cc_503 N_A_27_47#_M1036_s N_VGND_c_2301_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_c_304_n N_VGND_c_2301_n 0.00934473f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_c_306_n N_VGND_c_2301_n 0.00772301f $X=5.36 $Y=0.67 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_M1011_g N_VGND_c_2301_n 0.00565064f $X=8.43 $Y=0.415 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_310_n N_VGND_c_2301_n 0.00898615f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_339_n N_VGND_c_2301_n 0.00573594f $X=0.66 $Y=0.72 $X2=0
+ $Y2=0
cc_509 N_A_299_66#_M1004_g N_D_M1026_g 0.0104028f $X=3.825 $Y=2.215 $X2=0 $Y2=0
cc_510 N_A_299_66#_c_567_n N_D_M1018_g 0.0469999f $X=2.77 $Y=1.09 $X2=0 $Y2=0
cc_511 N_A_299_66#_c_568_n N_D_M1018_g 0.00693268f $X=3.825 $Y=1.685 $X2=0 $Y2=0
cc_512 N_A_299_66#_c_571_n N_D_M1018_g 0.00103624f $X=2.065 $Y=1.455 $X2=0 $Y2=0
cc_513 N_A_299_66#_c_572_n N_D_M1018_g 0.00378496f $X=2.915 $Y=1.09 $X2=0 $Y2=0
cc_514 N_A_299_66#_c_573_n N_D_M1018_g 0.0106539f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A_299_66#_c_574_n N_D_M1018_g 0.00295426f $X=3.68 $Y=0.34 $X2=0 $Y2=0
cc_516 N_A_299_66#_c_576_n N_D_M1018_g 7.55629e-19 $X=3.765 $Y=1.52 $X2=0 $Y2=0
cc_517 N_A_299_66#_c_577_n N_D_M1018_g 0.00427001f $X=2.385 $Y=1.29 $X2=0 $Y2=0
cc_518 N_A_299_66#_c_571_n D 0.00607625f $X=2.065 $Y=1.455 $X2=0 $Y2=0
cc_519 N_A_299_66#_c_572_n D 0.0246613f $X=2.915 $Y=1.09 $X2=0 $Y2=0
cc_520 N_A_299_66#_c_582_n D 0.0106084f $X=2.025 $Y=2.055 $X2=0 $Y2=0
cc_521 N_A_299_66#_c_577_n D 0.00301285f $X=2.385 $Y=1.29 $X2=0 $Y2=0
cc_522 N_A_299_66#_M1004_g N_D_c_710_n 0.00139776f $X=3.825 $Y=2.215 $X2=0 $Y2=0
cc_523 N_A_299_66#_c_572_n N_D_c_710_n 7.98046e-19 $X=2.915 $Y=1.09 $X2=0 $Y2=0
cc_524 N_A_299_66#_c_569_n N_SCE_M1025_g 0.014468f $X=2.055 $Y=0.815 $X2=0 $Y2=0
cc_525 N_A_299_66#_c_571_n N_SCE_M1025_g 0.00824697f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_526 N_A_299_66#_c_577_n N_SCE_M1025_g 0.0131f $X=2.385 $Y=1.29 $X2=0 $Y2=0
cc_527 N_A_299_66#_c_567_n N_SCE_c_751_n 0.0102879f $X=2.77 $Y=1.09 $X2=0 $Y2=0
cc_528 N_A_299_66#_c_569_n N_SCE_c_751_n 2.18848e-19 $X=2.055 $Y=0.815 $X2=0
+ $Y2=0
cc_529 N_A_299_66#_c_571_n N_SCE_c_751_n 0.001008f $X=2.065 $Y=1.455 $X2=0 $Y2=0
cc_530 N_A_299_66#_c_574_n N_SCE_c_751_n 0.00907768f $X=3.68 $Y=0.34 $X2=0 $Y2=0
cc_531 N_A_299_66#_c_575_n N_SCE_c_751_n 0.00370167f $X=3.085 $Y=0.34 $X2=0
+ $Y2=0
cc_532 N_A_299_66#_c_582_n N_SCE_c_756_n 0.0107883f $X=2.025 $Y=2.055 $X2=0
+ $Y2=0
cc_533 N_A_299_66#_c_615_p N_SCE_M1006_g 0.00391871f $X=1.985 $Y=2.22 $X2=0
+ $Y2=0
cc_534 N_A_299_66#_c_582_n N_SCE_M1006_g 0.0092899f $X=2.025 $Y=2.055 $X2=0
+ $Y2=0
cc_535 N_A_299_66#_c_572_n N_SCE_c_758_n 0.0019199f $X=2.915 $Y=1.09 $X2=0 $Y2=0
cc_536 N_A_299_66#_c_577_n N_SCE_c_758_n 0.00467364f $X=2.385 $Y=1.29 $X2=0
+ $Y2=0
cc_537 N_A_299_66#_c_582_n N_SCE_M1003_g 0.00170639f $X=2.025 $Y=2.055 $X2=0
+ $Y2=0
cc_538 N_A_299_66#_c_568_n N_SCE_c_753_n 0.00690009f $X=3.825 $Y=1.685 $X2=0
+ $Y2=0
cc_539 N_A_299_66#_c_573_n N_SCE_c_753_n 0.00163225f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_540 N_A_299_66#_c_574_n N_SCE_c_753_n 0.0153222f $X=3.68 $Y=0.34 $X2=0 $Y2=0
cc_541 N_A_299_66#_c_576_n N_SCE_c_753_n 0.0218997f $X=3.765 $Y=1.52 $X2=0 $Y2=0
cc_542 N_A_299_66#_c_571_n N_SCE_c_760_n 0.00752585f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_543 N_A_299_66#_c_582_n N_SCE_c_760_n 0.00484133f $X=2.025 $Y=2.055 $X2=0
+ $Y2=0
cc_544 N_A_299_66#_c_577_n N_SCE_c_760_n 0.021719f $X=2.385 $Y=1.29 $X2=0 $Y2=0
cc_545 N_A_299_66#_c_615_p N_SCE_c_761_n 0.0271281f $X=1.985 $Y=2.22 $X2=0 $Y2=0
cc_546 N_A_299_66#_c_569_n N_SCE_c_754_n 9.17465e-19 $X=2.055 $Y=0.815 $X2=0
+ $Y2=0
cc_547 N_A_299_66#_c_570_n N_SCE_c_754_n 0.00106256f $X=1.705 $Y=0.815 $X2=0
+ $Y2=0
cc_548 N_A_299_66#_c_571_n N_SCE_c_754_n 0.00265701f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_549 N_A_299_66#_c_615_p N_SCE_c_754_n 0.00266324f $X=1.985 $Y=2.22 $X2=0
+ $Y2=0
cc_550 N_A_299_66#_c_582_n N_SCE_c_754_n 0.00244193f $X=2.025 $Y=2.055 $X2=0
+ $Y2=0
cc_551 N_A_299_66#_c_569_n N_SCE_c_755_n 0.001843f $X=2.055 $Y=0.815 $X2=0 $Y2=0
cc_552 N_A_299_66#_c_570_n N_SCE_c_755_n 0.0143131f $X=1.705 $Y=0.815 $X2=0
+ $Y2=0
cc_553 N_A_299_66#_c_571_n N_SCE_c_755_n 0.0194368f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_554 N_A_299_66#_c_582_n N_SCE_c_755_n 0.0318889f $X=2.025 $Y=2.055 $X2=0
+ $Y2=0
cc_555 N_A_299_66#_c_577_n N_SCE_c_755_n 2.71658e-19 $X=2.385 $Y=1.29 $X2=0
+ $Y2=0
cc_556 N_A_299_66#_M1004_g N_SCD_M1035_g 0.0425828f $X=3.825 $Y=2.215 $X2=0
+ $Y2=0
cc_557 N_A_299_66#_c_568_n N_SCD_M1030_g 7.58826e-19 $X=3.825 $Y=1.685 $X2=0
+ $Y2=0
cc_558 N_A_299_66#_c_576_n N_SCD_M1030_g 0.00184558f $X=3.765 $Y=1.52 $X2=0
+ $Y2=0
cc_559 N_A_299_66#_c_568_n SCD 0.00265449f $X=3.825 $Y=1.685 $X2=0 $Y2=0
cc_560 N_A_299_66#_c_574_n SCD 0.010971f $X=3.68 $Y=0.34 $X2=0 $Y2=0
cc_561 N_A_299_66#_c_576_n SCD 0.0940519f $X=3.765 $Y=1.52 $X2=0 $Y2=0
cc_562 N_A_299_66#_c_568_n N_SCD_c_851_n 0.0141755f $X=3.825 $Y=1.685 $X2=0
+ $Y2=0
cc_563 N_A_299_66#_c_576_n N_SCD_c_851_n 2.87168e-19 $X=3.765 $Y=1.52 $X2=0
+ $Y2=0
cc_564 N_A_299_66#_c_646_p N_A_193_47#_c_894_n 0.00334973f $X=1.62 $Y=0.56 $X2=0
+ $Y2=0
cc_565 N_A_299_66#_c_570_n N_A_193_47#_c_894_n 0.0119534f $X=1.705 $Y=0.815
+ $X2=0 $Y2=0
cc_566 N_A_299_66#_c_646_p N_A_193_47#_c_900_n 0.0180018f $X=1.62 $Y=0.56 $X2=0
+ $Y2=0
cc_567 N_A_299_66#_c_568_n N_A_193_47#_c_912_n 9.25275e-19 $X=3.825 $Y=1.685
+ $X2=0 $Y2=0
cc_568 N_A_299_66#_M1004_g N_A_193_47#_c_912_n 0.00401957f $X=3.825 $Y=2.215
+ $X2=0 $Y2=0
cc_569 N_A_299_66#_c_571_n N_A_193_47#_c_912_n 0.00704301f $X=2.065 $Y=1.455
+ $X2=0 $Y2=0
cc_570 N_A_299_66#_c_572_n N_A_193_47#_c_912_n 0.00296925f $X=2.915 $Y=1.09
+ $X2=0 $Y2=0
cc_571 N_A_299_66#_c_576_n N_A_193_47#_c_912_n 0.00218994f $X=3.765 $Y=1.52
+ $X2=0 $Y2=0
cc_572 N_A_299_66#_c_615_p N_A_193_47#_c_912_n 0.00289777f $X=1.985 $Y=2.22
+ $X2=0 $Y2=0
cc_573 N_A_299_66#_c_582_n N_A_193_47#_c_912_n 0.0174959f $X=2.025 $Y=2.055
+ $X2=0 $Y2=0
cc_574 N_A_299_66#_c_577_n N_A_193_47#_c_912_n 7.16422e-19 $X=2.385 $Y=1.29
+ $X2=0 $Y2=0
cc_575 N_A_299_66#_c_571_n N_VPWR_c_1893_n 0.0022015f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_576 N_A_299_66#_c_577_n N_VPWR_c_1893_n 4.77202e-19 $X=2.385 $Y=1.29 $X2=0
+ $Y2=0
cc_577 N_A_299_66#_M1004_g N_VPWR_c_1894_n 0.00172182f $X=3.825 $Y=2.215 $X2=0
+ $Y2=0
cc_578 N_A_299_66#_c_615_p N_VPWR_c_1903_n 0.0106671f $X=1.985 $Y=2.22 $X2=0
+ $Y2=0
cc_579 N_A_299_66#_M1004_g N_VPWR_c_1908_n 0.00422112f $X=3.825 $Y=2.215 $X2=0
+ $Y2=0
cc_580 N_A_299_66#_M1006_s N_VPWR_c_1891_n 0.00338686f $X=1.77 $Y=1.945 $X2=0
+ $Y2=0
cc_581 N_A_299_66#_M1004_g N_VPWR_c_1891_n 0.00636449f $X=3.825 $Y=2.215 $X2=0
+ $Y2=0
cc_582 N_A_299_66#_c_615_p N_VPWR_c_1891_n 0.00425897f $X=1.985 $Y=2.22 $X2=0
+ $Y2=0
cc_583 N_A_299_66#_c_574_n N_A_620_389#_M1018_d 0.00577238f $X=3.68 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_584 N_A_299_66#_c_574_n N_A_620_389#_c_2129_n 0.00902749f $X=3.68 $Y=0.34
+ $X2=0 $Y2=0
cc_585 N_A_299_66#_c_576_n N_A_620_389#_c_2129_n 0.0179883f $X=3.765 $Y=1.52
+ $X2=0 $Y2=0
cc_586 N_A_299_66#_c_568_n N_A_620_389#_c_2098_n 0.00285088f $X=3.825 $Y=1.685
+ $X2=0 $Y2=0
cc_587 N_A_299_66#_M1004_g N_A_620_389#_c_2098_n 0.00418139f $X=3.825 $Y=2.215
+ $X2=0 $Y2=0
cc_588 N_A_299_66#_M1004_g N_A_620_389#_c_2133_n 0.00726498f $X=3.825 $Y=2.215
+ $X2=0 $Y2=0
cc_589 N_A_299_66#_c_568_n N_A_620_389#_c_2106_n 0.00194245f $X=3.825 $Y=1.685
+ $X2=0 $Y2=0
cc_590 N_A_299_66#_M1004_g N_A_620_389#_c_2106_n 0.0130365f $X=3.825 $Y=2.215
+ $X2=0 $Y2=0
cc_591 N_A_299_66#_c_576_n N_A_620_389#_c_2106_n 0.00719f $X=3.765 $Y=1.52 $X2=0
+ $Y2=0
cc_592 N_A_299_66#_c_572_n N_A_620_389#_c_2103_n 0.0137757f $X=2.915 $Y=1.09
+ $X2=0 $Y2=0
cc_593 N_A_299_66#_c_574_n N_A_620_389#_c_2103_n 0.001089f $X=3.68 $Y=0.34 $X2=0
+ $Y2=0
cc_594 N_A_299_66#_c_576_n N_A_620_389#_c_2103_n 0.0397275f $X=3.765 $Y=1.52
+ $X2=0 $Y2=0
cc_595 N_A_299_66#_c_569_n N_VGND_M1025_d 8.82396e-19 $X=2.055 $Y=0.815 $X2=0
+ $Y2=0
cc_596 N_A_299_66#_c_571_n N_VGND_M1025_d 0.00113622f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_597 N_A_299_66#_c_571_n N_VGND_M1009_s 3.82728e-19 $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_598 N_A_299_66#_c_572_n N_VGND_M1009_s 0.00178135f $X=2.915 $Y=1.09 $X2=0
+ $Y2=0
cc_599 N_A_299_66#_c_567_n N_VGND_c_2278_n 3.73754e-19 $X=2.77 $Y=1.09 $X2=0
+ $Y2=0
cc_600 N_A_299_66#_c_569_n N_VGND_c_2278_n 0.00904339f $X=2.055 $Y=0.815 $X2=0
+ $Y2=0
cc_601 N_A_299_66#_c_571_n N_VGND_c_2278_n 0.0126633f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_602 N_A_299_66#_c_571_n N_VGND_c_2279_n 3.29112e-19 $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_603 N_A_299_66#_c_567_n N_VGND_c_2280_n 0.00714612f $X=2.77 $Y=1.09 $X2=0
+ $Y2=0
cc_604 N_A_299_66#_c_571_n N_VGND_c_2280_n 0.0145653f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_605 N_A_299_66#_c_572_n N_VGND_c_2280_n 0.0147146f $X=2.915 $Y=1.09 $X2=0
+ $Y2=0
cc_606 N_A_299_66#_c_573_n N_VGND_c_2280_n 0.0274669f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_607 N_A_299_66#_c_575_n N_VGND_c_2280_n 0.0139003f $X=3.085 $Y=0.34 $X2=0
+ $Y2=0
cc_608 N_A_299_66#_c_577_n N_VGND_c_2280_n 0.00174383f $X=2.385 $Y=1.29 $X2=0
+ $Y2=0
cc_609 N_A_299_66#_c_574_n N_VGND_c_2281_n 8.32093e-19 $X=3.68 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_299_66#_c_574_n N_VGND_c_2287_n 0.049583f $X=3.68 $Y=0.34 $X2=0 $Y2=0
cc_611 N_A_299_66#_c_575_n N_VGND_c_2287_n 0.0115906f $X=3.085 $Y=0.34 $X2=0
+ $Y2=0
cc_612 N_A_299_66#_c_646_p N_VGND_c_2298_n 0.00594281f $X=1.62 $Y=0.56 $X2=0
+ $Y2=0
cc_613 N_A_299_66#_c_569_n N_VGND_c_2298_n 0.00195917f $X=2.055 $Y=0.815 $X2=0
+ $Y2=0
cc_614 N_A_299_66#_c_567_n N_VGND_c_2301_n 7.52198e-19 $X=2.77 $Y=1.09 $X2=0
+ $Y2=0
cc_615 N_A_299_66#_c_646_p N_VGND_c_2301_n 0.00591457f $X=1.62 $Y=0.56 $X2=0
+ $Y2=0
cc_616 N_A_299_66#_c_569_n N_VGND_c_2301_n 0.00455645f $X=2.055 $Y=0.815 $X2=0
+ $Y2=0
cc_617 N_A_299_66#_c_571_n N_VGND_c_2301_n 0.00116163f $X=2.065 $Y=1.455 $X2=0
+ $Y2=0
cc_618 N_A_299_66#_c_574_n N_VGND_c_2301_n 0.0254695f $X=3.68 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_299_66#_c_575_n N_VGND_c_2301_n 0.00576957f $X=3.085 $Y=0.34 $X2=0
+ $Y2=0
cc_620 N_A_299_66#_c_572_n A_569_119# 4.64076e-19 $X=2.915 $Y=1.09 $X2=-0.19
+ $Y2=-0.24
cc_621 N_A_299_66#_c_573_n A_569_119# 0.00382069f $X=3 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_622 N_D_M1018_g N_SCE_c_751_n 0.00900792f $X=3.13 $Y=0.805 $X2=0 $Y2=0
cc_623 D N_SCE_c_758_n 0.00218397f $X=2.795 $Y=1.445 $X2=0 $Y2=0
cc_624 N_D_c_710_n N_SCE_c_758_n 0.00980075f $X=3.035 $Y=1.62 $X2=0 $Y2=0
cc_625 N_D_M1026_g N_SCE_M1003_g 0.0395364f $X=3.025 $Y=2.215 $X2=0 $Y2=0
cc_626 D N_SCE_M1003_g 0.0082176f $X=2.925 $Y=2.125 $X2=0 $Y2=0
cc_627 N_D_M1018_g N_SCE_c_753_n 0.00950132f $X=3.13 $Y=0.805 $X2=0 $Y2=0
cc_628 D N_A_193_47#_c_912_n 0.00553465f $X=2.795 $Y=1.445 $X2=0 $Y2=0
cc_629 D N_A_193_47#_c_912_n 0.0237797f $X=2.925 $Y=2.125 $X2=0 $Y2=0
cc_630 N_D_c_710_n N_A_193_47#_c_912_n 0.0020276f $X=3.035 $Y=1.62 $X2=0 $Y2=0
cc_631 N_D_M1026_g N_VPWR_c_1908_n 0.00357668f $X=3.025 $Y=2.215 $X2=0 $Y2=0
cc_632 D N_VPWR_c_1908_n 0.0148222f $X=2.925 $Y=2.125 $X2=0 $Y2=0
cc_633 N_D_M1026_g N_VPWR_c_1891_n 0.00594623f $X=3.025 $Y=2.215 $X2=0 $Y2=0
cc_634 D N_VPWR_c_1891_n 0.00431744f $X=2.925 $Y=2.125 $X2=0 $Y2=0
cc_635 D A_538_389# 0.0064363f $X=2.925 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_636 N_D_M1026_g N_A_620_389#_c_2098_n 5.25693e-19 $X=3.025 $Y=2.215 $X2=0
+ $Y2=0
cc_637 N_D_M1018_g N_A_620_389#_c_2098_n 0.00974864f $X=3.13 $Y=0.805 $X2=0
+ $Y2=0
cc_638 D N_A_620_389#_c_2098_n 0.0433703f $X=2.795 $Y=1.445 $X2=0 $Y2=0
cc_639 N_D_M1026_g N_A_620_389#_c_2133_n 0.00141769f $X=3.025 $Y=2.215 $X2=0
+ $Y2=0
cc_640 N_D_M1026_g N_A_620_389#_c_2107_n 7.97227e-19 $X=3.025 $Y=2.215 $X2=0
+ $Y2=0
cc_641 D N_A_620_389#_c_2107_n 0.00782199f $X=2.925 $Y=2.125 $X2=0 $Y2=0
cc_642 N_D_M1018_g N_A_620_389#_c_2103_n 0.00367537f $X=3.13 $Y=0.805 $X2=0
+ $Y2=0
cc_643 N_D_M1018_g N_VGND_c_2280_n 2.94691e-19 $X=3.13 $Y=0.805 $X2=0 $Y2=0
cc_644 N_SCE_c_751_n N_SCD_M1030_g 0.041995f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_645 N_SCE_c_753_n SCD 0.0184489f $X=3.835 $Y=0.255 $X2=0 $Y2=0
cc_646 N_SCE_c_761_n N_A_193_47#_c_924_n 0.0271009f $X=1.597 $Y=2.117 $X2=0
+ $Y2=0
cc_647 N_SCE_c_755_n N_A_193_47#_c_924_n 0.00343293f $X=1.645 $Y=1.31 $X2=0
+ $Y2=0
cc_648 N_SCE_M1025_g N_A_193_47#_c_894_n 0.00514755f $X=1.83 $Y=0.54 $X2=0 $Y2=0
cc_649 N_SCE_c_754_n N_A_193_47#_c_894_n 0.00379441f $X=1.645 $Y=1.31 $X2=0
+ $Y2=0
cc_650 N_SCE_c_755_n N_A_193_47#_c_894_n 0.0487008f $X=1.645 $Y=1.31 $X2=0 $Y2=0
cc_651 N_SCE_M1025_g N_A_193_47#_c_900_n 9.91666e-19 $X=1.83 $Y=0.54 $X2=0 $Y2=0
cc_652 N_SCE_M1006_g N_A_193_47#_c_912_n 0.00380606f $X=2.195 $Y=2.215 $X2=0
+ $Y2=0
cc_653 N_SCE_c_758_n N_A_193_47#_c_912_n 0.00146367f $X=2.54 $Y=1.71 $X2=0 $Y2=0
cc_654 N_SCE_M1003_g N_A_193_47#_c_912_n 0.0063259f $X=2.615 $Y=2.215 $X2=0
+ $Y2=0
cc_655 N_SCE_c_761_n N_A_193_47#_c_912_n 7.97975e-19 $X=1.597 $Y=2.117 $X2=0
+ $Y2=0
cc_656 N_SCE_c_754_n N_A_193_47#_c_912_n 0.00668205f $X=1.645 $Y=1.31 $X2=0
+ $Y2=0
cc_657 N_SCE_c_755_n N_A_193_47#_c_912_n 0.0209535f $X=1.645 $Y=1.31 $X2=0 $Y2=0
cc_658 N_SCE_c_755_n N_A_193_47#_c_913_n 0.00162128f $X=1.645 $Y=1.31 $X2=0
+ $Y2=0
cc_659 N_SCE_c_755_n N_A_193_47#_c_919_n 0.0123906f $X=1.645 $Y=1.31 $X2=0 $Y2=0
cc_660 N_SCE_M1006_g N_VPWR_c_1893_n 0.0029521f $X=2.195 $Y=2.215 $X2=0 $Y2=0
cc_661 N_SCE_c_758_n N_VPWR_c_1893_n 0.00207809f $X=2.54 $Y=1.71 $X2=0 $Y2=0
cc_662 N_SCE_M1003_g N_VPWR_c_1893_n 0.0029521f $X=2.615 $Y=2.215 $X2=0 $Y2=0
cc_663 N_SCE_M1006_g N_VPWR_c_1903_n 0.00543919f $X=2.195 $Y=2.215 $X2=0 $Y2=0
cc_664 SCE N_VPWR_c_1903_n 0.0188207f $X=1.56 $Y=2.125 $X2=0 $Y2=0
cc_665 N_SCE_M1003_g N_VPWR_c_1908_n 0.00585385f $X=2.615 $Y=2.215 $X2=0 $Y2=0
cc_666 N_SCE_M1006_g N_VPWR_c_1891_n 0.00745913f $X=2.195 $Y=2.215 $X2=0 $Y2=0
cc_667 N_SCE_M1003_g N_VPWR_c_1891_n 0.00631707f $X=2.615 $Y=2.215 $X2=0 $Y2=0
cc_668 SCE N_VPWR_c_1891_n 0.00481824f $X=1.56 $Y=2.125 $X2=0 $Y2=0
cc_669 N_SCE_c_753_n N_A_620_389#_c_2129_n 0.00186401f $X=3.835 $Y=0.255 $X2=0
+ $Y2=0
cc_670 N_SCE_M1025_g N_VGND_c_2278_n 0.00716396f $X=1.83 $Y=0.54 $X2=0 $Y2=0
cc_671 N_SCE_c_751_n N_VGND_c_2278_n 0.015168f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_672 N_SCE_c_752_n N_VGND_c_2278_n 0.00414542f $X=1.905 $Y=0.18 $X2=0 $Y2=0
cc_673 N_SCE_c_751_n N_VGND_c_2279_n 0.00648503f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_674 N_SCE_M1025_g N_VGND_c_2280_n 0.00354677f $X=1.83 $Y=0.54 $X2=0 $Y2=0
cc_675 N_SCE_c_751_n N_VGND_c_2280_n 0.0230698f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_676 N_SCE_c_751_n N_VGND_c_2281_n 0.00262905f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_677 N_SCE_c_751_n N_VGND_c_2287_n 0.035035f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_678 N_SCE_c_752_n N_VGND_c_2298_n 0.00350026f $X=1.905 $Y=0.18 $X2=0 $Y2=0
cc_679 N_SCE_c_751_n N_VGND_c_2301_n 0.0526889f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_680 N_SCE_c_752_n N_VGND_c_2301_n 0.00563019f $X=1.905 $Y=0.18 $X2=0 $Y2=0
cc_681 N_SCD_M1035_g N_A_193_47#_c_912_n 0.004386f $X=4.255 $Y=2.215 $X2=0 $Y2=0
cc_682 SCD N_A_193_47#_c_912_n 0.00510982f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_683 N_SCD_c_851_n N_A_193_47#_c_912_n 0.00179125f $X=4.31 $Y=1.535 $X2=0
+ $Y2=0
cc_684 N_SCD_c_851_n N_A_193_47#_c_917_n 0.00101301f $X=4.31 $Y=1.535 $X2=0
+ $Y2=0
cc_685 N_SCD_M1035_g N_VPWR_c_1894_n 0.0105334f $X=4.255 $Y=2.215 $X2=0 $Y2=0
cc_686 N_SCD_M1035_g N_VPWR_c_1908_n 0.00337001f $X=4.255 $Y=2.215 $X2=0 $Y2=0
cc_687 N_SCD_M1035_g N_VPWR_c_1891_n 0.00379951f $X=4.255 $Y=2.215 $X2=0 $Y2=0
cc_688 SCD N_A_620_389#_c_2098_n 5.20671e-19 $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_689 N_SCD_M1035_g N_A_620_389#_c_2106_n 0.0129931f $X=4.255 $Y=2.215 $X2=0
+ $Y2=0
cc_690 SCD N_A_620_389#_c_2106_n 0.0178473f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_691 N_SCD_c_851_n N_A_620_389#_c_2106_n 0.00321619f $X=4.31 $Y=1.535 $X2=0
+ $Y2=0
cc_692 N_SCD_M1035_g N_A_620_389#_c_2099_n 0.00923383f $X=4.255 $Y=2.215 $X2=0
+ $Y2=0
cc_693 N_SCD_M1030_g N_A_620_389#_c_2099_n 0.0101759f $X=4.385 $Y=0.54 $X2=0
+ $Y2=0
cc_694 SCD N_A_620_389#_c_2099_n 0.0595722f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_695 N_SCD_M1030_g N_A_620_389#_c_2101_n 0.00185622f $X=4.385 $Y=0.54 $X2=0
+ $Y2=0
cc_696 SCD N_A_620_389#_c_2101_n 0.0150549f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_697 N_SCD_M1030_g N_A_620_389#_c_2102_n 0.00249829f $X=4.385 $Y=0.54 $X2=0
+ $Y2=0
cc_698 N_SCD_M1030_g N_VGND_c_2281_n 0.00852014f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_699 SCD N_VGND_c_2281_n 0.0113287f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_700 N_SCD_M1030_g N_VGND_c_2287_n 0.00405203f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_701 SCD N_VGND_c_2287_n 0.0167004f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_702 N_SCD_M1030_g N_VGND_c_2301_n 0.00614202f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_703 SCD N_VGND_c_2301_n 0.0121815f $X=4.075 $Y=1.445 $X2=0 $Y2=0
cc_704 N_A_193_47#_c_907_n N_A_1245_303#_M1021_d 3.72821e-19 $X=8.31 $Y=1.58
+ $X2=0 $Y2=0
cc_705 N_A_193_47#_c_908_n N_A_1245_303#_M1021_d 0.00157673f $X=8.095 $Y=1.58
+ $X2=0 $Y2=0
cc_706 N_A_193_47#_c_914_n N_A_1245_303#_M1021_d 0.00171601f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_707 N_A_193_47#_c_914_n N_A_1245_303#_M1038_g 0.00117999f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_708 N_A_193_47#_c_896_n N_A_1245_303#_M1010_g 0.00101776f $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_709 N_A_193_47#_c_901_n N_A_1245_303#_M1010_g 0.0284437f $X=5.8 $Y=0.705
+ $X2=0 $Y2=0
cc_710 N_A_193_47#_c_914_n N_A_1245_303#_c_1167_n 0.0203611f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_711 N_A_193_47#_c_914_n N_A_1245_303#_c_1168_n 0.00588349f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_712 N_A_193_47#_c_893_n N_A_1245_303#_c_1193_n 0.00348548f $X=7.885 $Y=0.705
+ $X2=0 $Y2=0
cc_713 N_A_193_47#_c_907_n N_A_1245_303#_c_1169_n 0.00289443f $X=8.31 $Y=1.58
+ $X2=0 $Y2=0
cc_714 N_A_193_47#_c_908_n N_A_1245_303#_c_1169_n 0.0119354f $X=8.095 $Y=1.58
+ $X2=0 $Y2=0
cc_715 N_A_193_47#_c_909_n N_A_1245_303#_c_1169_n 0.00834716f $X=8.415 $Y=1.58
+ $X2=0 $Y2=0
cc_716 N_A_193_47#_c_914_n N_A_1245_303#_c_1169_n 0.0183749f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_717 N_A_193_47#_c_916_n N_A_1245_303#_c_1169_n 0.00158802f $X=8.53 $Y=1.87
+ $X2=0 $Y2=0
cc_718 N_A_193_47#_c_898_n N_A_1245_303#_c_1181_n 0.0573468f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_719 N_A_193_47#_c_899_n N_A_1245_303#_c_1181_n 0.00348548f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_720 N_A_193_47#_c_909_n N_A_1245_303#_c_1171_n 0.00205198f $X=8.415 $Y=1.58
+ $X2=0 $Y2=0
cc_721 N_A_193_47#_c_914_n N_A_1245_303#_c_1171_n 0.0199108f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_722 N_A_193_47#_c_908_n N_A_1245_303#_c_1164_n 0.0120685f $X=8.095 $Y=1.58
+ $X2=0 $Y2=0
cc_723 N_A_193_47#_c_914_n N_RESET_B_M1033_g 0.0046833f $X=8.385 $Y=1.87 $X2=0
+ $Y2=0
cc_724 N_A_193_47#_c_898_n N_RESET_B_c_1282_n 0.0145517f $X=8.01 $Y=0.87 $X2=0
+ $Y2=0
cc_725 N_A_193_47#_c_899_n N_RESET_B_c_1282_n 0.00385878f $X=8.01 $Y=0.87 $X2=0
+ $Y2=0
cc_726 N_A_193_47#_c_893_n N_A_1079_413#_M1039_g 0.011215f $X=7.885 $Y=0.705
+ $X2=0 $Y2=0
cc_727 N_A_193_47#_c_898_n N_A_1079_413#_c_1451_n 7.85121e-19 $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_728 N_A_193_47#_c_899_n N_A_1079_413#_c_1451_n 0.00297112f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_729 N_A_193_47#_c_908_n N_A_1079_413#_c_1451_n 0.00170165f $X=8.095 $Y=1.58
+ $X2=0 $Y2=0
cc_730 N_A_193_47#_c_909_n N_A_1079_413#_c_1452_n 6.7969e-19 $X=8.415 $Y=1.58
+ $X2=0 $Y2=0
cc_731 N_A_193_47#_c_914_n N_A_1079_413#_c_1452_n 0.00270328f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_732 N_A_193_47#_c_895_n N_A_1079_413#_c_1479_n 4.06924e-19 $X=5.495 $Y=0.87
+ $X2=0 $Y2=0
cc_733 N_A_193_47#_c_896_n N_A_1079_413#_c_1479_n 0.023426f $X=5.8 $Y=0.87 $X2=0
+ $Y2=0
cc_734 N_A_193_47#_c_897_n N_A_1079_413#_c_1479_n 0.00243773f $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_735 N_A_193_47#_c_901_n N_A_1079_413#_c_1479_n 0.00884831f $X=5.8 $Y=0.705
+ $X2=0 $Y2=0
cc_736 N_A_193_47#_c_896_n N_A_1079_413#_c_1445_n 0.00859821f $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_737 N_A_193_47#_c_897_n N_A_1079_413#_c_1445_n 5.36138e-19 $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_738 N_A_193_47#_c_914_n N_A_1079_413#_c_1445_n 0.00508729f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_739 N_A_193_47#_c_896_n N_A_1079_413#_c_1446_n 0.0106449f $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_740 N_A_193_47#_c_897_n N_A_1079_413#_c_1446_n 9.03057e-19 $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_741 N_A_193_47#_c_902_n N_A_1079_413#_c_1446_n 0.012565f $X=5.37 $Y=1.575
+ $X2=0 $Y2=0
cc_742 N_A_193_47#_c_896_n N_A_1079_413#_c_1447_n 0.0245019f $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_743 N_A_193_47#_c_897_n N_A_1079_413#_c_1447_n 0.00103375f $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_744 N_A_193_47#_c_901_n N_A_1079_413#_c_1447_n 0.00463572f $X=5.8 $Y=0.705
+ $X2=0 $Y2=0
cc_745 N_A_193_47#_c_902_n N_A_1079_413#_c_1447_n 0.00379951f $X=5.37 $Y=1.575
+ $X2=0 $Y2=0
cc_746 N_A_193_47#_M1007_g N_A_1079_413#_c_1467_n 0.00376625f $X=5.32 $Y=2.275
+ $X2=0 $Y2=0
cc_747 N_A_193_47#_c_914_n N_A_1079_413#_c_1467_n 0.00363572f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_748 N_A_193_47#_c_915_n N_A_1079_413#_c_1467_n 0.00241651f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_749 N_A_193_47#_c_918_n N_A_1079_413#_c_1467_n 0.00151282f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_750 N_A_193_47#_M1007_g N_A_1079_413#_c_1455_n 0.00181645f $X=5.32 $Y=2.275
+ $X2=0 $Y2=0
cc_751 N_A_193_47#_c_914_n N_A_1079_413#_c_1455_n 0.0170929f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_752 N_A_193_47#_c_915_n N_A_1079_413#_c_1455_n 0.00294259f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_753 N_A_193_47#_c_917_n N_A_1079_413#_c_1455_n 0.00159864f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_754 N_A_193_47#_c_902_n N_A_1079_413#_c_1455_n 0.0410116f $X=5.37 $Y=1.575
+ $X2=0 $Y2=0
cc_755 N_A_193_47#_c_914_n N_A_1079_413#_c_1456_n 0.00155738f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_756 N_A_193_47#_c_899_n N_A_1079_413#_c_1450_n 0.011215f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_757 N_A_193_47#_c_914_n N_A_1079_413#_c_1450_n 3.00671e-19 $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_758 N_A_193_47#_M1031_g N_A_1767_21#_M1028_g 0.0350828f $X=8.715 $Y=2.275
+ $X2=0 $Y2=0
cc_759 N_A_193_47#_c_909_n N_A_1767_21#_M1028_g 3.42026e-19 $X=8.415 $Y=1.58
+ $X2=0 $Y2=0
cc_760 N_A_193_47#_c_910_n N_A_1767_21#_M1028_g 9.89492e-19 $X=8.69 $Y=1.805
+ $X2=0 $Y2=0
cc_761 N_A_193_47#_c_911_n N_A_1767_21#_M1028_g 0.0210643f $X=8.705 $Y=1.74
+ $X2=0 $Y2=0
cc_762 N_A_193_47#_c_898_n N_A_1592_47#_c_1783_n 0.0060004f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_763 N_A_193_47#_c_899_n N_A_1592_47#_c_1783_n 0.00264523f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_764 N_A_193_47#_M1031_g N_A_1592_47#_c_1779_n 0.0127238f $X=8.715 $Y=2.275
+ $X2=0 $Y2=0
cc_765 N_A_193_47#_c_909_n N_A_1592_47#_c_1779_n 0.0119715f $X=8.415 $Y=1.58
+ $X2=0 $Y2=0
cc_766 N_A_193_47#_c_910_n N_A_1592_47#_c_1779_n 0.0206842f $X=8.69 $Y=1.805
+ $X2=0 $Y2=0
cc_767 N_A_193_47#_c_911_n N_A_1592_47#_c_1779_n 3.21879e-19 $X=8.705 $Y=1.74
+ $X2=0 $Y2=0
cc_768 N_A_193_47#_c_914_n N_A_1592_47#_c_1779_n 2.92836e-19 $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_769 N_A_193_47#_c_916_n N_A_1592_47#_c_1779_n 0.00341459f $X=8.53 $Y=1.87
+ $X2=0 $Y2=0
cc_770 N_A_193_47#_c_898_n N_A_1592_47#_c_1775_n 0.00363555f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_771 N_A_193_47#_M1031_g N_A_1592_47#_c_1780_n 0.00160397f $X=8.715 $Y=2.275
+ $X2=0 $Y2=0
cc_772 N_A_193_47#_c_910_n N_A_1592_47#_c_1780_n 0.015723f $X=8.69 $Y=1.805
+ $X2=0 $Y2=0
cc_773 N_A_193_47#_c_911_n N_A_1592_47#_c_1780_n 4.32259e-19 $X=8.705 $Y=1.74
+ $X2=0 $Y2=0
cc_774 N_A_193_47#_c_916_n N_A_1592_47#_c_1780_n 0.00205399f $X=8.53 $Y=1.87
+ $X2=0 $Y2=0
cc_775 N_A_193_47#_c_898_n N_A_1592_47#_c_1781_n 0.00513856f $X=8.01 $Y=0.87
+ $X2=0 $Y2=0
cc_776 N_A_193_47#_c_909_n N_A_1592_47#_c_1781_n 0.00596879f $X=8.415 $Y=1.58
+ $X2=0 $Y2=0
cc_777 N_A_193_47#_c_910_n N_A_1592_47#_c_1781_n 0.0186201f $X=8.69 $Y=1.805
+ $X2=0 $Y2=0
cc_778 N_A_193_47#_c_911_n N_A_1592_47#_c_1781_n 0.00371643f $X=8.705 $Y=1.74
+ $X2=0 $Y2=0
cc_779 N_A_193_47#_c_914_n N_VPWR_M1021_s 2.16592e-19 $X=8.385 $Y=1.87 $X2=0
+ $Y2=0
cc_780 N_A_193_47#_c_912_n N_VPWR_c_1893_n 0.00399021f $X=5.265 $Y=1.87 $X2=0
+ $Y2=0
cc_781 N_A_193_47#_M1007_g N_VPWR_c_1894_n 0.00247529f $X=5.32 $Y=2.275 $X2=0
+ $Y2=0
cc_782 N_A_193_47#_c_912_n N_VPWR_c_1894_n 0.00117433f $X=5.265 $Y=1.87 $X2=0
+ $Y2=0
cc_783 N_A_193_47#_c_914_n N_VPWR_c_1895_n 0.00247761f $X=8.385 $Y=1.87 $X2=0
+ $Y2=0
cc_784 N_A_193_47#_c_924_n N_VPWR_c_1903_n 0.0116213f $X=1.12 $Y=1.96 $X2=0
+ $Y2=0
cc_785 N_A_193_47#_c_914_n N_VPWR_c_1905_n 0.00131518f $X=8.385 $Y=1.87 $X2=0
+ $Y2=0
cc_786 N_A_193_47#_M1007_g N_VPWR_c_1906_n 0.00541083f $X=5.32 $Y=2.275 $X2=0
+ $Y2=0
cc_787 N_A_193_47#_M1031_g N_VPWR_c_1910_n 0.00357877f $X=8.715 $Y=2.275 $X2=0
+ $Y2=0
cc_788 N_A_193_47#_M1041_d N_VPWR_c_1891_n 0.00222627f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_789 N_A_193_47#_M1007_g N_VPWR_c_1891_n 0.00731044f $X=5.32 $Y=2.275 $X2=0
+ $Y2=0
cc_790 N_A_193_47#_M1031_g N_VPWR_c_1891_n 0.00525625f $X=8.715 $Y=2.275 $X2=0
+ $Y2=0
cc_791 N_A_193_47#_c_924_n N_VPWR_c_1891_n 0.00290138f $X=1.12 $Y=1.96 $X2=0
+ $Y2=0
cc_792 N_A_193_47#_c_909_n N_VPWR_c_1891_n 2.9554e-19 $X=8.415 $Y=1.58 $X2=0
+ $Y2=0
cc_793 N_A_193_47#_c_912_n N_VPWR_c_1891_n 0.189767f $X=5.265 $Y=1.87 $X2=0
+ $Y2=0
cc_794 N_A_193_47#_c_913_n N_VPWR_c_1891_n 0.0157502f $X=1.27 $Y=1.87 $X2=0
+ $Y2=0
cc_795 N_A_193_47#_c_914_n N_VPWR_c_1891_n 0.129916f $X=8.385 $Y=1.87 $X2=0
+ $Y2=0
cc_796 N_A_193_47#_c_915_n N_VPWR_c_1891_n 0.01602f $X=5.555 $Y=1.87 $X2=0 $Y2=0
cc_797 N_A_193_47#_c_916_n N_VPWR_c_1891_n 0.0158836f $X=8.53 $Y=1.87 $X2=0
+ $Y2=0
cc_798 N_A_193_47#_c_918_n N_VPWR_c_1891_n 0.00217218f $X=5.33 $Y=1.74 $X2=0
+ $Y2=0
cc_799 N_A_193_47#_c_919_n N_VPWR_c_1891_n 7.75725e-19 $X=1.23 $Y=1.815 $X2=0
+ $Y2=0
cc_800 N_A_193_47#_c_912_n N_A_620_389#_c_2098_n 0.0132627f $X=5.265 $Y=1.87
+ $X2=0 $Y2=0
cc_801 N_A_193_47#_c_912_n N_A_620_389#_c_2133_n 2.97781e-19 $X=5.265 $Y=1.87
+ $X2=0 $Y2=0
cc_802 N_A_193_47#_c_912_n N_A_620_389#_c_2106_n 0.0327141f $X=5.265 $Y=1.87
+ $X2=0 $Y2=0
cc_803 N_A_193_47#_c_912_n N_A_620_389#_c_2107_n 0.0107741f $X=5.265 $Y=1.87
+ $X2=0 $Y2=0
cc_804 N_A_193_47#_M1007_g N_A_620_389#_c_2099_n 0.00829892f $X=5.32 $Y=2.275
+ $X2=0 $Y2=0
cc_805 N_A_193_47#_c_895_n N_A_620_389#_c_2099_n 0.00488629f $X=5.495 $Y=0.87
+ $X2=0 $Y2=0
cc_806 N_A_193_47#_c_912_n N_A_620_389#_c_2099_n 0.0385489f $X=5.265 $Y=1.87
+ $X2=0 $Y2=0
cc_807 N_A_193_47#_c_915_n N_A_620_389#_c_2099_n 0.00146664f $X=5.555 $Y=1.87
+ $X2=0 $Y2=0
cc_808 N_A_193_47#_c_917_n N_A_620_389#_c_2099_n 0.00491906f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_809 N_A_193_47#_c_918_n N_A_620_389#_c_2099_n 0.012343f $X=5.33 $Y=1.74 $X2=0
+ $Y2=0
cc_810 N_A_193_47#_c_902_n N_A_620_389#_c_2099_n 0.00662023f $X=5.37 $Y=1.575
+ $X2=0 $Y2=0
cc_811 N_A_193_47#_c_895_n N_A_620_389#_c_2100_n 0.014624f $X=5.495 $Y=0.87
+ $X2=0 $Y2=0
cc_812 N_A_193_47#_c_897_n N_A_620_389#_c_2100_n 2.34565e-19 $X=5.8 $Y=0.87
+ $X2=0 $Y2=0
cc_813 N_A_193_47#_c_895_n N_A_620_389#_c_2102_n 6.92432e-19 $X=5.495 $Y=0.87
+ $X2=0 $Y2=0
cc_814 N_A_193_47#_c_914_n N_A_1191_413#_c_2203_n 0.022443f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_815 N_A_193_47#_c_914_n N_A_1191_413#_c_2204_n 0.00700259f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_816 N_A_193_47#_c_914_n N_A_1191_413#_c_2205_n 0.00567047f $X=8.385 $Y=1.87
+ $X2=0 $Y2=0
cc_817 N_A_193_47#_c_900_n N_VGND_c_2278_n 0.00157059f $X=1.23 $Y=0.51 $X2=0
+ $Y2=0
cc_818 N_A_193_47#_c_893_n N_VGND_c_2289_n 0.0051118f $X=7.885 $Y=0.705 $X2=0
+ $Y2=0
cc_819 N_A_193_47#_c_898_n N_VGND_c_2289_n 0.00183172f $X=8.01 $Y=0.87 $X2=0
+ $Y2=0
cc_820 N_A_193_47#_c_899_n N_VGND_c_2289_n 2.13253e-19 $X=8.01 $Y=0.87 $X2=0
+ $Y2=0
cc_821 N_A_193_47#_c_900_n N_VGND_c_2298_n 0.0125774f $X=1.23 $Y=0.51 $X2=0
+ $Y2=0
cc_822 N_A_193_47#_c_895_n N_VGND_c_2299_n 0.00257694f $X=5.495 $Y=0.87 $X2=0
+ $Y2=0
cc_823 N_A_193_47#_c_901_n N_VGND_c_2299_n 0.00368123f $X=5.8 $Y=0.705 $X2=0
+ $Y2=0
cc_824 N_A_193_47#_M1022_d N_VGND_c_2301_n 0.00390713f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_825 N_A_193_47#_c_893_n N_VGND_c_2301_n 0.00649711f $X=7.885 $Y=0.705 $X2=0
+ $Y2=0
cc_826 N_A_193_47#_c_895_n N_VGND_c_2301_n 0.00403634f $X=5.495 $Y=0.87 $X2=0
+ $Y2=0
cc_827 N_A_193_47#_c_898_n N_VGND_c_2301_n 0.00150843f $X=8.01 $Y=0.87 $X2=0
+ $Y2=0
cc_828 N_A_193_47#_c_900_n N_VGND_c_2301_n 0.0107503f $X=1.23 $Y=0.51 $X2=0
+ $Y2=0
cc_829 N_A_193_47#_c_901_n N_VGND_c_2301_n 0.00574204f $X=5.8 $Y=0.705 $X2=0
+ $Y2=0
cc_830 N_A_1245_303#_M1038_g N_RESET_B_M1033_g 0.0200274f $X=6.3 $Y=2.275 $X2=0
+ $Y2=0
cc_831 N_A_1245_303#_M1010_g N_RESET_B_M1033_g 0.0156143f $X=6.39 $Y=0.445 $X2=0
+ $Y2=0
cc_832 N_A_1245_303#_c_1167_n N_RESET_B_M1033_g 0.0118675f $X=7.455 $Y=1.68
+ $X2=0 $Y2=0
cc_833 N_A_1245_303#_c_1168_n N_RESET_B_M1033_g 0.0229835f $X=6.45 $Y=1.68 $X2=0
+ $Y2=0
cc_834 N_A_1245_303#_c_1171_n N_RESET_B_M1033_g 0.00336641f $X=7.585 $Y=1.68
+ $X2=0 $Y2=0
cc_835 N_A_1245_303#_c_1164_n N_RESET_B_M1033_g 0.00114583f $X=7.585 $Y=1.595
+ $X2=0 $Y2=0
cc_836 N_A_1245_303#_M1010_g N_RESET_B_c_1280_n 0.0034695f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_837 N_A_1245_303#_M1010_g N_RESET_B_c_1281_n 0.00171689f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_838 N_A_1245_303#_c_1181_n N_RESET_B_c_1281_n 0.0017415f $X=7.585 $Y=0.835
+ $X2=0 $Y2=0
cc_839 N_A_1245_303#_c_1164_n N_RESET_B_c_1281_n 0.00429759f $X=7.585 $Y=1.595
+ $X2=0 $Y2=0
cc_840 N_A_1245_303#_c_1214_p N_RESET_B_c_1282_n 0.00176185f $X=7.62 $Y=0.36
+ $X2=0 $Y2=0
cc_841 N_A_1245_303#_c_1181_n N_RESET_B_c_1282_n 0.0120924f $X=7.585 $Y=0.835
+ $X2=0 $Y2=0
cc_842 N_A_1245_303#_c_1164_n N_RESET_B_c_1282_n 0.00688409f $X=7.585 $Y=1.595
+ $X2=0 $Y2=0
cc_843 N_A_1245_303#_c_1181_n N_RESET_B_c_1283_n 0.00169962f $X=7.585 $Y=0.835
+ $X2=0 $Y2=0
cc_844 N_A_1245_303#_c_1164_n N_RESET_B_c_1283_n 0.00124786f $X=7.585 $Y=1.595
+ $X2=0 $Y2=0
cc_845 N_A_1245_303#_M1010_g N_RESET_B_c_1286_n 0.0641839f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_846 N_A_1245_303#_c_1214_p N_RESET_B_c_1286_n 9.50035e-19 $X=7.62 $Y=0.36
+ $X2=0 $Y2=0
cc_847 N_A_1245_303#_c_1193_n N_A_1079_413#_M1039_g 0.00611564f $X=7.585
+ $Y=0.705 $X2=0 $Y2=0
cc_848 N_A_1245_303#_c_1214_p N_A_1079_413#_M1039_g 0.00225962f $X=7.62 $Y=0.36
+ $X2=0 $Y2=0
cc_849 N_A_1245_303#_c_1181_n N_A_1079_413#_M1039_g 0.003859f $X=7.585 $Y=0.835
+ $X2=0 $Y2=0
cc_850 N_A_1245_303#_c_1164_n N_A_1079_413#_M1039_g 0.0114806f $X=7.585 $Y=1.595
+ $X2=0 $Y2=0
cc_851 N_A_1245_303#_c_1169_n N_A_1079_413#_c_1451_n 4.11153e-19 $X=7.97 $Y=1.92
+ $X2=0 $Y2=0
cc_852 N_A_1245_303#_c_1181_n N_A_1079_413#_c_1451_n 8.88512e-19 $X=7.585
+ $Y=0.835 $X2=0 $Y2=0
cc_853 N_A_1245_303#_c_1164_n N_A_1079_413#_c_1451_n 0.0144527f $X=7.585
+ $Y=1.595 $X2=0 $Y2=0
cc_854 N_A_1245_303#_c_1169_n N_A_1079_413#_c_1452_n 0.0135494f $X=7.97 $Y=1.92
+ $X2=0 $Y2=0
cc_855 N_A_1245_303#_c_1170_n N_A_1079_413#_c_1452_n 0.00464109f $X=8.055 $Y=2.3
+ $X2=0 $Y2=0
cc_856 N_A_1245_303#_c_1171_n N_A_1079_413#_c_1452_n 0.00237614f $X=7.585
+ $Y=1.68 $X2=0 $Y2=0
cc_857 N_A_1245_303#_c_1164_n N_A_1079_413#_c_1452_n 0.00556533f $X=7.585
+ $Y=1.595 $X2=0 $Y2=0
cc_858 N_A_1245_303#_M1010_g N_A_1079_413#_c_1479_n 0.00572805f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_859 N_A_1245_303#_M1010_g N_A_1079_413#_c_1447_n 0.0186614f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_860 N_A_1245_303#_M1010_g N_A_1079_413#_c_1448_n 0.00932949f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_861 N_A_1245_303#_c_1167_n N_A_1079_413#_c_1448_n 0.0449153f $X=7.455 $Y=1.68
+ $X2=0 $Y2=0
cc_862 N_A_1245_303#_c_1168_n N_A_1079_413#_c_1448_n 0.00289824f $X=6.45 $Y=1.68
+ $X2=0 $Y2=0
cc_863 N_A_1245_303#_M1038_g N_A_1079_413#_c_1455_n 2.86579e-19 $X=6.3 $Y=2.275
+ $X2=0 $Y2=0
cc_864 N_A_1245_303#_M1010_g N_A_1079_413#_c_1455_n 6.14735e-19 $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_865 N_A_1245_303#_c_1167_n N_A_1079_413#_c_1455_n 0.00579774f $X=7.455
+ $Y=1.68 $X2=0 $Y2=0
cc_866 N_A_1245_303#_c_1168_n N_A_1079_413#_c_1455_n 0.00222517f $X=6.45 $Y=1.68
+ $X2=0 $Y2=0
cc_867 N_A_1245_303#_M1010_g N_A_1079_413#_c_1456_n 0.00333698f $X=6.39 $Y=0.445
+ $X2=0 $Y2=0
cc_868 N_A_1245_303#_c_1167_n N_A_1079_413#_c_1456_n 0.00280794f $X=7.455
+ $Y=1.68 $X2=0 $Y2=0
cc_869 N_A_1245_303#_c_1168_n N_A_1079_413#_c_1456_n 0.0029449f $X=6.45 $Y=1.68
+ $X2=0 $Y2=0
cc_870 N_A_1245_303#_c_1167_n N_A_1079_413#_c_1449_n 0.0096056f $X=7.455 $Y=1.68
+ $X2=0 $Y2=0
cc_871 N_A_1245_303#_c_1164_n N_A_1079_413#_c_1449_n 0.0266441f $X=7.585
+ $Y=1.595 $X2=0 $Y2=0
cc_872 N_A_1245_303#_c_1167_n N_A_1079_413#_c_1450_n 0.00625181f $X=7.455
+ $Y=1.68 $X2=0 $Y2=0
cc_873 N_A_1245_303#_c_1171_n N_A_1079_413#_c_1450_n 0.00421051f $X=7.585
+ $Y=1.68 $X2=0 $Y2=0
cc_874 N_A_1245_303#_c_1170_n N_A_1592_47#_c_1779_n 0.0254084f $X=8.055 $Y=2.3
+ $X2=0 $Y2=0
cc_875 N_A_1245_303#_c_1171_n N_VPWR_M1021_s 0.00330649f $X=7.585 $Y=1.68 $X2=0
+ $Y2=0
cc_876 N_A_1245_303#_c_1167_n N_VPWR_c_1895_n 0.00180429f $X=7.455 $Y=1.68 $X2=0
+ $Y2=0
cc_877 N_A_1245_303#_c_1169_n N_VPWR_c_1895_n 5.6212e-19 $X=7.97 $Y=1.92 $X2=0
+ $Y2=0
cc_878 N_A_1245_303#_c_1170_n N_VPWR_c_1895_n 0.0174112f $X=8.055 $Y=2.3 $X2=0
+ $Y2=0
cc_879 N_A_1245_303#_c_1171_n N_VPWR_c_1895_n 0.0173472f $X=7.585 $Y=1.68 $X2=0
+ $Y2=0
cc_880 N_A_1245_303#_M1038_g N_VPWR_c_1905_n 0.0039846f $X=6.3 $Y=2.275 $X2=0
+ $Y2=0
cc_881 N_A_1245_303#_M1038_g N_VPWR_c_1906_n 0.00422112f $X=6.3 $Y=2.275 $X2=0
+ $Y2=0
cc_882 N_A_1245_303#_c_1169_n N_VPWR_c_1910_n 0.00276762f $X=7.97 $Y=1.92 $X2=0
+ $Y2=0
cc_883 N_A_1245_303#_c_1170_n N_VPWR_c_1910_n 0.0117479f $X=8.055 $Y=2.3 $X2=0
+ $Y2=0
cc_884 N_A_1245_303#_M1021_d N_VPWR_c_1891_n 0.00287843f $X=7.885 $Y=1.645 $X2=0
+ $Y2=0
cc_885 N_A_1245_303#_M1038_g N_VPWR_c_1891_n 0.00581106f $X=6.3 $Y=2.275 $X2=0
+ $Y2=0
cc_886 N_A_1245_303#_c_1169_n N_VPWR_c_1891_n 0.00231913f $X=7.97 $Y=1.92 $X2=0
+ $Y2=0
cc_887 N_A_1245_303#_c_1170_n N_VPWR_c_1891_n 0.00306902f $X=8.055 $Y=2.3 $X2=0
+ $Y2=0
cc_888 N_A_1245_303#_c_1171_n N_VPWR_c_1891_n 7.10368e-19 $X=7.585 $Y=1.68 $X2=0
+ $Y2=0
cc_889 N_A_1245_303#_M1038_g N_A_1191_413#_c_2203_n 0.010597f $X=6.3 $Y=2.275
+ $X2=0 $Y2=0
cc_890 N_A_1245_303#_c_1167_n N_A_1191_413#_c_2203_n 0.0437915f $X=7.455 $Y=1.68
+ $X2=0 $Y2=0
cc_891 N_A_1245_303#_c_1168_n N_A_1191_413#_c_2203_n 0.00427615f $X=6.45 $Y=1.68
+ $X2=0 $Y2=0
cc_892 N_A_1245_303#_M1038_g N_A_1191_413#_c_2204_n 2.60163e-19 $X=6.3 $Y=2.275
+ $X2=0 $Y2=0
cc_893 N_A_1245_303#_c_1167_n N_A_1191_413#_c_2205_n 0.011083f $X=7.455 $Y=1.68
+ $X2=0 $Y2=0
cc_894 N_A_1245_303#_c_1171_n N_A_1191_413#_c_2205_n 0.0037013f $X=7.585 $Y=1.68
+ $X2=0 $Y2=0
cc_895 N_A_1245_303#_c_1214_p N_VGND_c_2282_n 0.0176707f $X=7.62 $Y=0.36 $X2=0
+ $Y2=0
cc_896 N_A_1245_303#_c_1214_p N_VGND_c_2289_n 0.0174179f $X=7.62 $Y=0.36 $X2=0
+ $Y2=0
cc_897 N_A_1245_303#_M1010_g N_VGND_c_2299_n 0.0055639f $X=6.39 $Y=0.445 $X2=0
+ $Y2=0
cc_898 N_A_1245_303#_M1039_d N_VGND_c_2301_n 0.00233415f $X=7.485 $Y=0.235 $X2=0
+ $Y2=0
cc_899 N_A_1245_303#_M1010_g N_VGND_c_2301_n 0.00962524f $X=6.39 $Y=0.445 $X2=0
+ $Y2=0
cc_900 N_A_1245_303#_c_1214_p N_VGND_c_2301_n 0.00575387f $X=7.62 $Y=0.36 $X2=0
+ $Y2=0
cc_901 N_RESET_B_c_1281_n N_A_1079_413#_M1039_g 0.00165023f $X=6.95 $Y=0.85
+ $X2=0 $Y2=0
cc_902 N_RESET_B_c_1282_n N_A_1079_413#_M1039_g 0.00521008f $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_903 N_RESET_B_c_1283_n N_A_1079_413#_M1039_g 0.00169797f $X=7.095 $Y=0.85
+ $X2=0 $Y2=0
cc_904 N_RESET_B_c_1285_n N_A_1079_413#_M1039_g 0.00740135f $X=6.81 $Y=0.96
+ $X2=0 $Y2=0
cc_905 N_RESET_B_c_1286_n N_A_1079_413#_M1039_g 0.0127085f $X=6.81 $Y=0.755
+ $X2=0 $Y2=0
cc_906 N_RESET_B_c_1286_n N_A_1079_413#_c_1479_n 4.85263e-19 $X=6.81 $Y=0.755
+ $X2=0 $Y2=0
cc_907 N_RESET_B_M1033_g N_A_1079_413#_c_1447_n 6.06578e-19 $X=6.87 $Y=2.275
+ $X2=0 $Y2=0
cc_908 N_RESET_B_c_1280_n N_A_1079_413#_c_1447_n 0.0076355f $X=6.98 $Y=0.85
+ $X2=0 $Y2=0
cc_909 N_RESET_B_c_1281_n N_A_1079_413#_c_1447_n 0.0189574f $X=6.95 $Y=0.85
+ $X2=0 $Y2=0
cc_910 N_RESET_B_c_1285_n N_A_1079_413#_c_1447_n 6.48617e-19 $X=6.81 $Y=0.96
+ $X2=0 $Y2=0
cc_911 N_RESET_B_c_1286_n N_A_1079_413#_c_1447_n 0.0012881f $X=6.81 $Y=0.755
+ $X2=0 $Y2=0
cc_912 N_RESET_B_M1033_g N_A_1079_413#_c_1448_n 0.00965887f $X=6.87 $Y=2.275
+ $X2=0 $Y2=0
cc_913 N_RESET_B_c_1280_n N_A_1079_413#_c_1448_n 0.00106869f $X=6.98 $Y=0.85
+ $X2=0 $Y2=0
cc_914 N_RESET_B_c_1281_n N_A_1079_413#_c_1448_n 0.0343562f $X=6.95 $Y=0.85
+ $X2=0 $Y2=0
cc_915 N_RESET_B_c_1282_n N_A_1079_413#_c_1448_n 5.4481e-19 $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_916 N_RESET_B_c_1283_n N_A_1079_413#_c_1448_n 2.36449e-19 $X=7.095 $Y=0.85
+ $X2=0 $Y2=0
cc_917 N_RESET_B_c_1285_n N_A_1079_413#_c_1448_n 0.00251038f $X=6.81 $Y=0.96
+ $X2=0 $Y2=0
cc_918 N_RESET_B_c_1281_n N_A_1079_413#_c_1449_n 0.00314358f $X=6.95 $Y=0.85
+ $X2=0 $Y2=0
cc_919 N_RESET_B_c_1282_n N_A_1079_413#_c_1449_n 0.0042685f $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_920 N_RESET_B_c_1285_n N_A_1079_413#_c_1449_n 0.00140529f $X=6.81 $Y=0.96
+ $X2=0 $Y2=0
cc_921 N_RESET_B_M1033_g N_A_1079_413#_c_1450_n 0.00817494f $X=6.87 $Y=2.275
+ $X2=0 $Y2=0
cc_922 N_RESET_B_c_1281_n N_A_1079_413#_c_1450_n 2.62214e-19 $X=6.95 $Y=0.85
+ $X2=0 $Y2=0
cc_923 N_RESET_B_c_1282_n N_A_1079_413#_c_1450_n 8.21109e-19 $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_924 N_RESET_B_c_1285_n N_A_1079_413#_c_1450_n 0.0219099f $X=6.81 $Y=0.96
+ $X2=0 $Y2=0
cc_925 N_RESET_B_M1000_g N_A_1767_21#_M1027_g 0.00832425f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_926 N_RESET_B_c_1282_n N_A_1767_21#_M1027_g 0.00153944f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_927 N_RESET_B_c_1276_n N_A_1767_21#_M1028_g 0.0473681f $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_928 N_RESET_B_c_1291_n N_A_1767_21#_M1028_g 0.0129297f $X=9.655 $Y=1.99 $X2=0
+ $Y2=0
cc_929 RESET_B N_A_1767_21#_M1028_g 0.00108111f $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_930 N_RESET_B_c_1276_n N_A_1767_21#_c_1589_n 3.89491e-19 $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_931 N_RESET_B_M1000_g N_A_1767_21#_c_1589_n 4.36318e-19 $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_932 RESET_B N_A_1767_21#_c_1589_n 0.00458036f $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_933 RESET_B N_A_1767_21#_c_1589_n 0.00341948f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_934 N_RESET_B_c_1282_n N_A_1767_21#_c_1589_n 0.00784735f $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_935 N_RESET_B_c_1284_n N_A_1767_21#_c_1589_n 0.0038541f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_936 N_RESET_B_c_1276_n N_A_1767_21#_c_1590_n 0.00387868f $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_937 N_RESET_B_M1000_g N_A_1767_21#_c_1590_n 0.0052827f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_938 RESET_B N_A_1767_21#_c_1590_n 0.00699765f $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_939 RESET_B N_A_1767_21#_c_1590_n 0.0124998f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_940 N_RESET_B_c_1282_n N_A_1767_21#_c_1590_n 0.0155247f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_941 N_RESET_B_c_1284_n N_A_1767_21#_c_1590_n 0.00226386f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_942 N_RESET_B_c_1282_n N_A_1767_21#_c_1591_n 0.00535772f $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_943 N_RESET_B_M1000_g N_A_1767_21#_c_1592_n 0.00686702f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_944 RESET_B N_A_1767_21#_c_1592_n 0.00441838f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_945 N_RESET_B_c_1276_n N_A_1767_21#_c_1593_n 8.95506e-19 $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_946 N_RESET_B_M1000_g N_A_1767_21#_c_1593_n 0.00556598f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_947 RESET_B N_A_1767_21#_c_1593_n 0.00153156f $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_948 RESET_B N_A_1767_21#_c_1593_n 0.0158276f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_949 N_RESET_B_c_1284_n N_A_1767_21#_c_1593_n 0.00476196f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_950 N_RESET_B_M1000_g N_A_1767_21#_c_1643_n 0.00391955f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_951 N_RESET_B_c_1292_n N_A_1767_21#_c_1605_n 0.0023084f $X=9.485 $Y=1.915
+ $X2=0 $Y2=0
cc_952 RESET_B N_A_1767_21#_c_1594_n 0.0177987f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_953 N_RESET_B_c_1284_n N_A_1767_21#_c_1594_n 0.00664316f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_954 RESET_B N_A_1767_21#_c_1596_n 0.00418829f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_955 N_RESET_B_c_1284_n N_A_1767_21#_c_1596_n 0.00288016f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_956 N_RESET_B_c_1287_n N_A_1767_21#_c_1596_n 0.0134093f $X=9.97 $Y=1.065
+ $X2=0 $Y2=0
cc_957 N_RESET_B_c_1276_n N_A_1767_21#_c_1597_n 0.0099528f $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_958 N_RESET_B_M1000_g N_A_1767_21#_c_1597_n 0.00976572f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_959 RESET_B N_A_1767_21#_c_1597_n 5.30274e-19 $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_960 N_RESET_B_c_1282_n N_A_1767_21#_c_1597_n 0.00565059f $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_961 N_RESET_B_c_1284_n N_A_1767_21#_c_1597_n 7.74628e-19 $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_962 N_RESET_B_M1000_g N_A_1592_47#_c_1773_n 0.0390661f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_963 RESET_B N_A_1592_47#_c_1773_n 0.00836902f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_964 N_RESET_B_c_1284_n N_A_1592_47#_c_1773_n 0.00134454f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_965 N_RESET_B_c_1290_n N_A_1592_47#_c_1776_n 0.0123371f $X=9.485 $Y=1.84
+ $X2=0 $Y2=0
cc_966 N_RESET_B_c_1284_n N_A_1592_47#_c_1776_n 4.36744e-19 $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_967 N_RESET_B_c_1287_n N_A_1592_47#_c_1776_n 0.00239709f $X=9.97 $Y=1.065
+ $X2=0 $Y2=0
cc_968 N_RESET_B_c_1290_n N_A_1592_47#_M1032_g 4.71931e-19 $X=9.485 $Y=1.84
+ $X2=0 $Y2=0
cc_969 N_RESET_B_c_1292_n N_A_1592_47#_M1032_g 0.019999f $X=9.485 $Y=1.915 $X2=0
+ $Y2=0
cc_970 N_RESET_B_c_1276_n N_A_1592_47#_c_1774_n 0.0263312f $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_971 N_RESET_B_c_1290_n N_A_1592_47#_c_1774_n 0.00185333f $X=9.485 $Y=1.84
+ $X2=0 $Y2=0
cc_972 N_RESET_B_M1000_g N_A_1592_47#_c_1774_n 0.0057628f $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_973 RESET_B N_A_1592_47#_c_1774_n 0.00464867f $X=9.945 $Y=0.765 $X2=0 $Y2=0
cc_974 N_RESET_B_c_1284_n N_A_1592_47#_c_1774_n 0.00238942f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_975 N_RESET_B_c_1287_n N_A_1592_47#_c_1774_n 0.00672376f $X=9.97 $Y=1.065
+ $X2=0 $Y2=0
cc_976 N_RESET_B_c_1282_n N_A_1592_47#_c_1783_n 0.0165715f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_977 N_RESET_B_c_1291_n N_A_1592_47#_c_1779_n 5.9045e-19 $X=9.655 $Y=1.99
+ $X2=0 $Y2=0
cc_978 N_RESET_B_M1000_g N_A_1592_47#_c_1775_n 2.70549e-19 $X=9.655 $Y=0.445
+ $X2=0 $Y2=0
cc_979 RESET_B N_A_1592_47#_c_1775_n 0.00424344f $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_980 N_RESET_B_c_1282_n N_A_1592_47#_c_1775_n 0.0214607f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_981 N_RESET_B_c_1290_n N_A_1592_47#_c_1780_n 0.00393349f $X=9.485 $Y=1.84
+ $X2=0 $Y2=0
cc_982 N_RESET_B_c_1291_n N_A_1592_47#_c_1780_n 3.26213e-19 $X=9.655 $Y=1.99
+ $X2=0 $Y2=0
cc_983 N_RESET_B_c_1276_n N_A_1592_47#_c_1781_n 0.00577456f $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_984 N_RESET_B_c_1282_n N_A_1592_47#_c_1781_n 0.00757576f $X=9.63 $Y=0.85
+ $X2=0 $Y2=0
cc_985 N_RESET_B_c_1276_n N_A_1592_47#_c_1782_n 0.00380276f $X=9.485 $Y=1.435
+ $X2=0 $Y2=0
cc_986 N_RESET_B_c_1290_n N_A_1592_47#_c_1782_n 0.0141248f $X=9.485 $Y=1.84
+ $X2=0 $Y2=0
cc_987 N_RESET_B_c_1292_n N_A_1592_47#_c_1782_n 0.00383937f $X=9.485 $Y=1.915
+ $X2=0 $Y2=0
cc_988 RESET_B N_A_1592_47#_c_1782_n 0.0114108f $X=9.825 $Y=1.105 $X2=0 $Y2=0
cc_989 N_RESET_B_c_1284_n N_A_1592_47#_c_1782_n 0.0101861f $X=9.775 $Y=0.965
+ $X2=0 $Y2=0
cc_990 N_RESET_B_c_1287_n N_A_1592_47#_c_1782_n 0.0127161f $X=9.97 $Y=1.065
+ $X2=0 $Y2=0
cc_991 N_RESET_B_M1033_g N_VPWR_c_1895_n 0.00347183f $X=6.87 $Y=2.275 $X2=0
+ $Y2=0
cc_992 N_RESET_B_c_1291_n N_VPWR_c_1896_n 0.00798618f $X=9.655 $Y=1.99 $X2=0
+ $Y2=0
cc_993 N_RESET_B_c_1292_n N_VPWR_c_1896_n 0.00452506f $X=9.485 $Y=1.915 $X2=0
+ $Y2=0
cc_994 N_RESET_B_c_1291_n N_VPWR_c_1897_n 7.21572e-19 $X=9.655 $Y=1.99 $X2=0
+ $Y2=0
cc_995 N_RESET_B_M1033_g N_VPWR_c_1905_n 0.00246816f $X=6.87 $Y=2.275 $X2=0
+ $Y2=0
cc_996 N_RESET_B_M1033_g N_VPWR_c_1909_n 0.00422112f $X=6.87 $Y=2.275 $X2=0
+ $Y2=0
cc_997 N_RESET_B_c_1291_n N_VPWR_c_1911_n 0.00466271f $X=9.655 $Y=1.99 $X2=0
+ $Y2=0
cc_998 N_RESET_B_M1033_g N_VPWR_c_1891_n 0.00721006f $X=6.87 $Y=2.275 $X2=0
+ $Y2=0
cc_999 N_RESET_B_c_1291_n N_VPWR_c_1891_n 0.00794889f $X=9.655 $Y=1.99 $X2=0
+ $Y2=0
cc_1000 N_RESET_B_M1033_g N_A_1191_413#_c_2203_n 0.0114021f $X=6.87 $Y=2.275
+ $X2=0 $Y2=0
cc_1001 N_RESET_B_M1033_g N_A_1191_413#_c_2205_n 0.00120854f $X=6.87 $Y=2.275
+ $X2=0 $Y2=0
cc_1002 N_RESET_B_c_1282_n N_VGND_M1013_d 0.00246367f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_1003 N_RESET_B_c_1283_n N_VGND_M1013_d 5.87293e-19 $X=7.095 $Y=0.85 $X2=0
+ $Y2=0
cc_1004 N_RESET_B_c_1280_n N_VGND_c_2282_n 0.00262628f $X=6.98 $Y=0.85 $X2=0
+ $Y2=0
cc_1005 N_RESET_B_c_1281_n N_VGND_c_2282_n 0.00640958f $X=6.95 $Y=0.85 $X2=0
+ $Y2=0
cc_1006 N_RESET_B_c_1282_n N_VGND_c_2282_n 0.0025629f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_1007 N_RESET_B_c_1285_n N_VGND_c_2282_n 5.41848e-19 $X=6.81 $Y=0.96 $X2=0
+ $Y2=0
cc_1008 N_RESET_B_c_1286_n N_VGND_c_2282_n 0.00852416f $X=6.81 $Y=0.755 $X2=0
+ $Y2=0
cc_1009 N_RESET_B_M1000_g N_VGND_c_2283_n 0.00368378f $X=9.655 $Y=0.445 $X2=0
+ $Y2=0
cc_1010 N_RESET_B_c_1282_n N_VGND_c_2283_n 0.0018919f $X=9.63 $Y=0.85 $X2=0
+ $Y2=0
cc_1011 N_RESET_B_M1000_g N_VGND_c_2291_n 0.0036601f $X=9.655 $Y=0.445 $X2=0
+ $Y2=0
cc_1012 N_RESET_B_c_1285_n N_VGND_c_2299_n 0.00111174f $X=6.81 $Y=0.96 $X2=0
+ $Y2=0
cc_1013 N_RESET_B_c_1286_n N_VGND_c_2299_n 0.00585385f $X=6.81 $Y=0.755 $X2=0
+ $Y2=0
cc_1014 N_RESET_B_M1000_g N_VGND_c_2301_n 0.00584295f $X=9.655 $Y=0.445 $X2=0
+ $Y2=0
cc_1015 N_RESET_B_c_1280_n N_VGND_c_2301_n 0.0354525f $X=6.98 $Y=0.85 $X2=0
+ $Y2=0
cc_1016 N_RESET_B_c_1281_n N_VGND_c_2301_n 0.00441112f $X=6.95 $Y=0.85 $X2=0
+ $Y2=0
cc_1017 N_RESET_B_c_1282_n N_VGND_c_2301_n 0.134033f $X=9.63 $Y=0.85 $X2=0 $Y2=0
cc_1018 N_RESET_B_c_1284_n N_VGND_c_2301_n 0.0147031f $X=9.775 $Y=0.965 $X2=0
+ $Y2=0
cc_1019 N_RESET_B_c_1285_n N_VGND_c_2301_n 5.47414e-19 $X=6.81 $Y=0.96 $X2=0
+ $Y2=0
cc_1020 N_RESET_B_c_1286_n N_VGND_c_2301_n 0.0060657f $X=6.81 $Y=0.755 $X2=0
+ $Y2=0
cc_1021 RESET_B A_1946_47# 0.00114648f $X=9.945 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_1022 N_A_1079_413#_c_1451_n N_VPWR_c_1895_n 5.04979e-19 $X=7.735 $Y=1.495
+ $X2=0 $Y2=0
cc_1023 N_A_1079_413#_c_1452_n N_VPWR_c_1895_n 0.00902097f $X=7.81 $Y=1.57 $X2=0
+ $Y2=0
cc_1024 N_A_1079_413#_c_1450_n N_VPWR_c_1895_n 4.01326e-19 $X=7.29 $Y=1.17 $X2=0
+ $Y2=0
cc_1025 N_A_1079_413#_c_1467_n N_VPWR_c_1906_n 0.0227585f $X=5.67 $Y=2.33 $X2=0
+ $Y2=0
cc_1026 N_A_1079_413#_c_1452_n N_VPWR_c_1910_n 0.00406603f $X=7.81 $Y=1.57 $X2=0
+ $Y2=0
cc_1027 N_A_1079_413#_M1007_d N_VPWR_c_1891_n 0.00289429f $X=5.395 $Y=2.065
+ $X2=0 $Y2=0
cc_1028 N_A_1079_413#_c_1452_n N_VPWR_c_1891_n 0.00451526f $X=7.81 $Y=1.57 $X2=0
+ $Y2=0
cc_1029 N_A_1079_413#_c_1467_n N_VPWR_c_1891_n 0.00635687f $X=5.67 $Y=2.33 $X2=0
+ $Y2=0
cc_1030 N_A_1079_413#_c_1467_n N_A_620_389#_c_2099_n 0.019896f $X=5.67 $Y=2.33
+ $X2=0 $Y2=0
cc_1031 N_A_1079_413#_c_1455_n N_A_620_389#_c_2099_n 0.00532808f $X=5.652
+ $Y=2.135 $X2=0 $Y2=0
cc_1032 N_A_1079_413#_c_1456_n N_A_1191_413#_c_2203_n 0.00204762f $X=6.25 $Y=1.3
+ $X2=0 $Y2=0
cc_1033 N_A_1079_413#_c_1445_n N_A_1191_413#_c_2204_n 0.00297929f $X=6.165
+ $Y=1.3 $X2=0 $Y2=0
cc_1034 N_A_1079_413#_c_1455_n N_A_1191_413#_c_2204_n 0.0205809f $X=5.652
+ $Y=2.135 $X2=0 $Y2=0
cc_1035 N_A_1079_413#_c_1452_n N_A_1191_413#_c_2205_n 0.00351626f $X=7.81
+ $Y=1.57 $X2=0 $Y2=0
cc_1036 N_A_1079_413#_M1039_g N_VGND_c_2282_n 0.00677972f $X=7.41 $Y=0.555 $X2=0
+ $Y2=0
cc_1037 N_A_1079_413#_c_1479_n N_VGND_c_2282_n 0.00530482f $X=6.165 $Y=0.39
+ $X2=0 $Y2=0
cc_1038 N_A_1079_413#_c_1447_n N_VGND_c_2282_n 0.00196456f $X=6.25 $Y=1.215
+ $X2=0 $Y2=0
cc_1039 N_A_1079_413#_c_1448_n N_VGND_c_2282_n 0.0020619f $X=7.205 $Y=1.3 $X2=0
+ $Y2=0
cc_1040 N_A_1079_413#_c_1449_n N_VGND_c_2282_n 6.81471e-19 $X=7.29 $Y=1.17 $X2=0
+ $Y2=0
cc_1041 N_A_1079_413#_c_1450_n N_VGND_c_2282_n 0.00132464f $X=7.29 $Y=1.17 $X2=0
+ $Y2=0
cc_1042 N_A_1079_413#_M1039_g N_VGND_c_2289_n 0.00542163f $X=7.41 $Y=0.555 $X2=0
+ $Y2=0
cc_1043 N_A_1079_413#_c_1479_n N_VGND_c_2299_n 0.0374514f $X=6.165 $Y=0.39 $X2=0
+ $Y2=0
cc_1044 N_A_1079_413#_M1023_d N_VGND_c_2301_n 0.0030735f $X=5.435 $Y=0.235 $X2=0
+ $Y2=0
cc_1045 N_A_1079_413#_M1039_g N_VGND_c_2301_n 0.00682459f $X=7.41 $Y=0.555 $X2=0
+ $Y2=0
cc_1046 N_A_1079_413#_c_1479_n N_VGND_c_2301_n 0.0300684f $X=6.165 $Y=0.39 $X2=0
+ $Y2=0
cc_1047 N_A_1079_413#_c_1479_n A_1187_47# 0.00955634f $X=6.165 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_1048 N_A_1079_413#_c_1447_n A_1187_47# 0.00216963f $X=6.25 $Y=1.215 $X2=-0.19
+ $Y2=-0.24
cc_1049 N_A_1767_21#_c_1592_n N_A_1592_47#_c_1773_n 9.88157e-19 $X=9.57 $Y=0.695
+ $X2=0 $Y2=0
cc_1050 N_A_1767_21#_c_1593_n N_A_1592_47#_c_1773_n 0.00903189f $X=10.345
+ $Y=0.38 $X2=0 $Y2=0
cc_1051 N_A_1767_21#_c_1594_n N_A_1592_47#_c_1773_n 0.0109288f $X=10.43 $Y=0.995
+ $X2=0 $Y2=0
cc_1052 N_A_1767_21#_c_1604_n N_A_1592_47#_c_1776_n 0.00224286f $X=10.375 $Y=2
+ $X2=0 $Y2=0
cc_1053 N_A_1767_21#_c_1605_n N_A_1592_47#_c_1776_n 0.00113085f $X=9.95 $Y=2
+ $X2=0 $Y2=0
cc_1054 N_A_1767_21#_c_1606_n N_A_1592_47#_c_1776_n 0.00403767f $X=10.46
+ $Y=1.915 $X2=0 $Y2=0
cc_1055 N_A_1767_21#_c_1604_n N_A_1592_47#_M1032_g 0.0124008f $X=10.375 $Y=2
+ $X2=0 $Y2=0
cc_1056 N_A_1767_21#_c_1606_n N_A_1592_47#_M1032_g 0.00287205f $X=10.46 $Y=1.915
+ $X2=0 $Y2=0
cc_1057 N_A_1767_21#_c_1606_n N_A_1592_47#_c_1774_n 0.00857906f $X=10.46
+ $Y=1.915 $X2=0 $Y2=0
cc_1058 N_A_1767_21#_c_1596_n N_A_1592_47#_c_1774_n 0.00447556f $X=10.345
+ $Y=0.995 $X2=0 $Y2=0
cc_1059 N_A_1767_21#_c_1598_n N_A_1592_47#_c_1774_n 0.00392382f $X=12.285
+ $Y=1.16 $X2=0 $Y2=0
cc_1060 N_A_1767_21#_M1027_g N_A_1592_47#_c_1783_n 0.00850482f $X=8.91 $Y=0.445
+ $X2=0 $Y2=0
cc_1061 N_A_1767_21#_c_1592_n N_A_1592_47#_c_1783_n 3.02597e-19 $X=9.57 $Y=0.695
+ $X2=0 $Y2=0
cc_1062 N_A_1767_21#_M1028_g N_A_1592_47#_c_1779_n 0.0139696f $X=9.125 $Y=2.275
+ $X2=0 $Y2=0
cc_1063 N_A_1767_21#_c_1605_n N_A_1592_47#_c_1779_n 0.00105649f $X=9.95 $Y=2
+ $X2=0 $Y2=0
cc_1064 N_A_1767_21#_M1027_g N_A_1592_47#_c_1775_n 0.00726792f $X=8.91 $Y=0.445
+ $X2=0 $Y2=0
cc_1065 N_A_1767_21#_c_1589_n N_A_1592_47#_c_1775_n 0.0161233f $X=9.21 $Y=0.98
+ $X2=0 $Y2=0
cc_1066 N_A_1767_21#_c_1591_n N_A_1592_47#_c_1775_n 0.0102727f $X=9.295 $Y=0.78
+ $X2=0 $Y2=0
cc_1067 N_A_1767_21#_c_1592_n N_A_1592_47#_c_1775_n 0.00439089f $X=9.57 $Y=0.695
+ $X2=0 $Y2=0
cc_1068 N_A_1767_21#_c_1597_n N_A_1592_47#_c_1775_n 0.00963909f $X=9.125 $Y=0.98
+ $X2=0 $Y2=0
cc_1069 N_A_1767_21#_M1028_g N_A_1592_47#_c_1780_n 0.00520507f $X=9.125 $Y=2.275
+ $X2=0 $Y2=0
cc_1070 N_A_1767_21#_c_1605_n N_A_1592_47#_c_1780_n 0.00429874f $X=9.95 $Y=2
+ $X2=0 $Y2=0
cc_1071 N_A_1767_21#_M1028_g N_A_1592_47#_c_1781_n 0.0146012f $X=9.125 $Y=2.275
+ $X2=0 $Y2=0
cc_1072 N_A_1767_21#_c_1589_n N_A_1592_47#_c_1781_n 0.00658052f $X=9.21 $Y=0.98
+ $X2=0 $Y2=0
cc_1073 N_A_1767_21#_c_1597_n N_A_1592_47#_c_1781_n 0.0043817f $X=9.125 $Y=0.98
+ $X2=0 $Y2=0
cc_1074 N_A_1767_21#_c_1589_n N_A_1592_47#_c_1782_n 0.00321233f $X=9.21 $Y=0.98
+ $X2=0 $Y2=0
cc_1075 N_A_1767_21#_c_1604_n N_A_1592_47#_c_1782_n 0.0177144f $X=10.375 $Y=2
+ $X2=0 $Y2=0
cc_1076 N_A_1767_21#_c_1605_n N_A_1592_47#_c_1782_n 0.0134553f $X=9.95 $Y=2
+ $X2=0 $Y2=0
cc_1077 N_A_1767_21#_c_1606_n N_A_1592_47#_c_1782_n 0.014187f $X=10.46 $Y=1.915
+ $X2=0 $Y2=0
cc_1078 N_A_1767_21#_c_1597_n N_A_1592_47#_c_1782_n 0.00192646f $X=9.125 $Y=0.98
+ $X2=0 $Y2=0
cc_1079 N_A_1767_21#_c_1604_n N_VPWR_M1032_d 0.00216549f $X=10.375 $Y=2 $X2=0
+ $Y2=0
cc_1080 N_A_1767_21#_M1028_g N_VPWR_c_1896_n 0.0046608f $X=9.125 $Y=2.275 $X2=0
+ $Y2=0
cc_1081 N_A_1767_21#_M1002_g N_VPWR_c_1897_n 9.67101e-19 $X=11.015 $Y=1.985
+ $X2=0 $Y2=0
cc_1082 N_A_1767_21#_c_1604_n N_VPWR_c_1897_n 0.0211796f $X=10.375 $Y=2 $X2=0
+ $Y2=0
cc_1083 N_A_1767_21#_c_1604_n N_VPWR_c_1898_n 0.0019191f $X=10.375 $Y=2 $X2=0
+ $Y2=0
cc_1084 N_A_1767_21#_M1002_g N_VPWR_c_1899_n 0.0168807f $X=11.015 $Y=1.985 $X2=0
+ $Y2=0
cc_1085 N_A_1767_21#_M1008_g N_VPWR_c_1899_n 0.00118718f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_1086 N_A_1767_21#_c_1604_n N_VPWR_c_1899_n 0.0141976f $X=10.375 $Y=2 $X2=0
+ $Y2=0
cc_1087 N_A_1767_21#_c_1606_n N_VPWR_c_1899_n 0.0312704f $X=10.46 $Y=1.915 $X2=0
+ $Y2=0
cc_1088 N_A_1767_21#_c_1595_n N_VPWR_c_1899_n 0.0181245f $X=10.935 $Y=1.16 $X2=0
+ $Y2=0
cc_1089 N_A_1767_21#_c_1598_n N_VPWR_c_1899_n 0.00308771f $X=12.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1090 N_A_1767_21#_M1008_g N_VPWR_c_1900_n 0.00528569f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_1091 N_A_1767_21#_M1024_g N_VPWR_c_1900_n 0.0155769f $X=11.865 $Y=1.985 $X2=0
+ $Y2=0
cc_1092 N_A_1767_21#_M1034_g N_VPWR_c_1900_n 0.00118f $X=12.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1093 N_A_1767_21#_c_1598_n N_VPWR_c_1900_n 0.00232957f $X=12.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1094 N_A_1767_21#_M1034_g N_VPWR_c_1902_n 0.00311793f $X=12.285 $Y=1.985
+ $X2=0 $Y2=0
cc_1095 N_A_1767_21#_M1028_g N_VPWR_c_1910_n 0.00361853f $X=9.125 $Y=2.275 $X2=0
+ $Y2=0
cc_1096 N_A_1767_21#_c_1702_p N_VPWR_c_1911_n 0.00701792f $X=9.865 $Y=2.21 $X2=0
+ $Y2=0
cc_1097 N_A_1767_21#_c_1604_n N_VPWR_c_1911_n 0.00243651f $X=10.375 $Y=2 $X2=0
+ $Y2=0
cc_1098 N_A_1767_21#_M1002_g N_VPWR_c_1912_n 0.0046653f $X=11.015 $Y=1.985 $X2=0
+ $Y2=0
cc_1099 N_A_1767_21#_M1008_g N_VPWR_c_1912_n 0.00533345f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_1100 N_A_1767_21#_M1024_g N_VPWR_c_1913_n 0.0046653f $X=11.865 $Y=1.985 $X2=0
+ $Y2=0
cc_1101 N_A_1767_21#_M1034_g N_VPWR_c_1913_n 0.00546688f $X=12.285 $Y=1.985
+ $X2=0 $Y2=0
cc_1102 N_A_1767_21#_M1012_d N_VPWR_c_1891_n 0.00416801f $X=9.73 $Y=2.065 $X2=0
+ $Y2=0
cc_1103 N_A_1767_21#_M1028_g N_VPWR_c_1891_n 0.00558649f $X=9.125 $Y=2.275 $X2=0
+ $Y2=0
cc_1104 N_A_1767_21#_M1002_g N_VPWR_c_1891_n 0.00796766f $X=11.015 $Y=1.985
+ $X2=0 $Y2=0
cc_1105 N_A_1767_21#_M1008_g N_VPWR_c_1891_n 0.00925272f $X=11.435 $Y=1.985
+ $X2=0 $Y2=0
cc_1106 N_A_1767_21#_M1024_g N_VPWR_c_1891_n 0.00796766f $X=11.865 $Y=1.985
+ $X2=0 $Y2=0
cc_1107 N_A_1767_21#_M1034_g N_VPWR_c_1891_n 0.0106176f $X=12.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1108 N_A_1767_21#_c_1702_p N_VPWR_c_1891_n 0.00608739f $X=9.865 $Y=2.21 $X2=0
+ $Y2=0
cc_1109 N_A_1767_21#_c_1604_n N_VPWR_c_1891_n 0.0086292f $X=10.375 $Y=2 $X2=0
+ $Y2=0
cc_1110 N_A_1767_21#_c_1585_n N_Q_c_2236_n 0.00232137f $X=11.015 $Y=0.995 $X2=0
+ $Y2=0
cc_1111 N_A_1767_21#_c_1586_n N_Q_c_2236_n 0.00514965f $X=11.435 $Y=0.995 $X2=0
+ $Y2=0
cc_1112 N_A_1767_21#_c_1594_n N_Q_c_2236_n 0.00559463f $X=10.43 $Y=0.995 $X2=0
+ $Y2=0
cc_1113 N_A_1767_21#_c_1598_n N_Q_c_2243_n 0.0598347f $X=12.285 $Y=1.16 $X2=0
+ $Y2=0
cc_1114 N_A_1767_21#_c_1587_n N_Q_c_2237_n 0.00235233f $X=11.865 $Y=0.995 $X2=0
+ $Y2=0
cc_1115 N_A_1767_21#_c_1588_n N_Q_c_2237_n 0.0253792f $X=12.285 $Y=0.995 $X2=0
+ $Y2=0
cc_1116 N_A_1767_21#_M1024_g N_Q_c_2238_n 0.00262852f $X=11.865 $Y=1.985 $X2=0
+ $Y2=0
cc_1117 N_A_1767_21#_M1034_g N_Q_c_2238_n 0.0193386f $X=12.285 $Y=1.985 $X2=0
+ $Y2=0
cc_1118 N_A_1767_21#_c_1586_n N_Q_c_2248_n 0.00252307f $X=11.435 $Y=0.995 $X2=0
+ $Y2=0
cc_1119 N_A_1767_21#_c_1598_n N_Q_c_2248_n 2.81601e-19 $X=12.285 $Y=1.16 $X2=0
+ $Y2=0
cc_1120 N_A_1767_21#_c_1598_n N_Q_c_2250_n 0.0269648f $X=12.285 $Y=1.16 $X2=0
+ $Y2=0
cc_1121 N_A_1767_21#_c_1586_n Q 0.00727483f $X=11.435 $Y=0.995 $X2=0 $Y2=0
cc_1122 N_A_1767_21#_c_1587_n Q 0.001414f $X=11.865 $Y=0.995 $X2=0 $Y2=0
cc_1123 N_A_1767_21#_M1008_g Q 0.00901955f $X=11.435 $Y=1.985 $X2=0 $Y2=0
cc_1124 N_A_1767_21#_M1002_g N_Q_c_2239_n 0.00238466f $X=11.015 $Y=1.985 $X2=0
+ $Y2=0
cc_1125 N_A_1767_21#_M1008_g N_Q_c_2239_n 0.00655045f $X=11.435 $Y=1.985 $X2=0
+ $Y2=0
cc_1126 N_A_1767_21#_M1024_g N_Q_c_2239_n 5.05521e-19 $X=11.865 $Y=1.985 $X2=0
+ $Y2=0
cc_1127 N_A_1767_21#_c_1606_n N_Q_c_2239_n 0.00499908f $X=10.46 $Y=1.915 $X2=0
+ $Y2=0
cc_1128 N_A_1767_21#_c_1595_n N_Q_c_2239_n 0.0277414f $X=10.935 $Y=1.16 $X2=0
+ $Y2=0
cc_1129 N_A_1767_21#_c_1598_n N_Q_c_2239_n 0.0155237f $X=12.285 $Y=1.16 $X2=0
+ $Y2=0
cc_1130 N_A_1767_21#_c_1592_n N_VGND_M1027_d 0.00273233f $X=9.57 $Y=0.695 $X2=0
+ $Y2=0
cc_1131 N_A_1767_21#_c_1643_n N_VGND_M1027_d 0.00230147f $X=9.655 $Y=0.38 $X2=0
+ $Y2=0
cc_1132 N_A_1767_21#_M1027_g N_VGND_c_2283_n 0.00382497f $X=8.91 $Y=0.445 $X2=0
+ $Y2=0
cc_1133 N_A_1767_21#_c_1591_n N_VGND_c_2283_n 0.0100722f $X=9.295 $Y=0.78 $X2=0
+ $Y2=0
cc_1134 N_A_1767_21#_c_1592_n N_VGND_c_2283_n 0.00345716f $X=9.57 $Y=0.695 $X2=0
+ $Y2=0
cc_1135 N_A_1767_21#_c_1643_n N_VGND_c_2283_n 0.0110509f $X=9.655 $Y=0.38 $X2=0
+ $Y2=0
cc_1136 N_A_1767_21#_c_1597_n N_VGND_c_2283_n 0.00205754f $X=9.125 $Y=0.98 $X2=0
+ $Y2=0
cc_1137 N_A_1767_21#_c_1585_n N_VGND_c_2284_n 0.00438629f $X=11.015 $Y=0.995
+ $X2=0 $Y2=0
cc_1138 N_A_1767_21#_c_1593_n N_VGND_c_2284_n 0.0123434f $X=10.345 $Y=0.38 $X2=0
+ $Y2=0
cc_1139 N_A_1767_21#_c_1594_n N_VGND_c_2284_n 0.00513747f $X=10.43 $Y=0.995
+ $X2=0 $Y2=0
cc_1140 N_A_1767_21#_c_1595_n N_VGND_c_2284_n 0.00669683f $X=10.935 $Y=1.16
+ $X2=0 $Y2=0
cc_1141 N_A_1767_21#_c_1598_n N_VGND_c_2284_n 0.00169434f $X=12.285 $Y=1.16
+ $X2=0 $Y2=0
cc_1142 N_A_1767_21#_c_1586_n N_VGND_c_2285_n 0.00395881f $X=11.435 $Y=0.995
+ $X2=0 $Y2=0
cc_1143 N_A_1767_21#_c_1587_n N_VGND_c_2285_n 0.00147955f $X=11.865 $Y=0.995
+ $X2=0 $Y2=0
cc_1144 N_A_1767_21#_c_1598_n N_VGND_c_2285_n 0.0019324f $X=12.285 $Y=1.16 $X2=0
+ $Y2=0
cc_1145 N_A_1767_21#_c_1588_n N_VGND_c_2286_n 0.00316354f $X=12.285 $Y=0.995
+ $X2=0 $Y2=0
cc_1146 N_A_1767_21#_M1027_g N_VGND_c_2289_n 0.00463936f $X=8.91 $Y=0.445 $X2=0
+ $Y2=0
cc_1147 N_A_1767_21#_c_1590_n N_VGND_c_2291_n 0.00305478f $X=9.485 $Y=0.78 $X2=0
+ $Y2=0
cc_1148 N_A_1767_21#_c_1591_n N_VGND_c_2291_n 6.89658e-19 $X=9.295 $Y=0.78 $X2=0
+ $Y2=0
cc_1149 N_A_1767_21#_c_1593_n N_VGND_c_2291_n 0.0403365f $X=10.345 $Y=0.38 $X2=0
+ $Y2=0
cc_1150 N_A_1767_21#_c_1643_n N_VGND_c_2291_n 0.00773128f $X=9.655 $Y=0.38 $X2=0
+ $Y2=0
cc_1151 N_A_1767_21#_c_1585_n N_VGND_c_2293_n 0.00585385f $X=11.015 $Y=0.995
+ $X2=0 $Y2=0
cc_1152 N_A_1767_21#_c_1586_n N_VGND_c_2293_n 0.00526721f $X=11.435 $Y=0.995
+ $X2=0 $Y2=0
cc_1153 N_A_1767_21#_c_1587_n N_VGND_c_2295_n 0.00585385f $X=11.865 $Y=0.995
+ $X2=0 $Y2=0
cc_1154 N_A_1767_21#_c_1588_n N_VGND_c_2295_n 0.00541763f $X=12.285 $Y=0.995
+ $X2=0 $Y2=0
cc_1155 N_A_1767_21#_M1015_d N_VGND_c_2301_n 0.00219929f $X=10.125 $Y=0.235
+ $X2=0 $Y2=0
cc_1156 N_A_1767_21#_M1027_g N_VGND_c_2301_n 0.00654514f $X=8.91 $Y=0.445 $X2=0
+ $Y2=0
cc_1157 N_A_1767_21#_c_1585_n N_VGND_c_2301_n 0.0119391f $X=11.015 $Y=0.995
+ $X2=0 $Y2=0
cc_1158 N_A_1767_21#_c_1586_n N_VGND_c_2301_n 0.00922259f $X=11.435 $Y=0.995
+ $X2=0 $Y2=0
cc_1159 N_A_1767_21#_c_1587_n N_VGND_c_2301_n 0.0106394f $X=11.865 $Y=0.995
+ $X2=0 $Y2=0
cc_1160 N_A_1767_21#_c_1588_n N_VGND_c_2301_n 0.0105952f $X=12.285 $Y=0.995
+ $X2=0 $Y2=0
cc_1161 N_A_1767_21#_c_1590_n N_VGND_c_2301_n 0.00219209f $X=9.485 $Y=0.78 $X2=0
+ $Y2=0
cc_1162 N_A_1767_21#_c_1591_n N_VGND_c_2301_n 8.93798e-19 $X=9.295 $Y=0.78 $X2=0
+ $Y2=0
cc_1163 N_A_1767_21#_c_1593_n N_VGND_c_2301_n 0.0204716f $X=10.345 $Y=0.38 $X2=0
+ $Y2=0
cc_1164 N_A_1767_21#_c_1643_n N_VGND_c_2301_n 0.00285745f $X=9.655 $Y=0.38 $X2=0
+ $Y2=0
cc_1165 N_A_1767_21#_c_1597_n N_VGND_c_2301_n 5.84978e-19 $X=9.125 $Y=0.98 $X2=0
+ $Y2=0
cc_1166 N_A_1767_21#_c_1593_n A_1946_47# 0.00282053f $X=10.345 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_1167 N_A_1592_47#_M1032_g N_VPWR_c_1896_n 7.34118e-19 $X=10.075 $Y=2.275
+ $X2=0 $Y2=0
cc_1168 N_A_1592_47#_c_1779_n N_VPWR_c_1896_n 0.0218074f $X=9.015 $Y=2.295 $X2=0
+ $Y2=0
cc_1169 N_A_1592_47#_c_1782_n N_VPWR_c_1896_n 0.00819386f $X=10.04 $Y=1.66 $X2=0
+ $Y2=0
cc_1170 N_A_1592_47#_M1032_g N_VPWR_c_1897_n 0.00837332f $X=10.075 $Y=2.275
+ $X2=0 $Y2=0
cc_1171 N_A_1592_47#_M1032_g N_VPWR_c_1899_n 0.00427541f $X=10.075 $Y=2.275
+ $X2=0 $Y2=0
cc_1172 N_A_1592_47#_c_1779_n N_VPWR_c_1910_n 0.0508194f $X=9.015 $Y=2.295 $X2=0
+ $Y2=0
cc_1173 N_A_1592_47#_M1032_g N_VPWR_c_1911_n 0.00339367f $X=10.075 $Y=2.275
+ $X2=0 $Y2=0
cc_1174 N_A_1592_47#_M1001_d N_VPWR_c_1891_n 0.00177113f $X=8.36 $Y=2.065 $X2=0
+ $Y2=0
cc_1175 N_A_1592_47#_M1032_g N_VPWR_c_1891_n 0.00401529f $X=10.075 $Y=2.275
+ $X2=0 $Y2=0
cc_1176 N_A_1592_47#_c_1779_n N_VPWR_c_1891_n 0.0247853f $X=9.015 $Y=2.295 $X2=0
+ $Y2=0
cc_1177 N_A_1592_47#_c_1779_n A_1758_413# 0.00405625f $X=9.015 $Y=2.295
+ $X2=-0.19 $Y2=-0.24
cc_1178 N_A_1592_47#_c_1783_n N_VGND_c_2283_n 0.0212216f $X=8.745 $Y=0.395 $X2=0
+ $Y2=0
cc_1179 N_A_1592_47#_c_1773_n N_VGND_c_2284_n 0.00231294f $X=10.05 $Y=0.73 $X2=0
+ $Y2=0
cc_1180 N_A_1592_47#_c_1783_n N_VGND_c_2289_n 0.05415f $X=8.745 $Y=0.395 $X2=0
+ $Y2=0
cc_1181 N_A_1592_47#_c_1773_n N_VGND_c_2291_n 0.00366111f $X=10.05 $Y=0.73 $X2=0
+ $Y2=0
cc_1182 N_A_1592_47#_M1014_d N_VGND_c_2301_n 0.00272411f $X=7.96 $Y=0.235 $X2=0
+ $Y2=0
cc_1183 N_A_1592_47#_c_1773_n N_VGND_c_2301_n 0.00642361f $X=10.05 $Y=0.73 $X2=0
+ $Y2=0
cc_1184 N_A_1592_47#_c_1783_n N_VGND_c_2301_n 0.0155364f $X=8.745 $Y=0.395 $X2=0
+ $Y2=0
cc_1185 N_A_1592_47#_c_1783_n A_1701_47# 0.00425471f $X=8.745 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_1186 N_A_1592_47#_c_1775_n A_1701_47# 0.00145404f $X=8.83 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_1187 N_VPWR_c_1891_n A_538_389# 0.00308654f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1188 N_VPWR_c_1891_n N_A_620_389#_M1026_d 0.00623687f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1891_n N_A_620_389#_M1007_s 0.00250496f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1894_n N_A_620_389#_c_2133_n 0.00469069f $X=4.465 $Y=2.36 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1908_n N_A_620_389#_c_2133_n 0.011287f $X=4.3 $Y=2.72 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1891_n N_A_620_389#_c_2133_n 0.00297981f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1193 N_VPWR_M1035_d N_A_620_389#_c_2106_n 0.00227835f $X=4.33 $Y=1.945 $X2=0
+ $Y2=0
cc_1194 N_VPWR_c_1894_n N_A_620_389#_c_2106_n 0.0143961f $X=4.465 $Y=2.36 $X2=0
+ $Y2=0
cc_1195 N_VPWR_c_1891_n N_A_620_389#_c_2106_n 7.21087e-19 $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1908_n N_A_620_389#_c_2107_n 0.0137161f $X=4.3 $Y=2.72 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1891_n N_A_620_389#_c_2107_n 0.00992616f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1198 N_VPWR_M1035_d N_A_620_389#_c_2099_n 8.75701e-19 $X=4.33 $Y=1.945 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1894_n N_A_620_389#_c_2099_n 0.0144588f $X=4.465 $Y=2.36 $X2=0
+ $Y2=0
cc_1200 N_VPWR_c_1906_n N_A_620_389#_c_2099_n 0.0247511f $X=6.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1201 N_VPWR_c_1891_n N_A_620_389#_c_2099_n 0.0102194f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1202 N_VPWR_c_1891_n A_780_389# 0.00241551f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1203 N_VPWR_c_1891_n N_A_1191_413#_M1005_d 0.00231077f $X=12.65 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_1204 N_VPWR_c_1891_n N_A_1191_413#_M1033_d 0.00218037f $X=12.65 $Y=2.72 $X2=0
+ $Y2=0
cc_1205 N_VPWR_M1038_d N_A_1191_413#_c_2203_n 0.00379929f $X=6.375 $Y=2.065
+ $X2=0 $Y2=0
cc_1206 N_VPWR_c_1905_n N_A_1191_413#_c_2203_n 0.0143155f $X=6.575 $Y=2.44 $X2=0
+ $Y2=0
cc_1207 N_VPWR_c_1906_n N_A_1191_413#_c_2203_n 0.00344259f $X=6.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1208 N_VPWR_c_1909_n N_A_1191_413#_c_2203_n 0.0036489f $X=7.375 $Y=2.72 $X2=0
+ $Y2=0
cc_1209 N_VPWR_c_1891_n N_A_1191_413#_c_2203_n 0.00664736f $X=12.65 $Y=2.72
+ $X2=0 $Y2=0
cc_1210 N_VPWR_c_1906_n N_A_1191_413#_c_2204_n 0.00699759f $X=6.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1211 N_VPWR_c_1891_n N_A_1191_413#_c_2204_n 0.00284468f $X=12.65 $Y=2.72
+ $X2=0 $Y2=0
cc_1212 N_VPWR_c_1895_n N_A_1191_413#_c_2205_n 0.0135177f $X=7.6 $Y=2.34 $X2=0
+ $Y2=0
cc_1213 N_VPWR_c_1909_n N_A_1191_413#_c_2205_n 0.00711582f $X=7.375 $Y=2.72
+ $X2=0 $Y2=0
cc_1214 N_VPWR_c_1891_n N_A_1191_413#_c_2205_n 0.00284468f $X=12.65 $Y=2.72
+ $X2=0 $Y2=0
cc_1215 N_VPWR_c_1891_n A_1758_413# 0.00208799f $X=12.65 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1216 N_VPWR_c_1891_n N_Q_M1002_s 0.00409194f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1217 N_VPWR_c_1891_n N_Q_M1024_s 0.00409194f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1218 N_VPWR_c_1900_n N_Q_c_2243_n 0.0177999f $X=11.655 $Y=1.66 $X2=0 $Y2=0
cc_1219 N_VPWR_c_1913_n N_Q_c_2238_n 0.00795791f $X=12.41 $Y=2.72 $X2=0 $Y2=0
cc_1220 N_VPWR_c_1891_n N_Q_c_2238_n 0.00867074f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1221 N_VPWR_c_1900_n Q 0.0548313f $X=11.655 $Y=1.66 $X2=0 $Y2=0
cc_1222 N_VPWR_c_1912_n Q 0.00830819f $X=11.57 $Y=2.72 $X2=0 $Y2=0
cc_1223 N_VPWR_c_1891_n Q 0.00897758f $X=12.65 $Y=2.72 $X2=0 $Y2=0
cc_1224 N_VPWR_c_1900_n N_Q_c_2239_n 0.0071282f $X=11.655 $Y=1.66 $X2=0 $Y2=0
cc_1225 N_A_620_389#_c_2106_n A_780_389# 0.00282776f $X=4.565 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_1226 N_A_620_389#_c_2100_n N_VGND_M1030_d 2.35236e-19 $X=4.975 $Y=0.805 $X2=0
+ $Y2=0
cc_1227 N_A_620_389#_c_2101_n N_VGND_M1030_d 0.00244143f $X=4.735 $Y=0.805 $X2=0
+ $Y2=0
cc_1228 N_A_620_389#_c_2100_n N_VGND_c_2281_n 0.0029069f $X=4.975 $Y=0.805 $X2=0
+ $Y2=0
cc_1229 N_A_620_389#_c_2101_n N_VGND_c_2281_n 0.0138829f $X=4.735 $Y=0.805 $X2=0
+ $Y2=0
cc_1230 N_A_620_389#_c_2102_n N_VGND_c_2281_n 0.00247574f $X=5.06 $Y=0.715 $X2=0
+ $Y2=0
cc_1231 N_A_620_389#_c_2104_n N_VGND_c_2281_n 0.0125584f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_1232 N_A_620_389#_c_2100_n N_VGND_c_2299_n 0.00310525f $X=4.975 $Y=0.805
+ $X2=0 $Y2=0
cc_1233 N_A_620_389#_c_2104_n N_VGND_c_2299_n 0.0132448f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_1234 N_A_620_389#_M1023_s N_VGND_c_2301_n 0.00216416f $X=5.025 $Y=0.235 $X2=0
+ $Y2=0
cc_1235 N_A_620_389#_c_2100_n N_VGND_c_2301_n 0.00552288f $X=4.975 $Y=0.805
+ $X2=0 $Y2=0
cc_1236 N_A_620_389#_c_2101_n N_VGND_c_2301_n 7.57107e-19 $X=4.735 $Y=0.805
+ $X2=0 $Y2=0
cc_1237 N_A_620_389#_c_2104_n N_VGND_c_2301_n 0.0118267f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_1238 N_Q_c_2243_n N_VGND_c_2285_n 0.00636507f $X=11.99 $Y=1.16 $X2=0 $Y2=0
cc_1239 Q N_VGND_c_2285_n 0.0202973f $X=11.17 $Y=0.425 $X2=0 $Y2=0
cc_1240 Q N_VGND_c_2293_n 0.0148631f $X=11.17 $Y=0.425 $X2=0 $Y2=0
cc_1241 N_Q_c_2237_n N_VGND_c_2295_n 0.0142742f $X=12.075 $Y=0.63 $X2=0 $Y2=0
cc_1242 N_Q_M1016_s N_VGND_c_2301_n 0.0039413f $X=11.09 $Y=0.235 $X2=0 $Y2=0
cc_1243 N_Q_M1037_s N_VGND_c_2301_n 0.0039413f $X=11.94 $Y=0.235 $X2=0 $Y2=0
cc_1244 N_Q_c_2237_n N_VGND_c_2301_n 0.00937227f $X=12.075 $Y=0.63 $X2=0 $Y2=0
cc_1245 Q N_VGND_c_2301_n 0.00969704f $X=11.17 $Y=0.425 $X2=0 $Y2=0
cc_1246 N_VGND_c_2301_n A_1187_47# 0.00309919f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1247 N_VGND_c_2301_n A_1293_47# 0.00214708f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1248 N_VGND_c_2301_n A_1701_47# 0.00217993f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1249 N_VGND_c_2301_n A_1946_47# 0.00161179f $X=12.65 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a311oi_1.spice
* Created: Thu Aug 27 14:04:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a311oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a311oi_1  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1009 A_109_47# N_A3_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.169 PD=0.925 PS=1.82 NRD=15.228 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002 A=0.0975 P=1.6 MULT=1
MM1002 A_194_47# N_A2_M1002_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.089375 PD=0.93 PS=0.925 NRD=15.684 NRS=15.228 M=1 R=4.33333 SA=75000.6
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_A1_M1005_g A_194_47# VNB NSHORT L=0.15 W=0.65 AD=0.115375
+ AS=0.091 PD=1.005 PS=0.93 NRD=14.76 NRS=15.684 M=1 R=4.33333 SA=75001
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.112125 AS=0.115375 PD=0.995 PS=1.005 NRD=4.608 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.112125 PD=1.82 PS=0.995 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75002 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1006 N_A_109_297#_M1006_d N_A3_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.26 PD=1.275 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_109_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1375 PD=1.28 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_109_297#_M1008_d N_A1_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.14 PD=1.33 PS=1.28 NRD=0 NRS=0.9653 M=1 R=6.66667 SA=75001
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1004 A_376_297# N_B1_M1004_g N_A_109_297#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1725 AS=0.165 PD=1.345 PS=1.33 NRD=23.1278 NRS=10.8153 M=1 R=6.66667
+ SA=75001.5 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g A_376_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.1725 PD=2.52 PS=1.345 NRD=0 NRS=23.1278 M=1 R=6.66667 SA=75002 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a311oi_1.pxi.spice"
*
.ends
*
*

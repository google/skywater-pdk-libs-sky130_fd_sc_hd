* File: sky130_fd_sc_hd__lpflow_decapkapwr_3.spice.pex
* Created: Thu Aug 27 14:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%VGND 1 7 9 12 15 25 28
r16 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r17 25 27 0.442563 $w=8.27e-07 $l=3e-08 $layer=LI1_cond $X=1.12 $Y=0.375
+ $X2=1.15 $Y2=0.375
r18 23 25 11.4329 $w=8.27e-07 $l=7.75e-07 $layer=LI1_cond $X=0.345 $Y=0.375
+ $X2=1.12 $Y2=0.375
r19 22 23 1.25393 $w=8.27e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.375
+ $X2=0.345 $Y2=0.375
r20 19 22 0.442563 $w=8.27e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.375
+ $X2=0.26 $Y2=0.375
r21 15 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r22 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r23 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.29 $X2=0.42 $Y2=1.29
r24 10 23 3.45185 $w=5.2e-07 $l=4.6e-07 $layer=LI1_cond $X=0.345 $Y=0.835
+ $X2=0.345 $Y2=0.375
r25 10 12 10.4657 $w=5.18e-07 $l=4.55e-07 $layer=LI1_cond $X=0.345 $Y=0.835
+ $X2=0.345 $Y2=1.29
r26 7 13 41.3046 $w=5.9e-07 $l=5.89746e-07 $layer=POLY_cond $X=0.69 $Y=1.76
+ $X2=0.42 $Y2=1.29
r27 7 9 23.6915 $w=5.9e-07 $l=2.9e-07 $layer=POLY_cond $X=0.69 $Y=1.76 $X2=0.69
+ $Y2=2.05
r28 1 25 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.485
r29 1 22 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=0.26 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%KAPWR 1 9 14 18 30 31 33 35
c19 31 0 7.9696e-20 $X=1.15 $Y=2.21
r20 33 35 0.0085136 $w=2.6e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.21
+ $X2=0.23 $Y2=2.21
r21 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.21
+ $X2=1.15 $Y2=2.21
r22 28 30 0.397826 $w=9.18e-07 $l=3e-08 $layer=LI1_cond $X=1.12 $Y=2.005
+ $X2=1.15 $Y2=2.005
r23 26 28 1.12717 $w=9.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=2.005
+ $X2=1.12 $Y2=2.005
r24 25 26 10.2772 $w=9.18e-07 $l=7.75e-07 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=1.035 $Y2=2.005
r25 21 25 0.397826 $w=9.18e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.005
+ $X2=0.26 $Y2=2.005
r26 21 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r27 14 33 0.0120192 $w=2.6e-07 $l=2.5e-08 $layer=MET1_cond $X=0.19 $Y=2.21
+ $X2=0.215 $Y2=2.21
r28 14 31 0.495491 $w=2.6e-07 $l=8.73e-07 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=1.15 $Y2=2.21
r29 14 35 0.0266759 $w=2.6e-07 $l=4.7e-08 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=0.23 $Y2=2.21
r30 10 18 54.7084 $w=5.11e-07 $l=6.72607e-07 $layer=POLY_cond $X=0.96 $Y=1.09
+ $X2=0.76 $Y2=0.51
r31 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.09 $X2=0.96 $Y2=1.09
r32 7 26 4.07606 $w=5.2e-07 $l=4.6e-07 $layer=LI1_cond $X=1.035 $Y=1.545
+ $X2=1.035 $Y2=2.005
r33 7 9 10.4657 $w=5.18e-07 $l=4.55e-07 $layer=LI1_cond $X=1.035 $Y=1.545
+ $X2=1.035 $Y2=1.09
r34 1 28 300 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.615 $X2=1.12 $Y2=1.865
r35 1 25 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.615 $X2=0.26 $Y2=1.865
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%VPWR 1 8 9
c10 8 0 7.9696e-20 $X=1.15 $Y=2.72
r11 8 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72 $X2=1.15
+ $Y2=2.72
r12 4 8 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=1.15
+ $Y2=2.72
r13 1 9 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=1.15
+ $Y2=2.72
r14 1 4 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends


* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s50_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
M1000 X a_390_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.491e+11p pd=1.55e+06u as=4.027e+11p ps=3.97e+06u
M1001 a_283_47# a_27_47# VGND VNB nshort w=650000u l=500000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1002 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=6.517e+11p pd=5.37e+06u as=2.7e+11p ps=2.54e+06u
M1004 VPWR a_283_47# a_390_47# VPB phighvt w=820000u l=500000u
+  ad=0p pd=0u as=2.173e+11p ps=2.17e+06u
M1005 a_283_47# a_27_47# VPWR VPB phighvt w=820000u l=500000u
+  ad=2.173e+11p pd=2.17e+06u as=0p ps=0u
M1006 VGND a_283_47# a_390_47# VNB nshort w=650000u l=500000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1007 X a_390_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.55e+11p pd=2.71e+06u as=0p ps=0u
.ends


* NGSPICE file created from sky130_fd_sc_hd__nor4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
M1000 a_297_297# B a_191_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=3.8e+11p ps=2.76e+06u
M1001 VGND A Y VNB nshort w=650000u l=150000u
+  ad=5.1675e+11p pd=5.49e+06u as=4.1275e+11p ps=3.87e+06u
M1002 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_191_297# C a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1005 a_109_297# D Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1006 VPWR A a_297_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1007 Y D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


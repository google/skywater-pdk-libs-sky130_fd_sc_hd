* File: sky130_fd_sc_hd__a31o_4.pex.spice
* Created: Thu Aug 27 14:04:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A31O_4%A3 3 6 10 13 15 19 20 22 23 27 28 29 32
c91 32 0 1.91119e-19 $X=2.69 $Y=0.995
c92 20 0 4.1943e-20 $X=2.69 $Y=1.16
c93 13 0 3.06607e-19 $X=2.63 $Y=1.985
r94 27 30 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.385 $Y2=1.325
r95 27 29 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.385 $Y2=0.995
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r97 22 23 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=0.337 $Y=1.19
+ $X2=0.337 $Y2=1.53
r98 22 28 0.921954 $w=3.73e-07 $l=3e-08 $layer=LI1_cond $X=0.337 $Y=1.19
+ $X2=0.337 $Y2=1.16
r99 20 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=1.325
r100 20 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=0.995
r101 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.16 $X2=2.69 $Y2=1.16
r102 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.69 $Y=1.445
+ $X2=2.69 $Y2=1.16
r103 16 23 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.525 $Y=1.53
+ $X2=0.337 $Y2=1.53
r104 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.525 $Y=1.53
+ $X2=2.69 $Y2=1.445
r105 15 16 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=2.525 $Y=1.53
+ $X2=0.525 $Y2=1.53
r106 13 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.63 $Y=1.985
+ $X2=2.63 $Y2=1.325
r107 10 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.63 $Y=0.56
+ $X2=2.63 $Y2=0.995
r108 6 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r109 3 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%A2 1 3 6 8 10 13 16 17 18 20 21 23 24 30 31
+ 32
c88 32 0 1.91119e-19 $X=2.077 $Y=0.905
c89 18 0 1.75522e-19 $X=0.975 $Y=0.82
r90 31 33 1.21796 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=2.077 $Y=1.175
+ $X2=2.077 $Y2=1.075
r91 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.16 $X2=2.15 $Y2=1.16
r92 24 31 0.110909 $w=1.98e-07 $l=2e-09 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=2.077 $Y2=1.175
r93 23 32 3.28106 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.077 $Y=0.82
+ $X2=2.077 $Y2=0.905
r94 23 33 9.29238 $w=1.83e-07 $l=1.55e-07 $layer=LI1_cond $X=2.077 $Y=0.92
+ $X2=2.077 $Y2=1.075
r95 23 32 0.899263 $w=1.83e-07 $l=1.5e-08 $layer=LI1_cond $X=2.077 $Y=0.92
+ $X2=2.077 $Y2=0.905
r96 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r97 17 23 3.55127 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=1.985 $Y=0.82
+ $X2=2.077 $Y2=0.82
r98 17 18 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.985 $Y=0.82
+ $X2=0.975 $Y2=0.82
r99 16 20 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=1.075
+ $X2=0.89 $Y2=1.16
r100 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.89 $Y=0.905
+ $X2=0.975 $Y2=0.82
r101 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.89 $Y=0.905
+ $X2=0.89 $Y2=1.075
r102 11 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r103 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r104 8 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r105 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
r106 4 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r107 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r108 1 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r109 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%A1 3 7 11 15 17 24
r45 22 24 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.73 $Y2=1.16
r46 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r47 19 22 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r48 17 23 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.52 $Y2=1.175
r49 13 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r50 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r51 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r52 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r53 5 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r54 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295 $X2=1.31
+ $Y2=1.985
r55 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r56 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%B1 1 3 6 8 10 13 15 19 20 24 35
r64 27 35 0.601528 $w=2.15e-07 $l=1.05e-07 $layer=LI1_cond $X=3.922 $Y=1.075
+ $X2=3.922 $Y2=1.18
r65 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.16 $X2=3.74 $Y2=1.16
r66 20 35 0.369697 $w=2.08e-07 $l=7e-09 $layer=LI1_cond $X=3.915 $Y=1.18
+ $X2=3.922 $Y2=1.18
r67 20 25 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=3.915 $Y=1.18
+ $X2=3.74 $Y2=1.18
r68 19 27 12.0604 $w=2.13e-07 $l=2.25e-07 $layer=LI1_cond $X=3.922 $Y=0.85
+ $X2=3.922 $Y2=1.075
r69 16 18 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.11 $Y=1.16
+ $X2=3.53 $Y2=1.16
r70 15 24 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=3.605 $Y=1.16
+ $X2=3.74 $Y2=1.16
r71 15 18 15.1926 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.605 $Y=1.16
+ $X2=3.53 $Y2=1.16
r72 11 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.16
r73 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.985
r74 8 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=1.16
r75 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=0.56
r76 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r77 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325 $X2=3.11
+ $Y2=1.985
r78 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=1.16
r79 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.11 $Y=0.995 $X2=3.11
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%A_277_47# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 38 42 46 49 52 54 56 61 62 64 68 69
c152 69 0 1.89237e-19 $X=3.32 $Y=1.54
c153 49 0 1.1737e-19 $X=3.25 $Y=1.455
r154 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.31 $Y=1.16
+ $X2=5.73 $Y2=1.16
r155 77 78 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.89 $Y=1.16
+ $X2=5.31 $Y2=1.16
r156 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.435 $Y=0.48
+ $X2=2.435 $Y2=0.785
r157 62 79 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.85 $Y=1.16
+ $X2=5.73 $Y2=1.16
r158 61 62 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.85
+ $Y=1.16 $X2=5.85 $Y2=1.16
r159 59 77 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=4.49 $Y=1.16 $X2=4.89
+ $Y2=1.16
r160 59 74 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.49 $Y=1.16 $X2=4.47
+ $Y2=1.16
r161 58 61 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=4.49 $Y=1.16
+ $X2=5.85 $Y2=1.16
r162 58 59 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.49
+ $Y=1.16 $X2=4.49 $Y2=1.16
r163 56 72 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.31 $Y=1.16
+ $X2=4.31 $Y2=1.54
r164 56 58 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.395 $Y=1.16
+ $X2=4.49 $Y2=1.16
r165 55 69 2.90867 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=1.54
+ $X2=3.32 $Y2=1.54
r166 54 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=1.54
+ $X2=4.31 $Y2=1.54
r167 54 55 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.225 $Y=1.54
+ $X2=3.485 $Y2=1.54
r168 50 69 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=1.625
+ $X2=3.32 $Y2=1.54
r169 50 52 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.32 $Y=1.625
+ $X2=3.32 $Y2=1.63
r170 49 69 3.58051 $w=2.6e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.25 $Y=1.455
+ $X2=3.32 $Y2=1.54
r171 48 68 3.58051 $w=2.6e-07 $l=2.1225e-07 $layer=LI1_cond $X=3.25 $Y=0.87
+ $X2=3.155 $Y2=0.7
r172 48 49 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=3.25 $Y=0.87
+ $X2=3.25 $Y2=1.455
r173 44 68 3.58051 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=0.7
+ $X2=3.155 $Y2=0.7
r174 44 46 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.32 $Y=0.7
+ $X2=3.32 $Y2=0.38
r175 43 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0.785
+ $X2=2.435 $Y2=0.785
r176 42 68 2.90867 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=0.785
+ $X2=3.155 $Y2=0.7
r177 42 43 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.155 $Y=0.785
+ $X2=2.52 $Y2=0.785
r178 38 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0.48
+ $X2=2.435 $Y2=0.48
r179 38 40 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.35 $Y=0.48
+ $X2=1.52 $Y2=0.48
r180 34 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.325
+ $X2=5.73 $Y2=1.16
r181 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.73 $Y=1.325
+ $X2=5.73 $Y2=1.985
r182 31 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=0.995
+ $X2=5.73 $Y2=1.16
r183 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.73 $Y=0.995
+ $X2=5.73 $Y2=0.56
r184 27 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.325
+ $X2=5.31 $Y2=1.16
r185 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.31 $Y=1.325
+ $X2=5.31 $Y2=1.985
r186 24 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=0.995
+ $X2=5.31 $Y2=1.16
r187 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.31 $Y=0.995
+ $X2=5.31 $Y2=0.56
r188 20 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.325
+ $X2=4.89 $Y2=1.16
r189 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.89 $Y=1.325
+ $X2=4.89 $Y2=1.985
r190 17 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=0.995
+ $X2=4.89 $Y2=1.16
r191 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.89 $Y=0.995
+ $X2=4.89 $Y2=0.56
r192 13 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.47 $Y=1.325
+ $X2=4.47 $Y2=1.16
r193 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.47 $Y=1.325
+ $X2=4.47 $Y2=1.985
r194 10 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=1.16
r195 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=0.56
r196 3 52 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=1.63
r197 2 46 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.185
+ $Y=0.235 $X2=3.32 $Y2=0.38
r198 1 40 182 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%A_27_297# 1 2 3 4 5 18 22 26 28 30 31 34 37
+ 39 41
c55 28 0 4.1943e-20 $X=2.9 $Y=1.955
r56 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.74 $Y=2.295
+ $X2=3.74 $Y2=1.96
r57 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=2.38
+ $X2=3.74 $Y2=2.295
r58 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.655 $Y=2.38
+ $X2=2.985 $Y2=2.38
r59 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.9 $Y=2.295
+ $X2=2.985 $Y2=2.38
r60 28 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=1.955 $X2=2.9
+ $Y2=1.87
r61 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.9 $Y=1.955 $X2=2.9
+ $Y2=2.295
r62 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.87
+ $X2=1.94 $Y2=1.87
r63 26 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=1.87 $X2=2.9
+ $Y2=1.87
r64 26 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.815 $Y=1.87
+ $X2=2.025 $Y2=1.87
r65 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.87 $X2=1.1
+ $Y2=1.87
r66 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=1.87
+ $X2=1.94 $Y2=1.87
r67 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=1.87
+ $X2=1.185 $Y2=1.87
r68 19 37 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.26 $Y2=1.87
r69 18 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=1.87 $X2=1.1
+ $Y2=1.87
r70 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=1.87
+ $X2=0.345 $Y2=1.87
r71 5 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.605
+ $Y=1.485 $X2=3.74 $Y2=1.96
r72 4 43 300 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=2 $X=2.705
+ $Y=1.485 $X2=2.9 $Y2=1.95
r73 3 41 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.95
r74 2 39 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.95
r75 1 37 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 53 54 56 57 58 60 85 86 89
r111 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r112 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r113 83 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r116 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r117 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r118 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r120 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r121 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 71 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r123 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r125 68 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r126 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 65 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r128 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r129 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r130 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r131 58 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 58 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r133 56 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.775 $Y=2.72
+ $X2=5.75 $Y2=2.72
r134 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=2.72
+ $X2=5.94 $Y2=2.72
r135 55 85 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.105 $Y=2.72
+ $X2=6.21 $Y2=2.72
r136 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=2.72
+ $X2=5.94 $Y2=2.72
r137 53 79 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=5.1 $Y2=2.72
r139 52 82 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.75 $Y2=2.72
r140 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.1 $Y2=2.72
r141 50 76 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=3.91 $Y2=2.72
r142 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=4.26 $Y2=2.72
r143 49 79 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.26 $Y2=2.72
r145 47 70 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r146 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.36 $Y2=2.72
r147 46 73 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.53 $Y2=2.72
r148 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.36 $Y2=2.72
r149 44 67 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.15 $Y2=2.72
r150 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.52 $Y2=2.72
r151 43 70 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=2.07 $Y2=2.72
r152 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.52 $Y2=2.72
r153 39 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.635
+ $X2=5.94 $Y2=2.72
r154 39 41 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.94 $Y=2.635
+ $X2=5.94 $Y2=2.21
r155 35 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=2.635 $X2=5.1
+ $Y2=2.72
r156 35 37 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.1 $Y=2.635
+ $X2=5.1 $Y2=2.21
r157 31 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=2.635
+ $X2=4.26 $Y2=2.72
r158 31 33 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.26 $Y=2.635
+ $X2=4.26 $Y2=2.21
r159 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r160 27 29 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.21
r161 23 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r162 23 25 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.21
r163 19 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r164 19 21 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.21
r165 6 41 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.94 $Y2=2.21
r166 5 37 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.485 $X2=5.1 $Y2=2.21
r167 4 33 600 $w=1.7e-07 $l=7.85016e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.26 $Y2=2.21
r168 3 29 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.21
r169 2 25 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.21
r170 1 21 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%X 1 2 3 4 15 20 23 24 25 26 27 36 39
r52 47 50 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.68 $Y=0.74
+ $X2=5.52 $Y2=0.74
r53 36 39 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.21 $Y=0.825
+ $X2=6.21 $Y2=0.85
r54 26 27 11.5225 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=6.21 $Y=1.53
+ $X2=6.21 $Y2=1.785
r55 25 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.21 $Y=1.19
+ $X2=6.21 $Y2=1.53
r56 24 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=0.74 $X2=6.21
+ $Y2=0.825
r57 24 50 31.122 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=6.125 $Y=0.74
+ $X2=5.52 $Y2=0.74
r58 24 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.21 $Y=0.88
+ $X2=6.21 $Y2=1.19
r59 24 39 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=6.21 $Y=0.88 $X2=6.21
+ $Y2=0.85
r60 21 27 19.0652 $w=3.38e-07 $l=5.2e-07 $layer=LI1_cond $X=5.605 $Y=1.87
+ $X2=6.125 $Y2=1.87
r61 21 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=1.87
+ $X2=5.52 $Y2=1.87
r62 16 20 3.40825 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.765 $Y=1.87
+ $X2=4.65 $Y2=1.87
r63 15 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=1.87
+ $X2=5.52 $Y2=1.87
r64 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.435 $Y=1.87
+ $X2=4.765 $Y2=1.87
r65 4 23 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.385
+ $Y=1.485 $X2=5.52 $Y2=1.95
r66 3 20 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.545
+ $Y=1.485 $X2=4.68 $Y2=1.95
r67 2 50 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.235 $X2=5.52 $Y2=0.74
r68 1 47 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_4%VGND 1 2 3 4 5 16 18 22 26 30 33 34 36 37 39
+ 40 41 50 62 63 70
r94 70 73 9.02701 $w=5.28e-07 $l=4e-07 $layer=LI1_cond $X=4 $Y=0 $X2=4 $Y2=0.4
r95 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r96 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r97 60 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r98 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r99 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r100 57 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r101 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r102 54 70 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4
+ $Y2=0
r103 54 56 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.83
+ $Y2=0
r104 53 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r105 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r106 50 70 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=4
+ $Y2=0
r107 50 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.45 $Y2=0
r108 49 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r109 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r110 46 49 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.53 $Y2=0
r111 45 48 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r112 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r113 43 66 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r114 43 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r115 41 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r116 41 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r117 39 59 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.75
+ $Y2=0
r118 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.94
+ $Y2=0
r119 38 62 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.105 $Y=0
+ $X2=6.21 $Y2=0
r120 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=5.94
+ $Y2=0
r121 36 56 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.935 $Y=0
+ $X2=4.83 $Y2=0
r122 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=5.1
+ $Y2=0
r123 35 59 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.265 $Y=0
+ $X2=5.75 $Y2=0
r124 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=0 $X2=5.1
+ $Y2=0
r125 33 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.53
+ $Y2=0
r126 33 34 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.842
+ $Y2=0
r127 32 52 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=3.45 $Y2=0
r128 32 34 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=2.842 $Y2=0
r129 28 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=0.085
+ $X2=5.94 $Y2=0
r130 28 30 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.94 $Y=0.085
+ $X2=5.94 $Y2=0.4
r131 24 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=0.085 $X2=5.1
+ $Y2=0
r132 24 26 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.1 $Y=0.085
+ $X2=5.1 $Y2=0.4
r133 20 34 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.842 $Y=0.085
+ $X2=2.842 $Y2=0
r134 20 22 11.3222 $w=2.83e-07 $l=2.8e-07 $layer=LI1_cond $X=2.842 $Y=0.085
+ $X2=2.842 $Y2=0.365
r135 16 66 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r136 16 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r137 5 30 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.235 $X2=5.94 $Y2=0.4
r138 4 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.1 $Y2=0.4
r139 3 73 91 $w=1.7e-07 $l=6.52304e-07 $layer=licon1_NDIFF $count=2 $X=3.605
+ $Y=0.235 $X2=4.18 $Y2=0.4
r140 2 22 182 $w=1.7e-07 $l=2.3103e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.235 $X2=2.88 $Y2=0.365
r141 1 18 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__or4bb_4.pex.spice
* Created: Thu Aug 27 14:44:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4BB_4%C_N 3 7 8 9 13 14 15
c33 3 0 1.33368e-19 $X=0.47 $Y=2.26
r34 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r35 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r37 8 9 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.53
r38 8 14 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.16
r39 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=0.675
+ $X2=0.505 $Y2=0.995
r40 3 16 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.47 $Y=2.26
+ $X2=0.47 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%D_N 3 6 8 11 13
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.16
+ $X2=1.03 $Y2=1.325
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.16
+ $X2=1.03 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.16 $X2=1.03 $Y2=1.16
r37 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.03
+ $Y2=1.16
r38 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.955 $Y=1.695
+ $X2=0.955 $Y2=1.325
r39 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.95 $Y=0.675
+ $X2=0.95 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%A_205_93# 1 2 7 9 12 14 15 16 23 25 28 30
c66 16 0 1.33368e-19 $X=1.405 $Y=1.61
r67 28 31 7.92688 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=1.16
+ $X2=1.55 $Y2=1.325
r68 28 30 7.92688 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=1.16
+ $X2=1.55 $Y2=0.995
r69 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r70 25 26 17.5021 $w=2.37e-07 $l=3.4e-07 $layer=LI1_cond $X=1.16 $Y=0.655
+ $X2=1.5 $Y2=0.655
r71 23 31 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=1.5 $Y=1.525 $X2=1.5
+ $Y2=1.325
r72 20 26 2.03416 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=1.5 $Y=0.825 $X2=1.5
+ $Y2=0.655
r73 20 30 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=1.5 $Y=0.825 $X2=1.5
+ $Y2=0.995
r74 16 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.405 $Y=1.61
+ $X2=1.5 $Y2=1.525
r75 16 18 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.405 $Y=1.61
+ $X2=1.165 $Y2=1.61
r76 14 29 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=1.61 $Y2=1.16
r77 14 15 5.03009 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=1.9 $Y2=1.16
r78 10 15 37.0704 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.91 $Y=1.325
+ $X2=1.9 $Y2=1.16
r79 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.91 $Y=1.325
+ $X2=1.91 $Y2=1.985
r80 7 15 37.0704 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.89 $Y=0.995
+ $X2=1.9 $Y2=1.16
r81 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.89 $Y=0.995 $X2=1.89
+ $Y2=0.56
r82 2 18 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.61
r83 1 25 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.465 $X2=1.16 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%A_27_410# 1 2 9 12 15 18 20 23 24 25 28 29
+ 34 36 38
r87 31 34 3.84148 $w=3.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.17 $Y=0.637
+ $X2=0.295 $Y2=0.637
r88 29 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.16
+ $X2=2.36 $Y2=1.325
r89 29 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.16
+ $X2=2.36 $Y2=0.995
r90 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r91 26 28 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.36 $Y=2.295
+ $X2=2.36 $Y2=1.16
r92 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.275 $Y=2.38
+ $X2=2.36 $Y2=2.295
r93 24 25 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.275 $Y=2.38
+ $X2=1.295 $Y2=2.38
r94 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.295
+ $X2=1.295 $Y2=2.38
r95 22 23 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.21 $Y=2.035
+ $X2=1.21 $Y2=2.295
r96 21 36 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.95
+ $X2=0.215 $Y2=1.95
r97 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.125 $Y=1.95
+ $X2=1.21 $Y2=2.035
r98 20 21 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.125 $Y=1.95
+ $X2=0.345 $Y2=1.95
r99 16 36 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=1.95
r100 16 18 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.29
r101 15 36 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.17 $Y=1.865
+ $X2=0.215 $Y2=1.95
r102 14 31 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.637
r103 14 15 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.865
r104 12 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.42 $Y=1.985
+ $X2=2.42 $Y2=1.325
r105 9 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.42 $Y=0.56
+ $X2=2.42 $Y2=0.995
r106 2 18 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r107 1 34 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.465 $X2=0.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%B 1 3 6 10 11 14 15 31
c39 11 0 5.72837e-20 $X=2.84 $Y=1.16
c40 6 0 2.99791e-19 $X=2.84 $Y=1.985
r41 21 31 2.70104 $w=3.18e-07 $l=7.5e-08 $layer=LI1_cond $X=2.955 $Y=1.945
+ $X2=2.955 $Y2=1.87
r42 14 31 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=2.955 $Y=1.865
+ $X2=2.955 $Y2=1.87
r43 14 15 9.3636 $w=3.18e-07 $l=2.6e-07 $layer=LI1_cond $X=2.955 $Y=1.95
+ $X2=2.955 $Y2=2.21
r44 14 21 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=2.955 $Y=1.95
+ $X2=2.955 $Y2=1.945
r45 13 14 14.2094 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.9 $Y=1.45 $X2=2.9
+ $Y2=1.785
r46 10 13 11.6456 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.84 $Y=1.16
+ $X2=2.84 $Y2=1.45
r47 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.16 $X2=2.84 $Y2=1.16
r48 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.325
+ $X2=2.84 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.84 $Y=1.325 $X2=2.84
+ $Y2=1.985
r50 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995 $X2=2.84
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%A 3 6 8 12 13 14
c41 13 0 1.24234e-19 $X=3.32 $Y=1.16
c42 8 0 1.75557e-19 $X=3.47 $Y=1.53
r43 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.32 $Y=1.16
+ $X2=3.32 $Y2=1.325
r44 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.32 $Y=1.16
+ $X2=3.32 $Y2=0.995
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.16 $X2=3.32 $Y2=1.16
r46 8 20 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.47 $Y=1.53 $X2=3.32
+ $Y2=1.53
r47 8 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=1.445
+ $X2=3.32 $Y2=1.53
r48 8 13 16.7846 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=3.32 $Y=1.445
+ $X2=3.32 $Y2=1.16
r49 6 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.26 $Y=1.985
+ $X2=3.26 $Y2=1.325
r50 3 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.26 $Y=0.56 $X2=3.26
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%A_315_380# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 43 46 48 49 52 54 57 58 63 69 76
c147 69 0 5.72837e-20 $X=3.05 $Y=0.74
c148 54 0 1.60701e-19 $X=3.575 $Y=0.74
r149 73 74 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.21 $Y=1.16
+ $X2=4.63 $Y2=1.16
r150 66 68 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.02 $Y=0.74
+ $X2=2.18 $Y2=0.74
r151 64 76 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.87 $Y=1.16
+ $X2=5.05 $Y2=1.16
r152 64 74 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.87 $Y=1.16
+ $X2=4.63 $Y2=1.16
r153 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.87
+ $Y=1.16 $X2=4.87 $Y2=1.16
r154 61 73 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.85 $Y=1.16
+ $X2=4.21 $Y2=1.16
r155 61 70 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.85 $Y=1.16 $X2=3.79
+ $Y2=1.16
r156 60 63 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=4.87 $Y2=1.16
r157 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.85
+ $Y=1.16 $X2=3.85 $Y2=1.16
r158 58 60 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.745 $Y=1.16
+ $X2=3.85 $Y2=1.16
r159 57 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.66 $Y=1.075
+ $X2=3.745 $Y2=1.16
r160 56 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.66 $Y=0.825
+ $X2=3.66 $Y2=1.075
r161 55 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=0.74
+ $X2=3.05 $Y2=0.74
r162 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.575 $Y=0.74
+ $X2=3.66 $Y2=0.825
r163 54 55 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.575 $Y=0.74
+ $X2=3.135 $Y2=0.74
r164 50 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=0.655
+ $X2=3.05 $Y2=0.74
r165 50 52 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0.655
+ $X2=3.05 $Y2=0.49
r166 49 68 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=0.74
+ $X2=2.18 $Y2=0.74
r167 48 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=0.74
+ $X2=3.05 $Y2=0.74
r168 48 49 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.965 $Y=0.74
+ $X2=2.265 $Y2=0.74
r169 44 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.655
+ $X2=2.18 $Y2=0.74
r170 44 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0.655
+ $X2=2.18 $Y2=0.49
r171 42 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.825
+ $X2=2.02 $Y2=0.74
r172 42 43 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.02 $Y=0.825
+ $X2=2.02 $Y2=1.955
r173 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.935 $Y=2.04
+ $X2=2.02 $Y2=1.955
r174 38 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.935 $Y=2.04
+ $X2=1.7 $Y2=2.04
r175 34 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.16
r176 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.985
r177 31 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=1.16
r178 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=0.56
r179 27 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=1.325
+ $X2=4.63 $Y2=1.16
r180 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.63 $Y=1.325
+ $X2=4.63 $Y2=1.985
r181 24 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.63 $Y2=1.16
r182 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.63 $Y2=0.56
r183 20 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.325
+ $X2=4.21 $Y2=1.16
r184 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.21 $Y=1.325
+ $X2=4.21 $Y2=1.985
r185 17 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=0.995
+ $X2=4.21 $Y2=1.16
r186 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.21 $Y=0.995
+ $X2=4.21 $Y2=0.56
r187 13 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=1.325
+ $X2=3.79 $Y2=1.16
r188 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.79 $Y=1.325
+ $X2=3.79 $Y2=1.985
r189 10 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=0.995
+ $X2=3.79 $Y2=1.16
r190 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.79 $Y=0.995
+ $X2=3.79 $Y2=0.56
r191 3 40 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.9 $X2=1.7 $Y2=2.04
r192 2 52 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.05 $Y2=0.49
r193 1 46 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.235 $X2=2.18 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%VPWR 1 2 3 4 15 19 21 25 27 29 31 33 38 43
+ 49 52 55 59
r73 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r74 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r75 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r77 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 47 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 47 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r80 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r81 44 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.42 $Y2=2.72
r82 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.83 $Y2=2.72
r83 43 58 3.98688 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.327 $Y2=2.72
r84 43 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=4.83 $Y2=2.72
r85 42 53 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 42 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r87 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 39 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r89 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r90 38 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.4 $Y=2.72
+ $X2=3.525 $Y2=2.72
r91 38 41 146.791 $w=1.68e-07 $l=2.25e-06 $layer=LI1_cond $X=3.4 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 33 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r93 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r94 31 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r96 27 58 3.15628 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=5.26 $Y=2.635
+ $X2=5.327 $Y2=2.72
r97 27 29 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.26 $Y=2.635
+ $X2=5.26 $Y2=1.96
r98 23 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.635
+ $X2=4.42 $Y2=2.72
r99 23 25 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.42 $Y=2.635
+ $X2=4.42 $Y2=1.96
r100 22 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.65 $Y=2.72
+ $X2=3.525 $Y2=2.72
r101 21 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.42 $Y2=2.72
r102 21 22 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=3.65 $Y2=2.72
r103 17 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.635
+ $X2=3.525 $Y2=2.72
r104 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.525 $Y=2.635
+ $X2=3.525 $Y2=1.96
r105 13 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r106 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.29
r107 4 29 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.485 $X2=5.26 $Y2=1.96
r108 3 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.285
+ $Y=1.485 $X2=4.42 $Y2=1.96
r109 2 19 300 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_PDIFF $count=2 $X=3.335
+ $Y=1.485 $X2=3.525 $Y2=1.96
r110 1 15 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=0.545 $Y=2.05
+ $X2=0.68 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%X 1 2 3 4 13 15 19 21 23 24 27 31 33 35 39
+ 41 43 46
r74 43 46 3.05086 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.32 $Y=0.815 $X2=5.32
+ $Y2=0.905
r75 43 46 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.32 $Y=0.92
+ $X2=5.32 $Y2=0.905
r76 42 43 26.8068 $w=2.28e-07 $l=5.35e-07 $layer=LI1_cond $X=5.32 $Y=1.455
+ $X2=5.32 $Y2=0.92
r77 36 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=0.815
+ $X2=4.84 $Y2=0.815
r78 35 43 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=5.205 $Y=0.815
+ $X2=5.32 $Y2=0.815
r79 35 36 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=5.205 $Y=0.815
+ $X2=5.005 $Y2=0.815
r80 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.965 $Y=1.54
+ $X2=4.84 $Y2=1.54
r81 33 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.205 $Y=1.54
+ $X2=5.32 $Y2=1.455
r82 33 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.205 $Y=1.54
+ $X2=4.965 $Y2=1.54
r83 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=1.625
+ $X2=4.84 $Y2=1.54
r84 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.84 $Y=1.625
+ $X2=4.84 $Y2=2.3
r85 25 39 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.84 $Y=0.725 $X2=4.84
+ $Y2=0.815
r86 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.84 $Y=0.725
+ $X2=4.84 $Y2=0.39
r87 23 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=0.815
+ $X2=4.84 $Y2=0.815
r88 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.675 $Y=0.815
+ $X2=4.165 $Y2=0.815
r89 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.125 $Y=1.54 $X2=4
+ $Y2=1.54
r90 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.715 $Y=1.54
+ $X2=4.84 $Y2=1.54
r91 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.715 $Y=1.54
+ $X2=4.125 $Y2=1.54
r92 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.04 $Y=0.725
+ $X2=4.165 $Y2=0.815
r93 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=4.04 $Y=0.725
+ $X2=4.04 $Y2=0.485
r94 13 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=1.625 $X2=4
+ $Y2=1.54
r95 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4 $Y=1.625 $X2=4
+ $Y2=2.3
r96 4 41 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.705
+ $Y=1.485 $X2=4.84 $Y2=1.62
r97 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.705
+ $Y=1.485 $X2=4.84 $Y2=2.3
r98 3 38 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.485 $X2=4 $Y2=1.62
r99 3 15 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.485 $X2=4 $Y2=2.3
r100 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.705
+ $Y=0.235 $X2=4.84 $Y2=0.39
r101 1 19 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=3.865
+ $Y=0.235 $X2=4 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_4%VGND 1 2 3 4 5 6 23 27 29 33 37 39 43 45 47
+ 49 51 56 61 67 70 73 76 79 83
c103 39 0 1.60701e-19 $X=4.335 $Y=0
r104 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r105 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r106 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r107 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r108 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r109 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r110 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r111 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r112 65 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r113 65 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r114 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r115 62 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.505 $Y=0 $X2=4.42
+ $Y2=0
r116 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=4.83 $Y2=0
r117 61 82 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.347 $Y2=0
r118 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=4.83
+ $Y2=0
r119 60 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r120 60 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r121 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r122 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r123 57 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=2.99 $Y2=0
r124 56 76 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.545
+ $Y2=0
r125 56 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.355 $Y=0
+ $X2=2.99 $Y2=0
r126 55 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r127 55 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r128 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r129 52 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.74
+ $Y2=0
r130 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=0
+ $X2=1.15 $Y2=0
r131 51 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.68
+ $Y2=0
r132 51 54 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=1.15 $Y2=0
r133 49 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r134 45 82 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=5.26 $Y=0.085
+ $X2=5.347 $Y2=0
r135 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.26 $Y=0.085
+ $X2=5.26 $Y2=0.39
r136 41 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=0.085
+ $X2=4.42 $Y2=0
r137 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.42 $Y=0.085
+ $X2=4.42 $Y2=0.39
r138 40 76 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.545
+ $Y2=0
r139 39 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.42
+ $Y2=0
r140 39 40 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=3.735
+ $Y2=0
r141 35 76 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0
r142 35 37 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0.4
r143 31 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r144 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.4
r145 30 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.68
+ $Y2=0
r146 29 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r147 29 30 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=1.845 $Y2=0
r148 25 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0
r149 25 27 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0.395
r150 21 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r151 21 23 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.66
r152 6 47 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.26 $Y2=0.39
r153 5 43 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.285
+ $Y=0.235 $X2=4.42 $Y2=0.39
r154 4 37 182 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.235 $X2=3.57 $Y2=0.4
r155 3 33 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.63 $Y2=0.4
r156 2 27 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.68 $Y2=0.395
r157 1 23 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.465 $X2=0.74 $Y2=0.66
.ends


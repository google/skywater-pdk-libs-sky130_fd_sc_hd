* File: sky130_fd_sc_hd__dlrtp_4.pex.spice
* Created: Thu Aug 27 14:17:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRTP_4%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%A_27_47# 1 2 9 13 17 19 20 23 27 30 34 35 36
+ 41 44 46 49 50 53 56 57 60 64
c145 57 0 7.61652e-20 $X=2.56 $Y=1.53
c146 13 0 2.6965e-20 $X=0.89 $Y=2.135
c147 9 0 2.6965e-20 $X=0.89 $Y=0.445
r148 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.52 $X2=2.675 $Y2=1.52
r149 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.56 $Y=1.53
+ $X2=2.56 $Y2=1.53
r150 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r151 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r152 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.415 $Y=1.53
+ $X2=2.56 $Y2=1.53
r153 49 50 1.94925 $w=1.4e-07 $l=1.575e-06 $layer=MET1_cond $X=2.415 $Y=1.53
+ $X2=0.84 $Y2=1.53
r154 48 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r155 47 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r156 45 64 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r157 44 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r158 44 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r159 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r160 38 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r161 37 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r162 36 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r163 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r164 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r165 34 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r166 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r167 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r168 26 60 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.675 $Y=1.55
+ $X2=2.675 $Y2=1.52
r169 26 27 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.675 $Y=1.55
+ $X2=2.675 $Y2=1.685
r170 25 60 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.675 $Y=1.395
+ $X2=2.675 $Y2=1.52
r171 21 23 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.225 $Y=1.245
+ $X2=3.225 $Y2=0.415
r172 20 25 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.81 $Y=1.32
+ $X2=2.675 $Y2=1.395
r173 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.15 $Y=1.32
+ $X2=3.225 $Y2=1.245
r174 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.15 $Y=1.32
+ $X2=2.81 $Y2=1.32
r175 17 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.685
r176 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r177 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r178 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r179 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r180 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r181 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.63 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.63 $Y=1.04
+ $X2=1.835 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.04 $X2=1.63 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.63 $Y=1.19 $X2=1.63
+ $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.205
+ $X2=1.835 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.835 $Y=1.205
+ $X2=1.835 $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=0.875
+ $X2=1.835 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.835 $Y=0.875
+ $X2=1.835 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%A_300_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c85 32 0 1.12109e-19 $X=2.26 $Y=0.93
c86 18 0 7.13094e-20 $X=1.975 $Y=0.7
r87 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.93
+ $X2=2.26 $Y2=1.095
r88 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.93
+ $X2=2.26 $Y2=0.765
r89 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=0.93 $X2=2.26 $Y2=0.93
r90 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.625 $Y=0.51
+ $X2=1.625 $Y2=0.7
r91 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.06 $Y=1.095
+ $X2=2.16 $Y2=0.93
r92 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.06 $Y=1.095 $X2=2.06
+ $Y2=1.495
r93 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.975 $Y=1.58
+ $X2=2.06 $Y2=1.495
r94 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=1.58
+ $X2=1.79 $Y2=1.58
r95 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.7
+ $X2=1.625 $Y2=0.7
r96 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.975 $Y=0.7
+ $X2=2.16 $Y2=0.93
r97 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.975 $Y=0.7
+ $X2=1.71 $Y2=0.7
r98 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.79 $Y2=1.58
r99 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.625 $Y2=1.99
r100 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.255 $Y=2.165
+ $X2=2.255 $Y2=1.095
r101 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.255 $Y=0.445
+ $X2=2.255 $Y2=0.765
r102 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.845 $X2=1.625 $Y2=1.99
r103 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.235 $X2=1.625 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%A_193_47# 1 2 9 12 16 20 24 26 28 29 32 35
+ 39 43 45 51
c122 45 0 7.61652e-20 $X=3.34 $Y=1.74
r123 43 51 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.1 $Y=1.74
+ $X2=3.1 $Y2=1.575
r124 42 45 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.185 $Y=1.74
+ $X2=3.34 $Y2=1.74
r125 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.74 $X2=3.185 $Y2=1.74
r126 35 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.02 $Y=1.87
+ $X2=3.02 $Y2=1.87
r127 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r128 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r129 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.875 $Y=1.87
+ $X2=3.02 $Y2=1.87
r130 28 29 1.94925 $w=1.4e-07 $l=1.575e-06 $layer=MET1_cond $X=2.875 $Y=1.87
+ $X2=1.3 $Y2=1.87
r131 24 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=0.87
+ $X2=2.805 $Y2=0.705
r132 23 26 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.805 $Y=0.87
+ $X2=3.015 $Y2=0.87
r133 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=0.87 $X2=2.805 $Y2=0.87
r134 20 32 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r135 20 21 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r136 18 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=1.035
+ $X2=3.015 $Y2=0.87
r137 18 51 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.015 $Y=1.035
+ $X2=3.015 $Y2=1.575
r138 16 21 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r139 10 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.34 $Y=1.875
+ $X2=3.34 $Y2=1.74
r140 10 12 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.34 $Y=1.875
+ $X2=3.34 $Y2=2.275
r141 9 39 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.795 $Y=0.415
+ $X2=2.795 $Y2=0.705
r142 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r143 1 16 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%A_725_21# 1 2 9 13 15 17 20 22 24 27 29 31
+ 34 36 38 41 43 46 50 52 53 56 58 63 66 75
c151 75 0 1.81835e-20 $X=6.89 $Y=1.16
r152 74 75 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=6.43 $Y=1.16
+ $X2=6.89 $Y2=1.16
r153 73 74 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=5.995 $Y=1.16
+ $X2=6.43 $Y2=1.16
r154 64 73 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=5.54 $Y=1.16
+ $X2=5.995 $Y2=1.16
r155 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.54
+ $Y=1.16 $X2=5.54 $Y2=1.16
r156 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.54 $Y=1.535
+ $X2=5.54 $Y2=1.16
r157 60 63 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.54 $Y=0.825
+ $X2=5.54 $Y2=1.16
r158 59 66 4.08801 $w=2.5e-07 $l=1.28938e-07 $layer=LI1_cond $X=4.945 $Y=1.62
+ $X2=4.85 $Y2=1.7
r159 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=1.62
+ $X2=5.54 $Y2=1.535
r160 58 59 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.455 $Y=1.62
+ $X2=4.945 $Y2=1.62
r161 54 66 2.34704 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=1.865
+ $X2=4.85 $Y2=1.7
r162 54 56 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=4.85 $Y=1.865
+ $X2=4.85 $Y2=2.27
r163 52 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=0.74
+ $X2=5.54 $Y2=0.825
r164 52 53 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.455 $Y=0.74
+ $X2=4.595 $Y2=0.74
r165 48 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.43 $Y=0.655
+ $X2=4.595 $Y2=0.74
r166 48 50 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.43 $Y=0.655
+ $X2=4.43 $Y2=0.4
r167 46 67 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.93 $Y=1.7 $X2=3.7
+ $Y2=1.7
r168 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.7 $X2=3.93 $Y2=1.7
r169 43 66 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.755 $Y=1.7
+ $X2=4.85 $Y2=1.7
r170 43 45 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.755 $Y=1.7
+ $X2=3.93 $Y2=1.7
r171 39 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.16
r172 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.985
r173 36 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=1.16
r174 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=0.56
r175 32 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.16
r176 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.985
r177 29 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=1.16
r178 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=0.56
r179 25 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.16
r180 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.985
r181 22 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=1.16
r182 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=0.56
r183 18 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=1.325
+ $X2=5.54 $Y2=1.16
r184 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.54 $Y=1.325
+ $X2=5.54 $Y2=1.985
r185 15 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=0.995
+ $X2=5.54 $Y2=1.16
r186 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.54 $Y=0.995
+ $X2=5.54 $Y2=0.56
r187 11 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.7 $Y=1.865
+ $X2=3.7 $Y2=1.7
r188 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.7 $Y=1.865
+ $X2=3.7 $Y2=2.275
r189 7 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.7 $Y=1.535
+ $X2=3.7 $Y2=1.7
r190 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.7 $Y=1.535 $X2=3.7
+ $Y2=0.445
r191 2 66 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=1.485 $X2=4.85 $Y2=1.755
r192 2 56 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=1.485 $X2=4.85 $Y2=2.27
r193 1 50 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.235 $X2=4.43 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%A_562_413# 1 2 9 13 15 16 17 21 26 27 28 31
c84 31 0 1.05688e-19 $X=4.15 $Y=1.16
c85 27 0 1.65126e-19 $X=3.57 $Y=1.325
r86 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.15
+ $Y=1.16 $X2=4.15 $Y2=1.16
r87 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.655 $Y=1.16
+ $X2=4.15 $Y2=1.16
r88 27 29 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.57 $Y=1.325
+ $X2=3.495 $Y2=1.16
r89 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=2.255
r90 26 29 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.42 $Y=0.995
+ $X2=3.495 $Y2=1.16
r91 25 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.42 $Y=0.535
+ $X2=3.42 $Y2=0.995
r92 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.485 $Y=2.34
+ $X2=3.57 $Y2=2.255
r93 21 23 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.485 $Y=2.34
+ $X2=3.07 $Y2=2.34
r94 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.45
+ $X2=3.42 $Y2=0.535
r95 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.335 $Y=0.45
+ $X2=3.01 $Y2=0.45
r96 15 32 92.2021 $w=2.7e-07 $l=4.15e-07 $layer=POLY_cond $X=4.565 $Y=1.16
+ $X2=4.15 $Y2=1.16
r97 15 16 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.565 $Y=1.16
+ $X2=4.64 $Y2=1.16
r98 11 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.64 $Y=1.295
+ $X2=4.64 $Y2=1.16
r99 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.64 $Y=1.295
+ $X2=4.64 $Y2=1.985
r100 7 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.64 $Y=1.025
+ $X2=4.64 $Y2=1.16
r101 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.64 $Y=1.025
+ $X2=4.64 $Y2=0.56
r102 2 23 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.065 $X2=3.07 $Y2=2.34
r103 1 19 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.01 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%RESET_B 1 3 6 8 11 12
c40 11 0 1.05688e-19 $X=5.06 $Y=1.16
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.06
+ $Y=1.16 $X2=5.06 $Y2=1.16
r42 8 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.88 $Y=1.16 $X2=5.06
+ $Y2=1.16
r43 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.325
+ $X2=5.06 $Y2=1.16
r44 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.06 $Y=1.325 $X2=5.06
+ $Y2=1.985
r45 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=0.995
+ $X2=5.06 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.06 $Y=0.995 $X2=5.06
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%VPWR 1 2 3 4 5 6 7 24 28 32 34 38 42 44 48
+ 52 54 58 60 65 70 78 83 89 92 95 98 101 104 108
c120 42 0 1.81835e-20 $X=5.3 $Y=2.02
r121 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r122 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r123 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r124 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r125 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r126 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r128 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r129 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 87 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r131 87 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r132 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r133 84 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.405 $Y=2.72
+ $X2=6.27 $Y2=2.72
r134 84 86 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=2.72
+ $X2=6.67 $Y2=2.72
r135 83 107 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=7.152 $Y2=2.72
r136 83 86 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=6.67 $Y2=2.72
r137 82 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r138 82 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r139 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r140 79 98 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.585 $Y=2.72
+ $X2=4.445 $Y2=2.72
r141 79 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.585 $Y=2.72
+ $X2=4.83 $Y2=2.72
r142 78 101 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.115 $Y=2.72
+ $X2=5.3 $Y2=2.72
r143 78 81 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.115 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 77 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r145 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r146 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r147 74 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r148 73 76 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r149 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r150 71 92 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.117 $Y2=2.72
r151 71 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.53 $Y2=2.72
r152 70 95 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.97 $Y2=2.72
r153 70 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.45 $Y2=2.72
r154 69 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r155 69 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r156 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r157 66 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r158 66 68 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r159 65 92 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.96 $Y=2.72
+ $X2=2.117 $Y2=2.72
r160 65 68 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.96 $Y=2.72
+ $X2=1.61 $Y2=2.72
r161 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r162 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r163 58 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r164 58 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r165 54 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.11 $Y=1.66
+ $X2=7.11 $Y2=2.34
r166 52 107 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.11 $Y=2.635
+ $X2=7.152 $Y2=2.72
r167 52 57 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.11 $Y=2.635
+ $X2=7.11 $Y2=2.34
r168 48 51 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.27 $Y=1.66
+ $X2=6.27 $Y2=2.34
r169 46 104 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=2.635
+ $X2=6.27 $Y2=2.72
r170 46 51 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.27 $Y=2.635
+ $X2=6.27 $Y2=2.34
r171 45 101 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.3 $Y2=2.72
r172 44 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.135 $Y=2.72
+ $X2=6.27 $Y2=2.72
r173 44 45 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.135 $Y=2.72
+ $X2=5.485 $Y2=2.72
r174 40 101 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r175 40 42 19.1555 $w=3.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.02
r176 36 98 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=2.635
+ $X2=4.445 $Y2=2.72
r177 36 38 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.445 $Y=2.635
+ $X2=4.445 $Y2=2.34
r178 35 95 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.115 $Y=2.72
+ $X2=3.97 $Y2=2.72
r179 34 98 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.445 $Y2=2.72
r180 34 35 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.115 $Y2=2.72
r181 30 95 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.72
r182 30 32 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.3
r183 26 92 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.117 $Y=2.635
+ $X2=2.117 $Y2=2.72
r184 26 28 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.117 $Y=2.635
+ $X2=2.117 $Y2=2
r185 22 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r186 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r187 7 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=2.34
r188 7 54 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=1.66
r189 6 51 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.22 $Y2=2.34
r190 6 48 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.22 $Y2=1.66
r191 5 42 300 $w=1.7e-07 $l=6.11964e-07 $layer=licon1_PDIFF $count=2 $X=5.135
+ $Y=1.485 $X2=5.3 $Y2=2.02
r192 4 38 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.485 $X2=4.43 $Y2=2.34
r193 3 32 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.775
+ $Y=2.065 $X2=3.91 $Y2=2.3
r194 2 28 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.91
+ $Y=1.845 $X2=2.045 $Y2=2
r195 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%Q 1 2 3 4 14 19 24 26 27 29 30 31 33 35 50
+ 56
r60 50 59 2.13585 $w=5.58e-07 $l=1e-07 $layer=LI1_cond $X=6.575 $Y=1.045
+ $X2=6.675 $Y2=1.045
r61 33 35 9.82493 $w=5.58e-07 $l=4.6e-07 $layer=LI1_cond $X=6.72 $Y=1.045
+ $X2=7.18 $Y2=1.045
r62 33 59 0.961134 $w=5.58e-07 $l=4.5e-08 $layer=LI1_cond $X=6.72 $Y=1.045
+ $X2=6.675 $Y2=1.045
r63 33 59 6.84897 $w=2e-07 $l=2.8e-07 $layer=LI1_cond $X=6.675 $Y=0.765
+ $X2=6.675 $Y2=1.045
r64 33 56 11.2591 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=6.675 $Y=0.765
+ $X2=6.675 $Y2=0.49
r65 31 50 6.72794 $w=5.58e-07 $l=3.15e-07 $layer=LI1_cond $X=6.26 $Y=1.045
+ $X2=6.575 $Y2=1.045
r66 30 48 3.63929 $w=2.83e-07 $l=9e-08 $layer=LI1_cond $X=5.822 $Y=2.21
+ $X2=5.822 $Y2=2.3
r67 28 31 6.30077 $w=5.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.965 $Y=1.045
+ $X2=6.26 $Y2=1.045
r68 28 29 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=1.045
+ $X2=5.88 $Y2=1.045
r69 26 30 7.80426 $w=2.83e-07 $l=1.93e-07 $layer=LI1_cond $X=5.822 $Y=2.017
+ $X2=5.822 $Y2=2.21
r70 26 27 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=5.822 $Y=2.017
+ $X2=5.822 $Y2=1.875
r71 22 24 5.26115 $w=2.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.775 $Y=0.37
+ $X2=5.88 $Y2=0.37
r72 17 59 6.84897 $w=2e-07 $l=2.8e-07 $layer=LI1_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=1.045
r73 17 19 35.2136 $w=1.98e-07 $l=6.35e-07 $layer=LI1_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=1.96
r74 15 29 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=5.88 $Y=1.325
+ $X2=5.88 $Y2=1.045
r75 15 27 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.88 $Y=1.325
+ $X2=5.88 $Y2=1.875
r76 14 29 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=5.88 $Y=0.765
+ $X2=5.88 $Y2=1.045
r77 13 24 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.88 $Y=0.485
+ $X2=5.88 $Y2=0.37
r78 13 14 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.88 $Y=0.485
+ $X2=5.88 $Y2=0.765
r79 4 19 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=6.505
+ $Y=1.485 $X2=6.66 $Y2=1.96
r80 3 48 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.615
+ $Y=1.485 $X2=5.765 $Y2=2.3
r81 2 56 182 $w=1.7e-07 $l=3.23342e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.66 $Y2=0.49
r82 1 22 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=5.615
+ $Y=0.235 $X2=5.775 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTP_4%VGND 1 2 3 4 5 6 21 25 29 33 35 39 41 43 45
+ 47 52 57 65 70 76 79 82 85 88 92
c126 92 0 2.71124e-20 $X=7.13 $Y=0
c127 2 0 7.13094e-20 $X=1.91 $Y=0.235
r128 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r129 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r130 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r131 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r132 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r133 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r134 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r135 74 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r136 74 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r137 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r138 71 88 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.27
+ $Y2=0
r139 71 73 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=0
+ $X2=6.67 $Y2=0
r140 70 91 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=7.152 $Y2=0
r141 70 73 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=6.67 $Y2=0
r142 69 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r143 69 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r144 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r145 66 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=0 $X2=3.91
+ $Y2=0
r146 66 68 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.075 $Y=0
+ $X2=4.83 $Y2=0
r147 65 85 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=5.27
+ $Y2=0
r148 65 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=4.83
+ $Y2=0
r149 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r150 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r151 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r152 61 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r153 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r154 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r155 58 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.045
+ $Y2=0
r156 58 60 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.53
+ $Y2=0
r157 57 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.91
+ $Y2=0
r158 57 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.45
+ $Y2=0
r159 56 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r160 56 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r161 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r162 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r163 53 55 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r164 52 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.045
+ $Y2=0
r165 52 55 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.61
+ $Y2=0
r166 47 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r167 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r168 45 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r169 45 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r170 41 91 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.11 $Y=0.085
+ $X2=7.152 $Y2=0
r171 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.11 $Y=0.085
+ $X2=7.11 $Y2=0.38
r172 37 88 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0
r173 37 39 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0.38
r174 36 85 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.27
+ $Y2=0
r175 35 88 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.135 $Y=0 $X2=6.27
+ $Y2=0
r176 35 36 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.135 $Y=0
+ $X2=5.44 $Y2=0
r177 31 85 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=0.085
+ $X2=5.27 $Y2=0
r178 31 33 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=5.27 $Y=0.085
+ $X2=5.27 $Y2=0.36
r179 27 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=0.085
+ $X2=3.91 $Y2=0
r180 27 29 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.91 $Y=0.085
+ $X2=3.91 $Y2=0.445
r181 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r182 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.36
r183 19 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r184 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r185 6 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.965
+ $Y=0.235 $X2=7.1 $Y2=0.38
r186 5 39 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.235 $X2=6.22 $Y2=0.38
r187 4 33 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.135
+ $Y=0.235 $X2=5.275 $Y2=0.36
r188 3 29 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.775
+ $Y=0.235 $X2=3.91 $Y2=0.445
r189 2 25 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.235 $X2=2.045 $Y2=0.36
r190 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


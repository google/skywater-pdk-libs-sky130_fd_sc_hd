* File: sky130_fd_sc_hd__nor3b_1.pxi.spice
* Created: Tue Sep  1 19:18:37 2020
* 
x_PM_SKY130_FD_SC_HD__NOR3B_1%A_91_199# N_A_91_199#_M1004_d N_A_91_199#_M1001_d
+ N_A_91_199#_M1006_g N_A_91_199#_M1003_g N_A_91_199#_c_48_n N_A_91_199#_c_49_n
+ N_A_91_199#_c_50_n N_A_91_199#_c_57_n N_A_91_199#_c_94_p N_A_91_199#_c_51_n
+ N_A_91_199#_c_52_n N_A_91_199#_c_53_n PM_SKY130_FD_SC_HD__NOR3B_1%A_91_199#
x_PM_SKY130_FD_SC_HD__NOR3B_1%B N_B_c_111_n N_B_M1000_g N_B_M1002_g B
+ N_B_c_113_n PM_SKY130_FD_SC_HD__NOR3B_1%B
x_PM_SKY130_FD_SC_HD__NOR3B_1%A N_A_M1007_g N_A_M1005_g A N_A_c_149_n
+ N_A_c_150_n PM_SKY130_FD_SC_HD__NOR3B_1%A
x_PM_SKY130_FD_SC_HD__NOR3B_1%C_N N_C_N_M1004_g N_C_N_M1001_g C_N N_C_N_c_183_n
+ N_C_N_c_184_n PM_SKY130_FD_SC_HD__NOR3B_1%C_N
x_PM_SKY130_FD_SC_HD__NOR3B_1%Y N_Y_M1006_s N_Y_M1000_d N_Y_M1003_s N_Y_c_216_n
+ N_Y_c_237_p N_Y_c_212_n Y Y PM_SKY130_FD_SC_HD__NOR3B_1%Y
x_PM_SKY130_FD_SC_HD__NOR3B_1%VPWR N_VPWR_M1005_d N_VPWR_c_251_n N_VPWR_c_252_n
+ N_VPWR_c_253_n VPWR N_VPWR_c_254_n N_VPWR_c_250_n
+ PM_SKY130_FD_SC_HD__NOR3B_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR3B_1%VGND N_VGND_M1006_d N_VGND_M1007_d N_VGND_c_277_n
+ N_VGND_c_278_n N_VGND_c_279_n N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n
+ VGND N_VGND_c_283_n N_VGND_c_284_n PM_SKY130_FD_SC_HD__NOR3B_1%VGND
cc_1 VNB N_A_91_199#_c_48_n 0.0040678f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.16
cc_2 VNB N_A_91_199#_c_49_n 0.0283018f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_3 VNB N_A_91_199#_c_50_n 3.54687e-19 $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.785
cc_4 VNB N_A_91_199#_c_51_n 0.0233028f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.785
cc_5 VNB N_A_91_199#_c_52_n 0.0206355f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=0.66
cc_6 VNB N_A_91_199#_c_53_n 0.019682f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.995
cc_7 VNB N_B_c_111_n 0.0162214f $X=-0.19 $Y=-0.24 $X2=2.13 $Y2=0.465
cc_8 VNB B 0.00271558f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_9 VNB N_B_c_113_n 0.0203512f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_10 VNB A 0.00611623f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_11 VNB N_A_c_149_n 0.0186156f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_12 VNB N_A_c_150_n 0.0185094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB C_N 0.00371265f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_14 VNB N_C_N_c_183_n 0.027206f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_15 VNB N_C_N_c_184_n 0.0203182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_212_n 0.0298186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB Y 0.0234854f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.87
cc_18 VNB N_VPWR_c_250_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.87
cc_19 VNB N_VGND_c_277_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_20 VNB N_VGND_c_278_n 0.00772861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_279_n 0.020151f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_22 VNB N_VGND_c_280_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_23 VNB N_VGND_c_281_n 0.0119183f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.245
cc_24 VNB N_VGND_c_282_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0.8 $Y2=1.785
cc_25 VNB N_VGND_c_283_n 0.0254957f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.995
cc_26 VNB N_VGND_c_284_n 0.173814f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.325
cc_27 VPB N_A_91_199#_M1003_g 0.0229082f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_28 VPB N_A_91_199#_c_49_n 0.00920264f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_29 VPB N_A_91_199#_c_50_n 0.00110724f $X=-0.19 $Y=1.305 $X2=0.8 $Y2=1.785
cc_30 VPB N_A_91_199#_c_57_n 0.017676f $X=-0.19 $Y=1.305 $X2=2.505 $Y2=1.87
cc_31 VPB N_A_91_199#_c_51_n 0.0234353f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.785
cc_32 VPB N_B_M1002_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB B 0.00212139f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_34 VPB N_B_c_113_n 0.00459538f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_35 VPB N_A_M1005_g 0.01942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB A 0.00221894f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_37 VPB N_A_c_149_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_38 VPB N_C_N_M1001_g 0.0367424f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB C_N 0.00489538f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_40 VPB N_C_N_c_183_n 0.00491111f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_41 VPB Y 0.0217075f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.87
cc_42 VPB Y 0.0392564f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.87
cc_43 VPB N_VPWR_c_251_n 0.0149263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_252_n 0.0482637f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_45 VPB N_VPWR_c_253_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.325
cc_46 VPB N_VPWR_c_254_n 0.0280782f $X=-0.19 $Y=1.305 $X2=2.505 $Y2=1.87
cc_47 VPB N_VPWR_c_250_n 0.0542793f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.87
cc_48 N_A_91_199#_c_53_n N_B_c_111_n 0.0260708f $X=0.63 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_49 N_A_91_199#_M1003_g N_B_M1002_g 0.0615749f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_91_199#_c_50_n N_B_M1002_g 0.00429358f $X=0.8 $Y=1.785 $X2=0 $Y2=0
cc_51 N_A_91_199#_c_57_n N_B_M1002_g 0.0115072f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_52 N_A_91_199#_M1003_g B 5.29605e-19 $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_53 N_A_91_199#_c_48_n B 0.0130107f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_54 N_A_91_199#_c_49_n B 7.60779e-19 $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_91_199#_c_50_n B 0.0219518f $X=0.8 $Y=1.785 $X2=0 $Y2=0
cc_56 N_A_91_199#_c_57_n B 0.0131145f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_57 N_A_91_199#_c_48_n N_B_c_113_n 0.00107792f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_91_199#_c_49_n N_B_c_113_n 0.02071f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_91_199#_c_50_n N_B_c_113_n 4.52901e-19 $X=0.8 $Y=1.785 $X2=0 $Y2=0
cc_60 N_A_91_199#_c_57_n N_B_c_113_n 9.49193e-19 $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_61 N_A_91_199#_c_57_n N_A_M1005_g 0.0116292f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_62 N_A_91_199#_c_57_n A 0.0203818f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_63 N_A_91_199#_c_57_n N_A_c_149_n 3.7381e-19 $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_64 N_A_91_199#_c_57_n N_C_N_M1001_g 0.00982299f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_65 N_A_91_199#_c_51_n N_C_N_M1001_g 0.00447475f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_66 N_A_91_199#_c_57_n C_N 0.0256345f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_67 N_A_91_199#_c_51_n C_N 0.0494531f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_68 N_A_91_199#_c_52_n C_N 0.0130216f $X=2.265 $Y=0.66 $X2=0 $Y2=0
cc_69 N_A_91_199#_c_57_n N_C_N_c_183_n 3.55624e-19 $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_70 N_A_91_199#_c_51_n N_C_N_c_183_n 0.00183894f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_71 N_A_91_199#_c_52_n N_C_N_c_183_n 0.00147244f $X=2.265 $Y=0.66 $X2=0 $Y2=0
cc_72 N_A_91_199#_c_51_n N_C_N_c_184_n 0.00424702f $X=2.59 $Y=1.785 $X2=0 $Y2=0
cc_73 N_A_91_199#_c_52_n N_C_N_c_184_n 0.00137912f $X=2.265 $Y=0.66 $X2=0 $Y2=0
cc_74 N_A_91_199#_c_48_n N_Y_c_216_n 0.0127182f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_91_199#_c_53_n N_Y_c_216_n 0.0125238f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_91_199#_c_48_n N_Y_c_212_n 0.0102716f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_91_199#_c_49_n N_Y_c_212_n 0.00360515f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_91_199#_M1003_g Y 0.0196026f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_91_199#_c_48_n Y 0.0223568f $X=0.715 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_91_199#_c_49_n Y 0.00832901f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_91_199#_c_50_n Y 0.0309037f $X=0.8 $Y=1.785 $X2=0 $Y2=0
cc_82 N_A_91_199#_c_53_n Y 0.00320726f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_91_199#_c_94_p Y 0.0143562f $X=0.885 $Y=1.87 $X2=0 $Y2=0
cc_84 N_A_91_199#_c_50_n A_161_297# 0.0031068f $X=0.8 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_91_199#_c_57_n A_161_297# 0.00741519f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_91_199#_c_94_p A_161_297# 4.90802e-19 $X=0.885 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_91_199#_c_57_n A_245_297# 0.00826124f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_91_199#_c_57_n N_VPWR_M1005_d 0.00757029f $X=2.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_91_199#_c_57_n N_VPWR_c_251_n 0.0205834f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_90 N_A_91_199#_M1003_g N_VPWR_c_252_n 0.00585385f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_91 N_A_91_199#_M1003_g N_VPWR_c_250_n 0.00912169f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_92 N_A_91_199#_c_57_n N_VPWR_c_250_n 0.0530816f $X=2.505 $Y=1.87 $X2=0 $Y2=0
cc_93 N_A_91_199#_c_94_p N_VPWR_c_250_n 0.0063769f $X=0.885 $Y=1.87 $X2=0 $Y2=0
cc_94 N_A_91_199#_c_53_n N_VGND_c_277_n 0.00853411f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_91_199#_c_52_n N_VGND_c_278_n 0.00374012f $X=2.265 $Y=0.66 $X2=0 $Y2=0
cc_96 N_A_91_199#_c_53_n N_VGND_c_279_n 0.00341689f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_91_199#_c_52_n N_VGND_c_283_n 0.0120161f $X=2.265 $Y=0.66 $X2=0 $Y2=0
cc_98 N_A_91_199#_c_52_n N_VGND_c_284_n 0.0152762f $X=2.265 $Y=0.66 $X2=0 $Y2=0
cc_99 N_A_91_199#_c_53_n N_VGND_c_284_n 0.0051968f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B_M1002_g N_A_M1005_g 0.0627989f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B_M1002_g A 5.5215e-19 $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_102 B A 0.0448494f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B_c_113_n A 0.00104218f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_104 B N_A_c_149_n 0.00189405f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_105 N_B_c_113_n N_A_c_149_n 0.0213684f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B_c_111_n N_A_c_150_n 0.0241358f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B_c_111_n N_Y_c_216_n 0.010671f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_108 B N_Y_c_216_n 0.0160356f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B_c_113_n N_Y_c_216_n 0.00114084f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_110 B A_245_297# 0.00135064f $X=1.065 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_111 N_B_M1002_g N_VPWR_c_251_n 0.00282002f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B_M1002_g N_VPWR_c_252_n 0.00585385f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B_M1002_g N_VPWR_c_250_n 0.00625469f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B_c_111_n N_VGND_c_277_n 0.00720306f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_111_n N_VGND_c_278_n 8.38908e-19 $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B_c_111_n N_VGND_c_281_n 0.00341689f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_111_n N_VGND_c_284_n 0.00405445f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_M1005_g N_C_N_M1001_g 0.0285585f $X=1.57 $Y=1.985 $X2=0 $Y2=0
cc_119 A N_C_N_M1001_g 0.00190954f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A_M1005_g C_N 2.82283e-19 $X=1.57 $Y=1.985 $X2=0 $Y2=0
cc_121 A C_N 0.0492394f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_c_149_n C_N 3.66689e-19 $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_123 A N_C_N_c_183_n 0.0018697f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_c_149_n N_C_N_c_183_n 0.0202813f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_150_n N_C_N_c_184_n 0.0125721f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_126 A N_VPWR_M1005_d 0.00233761f $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_127 N_A_M1005_g N_VPWR_c_251_n 0.0146914f $X=1.57 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_VPWR_c_252_n 0.0046653f $X=1.57 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1005_g N_VPWR_c_250_n 0.00427441f $X=1.57 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_c_150_n N_VGND_c_277_n 6.77973e-19 $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_131 A N_VGND_c_278_n 0.0147164f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A_c_149_n N_VGND_c_278_n 7.77033e-19 $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_c_150_n N_VGND_c_278_n 0.0118668f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_150_n N_VGND_c_281_n 0.0046653f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_150_n N_VGND_c_284_n 0.00799591f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_136 N_C_N_M1001_g N_VPWR_c_251_n 0.00214007f $X=2.055 $Y=1.86 $X2=0 $Y2=0
cc_137 N_C_N_M1001_g N_VPWR_c_254_n 0.00402388f $X=2.055 $Y=1.86 $X2=0 $Y2=0
cc_138 N_C_N_M1001_g N_VPWR_c_250_n 0.00459843f $X=2.055 $Y=1.86 $X2=0 $Y2=0
cc_139 N_C_N_c_184_n N_VGND_c_278_n 0.00441624f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_140 N_C_N_c_184_n N_VGND_c_283_n 0.00510437f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_141 N_C_N_c_184_n N_VGND_c_284_n 0.00512902f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_142 Y N_VPWR_c_252_n 0.0306029f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_143 N_Y_M1003_s N_VPWR_c_250_n 0.0064064f $X=0.335 $Y=1.485 $X2=0 $Y2=0
cc_144 Y N_VPWR_c_250_n 0.017555f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_145 N_Y_c_216_n N_VGND_M1006_d 0.00685192f $X=1.275 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_146 N_Y_c_216_n N_VGND_c_277_n 0.0160613f $X=1.275 $Y=0.74 $X2=0 $Y2=0
cc_147 N_Y_c_216_n N_VGND_c_279_n 0.0023303f $X=1.275 $Y=0.74 $X2=0 $Y2=0
cc_148 N_Y_c_212_n N_VGND_c_279_n 0.0362203f $X=0.44 $Y=0.39 $X2=0 $Y2=0
cc_149 N_Y_c_216_n N_VGND_c_281_n 0.00232396f $X=1.275 $Y=0.74 $X2=0 $Y2=0
cc_150 N_Y_c_237_p N_VGND_c_281_n 0.00825814f $X=1.36 $Y=0.495 $X2=0 $Y2=0
cc_151 N_Y_M1006_s N_VGND_c_284_n 0.00294593f $X=0.315 $Y=0.235 $X2=0 $Y2=0
cc_152 N_Y_M1000_d N_VGND_c_284_n 0.00415164f $X=1.225 $Y=0.235 $X2=0 $Y2=0
cc_153 N_Y_c_216_n N_VGND_c_284_n 0.009721f $X=1.275 $Y=0.74 $X2=0 $Y2=0
cc_154 N_Y_c_237_p N_VGND_c_284_n 0.00623764f $X=1.36 $Y=0.495 $X2=0 $Y2=0
cc_155 N_Y_c_212_n N_VGND_c_284_n 0.0198876f $X=0.44 $Y=0.39 $X2=0 $Y2=0
cc_156 A_161_297# N_VPWR_c_250_n 0.0036705f $X=0.805 $Y=1.485 $X2=0.885 $Y2=1.87
cc_157 A_245_297# N_VPWR_c_250_n 0.0036717f $X=1.225 $Y=1.485 $X2=0.885 $Y2=1.87

* File: sky130_fd_sc_hd__inv_1.pex.spice
* Created: Thu Aug 27 14:22:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_1%A 1 3 6 8 14
r22 11 14 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.485 $Y=1.16
+ $X2=0.675 $Y2=1.16
r23 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.16 $X2=0.485 $Y2=1.16
r24 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=1.325
+ $X2=0.675 $Y2=1.16
r25 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.675 $Y=1.325
+ $X2=0.675 $Y2=1.985
r26 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.675 $Y2=1.16
r27 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.675 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_1%VPWR 1 6 11 12 13 20 21
r14 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r15 13 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r16 13 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r17 11 16 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.34 $Y=2.72
+ $X2=0.23 $Y2=2.72
r18 11 12 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.34 $Y=2.72
+ $X2=0.445 $Y2=2.72
r19 10 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=1.15
+ $Y2=2.72
r20 10 12 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.55 $Y=2.72
+ $X2=0.445 $Y2=2.72
r21 6 9 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.445 $Y=1.66
+ $X2=0.445 $Y2=2.34
r22 4 12 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=2.635
+ $X2=0.445 $Y2=2.72
r23 4 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.445 $Y=2.635
+ $X2=0.445 $Y2=2.34
r24 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.485 $X2=0.465 $Y2=2.34
r25 1 6 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.485 $X2=0.465 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__INV_1%Y 1 2 9 13 18 19 20 29
r19 29 30 2.64191 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.885 $Y=1.53
+ $X2=0.885 $Y2=1.485
r20 20 29 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=0.885 $Y=1.55
+ $X2=0.885 $Y2=1.53
r21 20 30 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=0.935 $Y=1.465
+ $X2=0.935 $Y2=1.485
r22 19 20 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.935 $Y=1.19
+ $X2=0.935 $Y2=1.465
r23 18 19 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.935 $Y=0.885
+ $X2=0.935 $Y2=1.19
r24 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.885 $Y=1.66
+ $X2=0.885 $Y2=2.34
r25 11 20 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.885 $Y=1.65
+ $X2=0.885 $Y2=1.55
r26 11 13 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.885 $Y=1.65
+ $X2=0.885 $Y2=1.66
r27 7 18 6.83261 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0.72
+ $X2=0.885 $Y2=0.885
r28 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.885 $Y=0.72
+ $X2=0.885 $Y2=0.4
r29 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=1.485 $X2=0.885 $Y2=2.34
r30 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=1.485 $X2=0.885 $Y2=1.66
r31 1 9 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.75
+ $Y=0.235 $X2=0.885 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__INV_1%VGND 1 6 9 10 11 18 19
r14 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r15 11 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r16 11 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r17 9 14 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.23
+ $Y2=0
r18 9 10 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.435
+ $Y2=0
r19 8 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=1.15
+ $Y2=0
r20 8 10 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.435
+ $Y2=0
r21 4 10 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.435 $Y=0.085
+ $X2=0.435 $Y2=0
r22 4 6 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.435 $Y=0.085
+ $X2=0.435 $Y2=0.4
r23 1 6 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.34
+ $Y=0.235 $X2=0.465 $Y2=0.4
.ends


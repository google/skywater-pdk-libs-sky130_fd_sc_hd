# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__buf_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 2.485000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 0.255000  3.285000 0.260000 ;
        RECT 3.035000 0.260000  3.365000 0.735000 ;
        RECT 3.035000 0.735000 10.035000 0.905000 ;
        RECT 3.035000 1.445000 10.035000 1.615000 ;
        RECT 3.035000 1.615000  3.365000 2.465000 ;
        RECT 3.875000 0.260000  4.205000 0.735000 ;
        RECT 3.875000 1.615000  4.205000 2.465000 ;
        RECT 3.955000 0.255000  4.125000 0.260000 ;
        RECT 4.715000 0.260000  5.045000 0.735000 ;
        RECT 4.715000 1.615000  5.045000 2.465000 ;
        RECT 4.795000 0.255000  4.965000 0.260000 ;
        RECT 5.555000 0.260000  5.885000 0.735000 ;
        RECT 5.555000 1.615000  5.885000 2.465000 ;
        RECT 6.395000 0.260000  6.725000 0.735000 ;
        RECT 6.395000 1.615000  6.725000 2.465000 ;
        RECT 7.235000 0.260000  7.565000 0.735000 ;
        RECT 7.235000 1.615000  7.565000 2.465000 ;
        RECT 8.075000 0.260000  8.405000 0.735000 ;
        RECT 8.075000 1.615000  8.405000 2.465000 ;
        RECT 8.915000 0.260000  9.245000 0.735000 ;
        RECT 8.915000 1.615000  9.245000 2.465000 ;
        RECT 9.655000 0.905000 10.035000 1.445000 ;
        RECT 9.760000 0.365000 10.035000 0.735000 ;
        RECT 9.760000 1.615000 10.035000 2.360000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.175000  0.085000  0.345000 0.905000 ;
        RECT 1.015000  0.085000  1.185000 0.565000 ;
        RECT 1.855000  0.085000  2.025000 0.565000 ;
        RECT 2.695000  0.085000  2.865000 0.565000 ;
        RECT 3.535000  0.085000  3.705000 0.565000 ;
        RECT 4.375000  0.085000  4.545000 0.565000 ;
        RECT 5.215000  0.085000  5.385000 0.565000 ;
        RECT 6.055000  0.085000  6.225000 0.565000 ;
        RECT 6.895000  0.085000  7.065000 0.565000 ;
        RECT 7.735000  0.085000  7.905000 0.565000 ;
        RECT 8.575000  0.085000  8.745000 0.565000 ;
        RECT 9.415000  0.085000  9.585000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
        RECT 9.805000 -0.085000 9.975000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.175000 1.445000  0.345000 2.635000 ;
        RECT 1.015000 1.835000  1.185000 2.635000 ;
        RECT 1.855000 1.835000  2.025000 2.635000 ;
        RECT 2.695000 1.835000  2.865000 2.635000 ;
        RECT 3.535000 1.835000  3.705000 2.635000 ;
        RECT 4.375000 1.835000  4.545000 2.635000 ;
        RECT 5.215000 1.835000  5.385000 2.635000 ;
        RECT 6.055000 1.835000  6.225000 2.635000 ;
        RECT 6.895000 1.835000  7.065000 2.635000 ;
        RECT 7.735000 1.835000  7.905000 2.635000 ;
        RECT 8.575000 1.835000  8.745000 2.635000 ;
        RECT 9.415000 1.835000  9.585000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
        RECT 9.805000 2.635000 9.975000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 0.260000 0.845000 0.735000 ;
      RECT 0.515000 0.735000 2.865000 0.905000 ;
      RECT 0.515000 1.445000 2.865000 1.615000 ;
      RECT 0.515000 1.615000 0.845000 2.465000 ;
      RECT 1.355000 0.260000 1.685000 0.735000 ;
      RECT 1.355000 1.615000 1.685000 2.465000 ;
      RECT 2.195000 0.260000 2.525000 0.735000 ;
      RECT 2.195000 1.615000 2.525000 2.465000 ;
      RECT 2.690000 0.905000 2.865000 1.075000 ;
      RECT 2.690000 1.075000 9.410000 1.275000 ;
      RECT 2.690000 1.275000 2.865000 1.445000 ;
  END
END sky130_fd_sc_hd__buf_16

* File: sky130_fd_sc_hd__o32a_2.spice.pex
* Created: Thu Aug 27 14:40:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O32A_2%A_79_21# 1 2 7 9 12 14 16 19 23 24 26 27 30
+ 32 35 36 40
c84 36 0 1.52385e-19 $X=2.86 $Y=1.87
c85 23 0 4.0869e-20 $X=1.1 $Y=1.16
r86 42 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r87 38 40 3.2569 $w=2.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.36 $Y=0.71
+ $X2=3.425 $Y2=0.71
r88 34 40 1.55539 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=3.425 $Y=0.825
+ $X2=3.425 $Y2=0.71
r89 34 35 53.2364 $w=1.98e-07 $l=9.6e-07 $layer=LI1_cond $X=3.425 $Y=0.825
+ $X2=3.425 $Y2=1.785
r90 33 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=1.87
+ $X2=2.86 $Y2=1.87
r91 32 35 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.325 $Y=1.87
+ $X2=3.425 $Y2=1.785
r92 32 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.325 $Y=1.87
+ $X2=3.025 $Y2=1.87
r93 28 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=1.955
+ $X2=2.86 $Y2=1.87
r94 28 30 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.86 $Y=1.955
+ $X2=2.86 $Y2=2
r95 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=1.87
+ $X2=2.86 $Y2=1.87
r96 26 27 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=2.695 $Y=1.87
+ $X2=1.325 $Y2=1.87
r97 24 44 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=0.89
+ $Y2=1.16
r98 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r99 21 27 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=1.17 $Y=1.785
+ $X2=1.325 $Y2=1.87
r100 21 23 23.2347 $w=3.08e-07 $l=6.25e-07 $layer=LI1_cond $X=1.17 $Y=1.785
+ $X2=1.17 $Y2=1.16
r101 17 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r102 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r103 14 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r104 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r105 10 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r106 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r107 7 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r108 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r109 2 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.485 $X2=2.86 $Y2=2
r110 1 38 182 $w=1.7e-07 $l=5.82666e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.36 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%A1 3 6 8 11 13
r33 11 14 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.585 $Y2=1.325
r34 11 13 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.585 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.16 $X2=1.58 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.65 $Y=1.985
+ $X2=1.65 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.65 $Y=0.56 $X2=1.65
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%A2 1 3 6 8 11
c39 8 0 4.0869e-20 $X=2.075 $Y=1.19
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.16 $X2=2.07 $Y2=1.16
r41 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.325
+ $X2=2.07 $Y2=1.16
r42 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.07 $Y=1.325 $X2=2.07
+ $Y2=1.985
r43 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=0.995
+ $X2=2.07 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.07 $Y=0.995 $X2=2.07
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%A3 3 6 8 11 13
r38 11 14 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.57 $Y2=1.325
r39 11 13 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.57 $Y2=0.995
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.16 $X2=2.55 $Y2=1.16
r41 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.65 $Y=1.985
+ $X2=2.65 $Y2=1.325
r42 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.65 $Y=0.56 $X2=2.65
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%B2 1 3 6 8 11
c40 11 0 1.52385e-19 $X=3.07 $Y=1.16
r41 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.16 $X2=3.07 $Y2=1.16
r42 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.325
+ $X2=3.07 $Y2=1.16
r43 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.07 $Y=1.325 $X2=3.07
+ $Y2=1.985
r44 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=0.995
+ $X2=3.07 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.07 $Y=0.995 $X2=3.07
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%B1 3 7 9 14
r25 11 14 53.7814 $w=2.9e-07 $l=2.6e-07 $layer=POLY_cond $X=3.6 $Y=1.16 $X2=3.86
+ $Y2=1.16
r26 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.86
+ $Y=1.16 $X2=3.86 $Y2=1.16
r27 5 11 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.6 $Y=1.305 $X2=3.6
+ $Y2=1.16
r28 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.6 $Y=1.305 $X2=3.6
+ $Y2=1.985
r29 1 11 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.6 $Y=1.015 $X2=3.6
+ $Y2=1.16
r30 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.6 $Y=1.015 $X2=3.6
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%VPWR 1 2 3 10 12 16 18 22 24 29 41 49
r48 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r49 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 41 44 10.0846 $w=5.08e-07 $l=4.3e-07 $layer=LI1_cond $X=1.27 $Y=2.29
+ $X2=1.27 $Y2=2.72
r51 36 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r52 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 33 36 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 33 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 32 35 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 30 44 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.525 $Y=2.72
+ $X2=1.27 $Y2=2.72
r58 30 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 29 48 5.10352 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.917 $Y2=2.72
r60 29 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 28 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 25 38 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r64 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 24 44 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.27 $Y2=2.72
r66 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 18 21 21.7684 $w=3.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.875 $Y=1.66
+ $X2=3.875 $Y2=2.34
r70 16 48 2.91958 $w=3.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.875 $Y=2.635
+ $X2=3.917 $Y2=2.72
r71 16 21 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.875 $Y=2.635
+ $X2=3.875 $Y2=2.34
r72 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r73 10 38 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r74 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r75 3 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.81 $Y2=2.34
r76 3 18 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.81 $Y2=1.66
r77 2 41 300 $w=1.7e-07 $l=1.01509e-06 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.44 $Y2=2.29
r78 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r79 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%X 1 2 7 8 9 10 11 12 20
r13 12 37 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=2.21
+ $X2=0.68 $Y2=2.34
r14 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=2.21
r15 11 31 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=1.66
r16 10 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=1.53
+ $X2=0.68 $Y2=1.66
r17 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=1.19 $X2=0.68
+ $Y2=1.53
r18 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.85 $X2=0.68
+ $Y2=1.19
r19 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.51 $X2=0.68
+ $Y2=0.85
r20 7 20 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=0.51 $X2=0.68
+ $Y2=0.38
r21 2 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r22 2 31 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r23 1 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%VGND 1 2 3 10 12 14 18 22 25 26 27 37 38 44
r55 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r56 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r57 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r58 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r59 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r60 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r61 32 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r62 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 29 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.26
+ $Y2=0
r64 29 31 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=2.07
+ $Y2=0
r65 27 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r66 27 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r67 25 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.07
+ $Y2=0
r68 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.36
+ $Y2=0
r69 24 34 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.53
+ $Y2=0
r70 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.36
+ $Y2=0
r71 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r72 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.38
r73 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=0.085
+ $X2=1.26 $Y2=0
r74 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.26 $Y=0.085
+ $X2=1.26 $Y2=0.38
r75 15 41 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r76 14 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=0 $X2=1.26
+ $Y2=0
r77 14 15 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.095 $Y=0 $X2=0.345
+ $Y2=0
r78 10 41 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r79 10 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.38
r80 3 22 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.36 $Y2=0.38
r81 2 18 91 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.26 $Y2=0.38
r82 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_2%A_345_47# 1 2 3 12 14 15 16 17 18 25
r52 19 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=0.34
+ $X2=2.86 $Y2=0.34
r53 18 25 5.44966 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.875 $Y2=0.34
r54 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.025 $Y2=0.34
r55 16 23 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.425 $X2=2.86
+ $Y2=0.34
r56 16 17 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.86 $Y=0.425
+ $X2=2.86 $Y2=0.655
r57 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.695 $Y=0.74
+ $X2=2.86 $Y2=0.655
r58 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=0.74
+ $X2=2.025 $Y2=0.74
r59 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.86 $Y=0.655
+ $X2=2.025 $Y2=0.74
r60 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.86 $Y=0.655
+ $X2=1.86 $Y2=0.38
r61 3 25 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.675
+ $Y=0.235 $X2=3.81 $Y2=0.38
r62 2 23 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=0.235 $X2=2.86 $Y2=0.38
r63 1 12 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.725
+ $Y=0.235 $X2=1.86 $Y2=0.38
.ends


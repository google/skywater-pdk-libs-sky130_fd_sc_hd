* File: sky130_fd_sc_hd__o22ai_1.spice.SKY130_FD_SC_HD__O22AI_1.pxi
* Created: Thu Aug 27 14:37:52 2020
* 
x_PM_SKY130_FD_SC_HD__O22AI_1%B1 N_B1_c_44_n N_B1_M1007_g N_B1_M1006_g B1
+ N_B1_c_46_n PM_SKY130_FD_SC_HD__O22AI_1%B1
x_PM_SKY130_FD_SC_HD__O22AI_1%B2 N_B2_M1003_g N_B2_M1005_g N_B2_c_76_n
+ N_B2_c_77_n B2 N_B2_c_78_n PM_SKY130_FD_SC_HD__O22AI_1%B2
x_PM_SKY130_FD_SC_HD__O22AI_1%A2 N_A2_M1004_g N_A2_M1000_g N_A2_c_122_n
+ N_A2_c_123_n N_A2_c_124_n N_A2_c_129_n A2 N_A2_c_125_n
+ PM_SKY130_FD_SC_HD__O22AI_1%A2
x_PM_SKY130_FD_SC_HD__O22AI_1%A1 N_A1_M1001_g N_A1_M1002_g A1 N_A1_c_175_n
+ N_A1_c_176_n PM_SKY130_FD_SC_HD__O22AI_1%A1
x_PM_SKY130_FD_SC_HD__O22AI_1%VPWR N_VPWR_M1006_s N_VPWR_M1001_d N_VPWR_c_202_n
+ N_VPWR_c_203_n N_VPWR_c_204_n N_VPWR_c_205_n VPWR N_VPWR_c_206_n
+ N_VPWR_c_201_n PM_SKY130_FD_SC_HD__O22AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O22AI_1%Y N_Y_M1007_d N_Y_M1003_d N_Y_c_235_n N_Y_c_241_n
+ Y PM_SKY130_FD_SC_HD__O22AI_1%Y
x_PM_SKY130_FD_SC_HD__O22AI_1%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1005_d
+ N_A_27_47#_M1002_d N_A_27_47#_c_269_n N_A_27_47#_c_281_n N_A_27_47#_c_278_n
+ N_A_27_47#_c_270_n N_A_27_47#_c_271_n PM_SKY130_FD_SC_HD__O22AI_1%A_27_47#
x_PM_SKY130_FD_SC_HD__O22AI_1%VGND N_VGND_M1004_d N_VGND_c_311_n VGND
+ N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n
+ PM_SKY130_FD_SC_HD__O22AI_1%VGND
cc_1 VNB N_B1_c_44_n 0.0189108f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB B1 0.0242859f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B1_c_46_n 0.0351735f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B2_c_76_n 3.61466e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_5 VNB N_B2_c_77_n 0.0233554f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_6 VNB N_B2_c_78_n 0.0173583f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=0.85
cc_7 VNB N_A2_c_122_n 6.10894e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_123_n 0.0195481f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_9 VNB N_A2_c_124_n 0.00378985f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_10 VNB N_A2_c_125_n 0.017245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A1 0.0103792f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_12 VNB N_A1_c_175_n 0.0316454f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_13 VNB N_A1_c_176_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_201_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Y_c_235_n 0.00286868f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_16 VNB N_A_27_47#_c_269_n 0.00836668f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_17 VNB N_A_27_47#_c_270_n 0.00773281f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=0.85
cc_18 VNB N_A_27_47#_c_271_n 0.016608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_311_n 0.0046757f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_20 VNB N_VGND_c_312_n 0.0392944f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_21 VNB N_VGND_c_313_n 0.0173701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_314_n 0.142301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_315_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_B1_M1006_g 0.0206978f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_25 VPB B1 0.0270856f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_26 VPB N_B1_c_46_n 0.0116077f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_27 VPB N_B2_M1003_g 0.0194854f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_28 VPB N_B2_c_76_n 0.00106175f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_29 VPB N_B2_c_77_n 0.00486478f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_30 VPB B2 0.00387306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A2_M1000_g 0.0192402f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_32 VPB N_A2_c_122_n 0.00148417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A2_c_123_n 0.00602681f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_34 VPB N_A2_c_129_n 0.00259302f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.16
cc_35 VPB N_A1_M1001_g 0.0247168f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_36 VPB N_A1_c_175_n 0.00630501f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_37 VPB N_VPWR_c_202_n 0.0103382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_203_n 0.00495535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_204_n 0.0110416f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_40 VPB N_VPWR_c_205_n 0.0484563f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_206_n 0.0413545f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.16
cc_42 VPB N_VPWR_c_201_n 0.0428419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_Y_c_235_n 0.00104815f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_44 N_B1_M1006_g N_B2_M1003_g 0.0451122f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_45 N_B1_c_46_n N_B2_c_76_n 3.81697e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_46 N_B1_c_46_n N_B2_c_77_n 0.0451122f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_47 N_B1_M1006_g B2 2.26657e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_48 N_B1_c_44_n N_B2_c_78_n 0.0243847f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_49 B1 N_VPWR_M1006_s 0.011103f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_50 B1 N_VPWR_c_202_n 8.28574e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_51 N_B1_M1006_g N_VPWR_c_203_n 0.00444548f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_52 B1 N_VPWR_c_203_n 0.0151133f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_53 N_B1_M1006_g N_VPWR_c_206_n 0.00533841f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_54 N_B1_M1006_g N_VPWR_c_201_n 0.00986182f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_55 B1 N_VPWR_c_201_n 0.00223595f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_56 N_B1_c_44_n N_Y_c_235_n 0.00297647f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_57 N_B1_M1006_g N_Y_c_235_n 0.00899061f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_58 B1 N_Y_c_235_n 0.0723029f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_59 N_B1_c_46_n N_Y_c_235_n 0.00777743f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_60 N_B1_c_44_n N_Y_c_241_n 0.00365581f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_61 B1 N_Y_c_241_n 0.0121607f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_62 N_B1_M1006_g Y 0.0094833f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_63 B1 Y 0.0124824f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_64 B1 N_A_27_47#_M1007_s 0.00541864f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_65 N_B1_c_44_n N_A_27_47#_c_269_n 0.0112362f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_66 B1 N_A_27_47#_c_269_n 0.0168836f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_B1_c_46_n N_A_27_47#_c_269_n 0.0019308f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B1_c_44_n N_VGND_c_312_n 0.00366111f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B1_c_44_n N_VGND_c_314_n 0.00625137f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B2_M1003_g N_A2_M1000_g 0.0194981f $X=0.845 $Y=1.985 $X2=0 $Y2=0
cc_71 N_B2_c_76_n N_A2_M1000_g 6.0319e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_72 B2 N_A2_M1000_g 0.00213089f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_73 N_B2_c_76_n N_A2_c_122_n 0.00613421f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_74 N_B2_c_77_n N_A2_c_122_n 2.27495e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_75 B2 N_A2_c_122_n 0.00224479f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_76 N_B2_c_76_n N_A2_c_123_n 9.70263e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B2_c_77_n N_A2_c_123_n 0.0207332f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B2_c_76_n N_A2_c_124_n 0.0107814f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B2_c_77_n N_A2_c_124_n 0.00105604f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_80 B2 N_A2_c_124_n 0.00116357f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_81 B2 N_A2_c_129_n 0.0134013f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_82 N_B2_M1003_g A2 6.12942e-19 $X=0.845 $Y=1.985 $X2=0 $Y2=0
cc_83 B2 A2 0.00248342f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_84 N_B2_c_78_n N_A2_c_125_n 0.0182247f $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B2_M1003_g N_VPWR_c_206_n 0.00389338f $X=0.845 $Y=1.985 $X2=0 $Y2=0
cc_86 N_B2_M1003_g N_VPWR_c_201_n 0.005873f $X=0.845 $Y=1.985 $X2=0 $Y2=0
cc_87 B2 N_Y_M1003_d 0.00553586f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_88 N_B2_c_76_n N_Y_c_235_n 0.0300037f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B2_c_77_n N_Y_c_235_n 0.00763253f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_90 B2 N_Y_c_235_n 0.0187725f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_91 N_B2_c_78_n N_Y_c_235_n 0.0028752f $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B2_c_76_n N_Y_c_241_n 6.61482e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B2_c_77_n N_Y_c_241_n 0.00150271f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B2_c_78_n N_Y_c_241_n 0.00201612f $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B2_M1003_g Y 0.0203123f $X=0.845 $Y=1.985 $X2=0 $Y2=0
cc_96 B2 Y 0.0279522f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_97 N_B2_c_76_n N_A_27_47#_c_269_n 0.00434112f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_98 N_B2_c_78_n N_A_27_47#_c_269_n 0.0123138f $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_99 N_B2_c_77_n N_A_27_47#_c_278_n 9.61013e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_100 B2 N_A_27_47#_c_278_n 0.00662755f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_101 N_B2_c_78_n N_A_27_47#_c_278_n 4.59371e-19 $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B2_c_78_n N_VGND_c_312_n 0.00366111f $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B2_c_78_n N_VGND_c_314_n 0.00557587f $X=0.912 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A2_M1000_g N_A1_M1001_g 0.0489861f $X=1.46 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A2_c_129_n N_A1_M1001_g 9.03294e-19 $X=1.625 $Y=1.615 $X2=0 $Y2=0
cc_106 N_A2_c_122_n A1 0.00225656f $X=1.495 $Y=1.445 $X2=0 $Y2=0
cc_107 N_A2_c_123_n A1 2.18433e-19 $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A2_c_124_n A1 0.0138645f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A2_c_122_n N_A1_c_175_n 0.00366606f $X=1.495 $Y=1.445 $X2=0 $Y2=0
cc_110 N_A2_c_123_n N_A1_c_175_n 0.0489861f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A2_c_124_n N_A1_c_175_n 9.73585e-19 $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A2_c_125_n N_A1_c_176_n 0.0275253f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_129_n N_VPWR_c_205_n 0.00777738f $X=1.625 $Y=1.615 $X2=0 $Y2=0
cc_114 N_A2_M1000_g N_VPWR_c_206_n 0.00572457f $X=1.46 $Y=1.985 $X2=0 $Y2=0
cc_115 A2 N_VPWR_c_206_n 0.00775097f $X=1.525 $Y=1.785 $X2=0 $Y2=0
cc_116 N_A2_M1000_g N_VPWR_c_201_n 0.0107958f $X=1.46 $Y=1.985 $X2=0 $Y2=0
cc_117 A2 N_VPWR_c_201_n 0.00735105f $X=1.525 $Y=1.785 $X2=0 $Y2=0
cc_118 N_A2_c_123_n Y 0.00129776f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A2_c_124_n Y 0.0029507f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A2_c_129_n A_307_297# 2.83863e-19 $X=1.625 $Y=1.615 $X2=-0.19 $Y2=-0.24
cc_121 A2 A_307_297# 0.00134964f $X=1.525 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_122 N_A2_c_125_n N_A_27_47#_c_281_n 0.00181398f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A2_c_123_n N_A_27_47#_c_278_n 0.00152966f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A2_c_124_n N_A_27_47#_c_278_n 0.0062425f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A2_c_125_n N_A_27_47#_c_278_n 0.00352259f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_c_124_n N_A_27_47#_c_270_n 0.0123749f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A2_c_129_n N_A_27_47#_c_270_n 0.00389082f $X=1.625 $Y=1.615 $X2=0 $Y2=0
cc_128 N_A2_c_125_n N_A_27_47#_c_270_n 0.00962365f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_125_n N_A_27_47#_c_271_n 5.10226e-19 $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_125_n N_VGND_c_311_n 0.00268723f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_c_125_n N_VGND_c_312_n 0.00429196f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A2_c_125_n N_VGND_c_314_n 0.00601769f $X=1.4 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_M1001_g N_VPWR_c_205_n 0.00564336f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_134 A1 N_VPWR_c_205_n 0.0253819f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A1_c_175_n N_VPWR_c_205_n 0.00444551f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A1_M1001_g N_VPWR_c_206_n 0.00583607f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A1_M1001_g N_VPWR_c_201_n 0.0113033f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_c_176_n N_A_27_47#_c_278_n 4.35843e-19 $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_139 A1 N_A_27_47#_c_270_n 0.02808f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A1_c_175_n N_A_27_47#_c_270_n 0.0040271f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A1_c_176_n N_A_27_47#_c_270_n 0.00942444f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_176_n N_A_27_47#_c_271_n 0.00582398f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_176_n N_VGND_c_311_n 0.00268723f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_176_n N_VGND_c_313_n 0.00421028f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A1_c_176_n N_VGND_c_314_n 0.00663995f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_146 N_VPWR_c_201_n A_109_297# 0.00275535f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_147 N_VPWR_c_201_n N_Y_M1003_d 0.0054793f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_148 N_VPWR_c_206_n Y 0.037225f $X=1.895 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_c_201_n Y 0.027844f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_150 N_VPWR_c_201_n A_307_297# 0.00244669f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_151 A_109_297# N_Y_c_235_n 0.00336772f $X=0.545 $Y=1.485 $X2=0.24 $Y2=2.34
cc_152 A_109_297# Y 0.00394829f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_153 N_Y_M1007_d N_A_27_47#_c_269_n 0.00354591f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_154 N_Y_c_241_n N_A_27_47#_c_269_n 0.0160731f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_155 N_Y_c_235_n N_A_27_47#_c_278_n 0.0014108f $X=0.58 $Y=1.835 $X2=0 $Y2=0
cc_156 N_Y_M1007_d N_VGND_c_314_n 0.00231419f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_270_n N_VGND_M1004_d 0.00431108f $X=1.875 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_27_47#_c_270_n N_VGND_c_311_n 0.012114f $X=1.875 $Y=0.78 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_269_n N_VGND_c_312_n 0.0421545f $X=1.015 $Y=0.385 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_281_n N_VGND_c_312_n 0.0160422f $X=1.18 $Y=0.475 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_270_n N_VGND_c_312_n 0.00240491f $X=1.875 $Y=0.78 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_270_n N_VGND_c_313_n 0.00211912f $X=1.875 $Y=0.78 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_271_n N_VGND_c_313_n 0.01858f $X=2.04 $Y=0.39 $X2=0 $Y2=0
cc_164 N_A_27_47#_M1007_s N_VGND_c_314_n 0.00211652f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_M1005_d N_VGND_c_314_n 0.00287338f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_M1002_d N_VGND_c_314_n 0.00210425f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_269_n N_VGND_c_314_n 0.0323745f $X=1.015 $Y=0.385 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_281_n N_VGND_c_314_n 0.0122621f $X=1.18 $Y=0.475 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_270_n N_VGND_c_314_n 0.00901584f $X=1.875 $Y=0.78 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_271_n N_VGND_c_314_n 0.0125989f $X=2.04 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__mux2i_1.pxi.spice
* Created: Tue Sep  1 19:14:42 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2I_1%A0 N_A0_c_65_n N_A0_M1007_g N_A0_M1003_g A0
+ N_A0_c_67_n PM_SKY130_FD_SC_HD__MUX2I_1%A0
x_PM_SKY130_FD_SC_HD__MUX2I_1%A1 N_A1_M1005_g N_A1_M1001_g A1 A1 N_A1_c_91_n
+ N_A1_c_92_n N_A1_c_93_n A1 PM_SKY130_FD_SC_HD__MUX2I_1%A1
x_PM_SKY130_FD_SC_HD__MUX2I_1%A_283_205# N_A_283_205#_M1006_s
+ N_A_283_205#_M1000_s N_A_283_205#_M1004_g N_A_283_205#_M1009_g
+ N_A_283_205#_c_131_n N_A_283_205#_c_132_n N_A_283_205#_c_138_n
+ N_A_283_205#_c_133_n N_A_283_205#_c_134_n N_A_283_205#_c_135_n
+ PM_SKY130_FD_SC_HD__MUX2I_1%A_283_205#
x_PM_SKY130_FD_SC_HD__MUX2I_1%S N_S_M1008_g N_S_M1002_g N_S_c_195_n N_S_c_196_n
+ N_S_M1006_g N_S_M1000_g N_S_c_197_n S S S N_S_c_199_n
+ PM_SKY130_FD_SC_HD__MUX2I_1%S
x_PM_SKY130_FD_SC_HD__MUX2I_1%A_27_297# N_A_27_297#_M1003_s N_A_27_297#_M1008_d
+ N_A_27_297#_c_251_n N_A_27_297#_c_252_n N_A_27_297#_c_259_n
+ N_A_27_297#_c_265_n N_A_27_297#_c_253_n N_A_27_297#_c_263_n
+ N_A_27_297#_c_254_n N_A_27_297#_c_255_n PM_SKY130_FD_SC_HD__MUX2I_1%A_27_297#
x_PM_SKY130_FD_SC_HD__MUX2I_1%Y N_Y_M1007_d N_Y_M1003_d Y Y N_Y_c_292_n
+ PM_SKY130_FD_SC_HD__MUX2I_1%Y
x_PM_SKY130_FD_SC_HD__MUX2I_1%VPWR N_VPWR_M1004_d N_VPWR_M1000_d N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n VPWR
+ N_VPWR_c_322_n N_VPWR_c_316_n PM_SKY130_FD_SC_HD__MUX2I_1%VPWR
x_PM_SKY130_FD_SC_HD__MUX2I_1%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1009_s
+ N_A_27_47#_c_356_n N_A_27_47#_c_365_n N_A_27_47#_c_357_n N_A_27_47#_c_358_n
+ N_A_27_47#_c_364_n PM_SKY130_FD_SC_HD__MUX2I_1%A_27_47#
x_PM_SKY130_FD_SC_HD__MUX2I_1%A_193_47# N_A_193_47#_M1005_d N_A_193_47#_M1002_d
+ N_A_193_47#_c_382_n N_A_193_47#_c_383_n N_A_193_47#_c_384_n
+ N_A_193_47#_c_385_n PM_SKY130_FD_SC_HD__MUX2I_1%A_193_47#
x_PM_SKY130_FD_SC_HD__MUX2I_1%VGND N_VGND_M1009_d N_VGND_M1006_d N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n VGND N_VGND_c_418_n N_VGND_c_419_n
+ N_VGND_c_420_n N_VGND_c_421_n PM_SKY130_FD_SC_HD__MUX2I_1%VGND
cc_1 VNB N_A0_c_65_n 0.0221898f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A0 0.00925368f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A0_c_67_n 0.039606f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A1_c_91_n 0.0282278f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_5 VNB N_A1_c_92_n 0.0221895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A1_c_93_n 0.00279814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_283_205#_M1004_g 4.48114e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_283_205#_M1009_g 0.0240733f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_9 VNB N_A_283_205#_c_131_n 0.0131473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_283_205#_c_132_n 0.00856732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_283_205#_c_133_n 0.00282988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_283_205#_c_134_n 5.36744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_283_205#_c_135_n 0.042818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_S_M1002_g 0.0299549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_S_c_195_n 0.0291413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_S_c_196_n 0.0227703f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_17 VNB N_S_c_197_n 0.00507206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB S 0.0211218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_S_c_199_n 0.0361462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_292_n 0.0086171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_316_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_356_n 0.0176489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_357_n 0.00640165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_358_n 0.00921644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_c_382_n 0.0029015f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_26 VNB N_A_193_47#_c_383_n 0.0037308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_384_n 0.00239359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_385_n 0.00844407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_415_n 0.00466605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_416_n 0.0102534f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_31 VNB N_VGND_c_417_n 0.0160198f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_32 VNB N_VGND_c_418_n 0.0478121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_419_n 0.0309004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_420_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_421_n 0.210298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A0_M1003_g 0.0260553f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_37 VPB N_A0_c_67_n 0.0102093f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_38 VPB N_A1_M1001_g 0.0206808f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_39 VPB N_A1_c_91_n 0.00807244f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_40 VPB N_A1_c_93_n 0.00379723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_283_205#_M1004_g 0.0241837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_283_205#_c_131_n 0.00634988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_283_205#_c_138_n 0.00262368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_S_M1008_g 0.0242642f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_45 VPB N_S_c_195_n 0.0256471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_S_M1000_g 0.0247446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_S_c_197_n 0.00211602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB S 0.0126219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_S_c_199_n 0.0109066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_297#_c_251_n 0.00712721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_297#_c_252_n 0.0331813f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_253_n 0.00425745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_297#_c_254_n 0.00377351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_297#_c_255_n 0.00818989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB Y 0.00220261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_Y_c_292_n 0.00328556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_317_n 0.0050814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_318_n 0.0106178f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_59 VPB N_VPWR_c_319_n 0.0306458f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_60 VPB N_VPWR_c_320_n 0.0435345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_321_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_322_n 0.0366286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_316_n 0.0544872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 N_A0_M1003_g N_A1_M1001_g 0.0245475f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A0_c_67_n N_A1_c_91_n 0.0287631f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A0_c_65_n N_A1_c_92_n 0.0133018f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A0_M1003_g N_A_27_297#_c_252_n 0.00932467f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_68 A0 N_A_27_297#_c_252_n 0.0245948f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A0_c_67_n N_A_27_297#_c_252_n 0.00726508f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A0_M1003_g N_A_27_297#_c_259_n 0.0119907f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A0_M1003_g Y 0.00401017f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A0_c_65_n N_Y_c_292_n 0.00280474f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_73 A0 N_Y_c_292_n 0.0170715f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A0_c_67_n N_Y_c_292_n 0.00401017f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A0_M1003_g N_VPWR_c_320_n 0.0035787f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A0_M1003_g N_VPWR_c_316_n 0.00627709f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_77 A0 N_A_27_47#_c_356_n 0.0195144f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A0_c_67_n N_A_27_47#_c_356_n 0.00588963f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A0_c_65_n N_A_27_47#_c_358_n 0.00339071f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_80 A0 N_A_27_47#_c_358_n 0.00123148f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A0_c_67_n N_A_27_47#_c_358_n 7.09714e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A0_c_65_n N_A_27_47#_c_364_n 0.00904079f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A0_c_65_n N_VGND_c_418_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A0_c_65_n N_VGND_c_421_n 0.00620762f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A1_M1001_g N_A_283_205#_M1004_g 0.0336052f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_86 A1 N_A_283_205#_M1004_g 0.00197951f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_87 N_A1_c_93_n N_A_283_205#_M1004_g 0.00384556f $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_88 N_A1_c_91_n N_A_283_205#_M1009_g 6.59671e-19 $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A1_c_91_n N_A_283_205#_c_131_n 0.00115192f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A1_c_93_n N_A_283_205#_c_131_n 0.0175451f $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_91 N_A1_c_91_n N_A_283_205#_c_135_n 0.0166488f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A1_c_93_n N_A_283_205#_c_135_n 8.93471e-19 $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_93 N_A1_M1001_g N_A_27_297#_c_252_n 8.93484e-19 $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A1_M1001_g N_A_27_297#_c_259_n 0.0149514f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_95 A1 N_A_27_297#_c_259_n 0.0111209f $X=1.065 $Y=1.445 $X2=0 $Y2=0
cc_96 N_A1_c_93_n N_A_27_297#_c_263_n 0.00263799f $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_97 N_A1_M1001_g Y 2.48058e-19 $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A1_c_91_n Y 0.00120285f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A1_c_93_n Y 0.00207457f $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_100 N_A1_M1001_g N_Y_c_292_n 0.00103603f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A1_c_92_n N_Y_c_292_n 0.00531421f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A1_c_93_n N_Y_c_292_n 0.0311966f $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_103 A1 A_204_297# 0.0113841f $X=1.065 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_104 N_A1_c_93_n A_204_297# 8.53962e-19 $X=1.135 $Y=1.545 $X2=-0.19 $Y2=-0.24
cc_105 N_A1_M1001_g N_VPWR_c_320_n 0.00357877f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A1_M1001_g N_VPWR_c_316_n 0.00569486f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A1_c_92_n N_A_27_47#_c_365_n 0.00562452f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A1_c_92_n N_A_27_47#_c_364_n 0.0118771f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A1_c_91_n N_A_193_47#_c_384_n 0.00220841f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A1_c_92_n N_A_193_47#_c_384_n 0.0018135f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A1_c_93_n N_A_193_47#_c_384_n 0.0157579f $X=1.135 $Y=1.545 $X2=0 $Y2=0
cc_112 N_A1_c_92_n N_VGND_c_418_n 0.00357877f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A1_c_92_n N_VGND_c_421_n 0.00666937f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_283_205#_c_138_n N_S_M1008_g 0.00474138f $X=3 $Y=1.62 $X2=0 $Y2=0
cc_115 N_A_283_205#_M1009_g N_S_M1002_g 0.0287041f $X=1.85 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_283_205#_c_131_n N_S_M1002_g 0.00646483f $X=2.8 $Y=1.192 $X2=0 $Y2=0
cc_117 N_A_283_205#_c_132_n N_S_M1002_g 0.0057324f $X=3 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_283_205#_c_135_n N_S_M1002_g 0.00815798f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_283_205#_c_131_n N_S_c_195_n 0.0211205f $X=2.8 $Y=1.192 $X2=0 $Y2=0
cc_120 N_A_283_205#_c_138_n N_S_c_195_n 0.00760718f $X=3 $Y=1.62 $X2=0 $Y2=0
cc_121 N_A_283_205#_c_134_n N_S_c_195_n 0.0145751f $X=2.942 $Y=1.192 $X2=0 $Y2=0
cc_122 N_A_283_205#_c_132_n N_S_c_196_n 0.00470642f $X=3 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_283_205#_c_133_n N_S_c_196_n 0.00405253f $X=3 $Y=0.4 $X2=0 $Y2=0
cc_124 N_A_283_205#_c_138_n N_S_M1000_g 0.00299314f $X=3 $Y=1.62 $X2=0 $Y2=0
cc_125 N_A_283_205#_M1004_g N_S_c_197_n 0.0201695f $X=1.49 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_283_205#_c_131_n N_S_c_197_n 0.00680809f $X=2.8 $Y=1.192 $X2=0 $Y2=0
cc_127 N_A_283_205#_c_135_n N_S_c_197_n 0.00849063f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_283_205#_c_132_n S 0.0190326f $X=3 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_283_205#_c_138_n S 0.0178563f $X=3 $Y=1.62 $X2=0 $Y2=0
cc_130 N_A_283_205#_c_134_n S 0.0187515f $X=2.942 $Y=1.192 $X2=0 $Y2=0
cc_131 N_A_283_205#_c_134_n N_S_c_199_n 0.00257883f $X=2.942 $Y=1.192 $X2=0
+ $Y2=0
cc_132 N_A_283_205#_M1004_g N_A_27_297#_c_259_n 0.00775505f $X=1.49 $Y=1.985
+ $X2=0 $Y2=0
cc_133 N_A_283_205#_M1004_g N_A_27_297#_c_265_n 0.0182579f $X=1.49 $Y=1.985
+ $X2=0 $Y2=0
cc_134 N_A_283_205#_c_131_n N_A_27_297#_c_253_n 0.0538114f $X=2.8 $Y=1.192 $X2=0
+ $Y2=0
cc_135 N_A_283_205#_c_135_n N_A_27_297#_c_253_n 0.0025587f $X=1.85 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_283_205#_M1004_g N_A_27_297#_c_263_n 0.00870829f $X=1.49 $Y=1.985
+ $X2=0 $Y2=0
cc_137 N_A_283_205#_c_131_n N_A_27_297#_c_263_n 0.0134141f $X=2.8 $Y=1.192 $X2=0
+ $Y2=0
cc_138 N_A_283_205#_c_131_n N_A_27_297#_c_254_n 0.0270288f $X=2.8 $Y=1.192 $X2=0
+ $Y2=0
cc_139 N_A_283_205#_c_138_n N_A_27_297#_c_254_n 0.011079f $X=3 $Y=1.62 $X2=0
+ $Y2=0
cc_140 N_A_283_205#_c_138_n N_A_27_297#_c_255_n 0.0498445f $X=3 $Y=1.62 $X2=0
+ $Y2=0
cc_141 N_A_283_205#_M1004_g N_VPWR_c_317_n 0.00549893f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_283_205#_M1004_g N_VPWR_c_320_n 0.00357668f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_283_205#_c_138_n N_VPWR_c_322_n 0.0154725f $X=3 $Y=1.62 $X2=0 $Y2=0
cc_144 N_A_283_205#_M1000_s N_VPWR_c_316_n 0.00463037f $X=2.845 $Y=1.485 $X2=0
+ $Y2=0
cc_145 N_A_283_205#_M1004_g N_VPWR_c_316_n 0.00624492f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_283_205#_c_138_n N_VPWR_c_316_n 0.00858812f $X=3 $Y=1.62 $X2=0 $Y2=0
cc_147 N_A_283_205#_M1009_g N_A_27_47#_c_357_n 0.00292079f $X=1.85 $Y=0.56 $X2=0
+ $Y2=0
cc_148 N_A_283_205#_M1009_g N_A_193_47#_c_382_n 0.0139021f $X=1.85 $Y=0.56 $X2=0
+ $Y2=0
cc_149 N_A_283_205#_c_131_n N_A_193_47#_c_382_n 0.0175566f $X=2.8 $Y=1.192 $X2=0
+ $Y2=0
cc_150 N_A_283_205#_c_132_n N_A_193_47#_c_382_n 0.014291f $X=3 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_283_205#_c_133_n N_A_193_47#_c_383_n 0.0357313f $X=3 $Y=0.4 $X2=0
+ $Y2=0
cc_152 N_A_283_205#_M1009_g N_A_193_47#_c_385_n 0.00214388f $X=1.85 $Y=0.56
+ $X2=0 $Y2=0
cc_153 N_A_283_205#_c_131_n N_A_193_47#_c_385_n 0.0598351f $X=2.8 $Y=1.192 $X2=0
+ $Y2=0
cc_154 N_A_283_205#_c_135_n N_A_193_47#_c_385_n 0.00873518f $X=1.85 $Y=1.16
+ $X2=0 $Y2=0
cc_155 N_A_283_205#_M1009_g N_VGND_c_415_n 0.00268723f $X=1.85 $Y=0.56 $X2=0
+ $Y2=0
cc_156 N_A_283_205#_M1009_g N_VGND_c_418_n 0.00420765f $X=1.85 $Y=0.56 $X2=0
+ $Y2=0
cc_157 N_A_283_205#_c_133_n N_VGND_c_419_n 0.0234083f $X=3 $Y=0.4 $X2=0 $Y2=0
cc_158 N_A_283_205#_M1006_s N_VGND_c_421_n 0.00209319f $X=2.875 $Y=0.235 $X2=0
+ $Y2=0
cc_159 N_A_283_205#_M1009_g N_VGND_c_421_n 0.00705894f $X=1.85 $Y=0.56 $X2=0
+ $Y2=0
cc_160 N_A_283_205#_c_133_n N_VGND_c_421_n 0.0136987f $X=3 $Y=0.4 $X2=0 $Y2=0
cc_161 N_S_M1008_g N_A_27_297#_c_253_n 0.0119618f $X=2.24 $Y=1.985 $X2=0 $Y2=0
cc_162 N_S_M1008_g N_A_27_297#_c_254_n 8.99581e-19 $X=2.24 $Y=1.985 $X2=0 $Y2=0
cc_163 N_S_c_195_n N_A_27_297#_c_254_n 0.0047871f $X=3.135 $Y=1.257 $X2=0 $Y2=0
cc_164 N_S_M1008_g N_A_27_297#_c_255_n 0.0175042f $X=2.24 $Y=1.985 $X2=0 $Y2=0
cc_165 S N_VPWR_M1000_d 0.0029998f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_166 N_S_M1008_g N_VPWR_c_317_n 0.00917253f $X=2.24 $Y=1.985 $X2=0 $Y2=0
cc_167 N_S_M1000_g N_VPWR_c_319_n 0.00487552f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_168 S N_VPWR_c_319_n 0.018846f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_169 N_S_c_199_n N_VPWR_c_319_n 0.00109656f $X=3.21 $Y=1.17 $X2=0 $Y2=0
cc_170 N_S_M1008_g N_VPWR_c_322_n 0.00541359f $X=2.24 $Y=1.985 $X2=0 $Y2=0
cc_171 N_S_M1000_g N_VPWR_c_322_n 0.00585385f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_172 N_S_M1008_g N_VPWR_c_316_n 0.0116918f $X=2.24 $Y=1.985 $X2=0 $Y2=0
cc_173 N_S_M1000_g N_VPWR_c_316_n 0.012717f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_174 N_S_M1002_g N_A_193_47#_c_382_n 0.0129258f $X=2.27 $Y=0.56 $X2=0 $Y2=0
cc_175 N_S_c_195_n N_A_193_47#_c_382_n 0.00115948f $X=3.135 $Y=1.257 $X2=0 $Y2=0
cc_176 S N_VGND_M1006_d 0.00265397f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_177 N_S_M1002_g N_VGND_c_415_n 0.00268723f $X=2.27 $Y=0.56 $X2=0 $Y2=0
cc_178 S N_VGND_c_416_n 6.24443e-19 $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_179 N_S_c_196_n N_VGND_c_417_n 0.0044587f $X=3.21 $Y=0.99 $X2=0 $Y2=0
cc_180 S N_VGND_c_417_n 0.0150646f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_181 N_S_c_199_n N_VGND_c_417_n 0.0010142f $X=3.21 $Y=1.17 $X2=0 $Y2=0
cc_182 N_S_M1002_g N_VGND_c_419_n 0.00436487f $X=2.27 $Y=0.56 $X2=0 $Y2=0
cc_183 N_S_c_196_n N_VGND_c_419_n 0.00518482f $X=3.21 $Y=0.99 $X2=0 $Y2=0
cc_184 S N_VGND_c_419_n 6.78075e-19 $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_185 N_S_M1002_g N_VGND_c_421_n 0.00731071f $X=2.27 $Y=0.56 $X2=0 $Y2=0
cc_186 N_S_c_196_n N_VGND_c_421_n 0.0110721f $X=3.21 $Y=0.99 $X2=0 $Y2=0
cc_187 S N_VGND_c_421_n 0.00398521f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_188 N_A_27_297#_c_259_n N_Y_M1003_d 0.00382426f $X=1.405 $Y=2.38 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_252_n Y 0.0259326f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_190 N_A_27_297#_c_259_n Y 0.0145504f $X=1.405 $Y=2.38 $X2=0 $Y2=0
cc_191 N_A_27_297#_c_259_n A_204_297# 0.00938736f $X=1.405 $Y=2.38 $X2=-0.19
+ $Y2=1.305
cc_192 N_A_27_297#_c_253_n N_VPWR_M1004_d 0.0145345f $X=2.285 $Y=1.565 $X2=-0.19
+ $Y2=1.305
cc_193 N_A_27_297#_c_253_n N_VPWR_c_317_n 0.0174139f $X=2.285 $Y=1.565 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_255_n N_VPWR_c_317_n 0.0300045f $X=2.45 $Y=2.32 $X2=0 $Y2=0
cc_195 N_A_27_297#_c_251_n N_VPWR_c_320_n 0.0190876f $X=0.27 $Y=2.295 $X2=0
+ $Y2=0
cc_196 N_A_27_297#_c_259_n N_VPWR_c_320_n 0.0666676f $X=1.405 $Y=2.38 $X2=0
+ $Y2=0
cc_197 N_A_27_297#_c_255_n N_VPWR_c_322_n 0.0210382f $X=2.45 $Y=2.32 $X2=0 $Y2=0
cc_198 N_A_27_297#_M1003_s N_VPWR_c_316_n 0.00225715f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_M1008_d N_VPWR_c_316_n 0.00209319f $X=2.315 $Y=1.485 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_c_251_n N_VPWR_c_316_n 0.0114582f $X=0.27 $Y=2.295 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_c_259_n N_VPWR_c_316_n 0.0411989f $X=1.405 $Y=2.38 $X2=0
+ $Y2=0
cc_202 N_A_27_297#_c_255_n N_VPWR_c_316_n 0.0124268f $X=2.45 $Y=2.32 $X2=0 $Y2=0
cc_203 N_Y_M1003_d N_VPWR_c_316_n 0.00244941f $X=0.565 $Y=1.485 $X2=0 $Y2=0
cc_204 N_Y_M1007_d N_A_27_47#_c_364_n 0.00312348f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_205 N_Y_c_292_n N_A_27_47#_c_364_n 0.0118865f $X=0.68 $Y=0.76 $X2=0 $Y2=0
cc_206 N_Y_M1007_d N_VGND_c_421_n 0.00216833f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_207 A_204_297# N_VPWR_c_316_n 0.00317218f $X=1.02 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_365_n N_A_193_47#_M1005_d 0.00334172f $X=1.175 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_209 N_A_27_47#_c_357_n N_A_193_47#_M1005_d 0.00222246f $X=1.64 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_210 N_A_27_47#_M1009_s N_A_193_47#_c_382_n 0.00480511f $X=1.515 $Y=0.235
+ $X2=0 $Y2=0
cc_211 N_A_27_47#_c_357_n N_A_193_47#_c_382_n 0.0113937f $X=1.64 $Y=0.38 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_365_n N_A_193_47#_c_384_n 0.0163927f $X=1.175 $Y=0.36 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_364_n N_A_193_47#_c_384_n 4.37145e-19 $X=0.965 $Y=0.36 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1009_s N_A_193_47#_c_385_n 0.00100435f $X=1.515 $Y=0.235
+ $X2=0 $Y2=0
cc_215 N_A_27_47#_c_357_n N_A_193_47#_c_385_n 0.0163927f $X=1.64 $Y=0.38 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_358_n N_VGND_c_418_n 0.101535f $X=0.44 $Y=0.36 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1007_s N_VGND_c_421_n 0.00209344f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_M1009_s N_VGND_c_421_n 0.00209344f $X=1.515 $Y=0.235 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_358_n N_VGND_c_421_n 0.062612f $X=0.44 $Y=0.36 $X2=0 $Y2=0
cc_220 N_A_193_47#_c_382_n N_VGND_M1009_d 0.00335838f $X=2.385 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_193_47#_c_382_n N_VGND_c_415_n 0.012179f $X=2.385 $Y=0.8 $X2=0 $Y2=0
cc_222 N_A_193_47#_c_382_n N_VGND_c_418_n 0.00203142f $X=2.385 $Y=0.8 $X2=0
+ $Y2=0
cc_223 N_A_193_47#_c_382_n N_VGND_c_419_n 0.00275431f $X=2.385 $Y=0.8 $X2=0
+ $Y2=0
cc_224 N_A_193_47#_c_383_n N_VGND_c_419_n 0.0157611f $X=2.48 $Y=0.55 $X2=0 $Y2=0
cc_225 N_A_193_47#_M1005_d N_VGND_c_421_n 0.00226545f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_193_47#_M1002_d N_VGND_c_421_n 0.00228609f $X=2.345 $Y=0.235 $X2=0
+ $Y2=0
cc_227 N_A_193_47#_c_382_n N_VGND_c_421_n 0.0108006f $X=2.385 $Y=0.8 $X2=0 $Y2=0
cc_228 N_A_193_47#_c_383_n N_VGND_c_421_n 0.00895528f $X=2.48 $Y=0.55 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__or3_1.pex.spice
* Created: Thu Aug 27 14:43:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR3_1%C 3 7 9 15
r26 12 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.255 $Y=1.16
+ $X2=0.48 $Y2=1.16
r27 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r28 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r29 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.48 $Y=1.325 $X2=0.48
+ $Y2=1.695
r30 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r31 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.48 $Y=0.995 $X2=0.48
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_1%B 4 7 8 9 10 11 15 16
r41 15 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.9 $Y=2.28 $X2=0.9
+ $Y2=2.145
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.9
+ $Y=2.28 $X2=0.9 $Y2=2.28
r43 11 16 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=0.685 $Y=2.27
+ $X2=0.9 $Y2=2.27
r44 10 11 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.225 $Y=2.27
+ $X2=0.685 $Y2=2.27
r45 8 9 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=0.87 $Y=0.76 $X2=0.87
+ $Y2=0.91
r46 7 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.9 $Y=0.475 $X2=0.9
+ $Y2=0.76
r47 4 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.84 $Y=1.695
+ $X2=0.84 $Y2=2.145
r48 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.84 $Y=1.695
+ $X2=0.84 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_1%A 3 7 9 10 11 16 17 20
c52 20 0 1.12051e-19 $X=0.697 $Y=1.325
r53 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=1.16
+ $X2=1.305 $Y2=1.325
r54 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=1.16
+ $X2=1.305 $Y2=0.995
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.305
+ $Y=1.16 $X2=1.305 $Y2=1.16
r56 11 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.145 $Y=1.16
+ $X2=1.305 $Y2=1.16
r57 11 24 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.145 $Y=1.16
+ $X2=0.795 $Y2=1.16
r58 10 20 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.697 $Y=1.53
+ $X2=0.697 $Y2=1.325
r59 9 20 4.65494 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.697 $Y=1.16
+ $X2=0.697 $Y2=1.325
r60 9 24 2.76475 $w=3.3e-07 $l=9.8e-08 $layer=LI1_cond $X=0.697 $Y=1.16
+ $X2=0.795 $Y2=1.16
r61 7 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.32 $Y=1.695
+ $X2=1.32 $Y2=1.325
r62 3 18 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.32 $Y=0.475
+ $X2=1.32 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_1%A_29_53# 1 2 3 12 15 19 21 22 23 27 29 31 36
+ 38 42 43 48 49 50 53
c93 48 0 1.14153e-19 $X=1.785 $Y=1.16
c94 36 0 1.06604e-19 $X=1.68 $Y=1.495
r95 49 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.16
+ $X2=1.785 $Y2=1.325
r96 49 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.16
+ $X2=1.785 $Y2=0.995
r97 48 51 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.732 $Y=1.16
+ $X2=1.732 $Y2=1.325
r98 48 50 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.732 $Y=1.16
+ $X2=1.732 $Y2=0.995
r99 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=1.16 $X2=1.785 $Y2=1.16
r100 43 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.19 $Y=1.58
+ $X2=1.19 $Y2=1.87
r101 38 40 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=0.267 $Y=1.685
+ $X2=0.267 $Y2=1.87
r102 36 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=1.495
+ $X2=1.68 $Y2=1.325
r103 33 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=0.825
+ $X2=1.68 $Y2=0.995
r104 32 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.58
+ $X2=1.19 $Y2=1.58
r105 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.595 $Y=1.58
+ $X2=1.68 $Y2=1.495
r106 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.595 $Y=1.58
+ $X2=1.275 $Y2=1.58
r107 30 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.74
+ $X2=1.11 $Y2=0.74
r108 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.595 $Y=0.74
+ $X2=1.68 $Y2=0.825
r109 29 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.595 $Y=0.74
+ $X2=1.195 $Y2=0.74
r110 25 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=0.655
+ $X2=1.11 $Y2=0.74
r111 25 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.11 $Y=0.655
+ $X2=1.11 $Y2=0.47
r112 24 40 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.43 $Y=1.87
+ $X2=0.267 $Y2=1.87
r113 23 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=1.87
+ $X2=1.19 $Y2=1.87
r114 23 24 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.105 $Y=1.87
+ $X2=0.43 $Y2=1.87
r115 21 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.025 $Y=0.74
+ $X2=1.11 $Y2=0.74
r116 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=0.74
+ $X2=0.355 $Y2=0.74
r117 17 22 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.227 $Y=0.655
+ $X2=0.355 $Y2=0.74
r118 17 19 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=0.227 $Y=0.655
+ $X2=0.227 $Y2=0.47
r119 15 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.81 $Y=1.985
+ $X2=1.81 $Y2=1.325
r120 12 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.81 $Y=0.56
+ $X2=1.81 $Y2=0.995
r121 3 38 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.685
r122 2 27 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.265 $X2=1.11 $Y2=0.47
r123 1 19 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.265 $X2=0.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_1%VPWR 1 6 8 10 20 21 24 29
c26 1 0 1.06604e-19 $X=1.395 $Y=1.485
r27 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r29 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r30 18 24 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.725 $Y=2.72
+ $X2=1.585 $Y2=2.72
r31 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.725 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 17 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r33 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.23 $Y2=2.72
r34 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 12 16 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 12 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r37 10 24 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.585 $Y2=2.72
r38 10 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 8 29 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r40 4 24 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=2.635
+ $X2=1.585 $Y2=2.72
r41 4 6 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.585 $Y=2.635
+ $X2=1.585 $Y2=2
r42 1 6 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.395
+ $Y=1.485 $X2=1.595 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_1%X 1 2 12 14 15 16
r18 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=2.072 $Y=1.632
+ $X2=2.072 $Y2=1.845
r19 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.072 $Y=1.632
+ $X2=2.072 $Y2=1.495
r20 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=2.02 $Y=0.587
+ $X2=2.125 $Y2=0.587
r21 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.125 $Y=0.76
+ $X2=2.125 $Y2=0.587
r22 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.125 $Y=0.76
+ $X2=2.125 $Y2=1.495
r23 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=1.885
+ $Y=1.485 $X2=2.02 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.235 $X2=2.02 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_1%VGND 1 2 9 13 15 17 22 29 30 33 36 41
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r43 34 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r44 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r46 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r47 27 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.555
+ $Y2=0
r48 27 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=2.07
+ $Y2=0
r49 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r50 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r51 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r53 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.15
+ $Y2=0
r54 22 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.555
+ $Y2=0
r55 22 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.15
+ $Y2=0
r56 19 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r57 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r58 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r59 15 41 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r60 11 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=0.085
+ $X2=1.555 $Y2=0
r61 11 13 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.555 $Y=0.085
+ $X2=1.555 $Y2=0.4
r62 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r63 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.4
r64 2 13 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.395
+ $Y=0.265 $X2=1.58 $Y2=0.4
r65 1 9 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.265 $X2=0.69 $Y2=0.4
.ends


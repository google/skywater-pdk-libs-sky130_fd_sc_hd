* File: sky130_fd_sc_hd__o21ai_1.pxi.spice
* Created: Tue Sep  1 19:21:31 2020
* 
x_PM_SKY130_FD_SC_HD__O21AI_1%A1 N_A1_M1005_g N_A1_M1003_g A1 N_A1_c_39_n
+ N_A1_c_40_n N_A1_c_41_n PM_SKY130_FD_SC_HD__O21AI_1%A1
x_PM_SKY130_FD_SC_HD__O21AI_1%A2 N_A2_M1000_g N_A2_M1002_g A2 A2 A2 A2
+ N_A2_c_64_n N_A2_c_65_n N_A2_c_66_n PM_SKY130_FD_SC_HD__O21AI_1%A2
x_PM_SKY130_FD_SC_HD__O21AI_1%B1 N_B1_M1004_g N_B1_M1001_g B1 N_B1_c_108_n
+ PM_SKY130_FD_SC_HD__O21AI_1%B1
x_PM_SKY130_FD_SC_HD__O21AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1001_d N_VPWR_c_138_n
+ N_VPWR_c_139_n N_VPWR_c_140_n N_VPWR_c_141_n VPWR N_VPWR_c_142_n
+ N_VPWR_c_137_n PM_SKY130_FD_SC_HD__O21AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O21AI_1%Y N_Y_M1004_d N_Y_M1000_d N_Y_c_166_n N_Y_c_167_n
+ N_Y_c_168_n Y Y N_Y_c_169_n PM_SKY130_FD_SC_HD__O21AI_1%Y
x_PM_SKY130_FD_SC_HD__O21AI_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1002_d
+ N_A_27_47#_c_200_n N_A_27_47#_c_202_n N_A_27_47#_c_201_n N_A_27_47#_c_210_n
+ PM_SKY130_FD_SC_HD__O21AI_1%A_27_47#
x_PM_SKY130_FD_SC_HD__O21AI_1%VGND N_VGND_M1005_d N_VGND_c_223_n VGND
+ N_VGND_c_224_n N_VGND_c_225_n N_VGND_c_226_n N_VGND_c_227_n
+ PM_SKY130_FD_SC_HD__O21AI_1%VGND
cc_1 VNB N_A1_c_39_n 0.0307012f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_2 VNB N_A1_c_40_n 0.0115946f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_3 VNB N_A1_c_41_n 0.0227675f $X=-0.19 $Y=-0.24 $X2=0.367 $Y2=0.995
cc_4 VNB N_A2_c_64_n 0.0215419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A2_c_65_n 0.00348809f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_6 VNB N_A2_c_66_n 0.0167529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B1_M1004_g 0.0396748f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_8 VNB B1 0.00499959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_108_n 0.0088983f $X=-0.19 $Y=-0.24 $X2=0.367 $Y2=1.325
cc_10 VNB N_VPWR_c_137_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_166_n 0.0101911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_Y_c_167_n 0.00260201f $X=-0.19 $Y=-0.24 $X2=0.367 $Y2=1.16
cc_13 VNB N_Y_c_168_n 0.00308674f $X=-0.19 $Y=-0.24 $X2=0.367 $Y2=0.995
cc_14 VNB N_Y_c_169_n 0.0010487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_200_n 0.013695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_201_n 0.00894105f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_17 VNB N_VGND_c_223_n 0.00280453f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_18 VNB N_VGND_c_224_n 0.0168743f $X=-0.19 $Y=-0.24 $X2=0.367 $Y2=1.16
cc_19 VNB N_VGND_c_225_n 0.0269163f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_226_n 0.125064f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_21 VNB N_VGND_c_227_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A1_M1003_g 0.0247502f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_23 VPB N_A1_c_39_n 0.00656253f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_24 VPB N_A1_c_40_n 0.00105932f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_25 VPB N_A2_M1000_g 0.0186378f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_26 VPB A2 0.00193343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A2_c_64_n 0.00632341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A2_c_65_n 5.81142e-19 $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_29 VPB N_B1_M1001_g 0.0258776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB B1 0.0150543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_B1_c_108_n 0.0388746f $X=-0.19 $Y=1.305 $X2=0.367 $Y2=1.325
cc_32 VPB N_VPWR_c_138_n 0.0100471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_139_n 0.0428697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_140_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0.367 $Y2=0.995
cc_35 VPB N_VPWR_c_141_n 0.0299462f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_36 VPB N_VPWR_c_142_n 0.0287826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_137_n 0.0424607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_Y_c_169_n 0.0014021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 N_A1_M1003_g N_A2_M1000_g 0.0484572f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_40 N_A1_M1003_g A2 0.00674592f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_41 N_A1_c_39_n N_A2_c_64_n 0.0484572f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_42 N_A1_c_40_n N_A2_c_64_n 2.49008e-19 $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_43 N_A1_c_39_n N_A2_c_65_n 0.00250441f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_44 N_A1_c_40_n N_A2_c_65_n 0.0249818f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_45 N_A1_c_41_n N_A2_c_66_n 0.0223313f $X=0.367 $Y=0.995 $X2=0 $Y2=0
cc_46 N_A1_M1003_g N_VPWR_c_139_n 0.015979f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_47 N_A1_c_39_n N_VPWR_c_139_n 0.00460192f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_48 N_A1_c_40_n N_VPWR_c_139_n 0.0189139f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A1_M1003_g N_VPWR_c_142_n 0.00525069f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A1_M1003_g N_VPWR_c_137_n 0.00875452f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_51 N_A1_c_40_n N_A_27_47#_c_202_n 0.00137991f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A1_c_41_n N_A_27_47#_c_202_n 0.0173435f $X=0.367 $Y=0.995 $X2=0 $Y2=0
cc_53 N_A1_c_39_n N_A_27_47#_c_201_n 0.0041554f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_54 N_A1_c_40_n N_A_27_47#_c_201_n 0.0144129f $X=0.325 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A1_c_41_n N_VGND_c_223_n 0.00308386f $X=0.367 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A1_c_41_n N_VGND_c_224_n 0.00422112f $X=0.367 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A1_c_41_n N_VGND_c_226_n 0.00669273f $X=0.367 $Y=0.995 $X2=0 $Y2=0
cc_58 N_A2_c_64_n N_B1_M1004_g 0.0152559f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A2_c_65_n N_B1_M1004_g 2.95851e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A2_c_66_n N_B1_M1004_g 0.024222f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_61 N_A2_M1000_g N_B1_c_108_n 0.0239558f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_62 A2 N_B1_c_108_n 3.57443e-19 $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_63 N_A2_M1000_g N_VPWR_c_139_n 0.00211424f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_64 N_A2_M1000_g N_VPWR_c_142_n 0.00544863f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_65 A2 N_VPWR_c_142_n 0.00708237f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_66 N_A2_M1000_g N_VPWR_c_137_n 0.00992036f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_67 A2 N_VPWR_c_137_n 0.00694416f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_68 A2 A_109_297# 0.00112971f $X=0.61 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_69 N_A2_c_64_n N_Y_c_167_n 9.62723e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A2_c_65_n N_Y_c_167_n 0.0108085f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A2_c_66_n N_Y_c_167_n 0.00108806f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A2_M1000_g Y 0.00905894f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_73 A2 Y 0.0622575f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_74 N_A2_c_64_n Y 0.00307667f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A2_c_65_n Y 7.11027e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A2_M1000_g N_Y_c_169_n 0.0013736f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_77 A2 N_Y_c_169_n 0.00736847f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_78 N_A2_c_64_n N_Y_c_169_n 0.00131834f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A2_c_65_n N_Y_c_169_n 0.0151692f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A2_c_64_n N_A_27_47#_c_202_n 0.00293285f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A2_c_65_n N_A_27_47#_c_202_n 0.0224662f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A2_c_66_n N_A_27_47#_c_202_n 0.0125549f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A2_c_66_n N_VGND_c_223_n 0.00807643f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A2_c_66_n N_VGND_c_225_n 0.00337001f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A2_c_66_n N_VGND_c_226_n 0.00397658f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B1_M1001_g N_VPWR_c_141_n 0.00450113f $X=1.37 $Y=2.135 $X2=0 $Y2=0
cc_87 B1 N_VPWR_c_141_n 0.0205041f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_88 N_B1_c_108_n N_VPWR_c_141_n 0.00194789f $X=1.6 $Y=1.46 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_VPWR_c_142_n 0.00585385f $X=1.37 $Y=2.135 $X2=0 $Y2=0
cc_90 N_B1_M1001_g N_VPWR_c_137_n 0.0117852f $X=1.37 $Y=2.135 $X2=0 $Y2=0
cc_91 N_B1_M1004_g N_Y_c_166_n 0.0166042f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_92 B1 N_Y_c_166_n 0.0135548f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_93 N_B1_c_108_n N_Y_c_166_n 0.00360827f $X=1.6 $Y=1.46 $X2=0 $Y2=0
cc_94 N_B1_M1004_g N_Y_c_167_n 0.00216703f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_95 N_B1_M1004_g N_Y_c_168_n 0.00529249f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_96 N_B1_M1001_g Y 0.00901363f $X=1.37 $Y=2.135 $X2=0 $Y2=0
cc_97 N_B1_c_108_n Y 0.00359015f $X=1.6 $Y=1.46 $X2=0 $Y2=0
cc_98 N_B1_M1004_g N_Y_c_169_n 0.00787472f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_99 B1 N_Y_c_169_n 0.0235643f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_100 N_B1_c_108_n N_Y_c_169_n 0.0053408f $X=1.6 $Y=1.46 $X2=0 $Y2=0
cc_101 N_B1_M1004_g N_A_27_47#_c_202_n 0.00316982f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_102 N_B1_M1004_g N_A_27_47#_c_210_n 0.00559155f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_103 N_B1_M1004_g N_VGND_c_223_n 0.00134679f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_104 N_B1_M1004_g N_VGND_c_225_n 0.00572397f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_105 N_B1_M1004_g N_VGND_c_226_n 0.0114994f $X=1.37 $Y=0.56 $X2=0 $Y2=0
cc_106 N_VPWR_c_137_n A_109_297# 0.00333694f $X=1.61 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_107 N_VPWR_c_137_n N_Y_M1000_d 0.00524128f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_108 N_VPWR_c_139_n Y 0.00275664f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_109 N_VPWR_c_142_n Y 0.0211142f $X=1.495 $Y=2.72 $X2=0 $Y2=0
cc_110 N_VPWR_c_137_n Y 0.0126319f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_111 N_Y_c_167_n N_A_27_47#_c_202_n 0.0118288f $X=1.315 $Y=1.04 $X2=0 $Y2=0
cc_112 N_Y_c_168_n N_VGND_c_225_n 0.00617006f $X=1.58 $Y=0.555 $X2=0 $Y2=0
cc_113 N_Y_M1004_d N_VGND_c_226_n 0.00540557f $X=1.445 $Y=0.235 $X2=0 $Y2=0
cc_114 N_Y_c_168_n N_VGND_c_226_n 0.0059977f $X=1.58 $Y=0.555 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_202_n N_VGND_M1005_d 0.00456716f $X=1.075 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_27_47#_c_202_n N_VGND_c_223_n 0.0183914f $X=1.075 $Y=0.7 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_200_n N_VGND_c_224_n 0.0174379f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_202_n N_VGND_c_224_n 0.00301967f $X=1.075 $Y=0.7 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_202_n N_VGND_c_225_n 0.00255672f $X=1.075 $Y=0.7 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_210_n N_VGND_c_225_n 0.0100025f $X=1.16 $Y=0.475 $X2=0 $Y2=0
cc_121 N_A_27_47#_M1005_s N_VGND_c_226_n 0.00213527f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_M1002_d N_VGND_c_226_n 0.00235968f $X=1.025 $Y=0.235 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_200_n N_VGND_c_226_n 0.01096f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_202_n N_VGND_c_226_n 0.0105687f $X=1.075 $Y=0.7 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_210_n N_VGND_c_226_n 0.00839213f $X=1.16 $Y=0.475 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__lpflow_isobufsrc_1.pex.spice
* Created: Tue Sep  1 19:12:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1%A 3 7 9 10 11 12
r30 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r31 11 12 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r32 9 16 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=0.63 $Y=1.16 $X2=0.24
+ $Y2=1.16
r33 9 10 5.03009 $w=3.3e-07 $l=7.7e-08 $layer=POLY_cond $X=0.63 $Y=1.16
+ $X2=0.707 $Y2=1.16
r34 5 10 37.0704 $w=1.5e-07 $l=1.66493e-07 $layer=POLY_cond $X=0.71 $Y=1.325
+ $X2=0.707 $Y2=1.16
r35 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.71 $Y=1.325 $X2=0.71
+ $Y2=1.695
r36 1 10 37.0704 $w=1.5e-07 $l=1.65997e-07 $layer=POLY_cond $X=0.705 $Y=0.995
+ $X2=0.707 $Y2=1.16
r37 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.705 $Y=0.995
+ $X2=0.705 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1%SLEEP 3 6 8 11 13
r39 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=1.16 $Y2=1.325
r40 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=1.16 $Y2=0.995
r41 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.16 $X2=1.16 $Y2=1.16
r42 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.25 $Y=1.985
+ $X2=1.25 $Y2=1.325
r43 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.19 $Y=0.56 $X2=1.19
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1%A_74_47# 1 2 9 12 16 19 23 25 26
+ 32 33 36
r69 33 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.16 $X2=1.7
+ $Y2=1.325
r70 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.16 $X2=1.7
+ $Y2=0.995
r71 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.16 $X2=1.7 $Y2=1.16
r72 25 28 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.545 $Y=1.595
+ $X2=0.545 $Y2=1.73
r73 25 26 4.86943 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=1.595
+ $X2=0.545 $Y2=1.51
r74 21 23 5.7039 $w=1.73e-07 $l=9e-08 $layer=LI1_cond $X=0.495 $Y=0.457
+ $X2=0.585 $Y2=0.457
r75 18 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=1.245
+ $X2=1.62 $Y2=1.16
r76 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.62 $Y=1.245
+ $X2=1.62 $Y2=1.51
r77 17 25 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.675 $Y=1.595
+ $X2=0.545 $Y2=1.595
r78 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.535 $Y=1.595
+ $X2=1.62 $Y2=1.51
r79 16 17 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.535 $Y=1.595
+ $X2=0.675 $Y2=1.595
r80 14 23 0.543965 $w=1.8e-07 $l=8.8e-08 $layer=LI1_cond $X=0.585 $Y=0.545
+ $X2=0.585 $Y2=0.457
r81 14 26 59.4596 $w=1.78e-07 $l=9.65e-07 $layer=LI1_cond $X=0.585 $Y=0.545
+ $X2=0.585 $Y2=1.51
r82 12 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.61 $Y=1.985
+ $X2=1.61 $Y2=1.325
r83 9 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.61 $Y=0.56 $X2=1.61
+ $Y2=0.995
r84 2 28 600 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_PDIFF $count=1 $X=0.375
+ $Y=1.485 $X2=0.5 $Y2=1.73
r85 1 21 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.37
+ $Y=0.235 $X2=0.495 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1%VPWR 1 6 8 10 17 18 21
r24 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r26 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=2.72
+ $X2=1.04 $Y2=2.72
r28 15 17 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.205 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 13 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.04 $Y2=2.72
r32 10 12 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.04 $Y=2.635 $X2=1.04
+ $Y2=2.72
r35 4 6 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.04 $Y=2.635
+ $X2=1.04 $Y2=2
r36 1 6 300 $w=1.7e-07 $l=6.29722e-07 $layer=licon1_PDIFF $count=2 $X=0.785
+ $Y=1.485 $X2=1.04 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1%X 1 2 9 11 12 15 18 19
r39 18 19 9.16965 $w=5.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.935 $Y=2 $X2=1.935
+ $Y2=1.85
r40 15 18 4.48529 $w=5.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.935 $Y=2.21
+ $X2=1.935 $Y2=2
r41 13 19 58.8434 $w=1.78e-07 $l=9.55e-07 $layer=LI1_cond $X=2.125 $Y=0.895
+ $X2=2.125 $Y2=1.85
r42 11 13 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.035 $Y=0.81
+ $X2=2.125 $Y2=0.895
r43 11 12 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.035 $Y=0.81
+ $X2=1.565 $Y2=0.81
r44 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.4 $Y=0.725
+ $X2=1.565 $Y2=0.81
r45 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.4 $Y=0.725 $X2=1.4
+ $Y2=0.39
r46 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.485 $X2=1.82 $Y2=2
r47 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.265
+ $Y=0.235 $X2=1.4 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1%VGND 1 2 9 11 13 16 17 18 24 30
r35 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r36 27 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r37 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r38 24 29 5.08477 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=2.017
+ $Y2=0
r39 24 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.61
+ $Y2=0
r40 22 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r41 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r42 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 16 21 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r44 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.96
+ $Y2=0
r45 15 26 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.61
+ $Y2=0
r46 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.96
+ $Y2=0
r47 11 29 3.15544 $w=3.85e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.927 $Y=0.085
+ $X2=2.017 $Y2=0
r48 11 13 9.12974 $w=3.83e-07 $l=3.05e-07 $layer=LI1_cond $X=1.927 $Y=0.085
+ $X2=1.927 $Y2=0.39
r49 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0
r50 7 9 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0.39
r51 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.235 $X2=1.82 $Y2=0.39
r52 1 9 91 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_NDIFF $count=2 $X=0.78
+ $Y=0.235 $X2=0.98 $Y2=0.39
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
M1000 KAPWR a_75_212# X VPB phighvt w=790000u l=150000u
+  ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u
M1001 a_75_212# A VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u
M1002 a_75_212# A KAPWR VPB phighvt w=790000u l=150000u
+  ad=2.054e+11p pd=2.1e+06u as=0p ps=0u
M1003 VGND a_75_212# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
.ends

* File: sky130_fd_sc_hd__a2111oi_1.pxi.spice
* Created: Thu Aug 27 13:58:58 2020
* 
x_PM_SKY130_FD_SC_HD__A2111OI_1%D1 N_D1_M1003_g N_D1_M1006_g D1 D1 D1 D1
+ N_D1_c_52_n N_D1_c_53_n N_D1_c_54_n PM_SKY130_FD_SC_HD__A2111OI_1%D1
x_PM_SKY130_FD_SC_HD__A2111OI_1%C1 N_C1_M1000_g N_C1_M1001_g C1 C1 C1 C1
+ N_C1_c_83_n N_C1_c_84_n N_C1_c_87_n PM_SKY130_FD_SC_HD__A2111OI_1%C1
x_PM_SKY130_FD_SC_HD__A2111OI_1%B1 N_B1_M1004_g N_B1_M1008_g B1 B1 B1 B1
+ N_B1_c_114_n N_B1_c_115_n PM_SKY130_FD_SC_HD__A2111OI_1%B1
x_PM_SKY130_FD_SC_HD__A2111OI_1%A1 N_A1_c_151_n N_A1_M1007_g N_A1_c_152_n
+ N_A1_M1002_g A1 N_A1_c_153_n PM_SKY130_FD_SC_HD__A2111OI_1%A1
x_PM_SKY130_FD_SC_HD__A2111OI_1%A2 N_A2_M1009_g N_A2_M1005_g N_A2_c_185_n A2 A2
+ A2 N_A2_c_188_n N_A2_c_189_n PM_SKY130_FD_SC_HD__A2111OI_1%A2
x_PM_SKY130_FD_SC_HD__A2111OI_1%Y N_Y_M1003_d N_Y_M1004_d N_Y_M1006_s
+ N_Y_c_222_n N_Y_c_249_p N_Y_c_230_n N_Y_c_233_n N_Y_c_225_n Y Y Y Y Y
+ N_Y_c_219_n PM_SKY130_FD_SC_HD__A2111OI_1%Y
x_PM_SKY130_FD_SC_HD__A2111OI_1%A_420_297# N_A_420_297#_M1008_d
+ N_A_420_297#_M1005_d N_A_420_297#_c_271_n N_A_420_297#_c_275_n
+ N_A_420_297#_c_273_n N_A_420_297#_c_286_p
+ PM_SKY130_FD_SC_HD__A2111OI_1%A_420_297#
x_PM_SKY130_FD_SC_HD__A2111OI_1%VPWR N_VPWR_M1007_d N_VPWR_c_292_n VPWR
+ N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_291_n N_VPWR_c_296_n
+ PM_SKY130_FD_SC_HD__A2111OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A2111OI_1%VGND N_VGND_M1003_s N_VGND_M1000_d
+ N_VGND_M1009_d N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n
+ N_VGND_c_332_n N_VGND_c_333_n VGND N_VGND_c_334_n N_VGND_c_335_n
+ N_VGND_c_336_n N_VGND_c_337_n PM_SKY130_FD_SC_HD__A2111OI_1%VGND
cc_1 VNB N_D1_c_52_n 0.026549f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_2 VNB N_D1_c_53_n 0.00305419f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_3 VNB N_D1_c_54_n 0.0208756f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=0.995
cc_4 VNB C1 0.00182947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_C1_c_83_n 0.0260751f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.16
cc_6 VNB N_C1_c_84_n 0.0165609f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_7 VNB B1 0.0034363f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_8 VNB N_B1_c_114_n 0.022496f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_9 VNB N_B1_c_115_n 0.01738f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=0.995
cc_10 VNB N_A1_c_151_n 0.0362645f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=0.995
cc_11 VNB N_A1_c_152_n 0.0167252f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_12 VNB N_A1_c_153_n 0.00269603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_185_n 0.003896f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_14 VNB A2 0.00243859f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.785
cc_15 VNB A2 0.0151379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_188_n 0.0336031f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_17 VNB N_A2_c_189_n 0.0196629f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=0.995
cc_18 VNB Y 0.0259069f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.19
cc_19 VNB N_Y_c_219_n 0.00754103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_291_n 0.155873f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.16
cc_21 VNB N_VGND_c_328_n 0.00555947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_329_n 0.00281836f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.16
cc_23 VNB N_VGND_c_330_n 0.0122401f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_24 VNB N_VGND_c_331_n 0.00512364f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.325
cc_25 VNB N_VGND_c_332_n 0.0115062f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.19
cc_26 VNB N_VGND_c_333_n 0.00602956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_334_n 0.0227961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_335_n 0.0391205f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_336_n 0.00507571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_337_n 0.20333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_D1_M1006_g 0.0232188f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_32 VPB N_D1_c_52_n 0.00571602f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_33 VPB N_D1_c_53_n 0.00290804f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_34 VPB C1 0.00109916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_C1_c_83_n 0.00942528f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.16
cc_36 VPB N_C1_c_87_n 0.0170714f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=0.995
cc_37 VPB N_B1_M1008_g 0.0203294f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_38 VPB B1 0.00326245f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_39 VPB B1 0.00166411f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.445
cc_40 VPB N_B1_c_114_n 0.00551977f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_41 VPB N_A1_c_151_n 0.00747022f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=0.995
cc_42 VPB N_A1_M1007_g 0.0213769f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=0.56
cc_43 VPB N_A1_c_153_n 0.0028884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A2_M1005_g 0.0261219f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_45 VPB N_A2_c_188_n 0.00703033f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_46 VPB Y 0.0493032f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.19
cc_47 VPB N_VPWR_c_292_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_48 VPB N_VPWR_c_293_n 0.074782f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.785
cc_49 VPB N_VPWR_c_294_n 0.0168006f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.325
cc_50 VPB N_VPWR_c_291_n 0.0485688f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.16
cc_51 VPB N_VPWR_c_296_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_D1_c_52_n C1 0.00143164f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_53 N_D1_c_53_n C1 0.0994047f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_54 N_D1_c_52_n N_C1_c_83_n 0.0262828f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_55 N_D1_c_53_n N_C1_c_83_n 0.0098617f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_56 N_D1_c_54_n N_C1_c_84_n 0.0167393f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_57 N_D1_M1006_g N_C1_c_87_n 0.0262828f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_58 N_D1_c_53_n N_Y_M1006_s 0.0137012f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_59 N_D1_c_52_n N_Y_c_222_n 0.00250895f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_60 N_D1_c_53_n N_Y_c_222_n 0.0179416f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_61 N_D1_c_54_n N_Y_c_222_n 0.0125037f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_62 N_D1_c_53_n N_Y_c_225_n 0.0145432f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_63 N_D1_M1006_g Y 0.00606922f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_64 N_D1_c_52_n Y 0.00790701f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_65 N_D1_c_53_n Y 0.0868105f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_66 N_D1_c_54_n Y 0.00350517f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_67 N_D1_c_53_n A_217_297# 0.00990606f $X=0.95 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_68 N_D1_M1006_g N_VPWR_c_293_n 0.00359757f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_69 N_D1_c_53_n N_VPWR_c_293_n 0.025574f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_70 N_D1_M1006_g N_VPWR_c_291_n 0.0068514f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_71 N_D1_c_53_n N_VPWR_c_291_n 0.0164812f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_72 N_D1_c_54_n N_VGND_c_328_n 0.00916907f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_73 N_D1_c_54_n N_VGND_c_329_n 0.00101145f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_74 N_D1_c_54_n N_VGND_c_334_n 0.00434414f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_75 N_D1_c_54_n N_VGND_c_337_n 0.00765318f $X=0.935 $Y=0.995 $X2=0 $Y2=0
cc_76 N_C1_c_87_n N_B1_M1008_g 0.0392656f $X=1.585 $Y=1.38 $X2=0 $Y2=0
cc_77 C1 B1 0.0750618f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_78 N_C1_c_83_n B1 0.00101123f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C1_c_87_n B1 8.86077e-19 $X=1.585 $Y=1.38 $X2=0 $Y2=0
cc_80 C1 N_B1_c_114_n 0.0050621f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_81 N_C1_c_83_n N_B1_c_114_n 0.0271117f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C1_c_84_n N_B1_c_115_n 0.0215279f $X=1.585 $Y=0.97 $X2=0 $Y2=0
cc_83 C1 N_Y_c_230_n 0.0239196f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_84 N_C1_c_83_n N_Y_c_230_n 0.00397595f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_85 N_C1_c_84_n N_Y_c_230_n 0.013137f $X=1.585 $Y=0.97 $X2=0 $Y2=0
cc_86 N_C1_c_84_n N_Y_c_233_n 7.0363e-19 $X=1.585 $Y=0.97 $X2=0 $Y2=0
cc_87 C1 A_316_297# 0.0100836f $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_88 C1 N_VPWR_c_293_n 0.0198444f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_89 N_C1_c_87_n N_VPWR_c_293_n 0.00368782f $X=1.585 $Y=1.38 $X2=0 $Y2=0
cc_90 C1 N_VPWR_c_291_n 0.0121009f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_91 N_C1_c_87_n N_VPWR_c_291_n 0.00595926f $X=1.585 $Y=1.38 $X2=0 $Y2=0
cc_92 N_C1_c_84_n N_VGND_c_329_n 0.00883522f $X=1.585 $Y=0.97 $X2=0 $Y2=0
cc_93 N_C1_c_84_n N_VGND_c_334_n 0.00347311f $X=1.585 $Y=0.97 $X2=0 $Y2=0
cc_94 N_C1_c_84_n N_VGND_c_337_n 0.00442034f $X=1.585 $Y=0.97 $X2=0 $Y2=0
cc_95 B1 N_A1_c_151_n 8.53244e-19 $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_96 N_B1_c_114_n N_A1_c_151_n 0.0231304f $X=2.105 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_97 N_B1_M1008_g N_A1_M1007_g 0.0142346f $X=2.025 $Y=1.985 $X2=0 $Y2=0
cc_98 B1 N_A1_M1007_g 0.00350902f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_99 N_B1_c_114_n N_A1_M1007_g 2.31588e-19 $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B1_c_115_n N_A1_c_152_n 0.00897431f $X=2.097 $Y=0.96 $X2=0 $Y2=0
cc_101 B1 N_A1_c_153_n 0.0288686f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_102 N_B1_c_114_n N_A1_c_153_n 0.00203559f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_103 B1 N_Y_c_230_n 0.0238246f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_104 N_B1_c_114_n N_Y_c_230_n 0.00362838f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B1_c_115_n N_Y_c_230_n 0.0103858f $X=2.097 $Y=0.96 $X2=0 $Y2=0
cc_106 N_B1_c_115_n N_Y_c_233_n 0.00555039f $X=2.097 $Y=0.96 $X2=0 $Y2=0
cc_107 B1 N_A_420_297#_M1008_d 0.0105531f $X=1.985 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_108 N_B1_M1008_g N_A_420_297#_c_271_n 0.00230185f $X=2.025 $Y=1.985 $X2=0
+ $Y2=0
cc_109 B1 N_A_420_297#_c_271_n 0.0520084f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_110 N_B1_M1008_g N_A_420_297#_c_273_n 6.28479e-19 $X=2.025 $Y=1.985 $X2=0
+ $Y2=0
cc_111 B1 N_A_420_297#_c_273_n 0.0136956f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_112 N_B1_M1008_g N_VPWR_c_293_n 0.00359757f $X=2.025 $Y=1.985 $X2=0 $Y2=0
cc_113 B1 N_VPWR_c_293_n 0.0155738f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_114 N_B1_M1008_g N_VPWR_c_291_n 0.00616599f $X=2.025 $Y=1.985 $X2=0 $Y2=0
cc_115 B1 N_VPWR_c_291_n 0.00977353f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_116 N_B1_c_115_n N_VGND_c_329_n 0.00685284f $X=2.097 $Y=0.96 $X2=0 $Y2=0
cc_117 N_B1_c_115_n N_VGND_c_335_n 0.00432079f $X=2.097 $Y=0.96 $X2=0 $Y2=0
cc_118 N_B1_c_115_n N_VGND_c_337_n 0.00676703f $X=2.097 $Y=0.96 $X2=0 $Y2=0
cc_119 N_A1_M1007_g N_A2_M1005_g 0.0291443f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A1_c_153_n N_A2_M1005_g 3.74832e-19 $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A1_c_151_n N_A2_c_185_n 0.00233384f $X=2.755 $Y=1.32 $X2=0 $Y2=0
cc_122 N_A1_c_153_n N_A2_c_185_n 0.0215686f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A1_c_152_n A2 0.0087325f $X=2.765 $Y=0.965 $X2=0 $Y2=0
cc_124 N_A1_c_153_n A2 0.00169095f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A1_c_151_n N_A2_c_188_n 0.0282404f $X=2.755 $Y=1.32 $X2=0 $Y2=0
cc_126 N_A1_c_153_n N_A2_c_188_n 4.13532e-19 $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A1_c_152_n N_A2_c_189_n 0.025279f $X=2.765 $Y=0.965 $X2=0 $Y2=0
cc_128 N_A1_c_152_n N_Y_c_230_n 0.00196122f $X=2.765 $Y=0.965 $X2=0 $Y2=0
cc_129 N_A1_c_152_n N_Y_c_233_n 0.00480205f $X=2.765 $Y=0.965 $X2=0 $Y2=0
cc_130 N_A1_M1007_g N_A_420_297#_c_275_n 0.016258f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_c_153_n N_A_420_297#_c_275_n 0.00538961f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A1_c_151_n N_A_420_297#_c_273_n 0.00108923f $X=2.755 $Y=1.32 $X2=0
+ $Y2=0
cc_133 N_A1_c_153_n N_A_420_297#_c_273_n 0.0155304f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A1_M1007_g N_VPWR_c_292_n 0.0122572f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A1_M1007_g N_VPWR_c_293_n 0.0046653f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A1_M1007_g N_VPWR_c_291_n 0.00860455f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A1_c_152_n N_VGND_c_335_n 0.00585385f $X=2.765 $Y=0.965 $X2=0 $Y2=0
cc_138 N_A1_c_152_n N_VGND_c_337_n 0.0114653f $X=2.765 $Y=0.965 $X2=0 $Y2=0
cc_139 A2 N_Y_c_230_n 0.00616287f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_140 A2 N_Y_c_233_n 0.0125136f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_141 N_A2_M1005_g N_A_420_297#_c_275_n 0.0150949f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A2_c_185_n N_A_420_297#_c_275_n 0.00946266f $X=3.09 $Y=1.155 $X2=0
+ $Y2=0
cc_143 A2 N_A_420_297#_c_275_n 0.0193024f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A2_c_188_n N_A_420_297#_c_275_n 0.00298993f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A2_M1005_g N_VPWR_c_292_n 0.0119191f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A2_M1005_g N_VPWR_c_294_n 0.00486043f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A2_M1005_g N_VPWR_c_291_n 0.00929437f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_148 A2 N_VGND_c_331_n 0.0130907f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A2_c_188_n N_VGND_c_331_n 0.00391971f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_189_n N_VGND_c_331_n 0.00740284f $X=3.27 $Y=0.965 $X2=0 $Y2=0
cc_151 A2 N_VGND_c_335_n 0.0070098f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_152 N_A2_c_189_n N_VGND_c_335_n 0.00585385f $X=3.27 $Y=0.965 $X2=0 $Y2=0
cc_153 A2 N_VGND_c_337_n 0.00669655f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_154 N_A2_c_189_n N_VGND_c_337_n 0.0116398f $X=3.27 $Y=0.965 $X2=0 $Y2=0
cc_155 A2 A_568_47# 0.0122023f $X=2.905 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_156 Y N_VPWR_c_293_n 0.0261425f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_157 N_Y_M1006_s N_VPWR_c_291_n 0.0150849f $X=0.18 $Y=1.485 $X2=0 $Y2=0
cc_158 Y N_VPWR_c_291_n 0.0147154f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_159 N_Y_c_222_n N_VGND_M1003_s 0.0168743f $X=1.045 $Y=0.79 $X2=-0.19
+ $Y2=-0.24
cc_160 N_Y_c_219_n N_VGND_M1003_s 0.00920947f $X=0.337 $Y=0.88 $X2=-0.19
+ $Y2=-0.24
cc_161 N_Y_c_230_n N_VGND_M1000_d 0.00873972f $X=2.09 $Y=0.792 $X2=0 $Y2=0
cc_162 N_Y_c_222_n N_VGND_c_328_n 0.00750157f $X=1.045 $Y=0.79 $X2=0 $Y2=0
cc_163 N_Y_c_249_p N_VGND_c_328_n 0.0113813f $X=1.21 $Y=0.39 $X2=0 $Y2=0
cc_164 N_Y_c_219_n N_VGND_c_328_n 0.0179197f $X=0.337 $Y=0.88 $X2=0 $Y2=0
cc_165 N_Y_c_230_n N_VGND_c_329_n 0.0209552f $X=2.09 $Y=0.792 $X2=0 $Y2=0
cc_166 N_Y_c_233_n N_VGND_c_329_n 0.0151756f $X=2.255 $Y=0.39 $X2=0 $Y2=0
cc_167 N_Y_c_219_n N_VGND_c_332_n 0.00287051f $X=0.337 $Y=0.88 $X2=0 $Y2=0
cc_168 N_Y_c_222_n N_VGND_c_334_n 0.00576665f $X=1.045 $Y=0.79 $X2=0 $Y2=0
cc_169 N_Y_c_249_p N_VGND_c_334_n 0.0203048f $X=1.21 $Y=0.39 $X2=0 $Y2=0
cc_170 N_Y_c_230_n N_VGND_c_334_n 0.00212146f $X=2.09 $Y=0.792 $X2=0 $Y2=0
cc_171 N_Y_c_230_n N_VGND_c_335_n 0.00260851f $X=2.09 $Y=0.792 $X2=0 $Y2=0
cc_172 N_Y_c_233_n N_VGND_c_335_n 0.0157082f $X=2.255 $Y=0.39 $X2=0 $Y2=0
cc_173 N_Y_M1003_d N_VGND_c_337_n 0.00333431f $X=1.045 $Y=0.235 $X2=0 $Y2=0
cc_174 N_Y_M1004_d N_VGND_c_337_n 0.0142155f $X=2.1 $Y=0.235 $X2=0 $Y2=0
cc_175 N_Y_c_222_n N_VGND_c_337_n 0.0108715f $X=1.045 $Y=0.79 $X2=0 $Y2=0
cc_176 N_Y_c_249_p N_VGND_c_337_n 0.012566f $X=1.21 $Y=0.39 $X2=0 $Y2=0
cc_177 N_Y_c_230_n N_VGND_c_337_n 0.0103899f $X=2.09 $Y=0.792 $X2=0 $Y2=0
cc_178 N_Y_c_233_n N_VGND_c_337_n 0.0121249f $X=2.255 $Y=0.39 $X2=0 $Y2=0
cc_179 N_Y_c_219_n N_VGND_c_337_n 0.00589719f $X=0.337 $Y=0.88 $X2=0 $Y2=0
cc_180 A_217_297# N_VPWR_c_291_n 0.00957645f $X=1.085 $Y=1.485 $X2=1.01 $Y2=1.16
cc_181 A_316_297# N_VPWR_c_291_n 0.00894463f $X=1.58 $Y=1.485 $X2=0 $Y2=0
cc_182 N_A_420_297#_c_275_n N_VPWR_M1007_d 0.00434036f $X=3.31 $Y=1.665
+ $X2=2.025 $Y2=0.96
cc_183 N_A_420_297#_c_275_n N_VPWR_c_292_n 0.0170518f $X=3.31 $Y=1.665 $X2=2.025
+ $Y2=1.985
cc_184 N_A_420_297#_c_271_n N_VPWR_c_293_n 0.0155013f $X=2.54 $Y=1.84 $X2=1.985
+ $Y2=1.785
cc_185 N_A_420_297#_c_286_p N_VPWR_c_294_n 0.0131165f $X=3.395 $Y=1.89 $X2=2.097
+ $Y2=1.33
cc_186 N_A_420_297#_M1008_d N_VPWR_c_291_n 0.0129593f $X=2.1 $Y=1.485 $X2=2.077
+ $Y2=1.4
cc_187 N_A_420_297#_M1005_d N_VPWR_c_291_n 0.00571563f $X=3.255 $Y=1.485
+ $X2=2.077 $Y2=1.4
cc_188 N_A_420_297#_c_271_n N_VPWR_c_291_n 0.00875479f $X=2.54 $Y=1.84 $X2=2.077
+ $Y2=1.4
cc_189 N_A_420_297#_c_286_p N_VPWR_c_291_n 0.00741004f $X=3.395 $Y=1.89
+ $X2=2.077 $Y2=1.4
cc_190 N_VGND_c_337_n A_568_47# 0.00482665f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
M1000 VGND SLEEP a_68_297# VNB nshort w=420000u l=150000u
+  ad=3.097e+11p pd=3.33e+06u as=1.134e+11p ps=1.38e+06u
M1001 X a_68_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1002 VPWR SLEEP a_150_297# VPB phighvt w=420000u l=150000u
+  ad=2.915e+11p pd=2.67e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_68_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_150_297# A a_68_297# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 X a_68_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.4e+11p pd=2.68e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__nand3_2.pex.spice
* Created: Tue Sep  1 19:16:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND3_2%A 1 3 6 8 10 13 15 22
r42 21 22 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r43 18 21 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r44 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r45 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r47 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r49 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r51 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%B 3 7 11 15 17 18 19 27
r51 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.16 $X2=1.82 $Y2=1.16
r52 25 27 18.6166 $w=2.9e-07 $l=9e-08 $layer=POLY_cond $X=1.73 $Y=1.16 $X2=1.82
+ $Y2=1.16
r53 23 25 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r54 19 28 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=1.82 $Y2=1.175
r55 18 28 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.82 $Y2=1.175
r56 17 18 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.615 $Y2=1.175
r57 13 25 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.73 $Y=1.305
+ $X2=1.73 $Y2=1.16
r58 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.73 $Y=1.305
+ $X2=1.73 $Y2=1.985
r59 9 25 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.73 $Y=1.015
+ $X2=1.73 $Y2=1.16
r60 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.73 $Y=1.015
+ $X2=1.73 $Y2=0.56
r61 5 23 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.31 $Y=1.305
+ $X2=1.31 $Y2=1.16
r62 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.31 $Y=1.305 $X2=1.31
+ $Y2=1.985
r63 1 23 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.31 $Y=1.015
+ $X2=1.31 $Y2=1.16
r64 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.31 $Y=1.015
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%C 3 7 9 11 14 16 17 18 23
r40 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.18
+ $Y=1.16 $X2=3.18 $Y2=1.16
r41 23 25 14.6554 $w=2.96e-07 $l=9e-08 $layer=POLY_cond $X=3.09 $Y=1.162
+ $X2=3.18 $Y2=1.162
r42 18 26 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.47 $Y=1.175
+ $X2=3.18 $Y2=1.175
r43 17 26 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.18 $Y2=1.175
r44 16 17 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=3.015 $Y2=1.175
r45 12 23 18.6531 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=3.09 $Y=1.315
+ $X2=3.09 $Y2=1.162
r46 12 14 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.09 $Y=1.315
+ $X2=3.09 $Y2=1.985
r47 9 23 18.6531 $w=1.5e-07 $l=1.52e-07 $layer=POLY_cond $X=3.09 $Y=1.01
+ $X2=3.09 $Y2=1.162
r48 9 11 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.09 $Y=1.01 $X2=3.09
+ $Y2=0.56
r49 1 23 68.3919 $w=2.96e-07 $l=4.2e-07 $layer=POLY_cond $X=2.67 $Y=1.162
+ $X2=3.09 $Y2=1.162
r50 1 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.67 $Y=1.305 $X2=2.67
+ $Y2=1.985
r51 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.67 $Y=1.015
+ $X2=2.67 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%VPWR 1 2 3 4 5 16 18 24 28 31 33 38 39 40 46
+ 50 59 63
r50 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 54 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 54 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 51 59 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.2 $Y2=2.72
r56 51 53 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 50 62 5.29703 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.447 $Y2=2.72
r58 50 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 49 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 46 59 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=2.2 $Y2=2.72
r62 46 48 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 42 56 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r66 42 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 40 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 38 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72 $X2=1.1
+ $Y2=2.72
r71 37 48 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72 $X2=1.1
+ $Y2=2.72
r73 33 36 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.405 $Y=1.66
+ $X2=3.405 $Y2=2.34
r74 31 62 2.89966 $w=3.8e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.447 $Y2=2.72
r75 31 36 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.405 $Y2=2.34
r76 26 59 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.635 $X2=2.2
+ $Y2=2.72
r77 26 28 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=2.2 $Y=2.635
+ $X2=2.2 $Y2=2
r78 22 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r79 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r80 18 21 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r81 16 56 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r82 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r83 5 36 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.33 $Y2=2.34
r84 5 33 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.33 $Y2=1.66
r85 4 28 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=2
r86 3 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r87 2 24 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r88 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r89 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%Y 1 2 3 4 15 17 21 23 25 27 30 33 34 35 42
r61 34 35 7.48369 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=0.68 $Y=1.19
+ $X2=0.68 $Y2=1.445
r62 33 34 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.85
+ $X2=0.68 $Y2=1.19
r63 33 42 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=0.85
+ $X2=0.68 $Y2=0.72
r64 25 32 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=1.555
r65 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=2.34
r66 24 30 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.555
+ $X2=1.52 $Y2=1.555
r67 23 32 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=1.555
+ $X2=2.88 $Y2=1.555
r68 23 24 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=2.715 $Y=1.555
+ $X2=1.685 $Y2=1.555
r69 19 30 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.555
r70 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r71 18 35 2.83584 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.555
+ $X2=0.68 $Y2=1.555
r72 17 30 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=1.52 $Y2=1.555
r73 17 18 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=0.845 $Y2=1.555
r74 13 35 3.64284 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.555
r75 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r76 4 32 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.66
r77 4 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2.34
r78 3 30 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r79 3 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r80 2 35 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r81 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r82 1 42 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%A_27_47# 1 2 3 10 13 17
r25 15 17 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=0.38 $X2=1.94
+ $Y2=0.38
r26 13 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.345 $Y=0.38
+ $X2=1.1 $Y2=0.38
r27 10 13 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.345 $Y2=0.38
r28 10 12 2.15294 $w=2.55e-07 $l=4.5e-08 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.217 $Y2=0.51
r29 3 17 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r30 2 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r31 1 12 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%A_277_47# 1 2 11
r22 8 11 58.049 $w=2.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.52 $Y=0.77 $X2=2.88
+ $Y2=0.77
r23 2 11 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.72
r24 1 8 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_2%VGND 1 2 9 11 13 15 17 25 31 35
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r43 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r44 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r45 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r46 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.46
+ $Y2=0
r47 26 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.99
+ $Y2=0
r48 25 34 5.29703 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.447
+ $Y2=0
r49 25 28 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=2.99
+ $Y2=0
r50 24 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r51 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r52 19 23 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r53 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.46
+ $Y2=0
r54 17 23 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.07
+ $Y2=0
r55 15 24 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r56 15 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r57 11 34 2.89966 $w=3.8e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.405 $Y=0.085
+ $X2=3.447 $Y2=0
r58 11 13 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.405 $Y=0.085
+ $X2=3.405 $Y2=0.38
r59 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085 $X2=2.46
+ $Y2=0
r60 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.38
r61 2 13 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.165
+ $Y=0.235 $X2=3.33 $Y2=0.38
r62 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.38
.ends


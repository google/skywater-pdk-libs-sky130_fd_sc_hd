* File: sky130_fd_sc_hd__maj3_2.pxi.spice
* Created: Tue Sep  1 19:14:05 2020
* 
x_PM_SKY130_FD_SC_HD__MAJ3_2%C N_C_M1008_g N_C_M1009_g N_C_M1011_g N_C_M1010_g
+ N_C_c_78_n C C C N_C_c_73_n N_C_c_74_n N_C_c_82_n N_C_c_83_n N_C_c_84_n C
+ PM_SKY130_FD_SC_HD__MAJ3_2%C
x_PM_SKY130_FD_SC_HD__MAJ3_2%A N_A_M1013_g N_A_M1004_g N_A_M1001_g N_A_M1003_g A
+ A N_A_c_159_n PM_SKY130_FD_SC_HD__MAJ3_2%A
x_PM_SKY130_FD_SC_HD__MAJ3_2%B N_B_M1002_g N_B_M1005_g N_B_M1000_g N_B_M1014_g B
+ N_B_c_203_n PM_SKY130_FD_SC_HD__MAJ3_2%B
x_PM_SKY130_FD_SC_HD__MAJ3_2%A_47_47# N_A_47_47#_M1008_s N_A_47_47#_M1002_d
+ N_A_47_47#_M1009_s N_A_47_47#_M1005_d N_A_47_47#_M1012_g N_A_47_47#_M1006_g
+ N_A_47_47#_M1015_g N_A_47_47#_M1007_g N_A_47_47#_c_248_n N_A_47_47#_c_258_n
+ N_A_47_47#_c_273_n N_A_47_47#_c_249_n N_A_47_47#_c_250_n N_A_47_47#_c_251_n
+ N_A_47_47#_c_259_n N_A_47_47#_c_252_n N_A_47_47#_c_253_n N_A_47_47#_c_261_n
+ N_A_47_47#_c_254_n N_A_47_47#_c_255_n PM_SKY130_FD_SC_HD__MAJ3_2%A_47_47#
x_PM_SKY130_FD_SC_HD__MAJ3_2%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1007_d
+ N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n
+ N_VPWR_c_393_n VPWR N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n
+ N_VPWR_c_387_n PM_SKY130_FD_SC_HD__MAJ3_2%VPWR
x_PM_SKY130_FD_SC_HD__MAJ3_2%X N_X_M1012_d N_X_M1006_s N_X_c_453_n N_X_c_458_n
+ N_X_c_450_n N_X_c_451_n X N_X_c_471_n PM_SKY130_FD_SC_HD__MAJ3_2%X
x_PM_SKY130_FD_SC_HD__MAJ3_2%VGND N_VGND_M1013_d N_VGND_M1011_d N_VGND_M1015_s
+ N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n
+ N_VGND_c_489_n VGND N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n
+ N_VGND_c_493_n PM_SKY130_FD_SC_HD__MAJ3_2%VGND
cc_1 VNB N_C_M1008_g 0.032831f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=0.445
cc_2 VNB N_C_M1011_g 0.0472988f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.445
cc_3 VNB N_C_c_73_n 0.0223893f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_4 VNB N_C_c_74_n 0.00385856f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_5 VNB N_A_M1013_g 0.0249949f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=0.445
cc_6 VNB N_A_M1001_g 0.024996f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.445
cc_7 VNB A 0.0019514f $X=-0.19 $Y=-0.24 $X2=0.775 $Y2=1.58
cc_8 VNB N_A_c_159_n 0.0292712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_M1002_g 0.0252157f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=0.445
cc_10 VNB N_B_M1000_g 0.0252157f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.445
cc_11 VNB N_B_c_203_n 0.0293333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_47_47#_M1012_g 0.0201934f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=2.165
cc_13 VNB N_A_47_47#_M1006_g 5.57054e-19 $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.495
cc_14 VNB N_A_47_47#_M1015_g 0.023255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_47_47#_M1007_g 6.82813e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_16 VNB N_A_47_47#_c_248_n 0.0144365f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.325
cc_17 VNB N_A_47_47#_c_249_n 0.0134387f $X=-0.19 $Y=-0.24 $X2=2.577 $Y2=1.54
cc_18 VNB N_A_47_47#_c_250_n 0.0033001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_47_47#_c_251_n 0.0313974f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=1.54
cc_20 VNB N_A_47_47#_c_252_n 0.0226423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_47_47#_c_253_n 0.00286921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_47_47#_c_254_n 0.00230621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_47_47#_c_255_n 0.0623849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_387_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_450_n 0.00158665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_451_n 6.17454e-19 $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=1.58
cc_27 VNB N_VGND_c_484_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_485_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_486_n 0.0101024f $X=-0.19 $Y=-0.24 $X2=0.775 $Y2=1.58
cc_30 VNB N_VGND_c_487_n 0.0353247f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_31 VNB N_VGND_c_488_n 0.0336114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_489_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_490_n 0.026269f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_34 VNB N_VGND_c_491_n 0.0221243f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.19
cc_35 VNB N_VGND_c_492_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_493_n 0.218704f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=1.53
cc_37 VPB N_C_M1009_g 0.0426367f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=2.165
cc_38 VPB N_C_M1011_g 0.00483716f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.445
cc_39 VPB N_C_M1010_g 0.0226705f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=2.165
cc_40 VPB N_C_c_78_n 0.00345395f $X=-0.19 $Y=1.305 $X2=0.775 $Y2=1.58
cc_41 VPB C 0.00949675f $X=-0.19 $Y=1.305 $X2=2.9 $Y2=1.445
cc_42 VPB N_C_c_73_n 0.00477149f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_43 VPB N_C_c_74_n 0.00338512f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_44 VPB N_C_c_82_n 0.0282764f $X=-0.19 $Y=1.305 $X2=2.58 $Y2=1.52
cc_45 VPB N_C_c_83_n 9.20478e-19 $X=-0.19 $Y=1.305 $X2=2.54 $Y2=1.54
cc_46 VPB N_C_c_84_n 0.0265534f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=1.54
cc_47 VPB N_A_M1004_g 0.0337272f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=2.165
cc_48 VPB N_A_M1003_g 0.0337549f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=2.165
cc_49 VPB A 0.0019514f $X=-0.19 $Y=1.305 $X2=0.775 $Y2=1.58
cc_50 VPB N_A_c_159_n 0.00391365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_B_M1005_g 0.0339828f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=2.165
cc_52 VPB N_B_M1014_g 0.0340519f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=2.165
cc_53 VPB N_B_c_203_n 0.00391774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_47_47#_M1006_g 0.0224841f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.495
cc_55 VPB N_A_47_47#_M1007_g 0.0268951f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_56 VPB N_A_47_47#_c_258_n 0.00614851f $X=-0.19 $Y=1.305 $X2=2.58 $Y2=1.52
cc_57 VPB N_A_47_47#_c_259_n 0.0355743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_47_47#_c_252_n 0.0251463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_47_47#_c_261_n 0.00234947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_388_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_389_n 0.00510406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_390_n 0.0100765f $X=-0.19 $Y=1.305 $X2=0.775 $Y2=1.58
cc_63 VPB N_VPWR_c_391_n 0.043721f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_64 VPB N_VPWR_c_392_n 0.0319555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_393_n 0.00498265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_394_n 0.0256239f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_67 VPB N_VPWR_c_395_n 0.0260603f $X=-0.19 $Y=1.305 $X2=2.577 $Y2=1.54
cc_68 VPB N_VPWR_c_396_n 0.00436611f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=1.54
cc_69 VPB N_VPWR_c_387_n 0.0438828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_X_c_451_n 0.00126449f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=1.58
cc_71 N_C_M1008_g N_A_M1013_g 0.0520385f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_72 N_C_M1009_g N_A_M1004_g 0.0520385f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_73 N_C_c_84_n N_A_M1004_g 0.0122069f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_74 N_C_c_84_n N_A_M1003_g 0.00992836f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_75 N_C_c_73_n A 2.64217e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_76 N_C_c_74_n A 0.0220365f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_c_84_n A 0.0519418f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_78 N_C_c_73_n N_A_c_159_n 0.0520385f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C_c_74_n N_A_c_159_n 0.0071019f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_80 N_C_c_84_n N_A_c_159_n 0.00201785f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_81 N_C_c_84_n N_B_M1005_g 0.0112936f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_82 N_C_M1011_g N_B_M1000_g 0.0524142f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_83 N_C_M1010_g N_B_M1014_g 0.0524142f $X=2.49 $Y=2.165 $X2=0 $Y2=0
cc_84 N_C_c_83_n N_B_M1014_g 5.22213e-19 $X=2.54 $Y=1.54 $X2=0 $Y2=0
cc_85 N_C_c_84_n N_B_M1014_g 0.0143516f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_86 N_C_M1011_g B 0.00194394f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_87 N_C_c_84_n B 0.0214226f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_88 N_C_c_82_n N_B_c_203_n 0.0524142f $X=2.58 $Y=1.52 $X2=0 $Y2=0
cc_89 N_C_c_84_n N_B_c_203_n 0.00201785f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_90 N_C_M1011_g N_A_47_47#_M1012_g 0.0139602f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_91 N_C_M1011_g N_A_47_47#_M1006_g 0.00224384f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_92 N_C_M1010_g N_A_47_47#_M1006_g 0.0105969f $X=2.49 $Y=2.165 $X2=0 $Y2=0
cc_93 C N_A_47_47#_M1006_g 0.00361411f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_94 N_C_c_82_n N_A_47_47#_M1006_g 0.00654515f $X=2.58 $Y=1.52 $X2=0 $Y2=0
cc_95 N_C_M1008_g N_A_47_47#_c_248_n 0.00838569f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_96 N_C_c_74_n N_A_47_47#_c_248_n 0.0200117f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_97 N_C_c_84_n N_A_47_47#_c_248_n 0.00680892f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_98 N_C_M1009_g N_A_47_47#_c_258_n 0.00367116f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_99 N_C_c_78_n N_A_47_47#_c_258_n 0.0132022f $X=0.775 $Y=1.58 $X2=0 $Y2=0
cc_100 N_C_c_84_n N_A_47_47#_c_258_n 0.0705647f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_101 N_C_M1011_g N_A_47_47#_c_273_n 0.00152276f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_102 N_C_M1011_g N_A_47_47#_c_249_n 0.014581f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_103 N_C_c_82_n N_A_47_47#_c_249_n 0.00291106f $X=2.58 $Y=1.52 $X2=0 $Y2=0
cc_104 N_C_c_83_n N_A_47_47#_c_249_n 0.0146579f $X=2.54 $Y=1.54 $X2=0 $Y2=0
cc_105 N_C_c_84_n N_A_47_47#_c_249_n 0.00712919f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_106 N_C_M1011_g N_A_47_47#_c_250_n 0.0046356f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_107 N_C_M1008_g N_A_47_47#_c_251_n 0.0120523f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_108 N_C_c_73_n N_A_47_47#_c_251_n 0.00272381f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_109 N_C_c_74_n N_A_47_47#_c_251_n 0.0084508f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_110 N_C_M1009_g N_A_47_47#_c_259_n 0.0155322f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_111 N_C_c_78_n N_A_47_47#_c_259_n 0.0165181f $X=0.775 $Y=1.58 $X2=0 $Y2=0
cc_112 N_C_c_73_n N_A_47_47#_c_259_n 0.00180964f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_113 N_C_M1008_g N_A_47_47#_c_252_n 0.00379516f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_114 N_C_M1009_g N_A_47_47#_c_252_n 0.00583364f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_115 N_C_c_78_n N_A_47_47#_c_252_n 0.0143566f $X=0.775 $Y=1.58 $X2=0 $Y2=0
cc_116 N_C_c_73_n N_A_47_47#_c_252_n 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_117 N_C_c_74_n N_A_47_47#_c_252_n 0.0384102f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C_c_84_n N_A_47_47#_c_253_n 0.0032605f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_119 N_C_M1010_g N_A_47_47#_c_261_n 0.00172059f $X=2.49 $Y=2.165 $X2=0 $Y2=0
cc_120 N_C_c_84_n N_A_47_47#_c_261_n 0.0272027f $X=2.415 $Y=1.54 $X2=0 $Y2=0
cc_121 N_C_M1011_g N_A_47_47#_c_254_n 0.00333506f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_122 C N_A_47_47#_c_254_n 0.010775f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_123 N_C_M1011_g N_A_47_47#_c_255_n 0.00839435f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_124 C N_A_47_47#_c_255_n 0.0028814f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_125 C N_VPWR_M1010_d 0.00934441f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_126 N_C_M1009_g N_VPWR_c_388_n 0.0019774f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_127 N_C_M1010_g N_VPWR_c_389_n 0.0164756f $X=2.49 $Y=2.165 $X2=0 $Y2=0
cc_128 N_C_c_82_n N_VPWR_c_389_n 0.00139198f $X=2.58 $Y=1.52 $X2=0 $Y2=0
cc_129 N_C_c_83_n N_VPWR_c_389_n 0.0277316f $X=2.54 $Y=1.54 $X2=0 $Y2=0
cc_130 N_C_M1010_g N_VPWR_c_392_n 0.0046653f $X=2.49 $Y=2.165 $X2=0 $Y2=0
cc_131 N_C_M1009_g N_VPWR_c_394_n 0.0037495f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_132 N_C_M1009_g N_VPWR_c_387_n 0.00628054f $X=0.57 $Y=2.165 $X2=0 $Y2=0
cc_133 N_C_M1010_g N_VPWR_c_387_n 0.00783311f $X=2.49 $Y=2.165 $X2=0 $Y2=0
cc_134 C N_X_c_453_n 0.0116124f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_135 C N_X_c_451_n 0.00140415f $X=2.9 $Y=1.445 $X2=0 $Y2=0
cc_136 N_C_M1008_g N_VGND_c_484_n 0.00191424f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_137 N_C_M1011_g N_VGND_c_485_n 0.00746397f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_138 N_C_M1011_g N_VGND_c_488_n 0.00428022f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_139 N_C_M1008_g N_VGND_c_490_n 0.00416472f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_140 N_C_M1008_g N_VGND_c_493_n 0.00672809f $X=0.57 $Y=0.445 $X2=0 $Y2=0
cc_141 N_C_M1011_g N_VGND_c_493_n 0.00638372f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1001_g N_B_M1002_g 0.0528781f $X=1.35 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_M1003_g N_B_M1005_g 0.0528781f $X=1.35 $Y=2.165 $X2=0 $Y2=0
cc_144 A B 0.0261078f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_145 A N_B_c_203_n 0.0112868f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A_c_159_n N_B_c_203_n 0.0528781f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_M1013_g N_A_47_47#_c_248_n 0.0133608f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_M1001_g N_A_47_47#_c_248_n 0.0110822f $X=1.35 $Y=0.445 $X2=0 $Y2=0
cc_149 A N_A_47_47#_c_248_n 0.0519418f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A_c_159_n N_A_47_47#_c_248_n 0.00201785f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_M1004_g N_A_47_47#_c_258_n 0.011279f $X=0.93 $Y=2.165 $X2=0 $Y2=0
cc_152 N_A_M1003_g N_A_47_47#_c_258_n 0.011279f $X=1.35 $Y=2.165 $X2=0 $Y2=0
cc_153 N_A_M1001_g N_A_47_47#_c_273_n 0.00148749f $X=1.35 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A_M1013_g N_A_47_47#_c_251_n 0.00149485f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_M1004_g N_A_47_47#_c_259_n 0.0020623f $X=0.93 $Y=2.165 $X2=0 $Y2=0
cc_156 N_A_M1003_g N_A_47_47#_c_261_n 0.00165163f $X=1.35 $Y=2.165 $X2=0 $Y2=0
cc_157 N_A_M1004_g N_VPWR_c_388_n 0.00982588f $X=0.93 $Y=2.165 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_VPWR_c_388_n 0.010314f $X=1.35 $Y=2.165 $X2=0 $Y2=0
cc_159 N_A_M1003_g N_VPWR_c_392_n 0.00348405f $X=1.35 $Y=2.165 $X2=0 $Y2=0
cc_160 N_A_M1004_g N_VPWR_c_394_n 0.00348405f $X=0.93 $Y=2.165 $X2=0 $Y2=0
cc_161 N_A_M1004_g N_VPWR_c_387_n 0.00401101f $X=0.93 $Y=2.165 $X2=0 $Y2=0
cc_162 N_A_M1003_g N_VPWR_c_387_n 0.00401101f $X=1.35 $Y=2.165 $X2=0 $Y2=0
cc_163 N_A_M1013_g N_VGND_c_484_n 0.00938687f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_M1001_g N_VGND_c_484_n 0.00934722f $X=1.35 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_M1001_g N_VGND_c_488_n 0.00341689f $X=1.35 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_M1013_g N_VGND_c_490_n 0.00341689f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A_M1013_g N_VGND_c_493_n 0.00389164f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_M1001_g N_VGND_c_493_n 0.00389164f $X=1.35 $Y=0.445 $X2=0 $Y2=0
cc_169 N_B_M1002_g N_A_47_47#_c_248_n 0.00870428f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_170 N_B_M1005_g N_A_47_47#_c_258_n 0.00800193f $X=1.71 $Y=2.165 $X2=0 $Y2=0
cc_171 N_B_M1002_g N_A_47_47#_c_273_n 0.00808019f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_172 N_B_M1000_g N_A_47_47#_c_273_n 0.00845957f $X=2.13 $Y=0.445 $X2=0 $Y2=0
cc_173 N_B_M1000_g N_A_47_47#_c_249_n 0.00856756f $X=2.13 $Y=0.445 $X2=0 $Y2=0
cc_174 B N_A_47_47#_c_249_n 0.00496499f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_175 N_B_M1002_g N_A_47_47#_c_253_n 0.00332168f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_176 N_B_M1000_g N_A_47_47#_c_253_n 0.00285314f $X=2.13 $Y=0.445 $X2=0 $Y2=0
cc_177 B N_A_47_47#_c_253_n 0.0181557f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_178 N_B_c_203_n N_A_47_47#_c_253_n 0.00208238f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_M1005_g N_A_47_47#_c_261_n 0.00887855f $X=1.71 $Y=2.165 $X2=0 $Y2=0
cc_180 N_B_M1014_g N_A_47_47#_c_261_n 0.010889f $X=2.13 $Y=2.165 $X2=0 $Y2=0
cc_181 N_B_M1005_g N_VPWR_c_388_n 0.00202008f $X=1.71 $Y=2.165 $X2=0 $Y2=0
cc_182 N_B_M1014_g N_VPWR_c_389_n 0.00294882f $X=2.13 $Y=2.165 $X2=0 $Y2=0
cc_183 N_B_M1005_g N_VPWR_c_392_n 0.00422241f $X=1.71 $Y=2.165 $X2=0 $Y2=0
cc_184 N_B_M1014_g N_VPWR_c_392_n 0.00541359f $X=2.13 $Y=2.165 $X2=0 $Y2=0
cc_185 N_B_M1005_g N_VPWR_c_387_n 0.00572905f $X=1.71 $Y=2.165 $X2=0 $Y2=0
cc_186 N_B_M1014_g N_VPWR_c_387_n 0.00956562f $X=2.13 $Y=2.165 $X2=0 $Y2=0
cc_187 N_B_M1002_g N_VGND_c_484_n 0.00185594f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_188 N_B_M1002_g N_VGND_c_488_n 0.00415469f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_189 N_B_M1000_g N_VGND_c_488_n 0.00415469f $X=2.13 $Y=0.445 $X2=0 $Y2=0
cc_190 N_B_M1002_g N_VGND_c_493_n 0.00561067f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_191 N_B_M1000_g N_VGND_c_493_n 0.00561067f $X=2.13 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A_47_47#_c_258_n A_129_369# 0.0018249f $X=1.755 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_193 N_A_47_47#_c_258_n N_VPWR_M1004_d 0.00161592f $X=1.755 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_194 N_A_47_47#_c_258_n N_VPWR_c_388_n 0.0163351f $X=1.755 $Y=1.92 $X2=0 $Y2=0
cc_195 N_A_47_47#_c_259_n N_VPWR_c_388_n 0.0123624f $X=0.35 $Y=1.92 $X2=0 $Y2=0
cc_196 N_A_47_47#_c_261_n N_VPWR_c_388_n 0.00988691f $X=1.92 $Y=2 $X2=0 $Y2=0
cc_197 N_A_47_47#_M1006_g N_VPWR_c_389_n 0.00835802f $X=3.24 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_47_47#_c_261_n N_VPWR_c_389_n 0.021788f $X=1.92 $Y=2 $X2=0 $Y2=0
cc_199 N_A_47_47#_M1007_g N_VPWR_c_391_n 0.00451776f $X=3.66 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_47_47#_c_258_n N_VPWR_c_392_n 0.00559495f $X=1.755 $Y=1.92 $X2=0
+ $Y2=0
cc_201 N_A_47_47#_c_261_n N_VPWR_c_392_n 0.0188215f $X=1.92 $Y=2 $X2=0 $Y2=0
cc_202 N_A_47_47#_c_258_n N_VPWR_c_394_n 0.00436946f $X=1.755 $Y=1.92 $X2=0
+ $Y2=0
cc_203 N_A_47_47#_c_259_n N_VPWR_c_394_n 0.0349444f $X=0.35 $Y=1.92 $X2=0 $Y2=0
cc_204 N_A_47_47#_M1006_g N_VPWR_c_395_n 0.00541359f $X=3.24 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_47_47#_M1007_g N_VPWR_c_395_n 0.00541359f $X=3.66 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_47_47#_M1009_s N_VPWR_c_387_n 0.00209319f $X=0.235 $Y=1.845 $X2=0
+ $Y2=0
cc_207 N_A_47_47#_M1005_d N_VPWR_c_387_n 0.00215201f $X=1.785 $Y=1.845 $X2=0
+ $Y2=0
cc_208 N_A_47_47#_M1006_g N_VPWR_c_387_n 0.0103658f $X=3.24 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_47_47#_M1007_g N_VPWR_c_387_n 0.0104652f $X=3.66 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_47_47#_c_258_n N_VPWR_c_387_n 0.0209323f $X=1.755 $Y=1.92 $X2=0 $Y2=0
cc_211 N_A_47_47#_c_259_n N_VPWR_c_387_n 0.0196901f $X=0.35 $Y=1.92 $X2=0 $Y2=0
cc_212 N_A_47_47#_c_261_n N_VPWR_c_387_n 0.0121968f $X=1.92 $Y=2 $X2=0 $Y2=0
cc_213 N_A_47_47#_c_258_n A_285_369# 0.0018249f $X=1.755 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_47_47#_M1006_g N_X_c_453_n 0.00267339f $X=3.24 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_47_47#_M1007_g N_X_c_453_n 0.00181417f $X=3.66 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_47_47#_c_255_n N_X_c_453_n 0.00108933f $X=3.66 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_47_47#_M1006_g N_X_c_458_n 0.0187224f $X=3.24 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_47_47#_M1007_g N_X_c_458_n 0.00907982f $X=3.66 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_47_47#_M1012_g N_X_c_450_n 0.0028418f $X=3.24 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A_47_47#_M1015_g N_X_c_450_n 0.00203593f $X=3.66 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A_47_47#_c_250_n N_X_c_450_n 0.00566735f $X=3.015 $Y=1.075 $X2=0 $Y2=0
cc_222 N_A_47_47#_c_255_n N_X_c_450_n 0.00120248f $X=3.66 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_47_47#_M1012_g N_X_c_451_n 5.50891e-19 $X=3.24 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_47_47#_M1006_g N_X_c_451_n 0.00285149f $X=3.24 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_47_47#_M1015_g N_X_c_451_n 0.00618421f $X=3.66 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A_47_47#_M1007_g N_X_c_451_n 0.00988228f $X=3.66 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_47_47#_c_250_n N_X_c_451_n 0.00521937f $X=3.015 $Y=1.075 $X2=0 $Y2=0
cc_228 N_A_47_47#_c_254_n N_X_c_451_n 0.0121172f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_47_47#_c_255_n N_X_c_451_n 0.0223629f $X=3.66 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_47_47#_M1012_g N_X_c_471_n 0.0120424f $X=3.24 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_47_47#_M1015_g N_X_c_471_n 0.00556143f $X=3.66 $Y=0.56 $X2=0 $Y2=0
cc_232 N_A_47_47#_c_249_n N_X_c_471_n 0.0133942f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_47_47#_c_249_n N_VGND_M1011_d 0.00903141f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_47_47#_c_250_n N_VGND_M1011_d 0.00148529f $X=3.015 $Y=1.075 $X2=0
+ $Y2=0
cc_235 N_A_47_47#_c_248_n N_VGND_c_484_n 0.020154f $X=1.755 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_47_47#_c_273_n N_VGND_c_484_n 0.00784134f $X=1.92 $Y=0.36 $X2=0 $Y2=0
cc_237 N_A_47_47#_c_251_n N_VGND_c_484_n 0.00714625f $X=0.36 $Y=0.445 $X2=0
+ $Y2=0
cc_238 N_A_47_47#_M1012_g N_VGND_c_485_n 0.0052788f $X=3.24 $Y=0.56 $X2=0 $Y2=0
cc_239 N_A_47_47#_c_273_n N_VGND_c_485_n 0.00711496f $X=1.92 $Y=0.36 $X2=0 $Y2=0
cc_240 N_A_47_47#_c_249_n N_VGND_c_485_n 0.0256109f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A_47_47#_M1015_g N_VGND_c_487_n 0.00496233f $X=3.66 $Y=0.56 $X2=0 $Y2=0
cc_242 N_A_47_47#_c_248_n N_VGND_c_488_n 0.0074151f $X=1.755 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_47_47#_c_273_n N_VGND_c_488_n 0.018715f $X=1.92 $Y=0.36 $X2=0 $Y2=0
cc_244 N_A_47_47#_c_249_n N_VGND_c_488_n 0.00911064f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_47_47#_c_248_n N_VGND_c_490_n 0.00742144f $X=1.755 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_47_47#_c_251_n N_VGND_c_490_n 0.0247545f $X=0.36 $Y=0.445 $X2=0 $Y2=0
cc_247 N_A_47_47#_M1012_g N_VGND_c_491_n 0.00541359f $X=3.24 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_47_47#_M1015_g N_VGND_c_491_n 0.00541359f $X=3.66 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A_47_47#_c_249_n N_VGND_c_491_n 0.00249459f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_47_47#_M1008_s N_VGND_c_493_n 0.00211233f $X=0.235 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_47_47#_M1002_d N_VGND_c_493_n 0.00215201f $X=1.785 $Y=0.235 $X2=0
+ $Y2=0
cc_252 N_A_47_47#_M1012_g N_VGND_c_493_n 0.0103658f $X=3.24 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A_47_47#_M1015_g N_VGND_c_493_n 0.0104652f $X=3.66 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_47_47#_c_248_n N_VGND_c_493_n 0.0241551f $X=1.755 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_47_47#_c_273_n N_VGND_c_493_n 0.0121647f $X=1.92 $Y=0.36 $X2=0 $Y2=0
cc_256 N_A_47_47#_c_249_n N_VGND_c_493_n 0.0195526f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_47_47#_c_251_n N_VGND_c_493_n 0.0164556f $X=0.36 $Y=0.445 $X2=0 $Y2=0
cc_258 A_129_369# N_VPWR_c_387_n 0.00269901f $X=0.645 $Y=1.845 $X2=0.35 $Y2=1.92
cc_259 N_VPWR_c_387_n A_285_369# 0.00269901f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_260 N_VPWR_c_387_n A_441_369# 0.00897657f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_261 N_VPWR_c_387_n N_X_M1006_s 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_262 N_VPWR_c_389_n N_X_c_458_n 0.0241158f $X=2.7 $Y=2 $X2=0 $Y2=0
cc_263 N_VPWR_c_395_n N_X_c_458_n 0.0189039f $X=3.785 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_c_387_n N_X_c_458_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_265 N_VPWR_c_391_n N_VGND_c_487_n 0.00998764f $X=3.87 $Y=1.66 $X2=0 $Y2=0
cc_266 N_X_c_471_n N_VGND_c_485_n 0.0109935f $X=3.45 $Y=0.4 $X2=0 $Y2=0
cc_267 N_X_c_471_n N_VGND_c_487_n 0.0251189f $X=3.45 $Y=0.4 $X2=0 $Y2=0
cc_268 N_X_c_471_n N_VGND_c_491_n 0.0188807f $X=3.45 $Y=0.4 $X2=0 $Y2=0
cc_269 N_X_M1012_d N_VGND_c_493_n 0.00215201f $X=3.315 $Y=0.235 $X2=0 $Y2=0
cc_270 N_X_c_471_n N_VGND_c_493_n 0.0122146f $X=3.45 $Y=0.4 $X2=0 $Y2=0
cc_271 A_129_47# N_VGND_c_493_n 0.00251327f $X=0.645 $Y=0.235 $X2=3.91 $Y2=0
cc_272 N_VGND_c_493_n A_285_47# 0.00251327f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_273 N_VGND_c_493_n A_441_47# 0.00251327f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

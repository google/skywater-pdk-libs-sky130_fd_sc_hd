* File: sky130_fd_sc_hd__mux2i_4.spice
* Created: Thu Aug 27 14:28:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2i_4.spice.pex"
.subckt sky130_fd_sc_hd__mux2i_4  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1015 N_Y_M1015_d N_A0_M1015_g N_A_109_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_A0_M1018_g N_A_109_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1018_d N_A0_M1023_g N_A_109_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1033 N_Y_M1033_d N_A0_M1033_g N_A_109_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1019 N_A_445_47#_M1019_d N_A1_M1019_g N_Y_M1033_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1025 N_A_445_47#_M1019_d N_A1_M1025_g N_Y_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1028 N_A_445_47#_M1028_d N_A1_M1028_g N_Y_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1029 N_A_445_47#_M1028_d N_A1_M1029_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_445_47#_M1012_d N_S_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_445_47#_M1012_d N_S_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1020 N_A_445_47#_M1020_d N_S_M1020_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1026 N_A_445_47#_M1020_d N_S_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1026_s N_A_1191_21#_M1003_g N_A_109_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75002 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_1191_21#_M1009_g N_A_109_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1009_d N_A_1191_21#_M1013_g N_A_109_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.105625 PD=0.92 PS=0.975 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A_1191_21#_M1021_g N_A_109_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.102375 AS=0.105625 PD=0.965 PS=0.975 NRD=7.38 NRS=9.228 M=1
+ R=4.33333 SA=75003.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_1191_21#_M1010_d N_S_M1010_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.102375 PD=1.82 PS=0.965 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_109_297#_M1004_d N_A0_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1006 N_A_109_297#_M1004_d N_A0_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1024 N_A_109_297#_M1024_d N_A0_M1024_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1030 N_A_109_297#_M1024_d N_A0_M1030_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_A_445_297#_M1000_d N_A1_M1000_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 N_A_445_297#_M1000_d N_A1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1027 N_A_445_297#_M1027_d N_A1_M1027_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1031 N_A_445_297#_M1027_d N_A1_M1031_g N_Y_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_109_297#_M1001_d N_S_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1011 N_A_109_297#_M1001_d N_S_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_109_297#_M1014_d N_S_M1014_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1032 N_A_109_297#_M1014_d N_S_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1002 N_A_445_297#_M1002_d N_A_1191_21#_M1002_g N_VPWR_M1032_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75002 A=0.15 P=2.3 MULT=1
MM1005 N_A_445_297#_M1002_d N_A_1191_21#_M1005_g N_VPWR_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1008 N_A_445_297#_M1008_d N_A_1191_21#_M1008_g N_VPWR_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.1625 AS=0.135 PD=1.325 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1022 N_A_445_297#_M1008_d N_A_1191_21#_M1022_g N_VPWR_M1022_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.1625 AS=0.1575 PD=1.325 PS=1.315 NRD=9.8303 NRS=7.8603 M=1
+ R=6.66667 SA=75003.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_A_1191_21#_M1017_d N_S_M1017_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1575 PD=2.52 PS=1.315 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX34_noxref VNB VPB NWDIODE A=13.8993 P=20.53
c_60 VNB 0 1.39126e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__mux2i_4.spice.SKY130_FD_SC_HD__MUX2I_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__xor3_1.pxi.spice
* Created: Thu Aug 27 14:50:04 2020
* 
x_PM_SKY130_FD_SC_HD__XOR3_1%A_112_21# N_A_112_21#_M1019_d N_A_112_21#_M1004_d
+ N_A_112_21#_c_162_n N_A_112_21#_M1001_g N_A_112_21#_M1002_g
+ N_A_112_21#_c_163_n N_A_112_21#_c_170_n N_A_112_21#_c_177_p
+ N_A_112_21#_c_182_p N_A_112_21#_c_220_p N_A_112_21#_c_164_n
+ N_A_112_21#_c_171_n N_A_112_21#_c_165_n N_A_112_21#_c_172_n
+ N_A_112_21#_c_173_n N_A_112_21#_c_166_n N_A_112_21#_c_187_p
+ N_A_112_21#_c_167_n PM_SKY130_FD_SC_HD__XOR3_1%A_112_21#
x_PM_SKY130_FD_SC_HD__XOR3_1%C N_C_c_264_n N_C_M1005_g N_C_c_270_n N_C_M1003_g
+ N_C_c_265_n N_C_M1004_g N_C_c_266_n N_C_M1019_g N_C_c_267_n C N_C_c_268_n
+ N_C_c_269_n PM_SKY130_FD_SC_HD__XOR3_1%C
x_PM_SKY130_FD_SC_HD__XOR3_1%A_266_93# N_A_266_93#_M1005_d N_A_266_93#_M1003_d
+ N_A_266_93#_M1020_g N_A_266_93#_M1013_g N_A_266_93#_c_346_n
+ N_A_266_93#_c_332_n N_A_266_93#_c_338_n N_A_266_93#_c_339_n
+ N_A_266_93#_c_340_n N_A_266_93#_c_333_n N_A_266_93#_c_334_n
+ N_A_266_93#_c_335_n PM_SKY130_FD_SC_HD__XOR3_1%A_266_93#
x_PM_SKY130_FD_SC_HD__XOR3_1%A_827_297# N_A_827_297#_M1012_d
+ N_A_827_297#_M1000_d N_A_827_297#_M1018_g N_A_827_297#_M1015_g
+ N_A_827_297#_c_411_n N_A_827_297#_M1008_g N_A_827_297#_c_413_n
+ N_A_827_297#_M1010_g N_A_827_297#_c_414_n N_A_827_297#_c_415_n
+ N_A_827_297#_c_428_n N_A_827_297#_c_416_n N_A_827_297#_c_417_n
+ N_A_827_297#_c_432_p N_A_827_297#_c_418_n N_A_827_297#_c_419_n
+ N_A_827_297#_c_420_n N_A_827_297#_c_421_n N_A_827_297#_c_422_n
+ N_A_827_297#_c_423_n PM_SKY130_FD_SC_HD__XOR3_1%A_827_297#
x_PM_SKY130_FD_SC_HD__XOR3_1%B N_B_M1000_g N_B_M1012_g N_B_c_581_n N_B_c_582_n
+ N_B_M1016_g N_B_M1017_g N_B_c_591_n N_B_c_592_n N_B_M1021_g N_B_M1011_g
+ N_B_c_585_n N_B_c_586_n N_B_c_587_n N_B_c_596_n B N_B_c_588_n
+ PM_SKY130_FD_SC_HD__XOR3_1%B
x_PM_SKY130_FD_SC_HD__XOR3_1%A N_A_M1007_g N_A_M1014_g A N_A_c_701_n N_A_c_702_n
+ N_A_c_703_n PM_SKY130_FD_SC_HD__XOR3_1%A
x_PM_SKY130_FD_SC_HD__XOR3_1%A_931_365# N_A_931_365#_M1016_s
+ N_A_931_365#_M1010_d N_A_931_365#_M1017_s N_A_931_365#_M1008_d
+ N_A_931_365#_c_745_n N_A_931_365#_M1006_g N_A_931_365#_M1009_g
+ N_A_931_365#_c_746_n N_A_931_365#_c_755_n N_A_931_365#_c_747_n
+ N_A_931_365#_c_748_n N_A_931_365#_c_749_n N_A_931_365#_c_757_n
+ N_A_931_365#_c_750_n N_A_931_365#_c_768_n N_A_931_365#_c_751_n
+ N_A_931_365#_c_752_n N_A_931_365#_c_781_n N_A_931_365#_c_782_n
+ PM_SKY130_FD_SC_HD__XOR3_1%A_931_365#
x_PM_SKY130_FD_SC_HD__XOR3_1%X N_X_M1001_s N_X_M1002_s N_X_c_880_n N_X_c_882_n
+ N_X_c_881_n X PM_SKY130_FD_SC_HD__XOR3_1%X
x_PM_SKY130_FD_SC_HD__XOR3_1%VPWR N_VPWR_M1002_d N_VPWR_M1000_s N_VPWR_M1014_d
+ N_VPWR_c_905_n N_VPWR_c_906_n N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n
+ VPWR N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_904_n
+ N_VPWR_c_914_n N_VPWR_c_915_n PM_SKY130_FD_SC_HD__XOR3_1%VPWR
x_PM_SKY130_FD_SC_HD__XOR3_1%A_386_325# N_A_386_325#_M1013_d
+ N_A_386_325#_M1021_d N_A_386_325#_M1004_s N_A_386_325#_M1017_d
+ N_A_386_325#_c_1001_n N_A_386_325#_c_1022_n N_A_386_325#_c_999_n
+ N_A_386_325#_c_1003_n N_A_386_325#_c_1039_n N_A_386_325#_c_1004_n
+ N_A_386_325#_c_1000_n N_A_386_325#_c_1126_p N_A_386_325#_c_1050_n
+ N_A_386_325#_c_1070_n N_A_386_325#_c_1006_n N_A_386_325#_c_1007_n
+ N_A_386_325#_c_1008_n N_A_386_325#_c_1009_n
+ PM_SKY130_FD_SC_HD__XOR3_1%A_386_325#
x_PM_SKY130_FD_SC_HD__XOR3_1%A_404_49# N_A_404_49#_M1019_s N_A_404_49#_M1016_d
+ N_A_404_49#_M1020_d N_A_404_49#_M1011_d N_A_404_49#_c_1140_n
+ N_A_404_49#_c_1164_n N_A_404_49#_c_1141_n N_A_404_49#_c_1165_n
+ N_A_404_49#_c_1147_n N_A_404_49#_c_1148_n N_A_404_49#_c_1149_n
+ N_A_404_49#_c_1142_n N_A_404_49#_c_1143_n N_A_404_49#_c_1151_n
+ N_A_404_49#_c_1152_n N_A_404_49#_c_1153_n N_A_404_49#_c_1154_n
+ N_A_404_49#_c_1144_n N_A_404_49#_c_1156_n N_A_404_49#_c_1200_n
+ N_A_404_49#_c_1157_n N_A_404_49#_c_1145_n N_A_404_49#_c_1158_n
+ N_A_404_49#_c_1146_n N_A_404_49#_c_1159_n PM_SKY130_FD_SC_HD__XOR3_1%A_404_49#
x_PM_SKY130_FD_SC_HD__XOR3_1%A_1198_49# N_A_1198_49#_M1018_d
+ N_A_1198_49#_M1006_d N_A_1198_49#_M1015_d N_A_1198_49#_M1009_d
+ N_A_1198_49#_c_1321_n N_A_1198_49#_c_1333_n N_A_1198_49#_c_1325_n
+ N_A_1198_49#_c_1322_n N_A_1198_49#_c_1334_n N_A_1198_49#_c_1327_n
+ N_A_1198_49#_c_1323_n PM_SKY130_FD_SC_HD__XOR3_1%A_1198_49#
x_PM_SKY130_FD_SC_HD__XOR3_1%VGND N_VGND_M1001_d N_VGND_M1012_s N_VGND_M1007_d
+ N_VGND_c_1388_n N_VGND_c_1389_n N_VGND_c_1390_n N_VGND_c_1391_n
+ N_VGND_c_1392_n N_VGND_c_1393_n N_VGND_c_1394_n N_VGND_c_1395_n
+ N_VGND_c_1396_n VGND N_VGND_c_1397_n N_VGND_c_1398_n
+ PM_SKY130_FD_SC_HD__XOR3_1%VGND
cc_1 VNB N_A_112_21#_c_162_n 0.0242681f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_2 VNB N_A_112_21#_c_163_n 0.00258613f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.325
cc_3 VNB N_A_112_21#_c_164_n 0.00130544f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.695
cc_4 VNB N_A_112_21#_c_165_n 0.00246179f $X=-0.19 $Y=-0.24 $X2=1.35 $Y2=0.34
cc_5 VNB N_A_112_21#_c_166_n 0.0346379f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=1.16
cc_6 VNB N_A_112_21#_c_167_n 0.0169571f $X=-0.19 $Y=-0.24 $X2=2.39 $Y2=0.355
cc_7 VNB N_C_c_264_n 0.0196386f $X=-0.19 $Y=-0.24 $X2=2.44 $Y2=0.245
cc_8 VNB N_C_c_265_n 0.0529033f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_9 VNB N_C_c_266_n 0.0215718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_C_c_267_n 0.010199f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.78
cc_11 VNB N_C_c_268_n 0.0112837f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.425
cc_12 VNB N_C_c_269_n 0.00240757f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.695
cc_13 VNB N_A_266_93#_c_332_n 0.00257308f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.96
cc_14 VNB N_A_266_93#_c_333_n 0.00242149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_266_93#_c_334_n 0.0237186f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.78
cc_16 VNB N_A_266_93#_c_335_n 0.0215524f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=1.16
cc_17 VNB N_A_827_297#_M1018_g 0.0355962f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.56
cc_18 VNB N_A_827_297#_c_411_n 0.0259644f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.875
cc_19 VNB N_A_827_297#_M1008_g 0.00127227f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.78
cc_20 VNB N_A_827_297#_c_413_n 0.018065f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.96
cc_21 VNB N_A_827_297#_c_414_n 0.0291429f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=2.045
cc_22 VNB N_A_827_297#_c_415_n 0.0141001f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=2.235
cc_23 VNB N_A_827_297#_c_416_n 0.00221738f $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=0.37
cc_24 VNB N_A_827_297#_c_417_n 0.00809515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_827_297#_c_418_n 0.0124845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_827_297#_c_419_n 5.9975e-19 $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_27 VNB N_A_827_297#_c_420_n 0.00274838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_827_297#_c_421_n 9.00189e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_827_297#_c_422_n 0.00544296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_827_297#_c_423_n 0.00247748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_B_M1000_g 0.00410984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_B_M1012_g 0.0298477f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_33 VNB N_B_c_581_n 0.0515413f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.56
cc_34 VNB N_B_c_582_n 0.0167379f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.325
cc_35 VNB N_B_M1016_g 0.0285283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_B_M1017_g 0.00419891f $X=-0.19 $Y=-0.24 $X2=1.3 $Y2=1.96
cc_37 VNB N_B_c_585_n 0.00493047f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=1.16
cc_38 VNB N_B_c_586_n 7.60368e-19 $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=0.355
cc_39 VNB N_B_c_587_n 0.0267383f $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=0.37
cc_40 VNB N_B_c_588_n 0.0206335f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=1.16
cc_41 VNB N_A_c_701_n 0.0201493f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.985
cc_42 VNB N_A_c_702_n 0.00393727f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.985
cc_43 VNB N_A_c_703_n 0.0173356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_931_365#_c_745_n 0.0193901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_931_365#_c_746_n 0.00630737f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=2.045
cc_46 VNB N_A_931_365#_c_747_n 0.00264442f $X=-0.19 $Y=-0.24 $X2=2.58 $Y2=2.32
cc_47 VNB N_A_931_365#_c_748_n 0.00179065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_931_365#_c_749_n 0.00347802f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.78
cc_49 VNB N_A_931_365#_c_750_n 0.0235243f $X=-0.19 $Y=-0.24 $X2=2.39 $Y2=0.355
cc_50 VNB N_A_931_365#_c_751_n 0.00195542f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_51 VNB N_A_931_365#_c_752_n 0.00471664f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=1.16
cc_52 VNB N_X_c_880_n 0.0311326f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.325
cc_53 VNB N_X_c_881_n 0.0210474f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.78
cc_54 VNB N_VPWR_c_904_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_386_325#_c_999_n 0.00971866f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.695
cc_56 VNB N_A_386_325#_c_1000_n 0.00928634f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.78
cc_57 VNB N_A_404_49#_c_1140_n 0.0026153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_404_49#_c_1141_n 0.00844142f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.96
cc_59 VNB N_A_404_49#_c_1142_n 0.0137061f $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=2.32
cc_60 VNB N_A_404_49#_c_1143_n 0.00301265f $X=-0.19 $Y=-0.24 $X2=2.58 $Y2=2.32
cc_61 VNB N_A_404_49#_c_1144_n 0.00223087f $X=-0.19 $Y=-0.24 $X2=2.39 $Y2=0.355
cc_62 VNB N_A_404_49#_c_1145_n 0.0106987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_404_49#_c_1146_n 3.20957e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1198_49#_c_1321_n 0.00783929f $X=-0.19 $Y=-0.24 $X2=0.865
+ $Y2=1.875
cc_65 VNB N_A_1198_49#_c_1322_n 0.0307334f $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=2.32
cc_66 VNB N_A_1198_49#_c_1323_n 0.0135316f $X=-0.19 $Y=-0.24 $X2=2.39 $Y2=0.355
cc_67 VNB N_VGND_c_1388_n 0.00513547f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.985
cc_68 VNB N_VGND_c_1389_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.78
cc_69 VNB N_VGND_c_1390_n 0.00468014f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.425
cc_70 VNB N_VGND_c_1391_n 0.0223986f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=2.235
cc_71 VNB N_VGND_c_1392_n 0.00478003f $X=-0.19 $Y=-0.24 $X2=2.39 $Y2=0.34
cc_72 VNB N_VGND_c_1393_n 0.0685298f $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=2.32
cc_73 VNB N_VGND_c_1394_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.58 $Y2=2.32
cc_74 VNB N_VGND_c_1395_n 0.0990794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1396_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0.85 $Y2=0.78
cc_76 VNB N_VGND_c_1397_n 0.0189867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1398_n 0.444211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VPB N_A_112_21#_M1002_g 0.0273676f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.985
cc_79 VPB N_A_112_21#_c_163_n 0.00111888f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.325
cc_80 VPB N_A_112_21#_c_170_n 0.00272455f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.875
cc_81 VPB N_A_112_21#_c_171_n 0.00374454f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=2.235
cc_82 VPB N_A_112_21#_c_172_n 0.00112766f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=2.32
cc_83 VPB N_A_112_21#_c_173_n 0.0127396f $X=-0.19 $Y=1.305 $X2=2.58 $Y2=2.32
cc_84 VPB N_A_112_21#_c_166_n 0.00952188f $X=-0.19 $Y=1.305 $X2=0.835 $Y2=1.16
cc_85 VPB N_C_c_270_n 0.0341603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_C_c_265_n 0.0208673f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=0.995
cc_87 VPB N_C_M1004_g 0.0316695f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.985
cc_88 VPB N_C_c_267_n 6.57998e-19 $X=-0.19 $Y=1.305 $X2=1.18 $Y2=0.78
cc_89 VPB N_C_c_268_n 0.00399716f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.425
cc_90 VPB N_C_c_269_n 6.20084e-19 $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.695
cc_91 VPB N_A_266_93#_M1020_g 0.0309169f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=0.56
cc_92 VPB N_A_266_93#_c_332_n 0.00441629f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.96
cc_93 VPB N_A_266_93#_c_338_n 0.0163681f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.695
cc_94 VPB N_A_266_93#_c_339_n 0.00230347f $X=-0.19 $Y=1.305 $X2=2.39 $Y2=0.34
cc_95 VPB N_A_266_93#_c_340_n 0.00173244f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=0.34
cc_96 VPB N_A_266_93#_c_333_n 2.71647e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_266_93#_c_334_n 0.00512541f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=0.78
cc_98 VPB N_A_827_297#_M1015_g 0.0248305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_827_297#_M1008_g 0.0307087f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=0.78
cc_100 VPB N_A_827_297#_c_414_n 0.0105814f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=2.045
cc_101 VPB N_A_827_297#_c_415_n 9.09687e-19 $X=-0.19 $Y=1.305 $X2=1.385
+ $Y2=2.235
cc_102 VPB N_A_827_297#_c_428_n 0.0079496f $X=-0.19 $Y=1.305 $X2=2.58 $Y2=2.32
cc_103 VPB N_A_827_297#_c_423_n 0.00295841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_B_M1000_g 0.0262931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_B_M1017_g 0.0236365f $X=-0.19 $Y=1.305 $X2=1.3 $Y2=1.96
cc_106 VPB N_B_c_591_n 0.110749f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.96
cc_107 VPB N_B_c_592_n 0.0129123f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.425
cc_108 VPB N_B_M1011_g 0.0314866f $X=-0.19 $Y=1.305 $X2=2.58 $Y2=2.32
cc_109 VPB N_B_c_586_n 9.25804e-19 $X=-0.19 $Y=1.305 $X2=2.575 $Y2=0.355
cc_110 VPB N_B_c_587_n 0.00514585f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=0.37
cc_111 VPB N_B_c_596_n 0.00168086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB B 0.00780431f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_113 VPB N_A_M1014_g 0.0197671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_c_701_n 0.00439035f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.985
cc_115 VPB N_A_c_702_n 0.00141167f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.985
cc_116 VPB N_A_931_365#_M1009_g 0.0211416f $X=-0.19 $Y=1.305 $X2=1.3 $Y2=1.96
cc_117 VPB N_A_931_365#_c_746_n 0.00270427f $X=-0.19 $Y=1.305 $X2=1.385
+ $Y2=2.045
cc_118 VPB N_A_931_365#_c_755_n 0.00177722f $X=-0.19 $Y=1.305 $X2=2.39 $Y2=0.34
cc_119 VPB N_A_931_365#_c_749_n 2.70069e-19 $X=-0.19 $Y=1.305 $X2=0.85 $Y2=0.78
cc_120 VPB N_A_931_365#_c_757_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=1.16
cc_121 VPB N_A_931_365#_c_750_n 0.004813f $X=-0.19 $Y=1.305 $X2=2.39 $Y2=0.355
cc_122 VPB N_X_c_882_n 0.014777f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.875
cc_123 VPB N_X_c_881_n 0.00737692f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=0.78
cc_124 VPB X 0.0376478f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=0.78
cc_125 VPB N_VPWR_c_905_n 0.009518f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.985
cc_126 VPB N_VPWR_c_906_n 0.00798922f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=0.78
cc_127 VPB N_VPWR_c_907_n 4.89207e-19 $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.425
cc_128 VPB N_VPWR_c_908_n 0.0219184f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=2.235
cc_129 VPB N_VPWR_c_909_n 0.00640957f $X=-0.19 $Y=1.305 $X2=2.39 $Y2=0.34
cc_130 VPB N_VPWR_c_910_n 0.0626165f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=1.16
cc_131 VPB N_VPWR_c_911_n 0.0887551f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_132 VPB N_VPWR_c_912_n 0.0150434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_904_n 0.0721285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_914_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_915_n 0.00442675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_386_325#_c_1001_n 0.00305158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_386_325#_c_999_n 0.00162217f $X=-0.19 $Y=1.305 $X2=1.265
+ $Y2=0.695
cc_138 VPB N_A_386_325#_c_1003_n 0.00266445f $X=-0.19 $Y=1.305 $X2=1.385
+ $Y2=2.235
cc_139 VPB N_A_386_325#_c_1004_n 6.69494e-19 $X=-0.19 $Y=1.305 $X2=2.58 $Y2=2.32
cc_140 VPB N_A_386_325#_c_1000_n 0.00210227f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=0.78
cc_141 VPB N_A_386_325#_c_1006_n 0.0147473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_386_325#_c_1007_n 0.00318502f $X=-0.19 $Y=1.305 $X2=0.635
+ $Y2=1.16
cc_143 VPB N_A_386_325#_c_1008_n 0.00144605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_386_325#_c_1009_n 0.0214396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_404_49#_c_1147_n 0.00262503f $X=-0.19 $Y=1.305 $X2=1.385
+ $Y2=2.045
cc_146 VPB N_A_404_49#_c_1148_n 0.00579762f $X=-0.19 $Y=1.305 $X2=1.385
+ $Y2=2.235
cc_147 VPB N_A_404_49#_c_1149_n 8.62166e-19 $X=-0.19 $Y=1.305 $X2=2.39 $Y2=0.34
cc_148 VPB N_A_404_49#_c_1143_n 0.00842441f $X=-0.19 $Y=1.305 $X2=2.58 $Y2=2.32
cc_149 VPB N_A_404_49#_c_1151_n 0.00305847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_404_49#_c_1152_n 0.00297262f $X=-0.19 $Y=1.305 $X2=0.835 $Y2=1.16
cc_151 VPB N_A_404_49#_c_1153_n 0.0102984f $X=-0.19 $Y=1.305 $X2=0.835 $Y2=1.16
cc_152 VPB N_A_404_49#_c_1154_n 0.00185607f $X=-0.19 $Y=1.305 $X2=2.575
+ $Y2=0.355
cc_153 VPB N_A_404_49#_c_1144_n 0.00149669f $X=-0.19 $Y=1.305 $X2=2.39 $Y2=0.355
cc_154 VPB N_A_404_49#_c_1156_n 0.0239398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_404_49#_c_1157_n 0.00221054f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_404_49#_c_1158_n 2.86933e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_404_49#_c_1159_n 3.31954e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_1198_49#_c_1321_n 0.00467504f $X=-0.19 $Y=1.305 $X2=0.865
+ $Y2=1.875
cc_159 VPB N_A_1198_49#_c_1325_n 0.0147295f $X=-0.19 $Y=1.305 $X2=1.385
+ $Y2=2.235
cc_160 VPB N_A_1198_49#_c_1322_n 0.0229143f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=2.32
cc_161 VPB N_A_1198_49#_c_1327_n 0.0100871f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=1.16
cc_162 N_A_112_21#_c_162_n N_C_c_264_n 0.0121901f $X=0.635 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A_112_21#_c_163_n N_C_c_264_n 0.00133731f $X=0.865 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_164 N_A_112_21#_c_177_p N_C_c_264_n 0.0121231f $X=1.18 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_165 N_A_112_21#_c_164_n N_C_c_264_n 0.0102997f $X=1.265 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_112_21#_c_165_n N_C_c_264_n 0.00580453f $X=1.35 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_112_21#_M1002_g N_C_c_270_n 0.0204444f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_112_21#_c_170_n N_C_c_270_n 0.00686675f $X=0.865 $Y=1.875 $X2=0 $Y2=0
cc_169 N_A_112_21#_c_182_p N_C_c_270_n 0.0126643f $X=1.3 $Y=1.96 $X2=0 $Y2=0
cc_170 N_A_112_21#_c_171_n N_C_c_270_n 0.00679222f $X=1.385 $Y=2.235 $X2=0 $Y2=0
cc_171 N_A_112_21#_c_172_n N_C_c_270_n 0.00618407f $X=1.47 $Y=2.32 $X2=0 $Y2=0
cc_172 N_A_112_21#_c_167_n N_C_c_265_n 0.00939225f $X=2.39 $Y=0.355 $X2=0 $Y2=0
cc_173 N_A_112_21#_c_173_n N_C_M1004_g 0.0100647f $X=2.58 $Y=2.32 $X2=0 $Y2=0
cc_174 N_A_112_21#_c_187_p N_C_c_266_n 0.00326397f $X=2.575 $Y=0.37 $X2=0 $Y2=0
cc_175 N_A_112_21#_c_167_n N_C_c_266_n 0.00805634f $X=2.39 $Y=0.355 $X2=0 $Y2=0
cc_176 N_A_112_21#_c_163_n N_C_c_267_n 0.00155161f $X=0.865 $Y=1.325 $X2=0 $Y2=0
cc_177 N_A_112_21#_c_166_n N_C_c_267_n 0.0230234f $X=0.835 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_112_21#_c_167_n N_C_c_269_n 0.00331115f $X=2.39 $Y=0.355 $X2=0 $Y2=0
cc_179 N_A_112_21#_c_182_p N_A_266_93#_M1003_d 0.00430647f $X=1.3 $Y=1.96 $X2=0
+ $Y2=0
cc_180 N_A_112_21#_c_171_n N_A_266_93#_M1003_d 0.00261589f $X=1.385 $Y=2.235
+ $X2=0 $Y2=0
cc_181 N_A_112_21#_c_173_n N_A_266_93#_M1020_g 0.00829016f $X=2.58 $Y=2.32 $X2=0
+ $Y2=0
cc_182 N_A_112_21#_c_170_n N_A_266_93#_c_346_n 0.0102753f $X=0.865 $Y=1.875
+ $X2=0 $Y2=0
cc_183 N_A_112_21#_c_177_p N_A_266_93#_c_346_n 0.00345572f $X=1.18 $Y=0.78 $X2=0
+ $Y2=0
cc_184 N_A_112_21#_c_182_p N_A_266_93#_c_346_n 0.0165826f $X=1.3 $Y=1.96 $X2=0
+ $Y2=0
cc_185 N_A_112_21#_c_173_n N_A_266_93#_c_346_n 0.00160427f $X=2.58 $Y=2.32 $X2=0
+ $Y2=0
cc_186 N_A_112_21#_c_163_n N_A_266_93#_c_332_n 0.0125145f $X=0.865 $Y=1.325
+ $X2=0 $Y2=0
cc_187 N_A_112_21#_c_170_n N_A_266_93#_c_332_n 0.00659165f $X=0.865 $Y=1.875
+ $X2=0 $Y2=0
cc_188 N_A_112_21#_c_166_n N_A_266_93#_c_332_n 7.31438e-19 $X=0.835 $Y=1.16
+ $X2=0 $Y2=0
cc_189 N_A_112_21#_c_167_n N_A_266_93#_c_332_n 0.0130244f $X=2.39 $Y=0.355 $X2=0
+ $Y2=0
cc_190 N_A_112_21#_M1004_d N_A_266_93#_c_338_n 0.0030509f $X=2.4 $Y=1.625 $X2=0
+ $Y2=0
cc_191 N_A_112_21#_c_173_n N_A_266_93#_c_338_n 0.00614909f $X=2.58 $Y=2.32 $X2=0
+ $Y2=0
cc_192 N_A_112_21#_c_173_n N_A_266_93#_c_340_n 0.00632099f $X=2.58 $Y=2.32 $X2=0
+ $Y2=0
cc_193 N_A_112_21#_c_187_p N_A_266_93#_c_335_n 0.00171346f $X=2.575 $Y=0.37
+ $X2=0 $Y2=0
cc_194 N_A_112_21#_c_162_n N_X_c_880_n 0.0129344f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_112_21#_c_163_n N_X_c_880_n 0.0173722f $X=0.865 $Y=1.325 $X2=0 $Y2=0
cc_196 N_A_112_21#_c_164_n N_X_c_880_n 0.00448472f $X=1.265 $Y=0.695 $X2=0 $Y2=0
cc_197 N_A_112_21#_M1002_g N_X_c_882_n 0.00505101f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_112_21#_c_170_n N_X_c_882_n 0.0191384f $X=0.865 $Y=1.875 $X2=0 $Y2=0
cc_199 N_A_112_21#_c_166_n N_X_c_882_n 6.92625e-19 $X=0.835 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_112_21#_c_162_n N_X_c_881_n 0.00914182f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_112_21#_M1002_g N_X_c_881_n 0.0014005f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_112_21#_c_163_n N_X_c_881_n 0.0156273f $X=0.865 $Y=1.325 $X2=0 $Y2=0
cc_203 N_A_112_21#_c_170_n N_X_c_881_n 0.00291144f $X=0.865 $Y=1.875 $X2=0 $Y2=0
cc_204 N_A_112_21#_M1002_g X 0.0103319f $X=0.655 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_112_21#_c_170_n N_VPWR_M1002_d 0.00767127f $X=0.865 $Y=1.875
+ $X2=-0.19 $Y2=-0.24
cc_206 N_A_112_21#_c_182_p N_VPWR_M1002_d 0.00842351f $X=1.3 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_207 N_A_112_21#_c_220_p N_VPWR_M1002_d 0.00325153f $X=0.95 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_208 N_A_112_21#_M1002_g N_VPWR_c_905_n 0.00718896f $X=0.655 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_112_21#_c_182_p N_VPWR_c_905_n 0.0126462f $X=1.3 $Y=1.96 $X2=0 $Y2=0
cc_210 N_A_112_21#_c_220_p N_VPWR_c_905_n 0.0138637f $X=0.95 $Y=1.96 $X2=0 $Y2=0
cc_211 N_A_112_21#_c_171_n N_VPWR_c_905_n 0.00138743f $X=1.385 $Y=2.235 $X2=0
+ $Y2=0
cc_212 N_A_112_21#_c_172_n N_VPWR_c_905_n 0.0133932f $X=1.47 $Y=2.32 $X2=0 $Y2=0
cc_213 N_A_112_21#_M1002_g N_VPWR_c_908_n 0.00541359f $X=0.655 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_112_21#_c_182_p N_VPWR_c_910_n 0.00240851f $X=1.3 $Y=1.96 $X2=0 $Y2=0
cc_215 N_A_112_21#_c_172_n N_VPWR_c_910_n 0.00857493f $X=1.47 $Y=2.32 $X2=0
+ $Y2=0
cc_216 N_A_112_21#_c_173_n N_VPWR_c_910_n 0.0619991f $X=2.58 $Y=2.32 $X2=0 $Y2=0
cc_217 N_A_112_21#_M1002_g N_VPWR_c_904_n 0.0120447f $X=0.655 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_112_21#_c_182_p N_VPWR_c_904_n 0.00566226f $X=1.3 $Y=1.96 $X2=0 $Y2=0
cc_219 N_A_112_21#_c_220_p N_VPWR_c_904_n 7.91584e-19 $X=0.95 $Y=1.96 $X2=0
+ $Y2=0
cc_220 N_A_112_21#_c_172_n N_VPWR_c_904_n 0.00627734f $X=1.47 $Y=2.32 $X2=0
+ $Y2=0
cc_221 N_A_112_21#_c_173_n N_VPWR_c_904_n 0.0498596f $X=2.58 $Y=2.32 $X2=0 $Y2=0
cc_222 N_A_112_21#_c_173_n N_A_386_325#_M1004_s 0.00690533f $X=2.58 $Y=2.32
+ $X2=0 $Y2=0
cc_223 N_A_112_21#_M1004_d N_A_386_325#_c_1001_n 0.00585874f $X=2.4 $Y=1.625
+ $X2=0 $Y2=0
cc_224 N_A_112_21#_c_182_p N_A_386_325#_c_1001_n 0.00741315f $X=1.3 $Y=1.96
+ $X2=0 $Y2=0
cc_225 N_A_112_21#_c_171_n N_A_386_325#_c_1001_n 8.38378e-19 $X=1.385 $Y=2.235
+ $X2=0 $Y2=0
cc_226 N_A_112_21#_c_173_n N_A_386_325#_c_1001_n 0.0579338f $X=2.58 $Y=2.32
+ $X2=0 $Y2=0
cc_227 N_A_112_21#_c_167_n N_A_404_49#_M1019_s 0.00521002f $X=2.39 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_228 N_A_112_21#_M1019_d N_A_404_49#_c_1140_n 0.0113061f $X=2.44 $Y=0.245
+ $X2=0 $Y2=0
cc_229 N_A_112_21#_c_187_p N_A_404_49#_c_1140_n 0.017564f $X=2.575 $Y=0.37 $X2=0
+ $Y2=0
cc_230 N_A_112_21#_c_167_n N_A_404_49#_c_1140_n 0.0188825f $X=2.39 $Y=0.355
+ $X2=0 $Y2=0
cc_231 N_A_112_21#_c_187_p N_A_404_49#_c_1164_n 0.00213283f $X=2.575 $Y=0.37
+ $X2=0 $Y2=0
cc_232 N_A_112_21#_c_187_p N_A_404_49#_c_1165_n 0.0147712f $X=2.575 $Y=0.37
+ $X2=0 $Y2=0
cc_233 N_A_112_21#_c_173_n N_A_404_49#_c_1157_n 0.0117643f $X=2.58 $Y=2.32 $X2=0
+ $Y2=0
cc_234 N_A_112_21#_c_163_n N_VGND_M1001_d 0.0049093f $X=0.865 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_235 N_A_112_21#_c_177_p N_VGND_M1001_d 0.00907954f $X=1.18 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_236 N_A_112_21#_c_162_n N_VGND_c_1388_n 0.00766034f $X=0.635 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_112_21#_c_163_n N_VGND_c_1388_n 0.0151684f $X=0.865 $Y=1.325 $X2=0
+ $Y2=0
cc_238 N_A_112_21#_c_177_p N_VGND_c_1388_n 0.00454809f $X=1.18 $Y=0.78 $X2=0
+ $Y2=0
cc_239 N_A_112_21#_c_164_n N_VGND_c_1388_n 0.00720259f $X=1.265 $Y=0.695 $X2=0
+ $Y2=0
cc_240 N_A_112_21#_c_165_n N_VGND_c_1388_n 0.0140929f $X=1.35 $Y=0.34 $X2=0
+ $Y2=0
cc_241 N_A_112_21#_c_166_n N_VGND_c_1388_n 7.93989e-19 $X=0.835 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A_112_21#_c_162_n N_VGND_c_1391_n 0.0054505f $X=0.635 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_112_21#_c_177_p N_VGND_c_1393_n 0.0022086f $X=1.18 $Y=0.78 $X2=0
+ $Y2=0
cc_244 N_A_112_21#_c_165_n N_VGND_c_1393_n 0.0120884f $X=1.35 $Y=0.34 $X2=0
+ $Y2=0
cc_245 N_A_112_21#_c_167_n N_VGND_c_1393_n 0.0854399f $X=2.39 $Y=0.355 $X2=0
+ $Y2=0
cc_246 N_A_112_21#_c_162_n N_VGND_c_1398_n 0.0121255f $X=0.635 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_112_21#_c_163_n N_VGND_c_1398_n 7.71903e-19 $X=0.865 $Y=1.325 $X2=0
+ $Y2=0
cc_248 N_A_112_21#_c_177_p N_VGND_c_1398_n 0.00486519f $X=1.18 $Y=0.78 $X2=0
+ $Y2=0
cc_249 N_A_112_21#_c_165_n N_VGND_c_1398_n 0.00652842f $X=1.35 $Y=0.34 $X2=0
+ $Y2=0
cc_250 N_A_112_21#_c_167_n N_VGND_c_1398_n 0.0511191f $X=2.39 $Y=0.355 $X2=0
+ $Y2=0
cc_251 N_C_M1004_g N_A_266_93#_M1020_g 0.0343211f $X=2.325 $Y=2.045 $X2=0 $Y2=0
cc_252 N_C_c_268_n N_A_266_93#_M1020_g 9.62949e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_253 N_C_c_270_n N_A_266_93#_c_346_n 0.00943923f $X=1.255 $Y=1.325 $X2=0 $Y2=0
cc_254 N_C_c_265_n N_A_266_93#_c_346_n 0.00358164f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_255 N_C_c_264_n N_A_266_93#_c_332_n 0.00475343f $X=1.255 $Y=0.995 $X2=0 $Y2=0
cc_256 N_C_c_270_n N_A_266_93#_c_332_n 0.0038946f $X=1.255 $Y=1.325 $X2=0 $Y2=0
cc_257 N_C_c_265_n N_A_266_93#_c_332_n 0.0235777f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_258 N_C_c_266_n N_A_266_93#_c_332_n 0.00307699f $X=2.365 $Y=0.985 $X2=0 $Y2=0
cc_259 N_C_c_268_n N_A_266_93#_c_332_n 0.00478624f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_260 N_C_c_269_n N_A_266_93#_c_332_n 0.0248423f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_261 N_C_c_265_n N_A_266_93#_c_338_n 0.0126513f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_262 N_C_M1004_g N_A_266_93#_c_338_n 0.0133707f $X=2.325 $Y=2.045 $X2=0 $Y2=0
cc_263 N_C_c_268_n N_A_266_93#_c_338_n 0.00117647f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_264 N_C_c_269_n N_A_266_93#_c_338_n 0.0403344f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_265 N_C_M1004_g N_A_266_93#_c_339_n 0.00345696f $X=2.325 $Y=2.045 $X2=0 $Y2=0
cc_266 N_C_c_268_n N_A_266_93#_c_339_n 6.06227e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_267 N_C_c_268_n N_A_266_93#_c_333_n 9.73749e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_268 N_C_c_269_n N_A_266_93#_c_333_n 0.0286115f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_269 N_C_c_268_n N_A_266_93#_c_334_n 0.0153962f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_270 N_C_c_269_n N_A_266_93#_c_334_n 0.00111895f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_271 N_C_c_266_n N_A_266_93#_c_335_n 0.0223998f $X=2.365 $Y=0.985 $X2=0 $Y2=0
cc_272 N_C_c_268_n N_A_266_93#_c_335_n 3.54366e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_273 N_C_c_264_n N_X_c_880_n 6.48733e-19 $X=1.255 $Y=0.995 $X2=0 $Y2=0
cc_274 N_C_c_270_n X 9.14332e-19 $X=1.255 $Y=1.325 $X2=0 $Y2=0
cc_275 N_C_c_270_n N_VPWR_c_905_n 0.00211197f $X=1.255 $Y=1.325 $X2=0 $Y2=0
cc_276 N_C_c_270_n N_VPWR_c_910_n 0.00403219f $X=1.255 $Y=1.325 $X2=0 $Y2=0
cc_277 N_C_M1004_g N_VPWR_c_910_n 0.00356303f $X=2.325 $Y=2.045 $X2=0 $Y2=0
cc_278 N_C_c_270_n N_VPWR_c_904_n 0.00522107f $X=1.255 $Y=1.325 $X2=0 $Y2=0
cc_279 N_C_M1004_g N_VPWR_c_904_n 0.00649631f $X=2.325 $Y=2.045 $X2=0 $Y2=0
cc_280 N_C_c_270_n N_A_386_325#_c_1001_n 9.44709e-19 $X=1.255 $Y=1.325 $X2=0
+ $Y2=0
cc_281 N_C_M1004_g N_A_386_325#_c_1001_n 0.00901837f $X=2.325 $Y=2.045 $X2=0
+ $Y2=0
cc_282 N_C_c_265_n N_A_404_49#_c_1140_n 0.00531432f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_283 N_C_c_266_n N_A_404_49#_c_1140_n 0.00927259f $X=2.365 $Y=0.985 $X2=0
+ $Y2=0
cc_284 N_C_c_269_n N_A_404_49#_c_1140_n 0.0345339f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_285 N_C_c_266_n N_A_404_49#_c_1164_n 7.28465e-19 $X=2.365 $Y=0.985 $X2=0
+ $Y2=0
cc_286 N_C_c_264_n N_VGND_c_1388_n 0.00111462f $X=1.255 $Y=0.995 $X2=0 $Y2=0
cc_287 N_C_c_264_n N_VGND_c_1393_n 7.72982e-19 $X=1.255 $Y=0.995 $X2=0 $Y2=0
cc_288 N_C_c_266_n N_VGND_c_1393_n 0.00357877f $X=2.365 $Y=0.985 $X2=0 $Y2=0
cc_289 N_C_c_266_n N_VGND_c_1398_n 0.00696677f $X=2.365 $Y=0.985 $X2=0 $Y2=0
cc_290 N_A_266_93#_M1020_g N_VPWR_c_910_n 0.00369158f $X=2.855 $Y=2.045 $X2=0
+ $Y2=0
cc_291 N_A_266_93#_M1020_g N_VPWR_c_904_n 0.00664398f $X=2.855 $Y=2.045 $X2=0
+ $Y2=0
cc_292 N_A_266_93#_c_338_n N_A_386_325#_M1004_s 0.00354978f $X=2.665 $Y=1.62
+ $X2=0 $Y2=0
cc_293 N_A_266_93#_M1020_g N_A_386_325#_c_1001_n 0.0137617f $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_294 N_A_266_93#_c_338_n N_A_386_325#_c_1001_n 0.0526775f $X=2.665 $Y=1.62
+ $X2=0 $Y2=0
cc_295 N_A_266_93#_c_333_n N_A_386_325#_c_1001_n 0.00267573f $X=2.855 $Y=1.16
+ $X2=0 $Y2=0
cc_296 N_A_266_93#_c_334_n N_A_386_325#_c_1001_n 0.00111532f $X=2.855 $Y=1.16
+ $X2=0 $Y2=0
cc_297 N_A_266_93#_M1020_g N_A_386_325#_c_1022_n 0.00740594f $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_298 N_A_266_93#_c_338_n N_A_386_325#_c_1022_n 7.49507e-19 $X=2.665 $Y=1.62
+ $X2=0 $Y2=0
cc_299 N_A_266_93#_M1020_g N_A_386_325#_c_999_n 8.85667e-19 $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_300 N_A_266_93#_c_339_n N_A_386_325#_c_999_n 0.00180217f $X=2.75 $Y=1.535
+ $X2=0 $Y2=0
cc_301 N_A_266_93#_c_333_n N_A_386_325#_c_999_n 0.0155817f $X=2.855 $Y=1.16
+ $X2=0 $Y2=0
cc_302 N_A_266_93#_c_335_n N_A_386_325#_c_999_n 0.0134409f $X=2.855 $Y=0.995
+ $X2=0 $Y2=0
cc_303 N_A_266_93#_c_338_n N_A_386_325#_c_1007_n 4.43984e-19 $X=2.665 $Y=1.62
+ $X2=0 $Y2=0
cc_304 N_A_266_93#_c_339_n N_A_386_325#_c_1007_n 6.14306e-19 $X=2.75 $Y=1.535
+ $X2=0 $Y2=0
cc_305 N_A_266_93#_M1020_g N_A_386_325#_c_1009_n 0.00655666f $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_306 N_A_266_93#_c_338_n N_A_386_325#_c_1009_n 0.0135143f $X=2.665 $Y=1.62
+ $X2=0 $Y2=0
cc_307 N_A_266_93#_c_339_n N_A_386_325#_c_1009_n 0.00587493f $X=2.75 $Y=1.535
+ $X2=0 $Y2=0
cc_308 N_A_266_93#_c_332_n N_A_404_49#_c_1140_n 0.00977028f $X=1.605 $Y=0.76
+ $X2=0 $Y2=0
cc_309 N_A_266_93#_c_333_n N_A_404_49#_c_1140_n 0.0184041f $X=2.855 $Y=1.16
+ $X2=0 $Y2=0
cc_310 N_A_266_93#_c_334_n N_A_404_49#_c_1140_n 0.00280181f $X=2.855 $Y=1.16
+ $X2=0 $Y2=0
cc_311 N_A_266_93#_c_335_n N_A_404_49#_c_1140_n 0.0130512f $X=2.855 $Y=0.995
+ $X2=0 $Y2=0
cc_312 N_A_266_93#_c_335_n N_A_404_49#_c_1164_n 0.00862425f $X=2.855 $Y=0.995
+ $X2=0 $Y2=0
cc_313 N_A_266_93#_c_335_n N_A_404_49#_c_1165_n 0.00716742f $X=2.855 $Y=0.995
+ $X2=0 $Y2=0
cc_314 N_A_266_93#_M1020_g N_A_404_49#_c_1147_n 0.00447876f $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_315 N_A_266_93#_M1020_g N_A_404_49#_c_1149_n 7.78208e-19 $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_316 N_A_266_93#_c_335_n N_A_404_49#_c_1142_n 0.00103799f $X=2.855 $Y=0.995
+ $X2=0 $Y2=0
cc_317 N_A_266_93#_M1020_g N_A_404_49#_c_1157_n 0.00335543f $X=2.855 $Y=2.045
+ $X2=0 $Y2=0
cc_318 N_A_266_93#_c_335_n N_VGND_c_1393_n 0.00390499f $X=2.855 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_A_266_93#_c_335_n N_VGND_c_1398_n 0.00727536f $X=2.855 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_827_297#_c_428_n N_B_M1000_g 0.00527417f $X=4.4 $Y=1.58 $X2=0 $Y2=0
cc_321 N_A_827_297#_c_423_n N_B_M1000_g 0.00476142f $X=4.435 $Y=0.72 $X2=0 $Y2=0
cc_322 N_A_827_297#_c_432_p N_B_M1012_g 0.00360359f $X=4.515 $Y=0.85 $X2=0 $Y2=0
cc_323 N_A_827_297#_c_423_n N_B_M1012_g 0.0137047f $X=4.435 $Y=0.72 $X2=0 $Y2=0
cc_324 N_A_827_297#_c_417_n N_B_c_581_n 0.00436054f $X=5.605 $Y=0.85 $X2=0 $Y2=0
cc_325 N_A_827_297#_c_423_n N_B_c_581_n 0.0122014f $X=4.435 $Y=0.72 $X2=0 $Y2=0
cc_326 N_A_827_297#_c_428_n N_B_c_582_n 0.00335249f $X=4.4 $Y=1.58 $X2=0 $Y2=0
cc_327 N_A_827_297#_c_423_n N_B_c_582_n 0.00329164f $X=4.435 $Y=0.72 $X2=0 $Y2=0
cc_328 N_A_827_297#_M1018_g N_B_M1016_g 0.0114571f $X=5.915 $Y=0.455 $X2=0 $Y2=0
cc_329 N_A_827_297#_c_414_n N_B_M1016_g 0.0210118f $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_827_297#_c_416_n N_B_M1016_g 0.00170749f $X=5.727 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_827_297#_c_417_n N_B_M1016_g 7.57846e-19 $X=5.605 $Y=0.85 $X2=0 $Y2=0
cc_332 N_A_827_297#_c_419_n N_B_M1016_g 6.64234e-19 $X=5.895 $Y=0.85 $X2=0 $Y2=0
cc_333 N_A_827_297#_c_420_n N_B_M1016_g 0.00117063f $X=5.75 $Y=0.85 $X2=0 $Y2=0
cc_334 N_A_827_297#_M1015_g N_B_M1017_g 0.0137639f $X=5.915 $Y=1.805 $X2=0 $Y2=0
cc_335 N_A_827_297#_M1015_g N_B_c_591_n 0.00881703f $X=5.915 $Y=1.805 $X2=0
+ $Y2=0
cc_336 N_A_827_297#_M1008_g N_B_M1011_g 0.0403239f $X=7.305 $Y=2.065 $X2=0 $Y2=0
cc_337 N_A_827_297#_c_411_n N_B_c_586_n 0.00114568f $X=7.305 $Y=1.28 $X2=0 $Y2=0
cc_338 N_A_827_297#_c_418_n N_B_c_586_n 0.00555012f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_339 N_A_827_297#_c_422_n N_B_c_586_n 0.0211354f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_340 N_A_827_297#_c_411_n N_B_c_587_n 0.0189136f $X=7.305 $Y=1.28 $X2=0 $Y2=0
cc_341 N_A_827_297#_c_415_n N_B_c_587_n 0.00771356f $X=5.915 $Y=1.16 $X2=0 $Y2=0
cc_342 N_A_827_297#_c_418_n N_B_c_587_n 0.00134545f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_343 N_A_827_297#_c_422_n N_B_c_587_n 0.00169113f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_344 N_A_827_297#_c_411_n B 8.1069e-19 $X=7.305 $Y=1.28 $X2=0 $Y2=0
cc_345 N_A_827_297#_M1008_g B 0.00593518f $X=7.305 $Y=2.065 $X2=0 $Y2=0
cc_346 N_A_827_297#_c_418_n B 0.00414594f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_347 N_A_827_297#_c_421_n B 0.00235209f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_348 N_A_827_297#_c_422_n B 0.0183366f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_349 N_A_827_297#_M1018_g N_B_c_588_n 0.00771356f $X=5.915 $Y=0.455 $X2=0
+ $Y2=0
cc_350 N_A_827_297#_c_411_n N_B_c_588_n 0.00163786f $X=7.305 $Y=1.28 $X2=0 $Y2=0
cc_351 N_A_827_297#_c_413_n N_B_c_588_n 0.0180222f $X=7.31 $Y=0.945 $X2=0 $Y2=0
cc_352 N_A_827_297#_c_418_n N_B_c_588_n 0.00749482f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_353 N_A_827_297#_c_421_n N_B_c_588_n 0.00142159f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_354 N_A_827_297#_c_422_n N_B_c_588_n 0.00206701f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_355 N_A_827_297#_M1008_g N_A_M1014_g 0.0404776f $X=7.305 $Y=2.065 $X2=0 $Y2=0
cc_356 N_A_827_297#_c_411_n N_A_c_701_n 0.0176934f $X=7.305 $Y=1.28 $X2=0 $Y2=0
cc_357 N_A_827_297#_M1008_g N_A_c_701_n 0.00255062f $X=7.305 $Y=2.065 $X2=0
+ $Y2=0
cc_358 N_A_827_297#_c_422_n N_A_c_701_n 7.00021e-19 $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_359 N_A_827_297#_c_411_n N_A_c_702_n 0.00129629f $X=7.305 $Y=1.28 $X2=0 $Y2=0
cc_360 N_A_827_297#_M1008_g N_A_c_702_n 5.31842e-19 $X=7.305 $Y=2.065 $X2=0
+ $Y2=0
cc_361 N_A_827_297#_c_422_n N_A_c_702_n 0.016109f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_362 N_A_827_297#_c_413_n N_A_c_703_n 0.0225442f $X=7.31 $Y=0.945 $X2=0 $Y2=0
cc_363 N_A_827_297#_c_422_n N_A_c_703_n 2.68453e-19 $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_364 N_A_827_297#_c_417_n N_A_931_365#_M1016_s 8.44656e-19 $X=5.605 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_365 N_A_827_297#_c_428_n N_A_931_365#_c_746_n 0.019709f $X=4.4 $Y=1.58 $X2=0
+ $Y2=0
cc_366 N_A_827_297#_c_417_n N_A_931_365#_c_746_n 0.0123662f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_367 N_A_827_297#_c_432_p N_A_931_365#_c_746_n 6.70277e-19 $X=4.515 $Y=0.85
+ $X2=0 $Y2=0
cc_368 N_A_827_297#_c_423_n N_A_931_365#_c_746_n 0.0609172f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_369 N_A_827_297#_M1008_g N_A_931_365#_c_755_n 0.00235326f $X=7.305 $Y=2.065
+ $X2=0 $Y2=0
cc_370 N_A_827_297#_c_413_n N_A_931_365#_c_748_n 0.00164439f $X=7.31 $Y=0.945
+ $X2=0 $Y2=0
cc_371 N_A_827_297#_c_421_n N_A_931_365#_c_748_n 0.00485657f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_372 N_A_827_297#_c_422_n N_A_931_365#_c_748_n 0.00616889f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_373 N_A_827_297#_M1018_g N_A_931_365#_c_768_n 0.00602851f $X=5.915 $Y=0.455
+ $X2=0 $Y2=0
cc_374 N_A_827_297#_c_413_n N_A_931_365#_c_768_n 0.00716191f $X=7.31 $Y=0.945
+ $X2=0 $Y2=0
cc_375 N_A_827_297#_c_416_n N_A_931_365#_c_768_n 3.7129e-19 $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_376 N_A_827_297#_c_417_n N_A_931_365#_c_768_n 0.0490112f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_377 N_A_827_297#_c_418_n N_A_931_365#_c_768_n 0.0873524f $X=6.985 $Y=0.85
+ $X2=0 $Y2=0
cc_378 N_A_827_297#_c_419_n N_A_931_365#_c_768_n 0.0265257f $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_379 N_A_827_297#_c_420_n N_A_931_365#_c_768_n 0.00319269f $X=5.75 $Y=0.85
+ $X2=0 $Y2=0
cc_380 N_A_827_297#_c_421_n N_A_931_365#_c_768_n 0.0265508f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_381 N_A_827_297#_c_422_n N_A_931_365#_c_768_n 0.00472786f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_382 N_A_827_297#_c_417_n N_A_931_365#_c_751_n 0.0261136f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_383 N_A_827_297#_c_423_n N_A_931_365#_c_751_n 0.00675389f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_384 N_A_827_297#_c_417_n N_A_931_365#_c_752_n 0.00112331f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_385 N_A_827_297#_c_423_n N_A_931_365#_c_752_n 0.0117267f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_386 N_A_827_297#_c_413_n N_A_931_365#_c_781_n 0.00153367f $X=7.31 $Y=0.945
+ $X2=0 $Y2=0
cc_387 N_A_827_297#_c_413_n N_A_931_365#_c_782_n 0.0077529f $X=7.31 $Y=0.945
+ $X2=0 $Y2=0
cc_388 N_A_827_297#_M1008_g N_VPWR_c_907_n 0.00128985f $X=7.305 $Y=2.065 $X2=0
+ $Y2=0
cc_389 N_A_827_297#_M1008_g N_VPWR_c_911_n 0.00362032f $X=7.305 $Y=2.065 $X2=0
+ $Y2=0
cc_390 N_A_827_297#_M1000_d N_VPWR_c_904_n 0.00286702f $X=4.135 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_A_827_297#_M1008_g N_VPWR_c_904_n 0.00570414f $X=7.305 $Y=2.065 $X2=0
+ $Y2=0
cc_392 N_A_827_297#_c_418_n N_A_386_325#_M1021_d 0.00109392f $X=6.985 $Y=0.85
+ $X2=0 $Y2=0
cc_393 N_A_827_297#_c_421_n N_A_386_325#_M1021_d 7.4435e-19 $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_394 N_A_827_297#_c_422_n N_A_386_325#_M1021_d 0.00406077f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_395 N_A_827_297#_c_414_n N_A_386_325#_c_1003_n 0.00894291f $X=5.84 $Y=1.16
+ $X2=0 $Y2=0
cc_396 N_A_827_297#_c_416_n N_A_386_325#_c_1003_n 0.0270839f $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_397 N_A_827_297#_c_417_n N_A_386_325#_c_1003_n 5.63647e-19 $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_398 N_A_827_297#_M1015_g N_A_386_325#_c_1039_n 0.00368795f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_399 N_A_827_297#_M1015_g N_A_386_325#_c_1004_n 0.01555f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_400 N_A_827_297#_c_414_n N_A_386_325#_c_1004_n 7.42472e-19 $X=5.84 $Y=1.16
+ $X2=0 $Y2=0
cc_401 N_A_827_297#_c_416_n N_A_386_325#_c_1004_n 0.00152864f $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_402 N_A_827_297#_c_418_n N_A_386_325#_c_1004_n 0.00288457f $X=6.985 $Y=0.85
+ $X2=0 $Y2=0
cc_403 N_A_827_297#_c_419_n N_A_386_325#_c_1004_n 6.69145e-19 $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_827_297#_M1018_g N_A_386_325#_c_1000_n 0.0170984f $X=5.915 $Y=0.455
+ $X2=0 $Y2=0
cc_405 N_A_827_297#_c_416_n N_A_386_325#_c_1000_n 0.0210201f $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_406 N_A_827_297#_c_418_n N_A_386_325#_c_1000_n 0.0170211f $X=6.985 $Y=0.85
+ $X2=0 $Y2=0
cc_407 N_A_827_297#_c_419_n N_A_386_325#_c_1000_n 0.00240264f $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_408 N_A_827_297#_c_420_n N_A_386_325#_c_1000_n 0.0233729f $X=5.75 $Y=0.85
+ $X2=0 $Y2=0
cc_409 N_A_827_297#_c_413_n N_A_386_325#_c_1050_n 0.00328526f $X=7.31 $Y=0.945
+ $X2=0 $Y2=0
cc_410 N_A_827_297#_c_418_n N_A_386_325#_c_1050_n 0.00149151f $X=6.985 $Y=0.85
+ $X2=0 $Y2=0
cc_411 N_A_827_297#_c_421_n N_A_386_325#_c_1050_n 3.55136e-19 $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_412 N_A_827_297#_c_422_n N_A_386_325#_c_1050_n 0.00528249f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_413 N_A_827_297#_c_428_n N_A_386_325#_c_1006_n 0.0236641f $X=4.4 $Y=1.58
+ $X2=0 $Y2=0
cc_414 N_A_827_297#_c_416_n N_A_386_325#_c_1006_n 8.37577e-19 $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_415 N_A_827_297#_c_417_n N_A_386_325#_c_1006_n 0.0483476f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_416 N_A_827_297#_c_432_p N_A_386_325#_c_1006_n 0.0124517f $X=4.515 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_827_297#_c_423_n N_A_386_325#_c_1006_n 0.00191432f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_418 N_A_827_297#_M1015_g N_A_386_325#_c_1008_n 0.00414596f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_419 N_A_827_297#_c_414_n N_A_386_325#_c_1008_n 0.00431105f $X=5.84 $Y=1.16
+ $X2=0 $Y2=0
cc_420 N_A_827_297#_c_416_n N_A_386_325#_c_1008_n 0.00243787f $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_421 N_A_827_297#_c_419_n N_A_386_325#_c_1008_n 0.0153495f $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_422 N_A_827_297#_c_417_n N_A_404_49#_M1016_d 0.00139415f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_423 N_A_827_297#_c_419_n N_A_404_49#_M1016_d 5.07779e-19 $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_424 N_A_827_297#_c_420_n N_A_404_49#_M1016_d 0.00574398f $X=5.75 $Y=0.85
+ $X2=0 $Y2=0
cc_425 N_A_827_297#_c_432_p N_A_404_49#_c_1142_n 0.00244026f $X=4.515 $Y=0.85
+ $X2=0 $Y2=0
cc_426 N_A_827_297#_c_423_n N_A_404_49#_c_1142_n 0.00391248f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_427 N_A_827_297#_c_428_n N_A_404_49#_c_1143_n 0.0142825f $X=4.4 $Y=1.58 $X2=0
+ $Y2=0
cc_428 N_A_827_297#_c_423_n N_A_404_49#_c_1143_n 0.0100198f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_429 N_A_827_297#_M1000_d N_A_404_49#_c_1151_n 0.00530614f $X=4.135 $Y=1.485
+ $X2=0 $Y2=0
cc_430 N_A_827_297#_c_428_n N_A_404_49#_c_1151_n 0.0250069f $X=4.4 $Y=1.58 $X2=0
+ $Y2=0
cc_431 N_A_827_297#_M1000_d N_A_404_49#_c_1152_n 0.00285479f $X=4.135 $Y=1.485
+ $X2=0 $Y2=0
cc_432 N_A_827_297#_M1000_d N_A_404_49#_c_1154_n 0.00268234f $X=4.135 $Y=1.485
+ $X2=0 $Y2=0
cc_433 N_A_827_297#_M1015_g N_A_404_49#_c_1144_n 0.00176903f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_434 N_A_827_297#_c_414_n N_A_404_49#_c_1144_n 7.08656e-19 $X=5.84 $Y=1.16
+ $X2=0 $Y2=0
cc_435 N_A_827_297#_c_416_n N_A_404_49#_c_1144_n 0.0183299f $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_436 N_A_827_297#_c_417_n N_A_404_49#_c_1144_n 0.00613141f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_437 N_A_827_297#_c_419_n N_A_404_49#_c_1144_n 0.00108234f $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_438 N_A_827_297#_c_420_n N_A_404_49#_c_1144_n 0.00295805f $X=5.75 $Y=0.85
+ $X2=0 $Y2=0
cc_439 N_A_827_297#_M1015_g N_A_404_49#_c_1156_n 0.00215111f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_440 N_A_827_297#_M1008_g N_A_404_49#_c_1156_n 0.00693683f $X=7.305 $Y=2.065
+ $X2=0 $Y2=0
cc_441 N_A_827_297#_M1018_g N_A_404_49#_c_1200_n 0.00229256f $X=5.915 $Y=0.455
+ $X2=0 $Y2=0
cc_442 N_A_827_297#_c_420_n N_A_404_49#_c_1200_n 0.00181204f $X=5.75 $Y=0.85
+ $X2=0 $Y2=0
cc_443 N_A_827_297#_c_423_n N_A_404_49#_c_1145_n 0.00671983f $X=4.435 $Y=0.72
+ $X2=0 $Y2=0
cc_444 N_A_827_297#_c_414_n N_A_404_49#_c_1146_n 2.22283e-19 $X=5.84 $Y=1.16
+ $X2=0 $Y2=0
cc_445 N_A_827_297#_c_416_n N_A_404_49#_c_1146_n 0.00265833f $X=5.727 $Y=0.995
+ $X2=0 $Y2=0
cc_446 N_A_827_297#_c_417_n N_A_404_49#_c_1146_n 0.0156216f $X=5.605 $Y=0.85
+ $X2=0 $Y2=0
cc_447 N_A_827_297#_c_419_n N_A_404_49#_c_1146_n 0.00133614f $X=5.895 $Y=0.85
+ $X2=0 $Y2=0
cc_448 N_A_827_297#_c_420_n N_A_404_49#_c_1146_n 0.0141097f $X=5.75 $Y=0.85
+ $X2=0 $Y2=0
cc_449 N_A_827_297#_c_418_n N_A_1198_49#_M1018_d 0.00166227f $X=6.985 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_450 N_A_827_297#_M1015_g N_A_1198_49#_c_1321_n 0.00785518f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_451 N_A_827_297#_c_418_n N_A_1198_49#_c_1321_n 0.0179438f $X=6.985 $Y=0.85
+ $X2=0 $Y2=0
cc_452 N_A_827_297#_c_421_n N_A_1198_49#_c_1321_n 0.00214961f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_453 N_A_827_297#_c_422_n N_A_1198_49#_c_1321_n 0.00583126f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_454 N_A_827_297#_M1015_g N_A_1198_49#_c_1333_n 0.00421122f $X=5.915 $Y=1.805
+ $X2=0 $Y2=0
cc_455 N_A_827_297#_M1008_g N_A_1198_49#_c_1334_n 0.0138456f $X=7.305 $Y=2.065
+ $X2=0 $Y2=0
cc_456 N_A_827_297#_c_422_n N_A_1198_49#_c_1334_n 0.00161448f $X=7.13 $Y=0.85
+ $X2=0 $Y2=0
cc_457 N_A_827_297#_c_432_p N_VGND_c_1389_n 0.0038248f $X=4.515 $Y=0.85 $X2=0
+ $Y2=0
cc_458 N_A_827_297#_M1018_g N_VGND_c_1395_n 0.00575161f $X=5.915 $Y=0.455 $X2=0
+ $Y2=0
cc_459 N_A_827_297#_c_413_n N_VGND_c_1395_n 0.00585385f $X=7.31 $Y=0.945 $X2=0
+ $Y2=0
cc_460 N_A_827_297#_c_420_n N_VGND_c_1395_n 0.00316593f $X=5.75 $Y=0.85 $X2=0
+ $Y2=0
cc_461 N_A_827_297#_c_422_n N_VGND_c_1395_n 7.70543e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_462 N_A_827_297#_c_423_n N_VGND_c_1395_n 0.0072215f $X=4.435 $Y=0.72 $X2=0
+ $Y2=0
cc_463 N_A_827_297#_M1012_d N_VGND_c_1398_n 0.00194539f $X=4.3 $Y=0.235 $X2=0
+ $Y2=0
cc_464 N_A_827_297#_M1018_g N_VGND_c_1398_n 0.00663327f $X=5.915 $Y=0.455 $X2=0
+ $Y2=0
cc_465 N_A_827_297#_c_413_n N_VGND_c_1398_n 0.00607914f $X=7.31 $Y=0.945 $X2=0
+ $Y2=0
cc_466 N_A_827_297#_c_417_n N_VGND_c_1398_n 0.00899211f $X=5.605 $Y=0.85 $X2=0
+ $Y2=0
cc_467 N_A_827_297#_c_432_p N_VGND_c_1398_n 0.0148507f $X=4.515 $Y=0.85 $X2=0
+ $Y2=0
cc_468 N_A_827_297#_c_423_n N_VGND_c_1398_n 0.00376241f $X=4.435 $Y=0.72 $X2=0
+ $Y2=0
cc_469 B N_A_M1014_g 2.12214e-19 $X=7.045 $Y=1.445 $X2=0 $Y2=0
cc_470 N_B_c_586_n N_A_c_702_n 0.00135728f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_471 N_B_M1000_g N_A_931_365#_c_746_n 0.00405425f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_472 N_B_M1012_g N_A_931_365#_c_746_n 0.00120086f $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_473 N_B_c_581_n N_A_931_365#_c_746_n 0.014531f $X=5.08 $Y=1.16 $X2=0 $Y2=0
cc_474 N_B_M1016_g N_A_931_365#_c_746_n 0.00465425f $X=5.155 $Y=0.565 $X2=0
+ $Y2=0
cc_475 N_B_M1017_g N_A_931_365#_c_746_n 0.00542523f $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_476 B N_A_931_365#_c_755_n 0.0103993f $X=7.045 $Y=1.445 $X2=0 $Y2=0
cc_477 N_B_M1016_g N_A_931_365#_c_768_n 0.00165623f $X=5.155 $Y=0.565 $X2=0
+ $Y2=0
cc_478 N_B_c_588_n N_A_931_365#_c_768_n 0.00325031f $X=6.77 $Y=0.995 $X2=0 $Y2=0
cc_479 N_B_M1012_g N_A_931_365#_c_751_n 4.1997e-19 $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_480 N_B_M1016_g N_A_931_365#_c_751_n 9.47409e-19 $X=5.155 $Y=0.565 $X2=0
+ $Y2=0
cc_481 N_B_M1012_g N_A_931_365#_c_752_n 0.00326325f $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_482 N_B_c_581_n N_A_931_365#_c_752_n 0.00234074f $X=5.08 $Y=1.16 $X2=0 $Y2=0
cc_483 N_B_M1016_g N_A_931_365#_c_752_n 0.00457137f $X=5.155 $Y=0.565 $X2=0
+ $Y2=0
cc_484 N_B_M1000_g N_VPWR_c_906_n 0.0112156f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_485 N_B_M1000_g N_VPWR_c_911_n 0.00341689f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_486 N_B_c_592_n N_VPWR_c_911_n 0.038174f $X=5.23 $Y=2.54 $X2=0 $Y2=0
cc_487 N_B_M1000_g N_VPWR_c_904_n 0.00540327f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_488 N_B_c_591_n N_VPWR_c_904_n 0.0391964f $X=6.715 $Y=2.54 $X2=0 $Y2=0
cc_489 N_B_c_592_n N_VPWR_c_904_n 0.00592495f $X=5.23 $Y=2.54 $X2=0 $Y2=0
cc_490 N_B_c_582_n N_A_386_325#_c_999_n 4.45781e-19 $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_491 N_B_M1017_g N_A_386_325#_c_1003_n 0.00135024f $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_492 N_B_M1017_g N_A_386_325#_c_1039_n 0.00408716f $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_493 N_B_c_588_n N_A_386_325#_c_1000_n 0.0026019f $X=6.77 $Y=0.995 $X2=0 $Y2=0
cc_494 N_B_c_586_n N_A_386_325#_c_1050_n 0.00216976f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_495 N_B_c_587_n N_A_386_325#_c_1050_n 0.00134398f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_496 N_B_c_588_n N_A_386_325#_c_1050_n 0.00498906f $X=6.77 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_B_c_588_n N_A_386_325#_c_1070_n 0.00521263f $X=6.77 $Y=0.995 $X2=0
+ $Y2=0
cc_498 N_B_M1000_g N_A_386_325#_c_1006_n 0.00514339f $X=4.06 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_B_c_581_n N_A_386_325#_c_1006_n 0.0041572f $X=5.08 $Y=1.16 $X2=0 $Y2=0
cc_500 N_B_M1017_g N_A_386_325#_c_1006_n 0.00291393f $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_501 N_B_M1017_g N_A_386_325#_c_1008_n 4.42823e-19 $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_502 N_B_M1000_g N_A_404_49#_c_1147_n 0.00287704f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_503 N_B_M1012_g N_A_404_49#_c_1142_n 0.00331221f $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_504 N_B_c_582_n N_A_404_49#_c_1143_n 0.0176462f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_505 N_B_M1000_g N_A_404_49#_c_1151_n 0.0156612f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_506 N_B_M1000_g N_A_404_49#_c_1152_n 0.00631689f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_507 N_B_M1017_g N_A_404_49#_c_1152_n 9.06836e-19 $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_508 N_B_M1000_g N_A_404_49#_c_1154_n 0.00361658f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_509 N_B_c_581_n N_A_404_49#_c_1144_n 0.00266058f $X=5.08 $Y=1.16 $X2=0 $Y2=0
cc_510 N_B_M1016_g N_A_404_49#_c_1144_n 0.00664131f $X=5.155 $Y=0.565 $X2=0
+ $Y2=0
cc_511 N_B_M1017_g N_A_404_49#_c_1144_n 0.0375467f $X=5.155 $Y=1.905 $X2=0 $Y2=0
cc_512 N_B_c_585_n N_A_404_49#_c_1144_n 0.0026181f $X=5.155 $Y=1.16 $X2=0 $Y2=0
cc_513 N_B_M1017_g N_A_404_49#_c_1156_n 0.00571676f $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_514 N_B_c_591_n N_A_404_49#_c_1156_n 0.0278445f $X=6.715 $Y=2.54 $X2=0 $Y2=0
cc_515 N_B_M1011_g N_A_404_49#_c_1156_n 0.0122992f $X=6.79 $Y=1.965 $X2=0 $Y2=0
cc_516 N_B_M1016_g N_A_404_49#_c_1200_n 5.18677e-19 $X=5.155 $Y=0.565 $X2=0
+ $Y2=0
cc_517 N_B_M1012_g N_A_404_49#_c_1145_n 9.41344e-19 $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_518 N_B_c_582_n N_A_404_49#_c_1145_n 0.00378888f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_519 N_B_M1016_g N_A_404_49#_c_1146_n 0.0115325f $X=5.155 $Y=0.565 $X2=0 $Y2=0
cc_520 N_B_M1017_g N_A_404_49#_c_1159_n 0.00727105f $X=5.155 $Y=1.905 $X2=0
+ $Y2=0
cc_521 N_B_M1011_g N_A_1198_49#_c_1321_n 0.0107026f $X=6.79 $Y=1.965 $X2=0 $Y2=0
cc_522 N_B_c_586_n N_A_1198_49#_c_1321_n 0.0325983f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_523 N_B_c_596_n N_A_1198_49#_c_1321_n 0.0141708f $X=6.855 $Y=1.53 $X2=0 $Y2=0
cc_524 N_B_c_588_n N_A_1198_49#_c_1321_n 0.0103225f $X=6.77 $Y=0.995 $X2=0 $Y2=0
cc_525 N_B_M1011_g N_A_1198_49#_c_1334_n 0.0096343f $X=6.79 $Y=1.965 $X2=0 $Y2=0
cc_526 N_B_c_587_n N_A_1198_49#_c_1334_n 0.00103367f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_527 N_B_c_596_n N_A_1198_49#_c_1334_n 0.00720786f $X=6.855 $Y=1.53 $X2=0
+ $Y2=0
cc_528 B N_A_1198_49#_c_1334_n 0.0164129f $X=7.045 $Y=1.445 $X2=0 $Y2=0
cc_529 N_B_M1012_g N_VGND_c_1389_n 0.00438629f $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_530 N_B_c_582_n N_VGND_c_1389_n 0.00508944f $X=4.3 $Y=1.16 $X2=0 $Y2=0
cc_531 N_B_M1012_g N_VGND_c_1395_n 0.00560495f $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_532 N_B_M1016_g N_VGND_c_1395_n 0.00414252f $X=5.155 $Y=0.565 $X2=0 $Y2=0
cc_533 N_B_c_588_n N_VGND_c_1395_n 0.00357877f $X=6.77 $Y=0.995 $X2=0 $Y2=0
cc_534 N_B_M1012_g N_VGND_c_1398_n 0.0109355f $X=4.225 $Y=0.56 $X2=0 $Y2=0
cc_535 N_B_M1016_g N_VGND_c_1398_n 0.00707752f $X=5.155 $Y=0.565 $X2=0 $Y2=0
cc_536 N_B_c_588_n N_VGND_c_1398_n 0.00596272f $X=6.77 $Y=0.995 $X2=0 $Y2=0
cc_537 N_A_c_703_n N_A_931_365#_c_745_n 0.0247826f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_538 N_A_M1014_g N_A_931_365#_M1009_g 0.0453081f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_539 N_A_M1014_g N_A_931_365#_c_755_n 0.00974519f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_540 N_A_c_701_n N_A_931_365#_c_755_n 0.00302292f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_541 N_A_c_702_n N_A_931_365#_c_755_n 0.0269201f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_542 N_A_c_702_n N_A_931_365#_c_747_n 0.0106752f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_543 N_A_c_703_n N_A_931_365#_c_747_n 0.00845772f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_544 N_A_c_701_n N_A_931_365#_c_748_n 0.00357599f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_545 N_A_c_702_n N_A_931_365#_c_748_n 0.0204454f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_546 N_A_c_703_n N_A_931_365#_c_748_n 0.00178341f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_547 N_A_c_701_n N_A_931_365#_c_749_n 7.09491e-19 $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_548 N_A_c_702_n N_A_931_365#_c_749_n 0.0206309f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_549 N_A_c_703_n N_A_931_365#_c_749_n 0.00347974f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_550 N_A_M1014_g N_A_931_365#_c_757_n 0.00333575f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_551 N_A_c_701_n N_A_931_365#_c_750_n 0.0211645f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_552 N_A_c_702_n N_A_931_365#_c_750_n 8.25692e-19 $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_553 N_A_c_702_n N_A_931_365#_c_781_n 9.51454e-19 $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_554 N_A_c_703_n N_A_931_365#_c_782_n 0.00774108f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_555 N_A_M1014_g N_VPWR_c_907_n 0.00873272f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_556 N_A_M1014_g N_VPWR_c_911_n 0.00337001f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_557 N_A_M1014_g N_VPWR_c_904_n 0.00417888f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_558 N_A_M1014_g N_A_404_49#_c_1156_n 0.00145186f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_559 N_A_M1014_g N_A_1198_49#_c_1334_n 0.0121115f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_560 N_A_M1014_g N_A_1198_49#_c_1327_n 3.59394e-19 $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_561 N_A_c_703_n N_VGND_c_1390_n 0.00268723f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_562 N_A_c_703_n N_VGND_c_1395_n 0.0042601f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_563 N_A_c_703_n N_VGND_c_1398_n 0.00602447f $X=7.74 $Y=0.995 $X2=0 $Y2=0
cc_564 N_A_931_365#_c_755_n N_VPWR_M1014_d 0.00452045f $X=8.085 $Y=1.6 $X2=0
+ $Y2=0
cc_565 N_A_931_365#_M1009_g N_VPWR_c_907_n 0.00837913f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_566 N_A_931_365#_M1009_g N_VPWR_c_912_n 0.00322931f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_567 N_A_931_365#_M1008_d N_VPWR_c_904_n 0.00382772f $X=7.38 $Y=1.645 $X2=0
+ $Y2=0
cc_568 N_A_931_365#_M1009_g N_VPWR_c_904_n 0.00475509f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_569 N_A_931_365#_c_768_n N_A_386_325#_M1021_d 0.00332817f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_570 N_A_931_365#_c_768_n N_A_386_325#_c_1000_n 0.0145847f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_571 N_A_931_365#_c_768_n N_A_386_325#_c_1050_n 0.0145995f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_572 N_A_931_365#_c_781_n N_A_386_325#_c_1050_n 0.00126391f $X=7.59 $Y=0.51
+ $X2=0 $Y2=0
cc_573 N_A_931_365#_c_782_n N_A_386_325#_c_1050_n 0.00765914f $X=7.59 $Y=0.51
+ $X2=0 $Y2=0
cc_574 N_A_931_365#_c_768_n N_A_386_325#_c_1070_n 0.0119237f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_575 N_A_931_365#_M1017_s N_A_386_325#_c_1006_n 0.00764502f $X=4.655 $Y=1.825
+ $X2=0 $Y2=0
cc_576 N_A_931_365#_c_746_n N_A_386_325#_c_1006_n 0.0182772f $X=4.78 $Y=1.94
+ $X2=0 $Y2=0
cc_577 N_A_931_365#_c_768_n N_A_404_49#_M1016_d 0.00519015f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_578 N_A_931_365#_c_746_n N_A_404_49#_c_1151_n 0.0138372f $X=4.78 $Y=1.94
+ $X2=0 $Y2=0
cc_579 N_A_931_365#_c_746_n N_A_404_49#_c_1152_n 0.0028603f $X=4.78 $Y=1.94
+ $X2=0 $Y2=0
cc_580 N_A_931_365#_M1017_s N_A_404_49#_c_1153_n 0.0100815f $X=4.655 $Y=1.825
+ $X2=0 $Y2=0
cc_581 N_A_931_365#_c_746_n N_A_404_49#_c_1153_n 0.0128549f $X=4.78 $Y=1.94
+ $X2=0 $Y2=0
cc_582 N_A_931_365#_c_746_n N_A_404_49#_c_1144_n 0.0675743f $X=4.78 $Y=1.94
+ $X2=0 $Y2=0
cc_583 N_A_931_365#_M1008_d N_A_404_49#_c_1156_n 0.00239642f $X=7.38 $Y=1.645
+ $X2=0 $Y2=0
cc_584 N_A_931_365#_c_768_n N_A_404_49#_c_1200_n 0.0121773f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_585 N_A_931_365#_c_751_n N_A_404_49#_c_1200_n 0.001476f $X=4.975 $Y=0.51
+ $X2=0 $Y2=0
cc_586 N_A_931_365#_c_752_n N_A_404_49#_c_1200_n 0.00942559f $X=4.83 $Y=0.51
+ $X2=0 $Y2=0
cc_587 N_A_931_365#_c_746_n N_A_404_49#_c_1146_n 0.0120431f $X=4.78 $Y=1.94
+ $X2=0 $Y2=0
cc_588 N_A_931_365#_c_768_n N_A_404_49#_c_1146_n 0.00300418f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_589 N_A_931_365#_c_752_n N_A_404_49#_c_1146_n 0.00248625f $X=4.83 $Y=0.51
+ $X2=0 $Y2=0
cc_590 N_A_931_365#_c_768_n N_A_1198_49#_M1018_d 0.00653094f $X=7.445 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_591 N_A_931_365#_c_768_n N_A_1198_49#_c_1321_n 0.00162336f $X=7.445 $Y=0.51
+ $X2=0 $Y2=0
cc_592 N_A_931_365#_c_745_n N_A_1198_49#_c_1322_n 0.00964261f $X=8.23 $Y=0.995
+ $X2=0 $Y2=0
cc_593 N_A_931_365#_M1009_g N_A_1198_49#_c_1322_n 0.0113295f $X=8.23 $Y=1.985
+ $X2=0 $Y2=0
cc_594 N_A_931_365#_c_755_n N_A_1198_49#_c_1322_n 0.0130585f $X=8.085 $Y=1.6
+ $X2=0 $Y2=0
cc_595 N_A_931_365#_c_749_n N_A_1198_49#_c_1322_n 0.040001f $X=8.17 $Y=1.325
+ $X2=0 $Y2=0
cc_596 N_A_931_365#_c_757_n N_A_1198_49#_c_1322_n 0.00963537f $X=8.17 $Y=1.495
+ $X2=0 $Y2=0
cc_597 N_A_931_365#_c_750_n N_A_1198_49#_c_1322_n 0.00752814f $X=8.23 $Y=1.16
+ $X2=0 $Y2=0
cc_598 N_A_931_365#_M1008_d N_A_1198_49#_c_1334_n 0.00689243f $X=7.38 $Y=1.645
+ $X2=0 $Y2=0
cc_599 N_A_931_365#_M1009_g N_A_1198_49#_c_1334_n 0.00253441f $X=8.23 $Y=1.985
+ $X2=0 $Y2=0
cc_600 N_A_931_365#_c_755_n N_A_1198_49#_c_1334_n 0.0324094f $X=8.085 $Y=1.6
+ $X2=0 $Y2=0
cc_601 N_A_931_365#_M1009_g N_A_1198_49#_c_1327_n 0.0090064f $X=8.23 $Y=1.985
+ $X2=0 $Y2=0
cc_602 N_A_931_365#_c_755_n N_A_1198_49#_c_1327_n 0.00661258f $X=8.085 $Y=1.6
+ $X2=0 $Y2=0
cc_603 N_A_931_365#_c_749_n N_A_1198_49#_c_1327_n 0.00152532f $X=8.17 $Y=1.325
+ $X2=0 $Y2=0
cc_604 N_A_931_365#_c_750_n N_A_1198_49#_c_1327_n 7.17833e-19 $X=8.23 $Y=1.16
+ $X2=0 $Y2=0
cc_605 N_A_931_365#_c_750_n N_A_1198_49#_c_1323_n 2.03932e-19 $X=8.23 $Y=1.16
+ $X2=0 $Y2=0
cc_606 N_A_931_365#_c_781_n N_A_1198_49#_c_1323_n 4.91816e-19 $X=7.59 $Y=0.51
+ $X2=0 $Y2=0
cc_607 N_A_931_365#_c_747_n N_VGND_M1007_d 0.00147467f $X=8.085 $Y=0.82 $X2=0
+ $Y2=0
cc_608 N_A_931_365#_c_751_n N_VGND_c_1389_n 7.53702e-19 $X=4.975 $Y=0.51 $X2=0
+ $Y2=0
cc_609 N_A_931_365#_c_745_n N_VGND_c_1390_n 0.00268723f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_610 N_A_931_365#_c_747_n N_VGND_c_1390_n 0.0111874f $X=8.085 $Y=0.82 $X2=0
+ $Y2=0
cc_611 N_A_931_365#_c_749_n N_VGND_c_1390_n 0.00112709f $X=8.17 $Y=1.325 $X2=0
+ $Y2=0
cc_612 N_A_931_365#_c_781_n N_VGND_c_1390_n 0.00115239f $X=7.59 $Y=0.51 $X2=0
+ $Y2=0
cc_613 N_A_931_365#_c_747_n N_VGND_c_1395_n 0.00193763f $X=8.085 $Y=0.82 $X2=0
+ $Y2=0
cc_614 N_A_931_365#_c_768_n N_VGND_c_1395_n 0.00505812f $X=7.445 $Y=0.51 $X2=0
+ $Y2=0
cc_615 N_A_931_365#_c_751_n N_VGND_c_1395_n 2.49898e-19 $X=4.975 $Y=0.51 $X2=0
+ $Y2=0
cc_616 N_A_931_365#_c_752_n N_VGND_c_1395_n 0.024795f $X=4.83 $Y=0.51 $X2=0
+ $Y2=0
cc_617 N_A_931_365#_c_781_n N_VGND_c_1395_n 3.63685e-19 $X=7.59 $Y=0.51 $X2=0
+ $Y2=0
cc_618 N_A_931_365#_c_782_n N_VGND_c_1395_n 0.0143515f $X=7.59 $Y=0.51 $X2=0
+ $Y2=0
cc_619 N_A_931_365#_c_745_n N_VGND_c_1397_n 0.00487842f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_620 N_A_931_365#_c_749_n N_VGND_c_1397_n 0.00181647f $X=8.17 $Y=1.325 $X2=0
+ $Y2=0
cc_621 N_A_931_365#_M1010_d N_VGND_c_1398_n 0.00190368f $X=7.385 $Y=0.235 $X2=0
+ $Y2=0
cc_622 N_A_931_365#_c_745_n N_VGND_c_1398_n 0.00845884f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_623 N_A_931_365#_c_747_n N_VGND_c_1398_n 0.00437041f $X=8.085 $Y=0.82 $X2=0
+ $Y2=0
cc_624 N_A_931_365#_c_749_n N_VGND_c_1398_n 0.00372241f $X=8.17 $Y=1.325 $X2=0
+ $Y2=0
cc_625 N_A_931_365#_c_768_n N_VGND_c_1398_n 0.215427f $X=7.445 $Y=0.51 $X2=0
+ $Y2=0
cc_626 N_A_931_365#_c_751_n N_VGND_c_1398_n 0.0285546f $X=4.975 $Y=0.51 $X2=0
+ $Y2=0
cc_627 N_A_931_365#_c_752_n N_VGND_c_1398_n 0.00391709f $X=4.83 $Y=0.51 $X2=0
+ $Y2=0
cc_628 N_A_931_365#_c_781_n N_VGND_c_1398_n 0.0285254f $X=7.59 $Y=0.51 $X2=0
+ $Y2=0
cc_629 N_A_931_365#_c_782_n N_VGND_c_1398_n 0.00348354f $X=7.59 $Y=0.51 $X2=0
+ $Y2=0
cc_630 X N_VPWR_c_908_n 0.0349912f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_631 N_X_M1002_s N_VPWR_c_904_n 0.00225715f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_632 X N_VPWR_c_904_n 0.0199366f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_633 N_X_c_880_n N_VGND_c_1391_n 0.0208342f $X=0.425 $Y=0.56 $X2=0 $Y2=0
cc_634 N_X_M1001_s N_VGND_c_1398_n 0.00219466f $X=0.3 $Y=0.235 $X2=0 $Y2=0
cc_635 N_X_c_880_n N_VGND_c_1398_n 0.0182278f $X=0.425 $Y=0.56 $X2=0 $Y2=0
cc_636 N_VPWR_c_910_n N_A_386_325#_c_1001_n 0.00328201f $X=3.685 $Y=2.72 $X2=0
+ $Y2=0
cc_637 N_VPWR_c_904_n N_A_386_325#_c_1001_n 0.00795134f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_638 N_VPWR_M1000_s N_A_386_325#_c_1006_n 0.00100785f $X=3.725 $Y=1.485 $X2=0
+ $Y2=0
cc_639 N_VPWR_c_904_n N_A_404_49#_M1011_d 0.00233026f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_640 N_VPWR_c_906_n N_A_404_49#_c_1148_n 0.00147971f $X=3.85 $Y=2.32 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_910_n N_A_404_49#_c_1148_n 0.00296166f $X=3.685 $Y=2.72 $X2=0
+ $Y2=0
cc_642 N_VPWR_c_904_n N_A_404_49#_c_1148_n 0.00485654f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_643 N_VPWR_M1000_s N_A_404_49#_c_1143_n 0.00648805f $X=3.725 $Y=1.485 $X2=0
+ $Y2=0
cc_644 N_VPWR_M1000_s N_A_404_49#_c_1151_n 0.00130442f $X=3.725 $Y=1.485 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_906_n N_A_404_49#_c_1151_n 0.00607843f $X=3.85 $Y=2.32 $X2=0
+ $Y2=0
cc_646 N_VPWR_c_911_n N_A_404_49#_c_1151_n 0.00503515f $X=7.855 $Y=2.72 $X2=0
+ $Y2=0
cc_647 N_VPWR_c_904_n N_A_404_49#_c_1151_n 0.00935628f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_648 N_VPWR_c_906_n N_A_404_49#_c_1152_n 0.00173147f $X=3.85 $Y=2.32 $X2=0
+ $Y2=0
cc_649 N_VPWR_c_911_n N_A_404_49#_c_1153_n 0.0294498f $X=7.855 $Y=2.72 $X2=0
+ $Y2=0
cc_650 N_VPWR_c_904_n N_A_404_49#_c_1153_n 0.0189426f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_651 N_VPWR_c_906_n N_A_404_49#_c_1154_n 0.00833535f $X=3.85 $Y=2.32 $X2=0
+ $Y2=0
cc_652 N_VPWR_c_911_n N_A_404_49#_c_1154_n 0.0105745f $X=7.855 $Y=2.72 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_904_n N_A_404_49#_c_1154_n 0.00644066f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_907_n N_A_404_49#_c_1156_n 0.00704283f $X=8.02 $Y=2.36 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_911_n N_A_404_49#_c_1156_n 0.124148f $X=7.855 $Y=2.72 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_904_n N_A_404_49#_c_1156_n 0.074875f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_657 N_VPWR_c_906_n N_A_404_49#_c_1157_n 0.0142739f $X=3.85 $Y=2.32 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_910_n N_A_404_49#_c_1157_n 0.0186431f $X=3.685 $Y=2.72 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_904_n N_A_404_49#_c_1157_n 0.0145279f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_660 N_VPWR_M1000_s N_A_404_49#_c_1158_n 0.00234468f $X=3.725 $Y=1.485 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_906_n N_A_404_49#_c_1158_n 0.0143988f $X=3.85 $Y=2.32 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_904_n N_A_404_49#_c_1158_n 8.22076e-19 $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_911_n N_A_404_49#_c_1159_n 0.0103342f $X=7.855 $Y=2.72 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_904_n N_A_404_49#_c_1159_n 0.00589464f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_665 N_VPWR_c_904_n N_A_1198_49#_M1009_d 0.00248304f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_912_n N_A_1198_49#_c_1325_n 0.0197307f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_904_n N_A_1198_49#_c_1325_n 0.0111012f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_668 N_VPWR_M1014_d N_A_1198_49#_c_1334_n 0.00343874f $X=7.885 $Y=1.485 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_907_n N_A_1198_49#_c_1334_n 0.0162117f $X=8.02 $Y=2.36 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_911_n N_A_1198_49#_c_1334_n 0.00690051f $X=7.855 $Y=2.72 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_904_n N_A_1198_49#_c_1334_n 0.0144976f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_912_n N_A_1198_49#_c_1327_n 0.00258024f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_904_n N_A_1198_49#_c_1327_n 0.00441029f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_674 N_A_386_325#_c_1001_n N_A_404_49#_M1020_d 0.00597024f $X=3.005 $Y=1.98
+ $X2=0 $Y2=0
cc_675 N_A_386_325#_c_1022_n N_A_404_49#_M1020_d 0.00664959f $X=3.09 $Y=1.895
+ $X2=0 $Y2=0
cc_676 N_A_386_325#_c_1009_n N_A_404_49#_M1020_d 0.00687512f $X=3.335 $Y=1.535
+ $X2=0 $Y2=0
cc_677 N_A_386_325#_M1013_d N_A_404_49#_c_1140_n 0.00334341f $X=2.99 $Y=0.245
+ $X2=0 $Y2=0
cc_678 N_A_386_325#_c_999_n N_A_404_49#_c_1140_n 0.0138308f $X=3.335 $Y=0.76
+ $X2=0 $Y2=0
cc_679 N_A_386_325#_M1013_d N_A_404_49#_c_1164_n 0.00347935f $X=2.99 $Y=0.245
+ $X2=0 $Y2=0
cc_680 N_A_386_325#_c_999_n N_A_404_49#_c_1164_n 0.00432164f $X=3.335 $Y=0.76
+ $X2=0 $Y2=0
cc_681 N_A_386_325#_M1013_d N_A_404_49#_c_1141_n 0.0175141f $X=2.99 $Y=0.245
+ $X2=0 $Y2=0
cc_682 N_A_386_325#_c_999_n N_A_404_49#_c_1141_n 0.0128008f $X=3.335 $Y=0.76
+ $X2=0 $Y2=0
cc_683 N_A_386_325#_M1013_d N_A_404_49#_c_1165_n 3.2099e-19 $X=2.99 $Y=0.245
+ $X2=0 $Y2=0
cc_684 N_A_386_325#_c_1006_n N_A_404_49#_c_1148_n 0.00437461f $X=5.605 $Y=1.53
+ $X2=0 $Y2=0
cc_685 N_A_386_325#_c_1007_n N_A_404_49#_c_1148_n 0.00277011f $X=3.595 $Y=1.53
+ $X2=0 $Y2=0
cc_686 N_A_386_325#_c_1009_n N_A_404_49#_c_1148_n 0.00125154f $X=3.335 $Y=1.535
+ $X2=0 $Y2=0
cc_687 N_A_386_325#_c_1001_n N_A_404_49#_c_1149_n 0.0153275f $X=3.005 $Y=1.98
+ $X2=0 $Y2=0
cc_688 N_A_386_325#_c_1007_n N_A_404_49#_c_1149_n 0.00119193f $X=3.595 $Y=1.53
+ $X2=0 $Y2=0
cc_689 N_A_386_325#_c_1009_n N_A_404_49#_c_1149_n 0.0114314f $X=3.335 $Y=1.535
+ $X2=0 $Y2=0
cc_690 N_A_386_325#_c_999_n N_A_404_49#_c_1142_n 0.0327455f $X=3.335 $Y=0.76
+ $X2=0 $Y2=0
cc_691 N_A_386_325#_c_1022_n N_A_404_49#_c_1143_n 0.00649967f $X=3.09 $Y=1.895
+ $X2=0 $Y2=0
cc_692 N_A_386_325#_c_999_n N_A_404_49#_c_1143_n 0.00891656f $X=3.335 $Y=0.76
+ $X2=0 $Y2=0
cc_693 N_A_386_325#_c_1006_n N_A_404_49#_c_1143_n 0.0161183f $X=5.605 $Y=1.53
+ $X2=0 $Y2=0
cc_694 N_A_386_325#_c_1007_n N_A_404_49#_c_1143_n 0.00275249f $X=3.595 $Y=1.53
+ $X2=0 $Y2=0
cc_695 N_A_386_325#_c_1009_n N_A_404_49#_c_1143_n 0.0233324f $X=3.335 $Y=1.535
+ $X2=0 $Y2=0
cc_696 N_A_386_325#_c_1006_n N_A_404_49#_c_1151_n 0.0108493f $X=5.605 $Y=1.53
+ $X2=0 $Y2=0
cc_697 N_A_386_325#_c_1003_n N_A_404_49#_c_1144_n 0.010588f $X=5.602 $Y=1.615
+ $X2=0 $Y2=0
cc_698 N_A_386_325#_c_1039_n N_A_404_49#_c_1144_n 0.0296035f $X=5.57 $Y=1.62
+ $X2=0 $Y2=0
cc_699 N_A_386_325#_c_1006_n N_A_404_49#_c_1144_n 0.0192106f $X=5.605 $Y=1.53
+ $X2=0 $Y2=0
cc_700 N_A_386_325#_c_1008_n N_A_404_49#_c_1144_n 0.0013191f $X=5.75 $Y=1.53
+ $X2=0 $Y2=0
cc_701 N_A_386_325#_M1017_d N_A_404_49#_c_1156_n 0.00904513f $X=5.23 $Y=1.485
+ $X2=0 $Y2=0
cc_702 N_A_386_325#_c_1039_n N_A_404_49#_c_1156_n 0.0235166f $X=5.57 $Y=1.62
+ $X2=0 $Y2=0
cc_703 N_A_386_325#_c_1004_n N_A_404_49#_c_1156_n 0.00873322f $X=6.005 $Y=1.53
+ $X2=0 $Y2=0
cc_704 N_A_386_325#_c_1000_n N_A_404_49#_c_1200_n 0.0028148f $X=6.09 $Y=1.445
+ $X2=0 $Y2=0
cc_705 N_A_386_325#_c_1001_n N_A_404_49#_c_1157_n 0.0049241f $X=3.005 $Y=1.98
+ $X2=0 $Y2=0
cc_706 N_A_386_325#_c_1007_n N_A_404_49#_c_1157_n 2.48159e-19 $X=3.595 $Y=1.53
+ $X2=0 $Y2=0
cc_707 N_A_386_325#_c_1009_n N_A_404_49#_c_1157_n 0.00535873f $X=3.335 $Y=1.535
+ $X2=0 $Y2=0
cc_708 N_A_386_325#_c_999_n N_A_404_49#_c_1145_n 0.0132287f $X=3.335 $Y=0.76
+ $X2=0 $Y2=0
cc_709 N_A_386_325#_c_1006_n N_A_404_49#_c_1145_n 0.0052436f $X=5.605 $Y=1.53
+ $X2=0 $Y2=0
cc_710 N_A_386_325#_c_1007_n N_A_404_49#_c_1145_n 2.29009e-19 $X=3.595 $Y=1.53
+ $X2=0 $Y2=0
cc_711 N_A_386_325#_c_1003_n N_A_404_49#_c_1146_n 2.53366e-19 $X=5.602 $Y=1.615
+ $X2=0 $Y2=0
cc_712 N_A_386_325#_c_1006_n N_A_404_49#_c_1146_n 4.20548e-19 $X=5.605 $Y=1.53
+ $X2=0 $Y2=0
cc_713 N_A_386_325#_c_1000_n N_A_1198_49#_M1018_d 0.00729398f $X=6.09 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_714 N_A_386_325#_c_1126_p N_A_1198_49#_M1018_d 0.0024562f $X=6.175 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_715 N_A_386_325#_c_1070_n N_A_1198_49#_M1018_d 0.0107136f $X=6.685 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_716 N_A_386_325#_c_1004_n N_A_1198_49#_M1015_d 0.00414782f $X=6.005 $Y=1.53
+ $X2=0 $Y2=0
cc_717 N_A_386_325#_c_1039_n N_A_1198_49#_c_1321_n 0.00487817f $X=5.57 $Y=1.62
+ $X2=0 $Y2=0
cc_718 N_A_386_325#_c_1004_n N_A_1198_49#_c_1321_n 0.0134336f $X=6.005 $Y=1.53
+ $X2=0 $Y2=0
cc_719 N_A_386_325#_c_1000_n N_A_1198_49#_c_1321_n 0.0622566f $X=6.09 $Y=1.445
+ $X2=0 $Y2=0
cc_720 N_A_386_325#_c_1070_n N_A_1198_49#_c_1321_n 0.0106102f $X=6.685 $Y=0.36
+ $X2=0 $Y2=0
cc_721 N_A_386_325#_c_1008_n N_A_1198_49#_c_1321_n 0.0013871f $X=5.75 $Y=1.53
+ $X2=0 $Y2=0
cc_722 N_A_386_325#_c_1006_n N_VGND_c_1389_n 0.00555354f $X=5.605 $Y=1.53 $X2=0
+ $Y2=0
cc_723 N_A_386_325#_c_1126_p N_VGND_c_1395_n 0.0104913f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_724 N_A_386_325#_c_1070_n N_VGND_c_1395_n 0.0586043f $X=6.685 $Y=0.36 $X2=0
+ $Y2=0
cc_725 N_A_386_325#_M1021_d N_VGND_c_1398_n 0.00184103f $X=6.785 $Y=0.245 $X2=0
+ $Y2=0
cc_726 N_A_386_325#_c_1126_p N_VGND_c_1398_n 0.00184693f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_727 N_A_386_325#_c_1070_n N_VGND_c_1398_n 0.0092581f $X=6.685 $Y=0.36 $X2=0
+ $Y2=0
cc_728 N_A_404_49#_c_1156_n N_A_1198_49#_M1015_d 0.0055303f $X=7.085 $Y=2.36
+ $X2=0 $Y2=0
cc_729 N_A_404_49#_c_1156_n N_A_1198_49#_c_1333_n 0.0129278f $X=7.085 $Y=2.36
+ $X2=0 $Y2=0
cc_730 N_A_404_49#_M1011_d N_A_1198_49#_c_1334_n 0.00612338f $X=6.865 $Y=1.645
+ $X2=0 $Y2=0
cc_731 N_A_404_49#_c_1156_n N_A_1198_49#_c_1334_n 0.0467387f $X=7.085 $Y=2.36
+ $X2=0 $Y2=0
cc_732 N_A_404_49#_c_1141_n N_VGND_c_1389_n 0.0141315f $X=3.59 $Y=0.34 $X2=0
+ $Y2=0
cc_733 N_A_404_49#_c_1142_n N_VGND_c_1389_n 0.0321143f $X=3.675 $Y=1.035 $X2=0
+ $Y2=0
cc_734 N_A_404_49#_c_1140_n N_VGND_c_1393_n 0.00233735f $X=2.91 $Y=0.74 $X2=0
+ $Y2=0
cc_735 N_A_404_49#_c_1141_n N_VGND_c_1393_n 0.0445697f $X=3.59 $Y=0.34 $X2=0
+ $Y2=0
cc_736 N_A_404_49#_c_1165_n N_VGND_c_1393_n 0.0096984f $X=3.08 $Y=0.34 $X2=0
+ $Y2=0
cc_737 N_A_404_49#_c_1200_n N_VGND_c_1395_n 0.00800682f $X=5.365 $Y=0.545 $X2=0
+ $Y2=0
cc_738 N_A_404_49#_c_1146_n N_VGND_c_1395_n 0.00224122f $X=5.12 $Y=0.772 $X2=0
+ $Y2=0
cc_739 N_A_404_49#_c_1140_n N_VGND_c_1398_n 0.00612861f $X=2.91 $Y=0.74 $X2=0
+ $Y2=0
cc_740 N_A_404_49#_c_1141_n N_VGND_c_1398_n 0.0255342f $X=3.59 $Y=0.34 $X2=0
+ $Y2=0
cc_741 N_A_404_49#_c_1165_n N_VGND_c_1398_n 0.00615131f $X=3.08 $Y=0.34 $X2=0
+ $Y2=0
cc_742 N_A_404_49#_c_1200_n N_VGND_c_1398_n 0.0018012f $X=5.365 $Y=0.545 $X2=0
+ $Y2=0
cc_743 N_A_1198_49#_c_1323_n N_VGND_c_1397_n 0.0197576f $X=8.57 $Y=0.42 $X2=0
+ $Y2=0
cc_744 N_A_1198_49#_M1006_d N_VGND_c_1398_n 0.00399944f $X=8.305 $Y=0.235 $X2=0
+ $Y2=0
cc_745 N_A_1198_49#_c_1323_n N_VGND_c_1398_n 0.0113402f $X=8.57 $Y=0.42 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__clkinv_1.pex.spice
* Created: Thu Aug 27 14:12:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINV_1%A 3 7 11 13 14 15 23
r30 23 24 0.678873 $w=3.55e-07 $l=5e-09 $layer=POLY_cond $X=0.885 $Y=1.16
+ $X2=0.89 $Y2=1.16
r31 22 23 56.3465 $w=3.55e-07 $l=4.15e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.885 $Y2=1.16
r32 20 22 31.2282 $w=3.55e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r33 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r34 14 15 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.205 $Y=0.85
+ $X2=0.205 $Y2=1.16
r35 13 14 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.205 $Y=0.51
+ $X2=0.205 $Y2=0.85
r36 9 24 22.9692 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.89 $Y=1.345
+ $X2=0.89 $Y2=1.16
r37 9 11 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.89 $Y=1.345
+ $X2=0.89 $Y2=2.065
r38 5 23 22.9692 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.885 $Y=0.975
+ $X2=0.885 $Y2=1.16
r39 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.885 $Y=0.975
+ $X2=0.885 $Y2=0.445
r40 1 22 22.9692 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.47 $Y=1.345
+ $X2=0.47 $Y2=1.16
r41 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.47 $Y=1.345 $X2=0.47
+ $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_1%VPWR 1 2 7 9 11 13 15 17 27
r19 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r20 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r21 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r22 18 23 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r23 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r24 17 26 4.33505 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.197 $Y2=2.72
r25 17 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r26 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r27 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r28 11 26 3.02501 $w=2.8e-07 $l=1.03899e-07 $layer=LI1_cond $X=1.155 $Y=2.635
+ $X2=1.197 $Y2=2.72
r29 11 13 33.1327 $w=2.78e-07 $l=8.05e-07 $layer=LI1_cond $X=1.155 $Y=2.635
+ $X2=1.155 $Y2=1.83
r30 7 23 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r31 7 9 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=1.83
r32 2 13 300 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.645 $X2=1.1 $Y2=1.83
r33 1 9 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.645 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_1%Y 1 2 9 11 13 14
r22 27 29 0.0677026 $w=5.28e-07 $l=3e-09 $layer=LI1_cond $X=0.677 $Y=1.025
+ $X2=0.68 $Y2=1.025
r23 21 29 3.50913 $w=3.3e-07 $l=2.65e-07 $layer=LI1_cond $X=0.68 $Y=1.29
+ $X2=0.68 $Y2=1.025
r24 13 25 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.68 $Y=1.53 $X2=0.68
+ $Y2=1.83
r25 13 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.68 $Y=1.53 $X2=0.68
+ $Y2=1.29
r26 11 14 10.3811 $w=5.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=1.15 $Y2=1.025
r27 11 29 0.225675 $w=5.28e-07 $l=1e-08 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.68 $Y2=1.025
r28 7 27 3.60987 $w=3.25e-07 $l=2.65e-07 $layer=LI1_cond $X=0.677 $Y=0.76
+ $X2=0.677 $Y2=1.025
r29 7 9 11.5244 $w=3.23e-07 $l=3.25e-07 $layer=LI1_cond $X=0.677 $Y=0.76
+ $X2=0.677 $Y2=0.435
r30 2 25 300 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.645 $X2=0.68 $Y2=1.83
r31 1 9 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.675 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_1%VGND 1 4 6 8 10 17
r15 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r16 13 17 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r17 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r18 10 16 4.37302 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.195
+ $Y2=0
r19 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.69
+ $Y2=0
r20 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r21 4 16 3.02565 $w=2.85e-07 $l=1.04307e-07 $layer=LI1_cond $X=1.152 $Y=0.085
+ $X2=1.195 $Y2=0
r22 4 6 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.152 $Y=0.085
+ $X2=1.152 $Y2=0.425
r23 1 6 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.235 $X2=1.095 $Y2=0.425
.ends


* File: sky130_fd_sc_hd__o31ai_4.spice.SKY130_FD_SC_HD__O31AI_4.pxi
* Created: Thu Aug 27 14:40:37 2020
* 
x_PM_SKY130_FD_SC_HD__O31AI_4%A1 N_A1_M1008_g N_A1_M1007_g N_A1_M1012_g
+ N_A1_M1022_g N_A1_M1019_g N_A1_M1026_g N_A1_M1020_g N_A1_M1031_g A1 A1 A1 A1
+ N_A1_c_125_n PM_SKY130_FD_SC_HD__O31AI_4%A1
x_PM_SKY130_FD_SC_HD__O31AI_4%A2 N_A2_M1016_g N_A2_M1005_g N_A2_M1021_g
+ N_A2_M1017_g N_A2_M1023_g N_A2_M1018_g N_A2_M1029_g N_A2_M1027_g A2 A2 A2 A2
+ N_A2_c_216_n PM_SKY130_FD_SC_HD__O31AI_4%A2
x_PM_SKY130_FD_SC_HD__O31AI_4%A3 N_A3_M1001_g N_A3_M1004_g N_A3_M1002_g
+ N_A3_M1009_g N_A3_M1013_g N_A3_M1028_g N_A3_M1024_g N_A3_M1030_g N_A3_c_307_n
+ A3 A3 A3 A3 A3 N_A3_c_309_n N_A3_c_310_n PM_SKY130_FD_SC_HD__O31AI_4%A3
x_PM_SKY130_FD_SC_HD__O31AI_4%B1 N_B1_M1003_g N_B1_M1000_g N_B1_M1006_g
+ N_B1_M1010_g N_B1_M1011_g N_B1_M1015_g N_B1_M1014_g N_B1_M1025_g B1 B1 B1
+ N_B1_c_384_n PM_SKY130_FD_SC_HD__O31AI_4%B1
x_PM_SKY130_FD_SC_HD__O31AI_4%A_27_297# N_A_27_297#_M1007_s N_A_27_297#_M1022_s
+ N_A_27_297#_M1031_s N_A_27_297#_M1017_d N_A_27_297#_M1027_d
+ N_A_27_297#_c_449_n N_A_27_297#_c_450_n N_A_27_297#_c_456_n
+ N_A_27_297#_c_460_n N_A_27_297#_c_464_n N_A_27_297#_c_468_n
+ N_A_27_297#_c_469_n N_A_27_297#_c_479_n N_A_27_297#_c_451_n
+ N_A_27_297#_c_471_n N_A_27_297#_c_483_n PM_SKY130_FD_SC_HD__O31AI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__O31AI_4%VPWR N_VPWR_M1007_d N_VPWR_M1026_d N_VPWR_M1000_s
+ N_VPWR_M1015_s N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n
+ VPWR N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n
+ N_VPWR_c_522_n N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n
+ PM_SKY130_FD_SC_HD__O31AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O31AI_4%A_449_297# N_A_449_297#_M1005_s
+ N_A_449_297#_M1018_s N_A_449_297#_M1004_s N_A_449_297#_M1028_s
+ N_A_449_297#_c_627_n N_A_449_297#_c_637_n N_A_449_297#_c_628_n
+ N_A_449_297#_c_630_n N_A_449_297#_c_634_n N_A_449_297#_c_626_n
+ PM_SKY130_FD_SC_HD__O31AI_4%A_449_297#
x_PM_SKY130_FD_SC_HD__O31AI_4%Y N_Y_M1003_s N_Y_M1011_s N_Y_M1004_d N_Y_M1009_d
+ N_Y_M1030_d N_Y_M1010_d N_Y_M1025_d N_Y_c_716_n N_Y_c_718_n Y Y Y Y Y Y Y Y Y
+ Y Y Y Y N_Y_c_671_n Y N_Y_c_696_n N_Y_c_672_n N_Y_c_673_n N_Y_c_674_n
+ N_Y_c_706_n PM_SKY130_FD_SC_HD__O31AI_4%Y
x_PM_SKY130_FD_SC_HD__O31AI_4%A_31_47# N_A_31_47#_M1008_s N_A_31_47#_M1012_s
+ N_A_31_47#_M1020_s N_A_31_47#_M1021_d N_A_31_47#_M1029_d N_A_31_47#_M1002_d
+ N_A_31_47#_M1024_d N_A_31_47#_M1006_d N_A_31_47#_M1014_d N_A_31_47#_c_741_n
+ N_A_31_47#_c_753_n N_A_31_47#_c_742_n N_A_31_47#_c_759_n N_A_31_47#_c_763_n
+ N_A_31_47#_c_767_n N_A_31_47#_c_776_n N_A_31_47#_c_780_n N_A_31_47#_c_784_n
+ N_A_31_47#_c_788_n N_A_31_47#_c_799_n N_A_31_47#_c_845_p N_A_31_47#_c_743_n
+ N_A_31_47#_c_811_n N_A_31_47#_c_849_p N_A_31_47#_c_744_n N_A_31_47#_c_745_n
+ N_A_31_47#_c_746_n N_A_31_47#_c_747_n N_A_31_47#_c_748_n N_A_31_47#_c_749_n
+ N_A_31_47#_c_750_n PM_SKY130_FD_SC_HD__O31AI_4%A_31_47#
x_PM_SKY130_FD_SC_HD__O31AI_4%VGND N_VGND_M1008_d N_VGND_M1019_d N_VGND_M1016_s
+ N_VGND_M1023_s N_VGND_M1001_s N_VGND_M1013_s N_VGND_c_882_n N_VGND_c_883_n
+ N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n VGND
+ N_VGND_c_893_n N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n
+ N_VGND_c_898_n N_VGND_c_899_n PM_SKY130_FD_SC_HD__O31AI_4%VGND
cc_1 VNB N_A1_M1008_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_2 VNB N_A1_M1007_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_3 VNB N_A1_M1012_g 0.017456f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_4 VNB N_A1_M1022_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_5 VNB N_A1_M1019_g 0.017456f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_6 VNB N_A1_M1026_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_7 VNB N_A1_M1020_g 0.0177503f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_8 VNB N_A1_M1031_g 4.2554e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_9 VNB A1 0.0144966f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_10 VNB N_A1_c_125_n 0.0681838f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_11 VNB N_A2_M1016_g 0.0177503f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_12 VNB N_A2_M1005_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_13 VNB N_A2_M1021_g 0.017456f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_14 VNB N_A2_M1017_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_15 VNB N_A2_M1023_g 0.017456f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_16 VNB N_A2_M1018_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_17 VNB N_A2_M1029_g 0.0177503f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_18 VNB N_A2_M1027_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_19 VNB A2 0.00575743f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_20 VNB N_A2_c_216_n 0.0617935f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_21 VNB N_A3_M1001_g 0.0211443f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_22 VNB N_A3_M1004_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_23 VNB N_A3_M1002_g 0.0204855f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_24 VNB N_A3_M1009_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_25 VNB N_A3_M1013_g 0.0184397f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_26 VNB N_A3_M1028_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_27 VNB N_A3_M1024_g 0.0187228f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_28 VNB N_A3_M1030_g 4.65066e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_29 VNB N_A3_c_307_n 0.0120068f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_30 VNB A3 0.00698319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A3_c_309_n 0.0270143f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_32 VNB N_A3_c_310_n 0.0639108f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.24
cc_33 VNB N_B1_M1003_g 0.0172035f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_34 VNB N_B1_M1000_g 4.28089e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_35 VNB N_B1_M1006_g 0.0174197f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_36 VNB N_B1_M1010_g 4.47843e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_37 VNB N_B1_M1011_g 0.0174522f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_38 VNB N_B1_M1015_g 4.49965e-19 $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_39 VNB N_B1_M1014_g 0.0243627f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_40 VNB N_B1_M1025_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_41 VNB B1 0.0143034f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_42 VNB N_B1_c_384_n 0.0740056f $X=-0.19 $Y=-0.24 $X2=1.275 $Y2=1.16
cc_43 VNB N_VPWR_c_522_n 0.326667f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.16
cc_44 VNB Y 0.00139886f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_45 VNB N_A_31_47#_c_741_n 0.0188118f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_46 VNB N_A_31_47#_c_742_n 0.00983636f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_47 VNB N_A_31_47#_c_743_n 0.001463f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.24
cc_48 VNB N_A_31_47#_c_744_n 0.0101084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_31_47#_c_745_n 0.0186289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_31_47#_c_746_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_31_47#_c_747_n 0.00356912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_31_47#_c_748_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_31_47#_c_749_n 0.00496288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_31_47#_c_750_n 0.00115893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_882_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_56 VNB N_VGND_c_883_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_57 VNB N_VGND_c_884_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_58 VNB N_VGND_c_885_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_59 VNB N_VGND_c_886_n 5.61194e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_887_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_888_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_62 VNB N_VGND_c_889_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_63 VNB N_VGND_c_890_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_64 VNB N_VGND_c_891_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=1.275 $Y2=1.16
cc_65 VNB N_VGND_c_892_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=1.275 $Y2=1.16
cc_66 VNB N_VGND_c_893_n 0.0115586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_894_n 0.0521194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_895_n 0.371379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_896_n 0.0208501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_897_n 0.0172004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_898_n 0.0156478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_899_n 0.00614073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VPB N_A1_M1007_g 0.0249717f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_74 VPB N_A1_M1022_g 0.0185598f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_75 VPB N_A1_M1026_g 0.0185598f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_76 VPB N_A1_M1031_g 0.0193917f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_77 VPB A1 0.0160415f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_78 VPB N_A2_M1005_g 0.0187304f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_79 VPB N_A2_M1017_g 0.0185598f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_80 VPB N_A2_M1018_g 0.0185595f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_81 VPB N_A2_M1027_g 0.0240633f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_82 VPB A2 0.0168232f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_83 VPB N_A3_M1004_g 0.0267252f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_84 VPB N_A3_M1009_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_85 VPB N_A3_M1028_g 0.0191885f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_86 VPB N_A3_M1030_g 0.0194609f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_87 VPB N_B1_M1000_g 0.0186603f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_88 VPB N_B1_M1010_g 0.0189074f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_89 VPB N_B1_M1015_g 0.0189404f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_90 VPB N_B1_M1025_g 0.026498f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_91 VPB N_A_27_297#_c_449_n 0.0131401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_297#_c_450_n 0.0226427f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_93 VPB N_A_27_297#_c_451_n 0.00449223f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_94 VPB N_VPWR_c_523_n 0.00410835f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.025
cc_95 VPB N_VPWR_c_524_n 0.00410284f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.295
cc_96 VPB N_VPWR_c_525_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.025
cc_97 VPB N_VPWR_c_526_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.295
cc_98 VPB N_VPWR_c_527_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_99 VPB N_VPWR_c_528_n 0.104184f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_529_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_101 VPB N_VPWR_c_530_n 0.015618f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_102 VPB N_VPWR_c_522_n 0.0477745f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.16
cc_103 VPB N_VPWR_c_532_n 0.0214916f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_104 VPB N_VPWR_c_533_n 0.00323699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_534_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.24
cc_106 VPB N_VPWR_c_535_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_449_297#_c_626_n 0.00804166f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_108 VPB Y 0.00175406f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_109 VPB Y 0.00375323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB Y 0.0012991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB Y 0.0307929f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_112 VPB N_Y_c_671_n 0.0174025f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.24
cc_113 VPB N_Y_c_672_n 0.00186725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_Y_c_673_n 0.00295125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_Y_c_674_n 0.013547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 N_A1_M1020_g N_A2_M1016_g 0.0143105f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_117 N_A1_M1031_g N_A2_M1005_g 0.0143105f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_118 A1 A2 0.0327645f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_119 N_A1_c_125_n A2 0.00288484f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_120 A1 N_A2_c_216_n 3.34444e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A1_c_125_n N_A2_c_216_n 0.0143105f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A1_M1007_g N_A_27_297#_c_449_n 0.00123961f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_123 A1 N_A_27_297#_c_449_n 0.0283057f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A1_M1007_g N_A_27_297#_c_450_n 0.00735265f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A1_M1022_g N_A_27_297#_c_450_n 6.15622e-19 $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A1_M1007_g N_A_27_297#_c_456_n 0.0114894f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A1_M1022_g N_A_27_297#_c_456_n 0.0114894f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_128 A1 N_A_27_297#_c_456_n 0.035571f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_129 N_A1_c_125_n N_A_27_297#_c_456_n 4.81973e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_M1007_g N_A_27_297#_c_460_n 6.16084e-19 $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_M1022_g N_A_27_297#_c_460_n 0.00735265f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A1_M1026_g N_A_27_297#_c_460_n 0.00735265f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A1_M1031_g N_A_27_297#_c_460_n 6.16084e-19 $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A1_M1026_g N_A_27_297#_c_464_n 0.0114894f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A1_M1031_g N_A_27_297#_c_464_n 0.0119542f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_136 A1 N_A_27_297#_c_464_n 0.0344805f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A1_c_125_n N_A_27_297#_c_464_n 4.81973e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_M1031_g N_A_27_297#_c_468_n 0.00232477f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_M1026_g N_A_27_297#_c_469_n 5.39159e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_M1031_g N_A_27_297#_c_469_n 0.00736261f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_M1022_g N_A_27_297#_c_471_n 0.00123961f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A1_M1026_g N_A_27_297#_c_471_n 0.00123961f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_143 A1 N_A_27_297#_c_471_n 0.0232321f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A1_c_125_n N_A_27_297#_c_471_n 5.20942e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A1_M1007_g N_VPWR_c_523_n 0.00301669f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1022_g N_VPWR_c_523_n 0.00179394f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_M1026_g N_VPWR_c_524_n 0.00179394f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A1_M1031_g N_VPWR_c_524_n 0.00301669f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A1_M1022_g N_VPWR_c_527_n 0.00541359f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A1_M1026_g N_VPWR_c_527_n 0.00541359f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A1_M1031_g N_VPWR_c_528_n 0.00539841f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1007_g N_VPWR_c_522_n 0.00688717f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A1_M1022_g N_VPWR_c_522_n 0.00591429f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A1_M1026_g N_VPWR_c_522_n 0.00591429f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A1_M1031_g N_VPWR_c_522_n 0.00595057f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A1_M1007_g N_VPWR_c_532_n 0.00541359f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A1_M1008_g N_A_31_47#_c_741_n 0.00620543f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_158 N_A1_M1012_g N_A_31_47#_c_741_n 5.18879e-19 $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A1_M1008_g N_A_31_47#_c_753_n 0.00844123f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A1_M1012_g N_A_31_47#_c_753_n 0.00844123f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_161 A1 N_A_31_47#_c_753_n 0.0332055f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A1_c_125_n N_A_31_47#_c_753_n 0.0020061f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A1_M1008_g N_A_31_47#_c_742_n 8.68782e-19 $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_164 A1 N_A_31_47#_c_742_n 0.0281907f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A1_M1008_g N_A_31_47#_c_759_n 5.19281e-19 $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A1_M1012_g N_A_31_47#_c_759_n 0.00620543f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A1_M1019_g N_A_31_47#_c_759_n 0.00620543f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A1_M1020_g N_A_31_47#_c_759_n 5.19281e-19 $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A1_M1019_g N_A_31_47#_c_763_n 0.00844123f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_170 N_A1_M1020_g N_A_31_47#_c_763_n 0.00886881f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_171 A1 N_A_31_47#_c_763_n 0.0321583f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A1_c_125_n N_A_31_47#_c_763_n 0.0020061f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A1_M1019_g N_A_31_47#_c_767_n 5.19281e-19 $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A1_M1020_g N_A_31_47#_c_767_n 0.00620543f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A1_M1012_g N_A_31_47#_c_746_n 8.68782e-19 $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A1_M1019_g N_A_31_47#_c_746_n 8.68782e-19 $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_177 A1 N_A_31_47#_c_746_n 0.0219994f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A1_c_125_n N_A_31_47#_c_746_n 0.00208088f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A1_M1020_g N_A_31_47#_c_747_n 0.00190519f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A1_M1008_g N_VGND_c_882_n 0.00268723f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A1_M1012_g N_VGND_c_882_n 0.00146448f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A1_M1019_g N_VGND_c_883_n 0.00146448f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A1_M1020_g N_VGND_c_883_n 0.00146448f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A1_M1012_g N_VGND_c_887_n 0.00422241f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A1_M1019_g N_VGND_c_887_n 0.00422241f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A1_M1020_g N_VGND_c_889_n 0.00422241f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A1_M1008_g N_VGND_c_895_n 0.00666944f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A1_M1012_g N_VGND_c_895_n 0.00569656f $X=0.91 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A1_M1019_g N_VGND_c_895_n 0.00569656f $X=1.33 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A1_M1020_g N_VGND_c_895_n 0.00572376f $X=1.75 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A1_M1008_g N_VGND_c_896_n 0.00422241f $X=0.49 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A2_M1029_g N_A3_M1001_g 0.0137836f $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_193 A2 N_A3_c_307_n 0.00146591f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_194 N_A2_c_216_n N_A3_c_307_n 0.0137836f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_195 A2 A3 0.0194357f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_196 N_A2_c_216_n A3 2.27279e-19 $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A2_M1005_g N_A_27_297#_c_468_n 0.00355506f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_198 A2 N_A_27_297#_c_468_n 0.0124903f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A2_M1005_g N_A_27_297#_c_469_n 0.00534917f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A2_M1017_g N_A_27_297#_c_469_n 5.39159e-19 $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A2_M1005_g N_A_27_297#_c_479_n 0.0124301f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A2_M1017_g N_A_27_297#_c_479_n 0.0105223f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A2_M1018_g N_A_27_297#_c_451_n 0.0105223f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A2_M1027_g N_A_27_297#_c_451_n 0.00996642f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A2_M1005_g N_A_27_297#_c_483_n 6.5188e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A2_M1017_g N_A_27_297#_c_483_n 0.00610524f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A2_M1018_g N_A_27_297#_c_483_n 0.00631336f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_M1027_g N_A_27_297#_c_483_n 0.00103389f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_M1005_g N_VPWR_c_528_n 0.00357835f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1017_g N_VPWR_c_528_n 0.00359354f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A2_M1018_g N_VPWR_c_528_n 0.00359354f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A2_M1027_g N_VPWR_c_528_n 0.00357877f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A2_M1005_g N_VPWR_c_522_n 0.00525234f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A2_M1017_g N_VPWR_c_522_n 0.00521606f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A2_M1018_g N_VPWR_c_522_n 0.00521606f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A2_M1027_g N_VPWR_c_522_n 0.00655123f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A2_M1027_g N_A_449_297#_c_627_n 0.00415651f $X=3.43 $Y=1.985 $X2=0
+ $Y2=0
cc_218 A2 N_A_449_297#_c_628_n 0.0137102f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_219 N_A2_c_216_n N_A_449_297#_c_628_n 4.98274e-19 $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A2_M1017_g N_A_449_297#_c_630_n 0.00948336f $X=2.59 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A2_M1018_g N_A_449_297#_c_630_n 0.00943921f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_222 A2 N_A_449_297#_c_630_n 0.0763505f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_223 N_A2_c_216_n N_A_449_297#_c_630_n 4.60517e-19 $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A2_M1027_g N_A_449_297#_c_634_n 0.0195317f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A2_c_216_n N_A_449_297#_c_634_n 4.9805e-19 $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A2_M1027_g N_Y_c_671_n 0.00614957f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A2_M1016_g N_A_31_47#_c_767_n 0.00620543f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A2_M1021_g N_A_31_47#_c_767_n 5.19281e-19 $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A2_M1016_g N_A_31_47#_c_776_n 0.00844123f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A2_M1021_g N_A_31_47#_c_776_n 0.00844123f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_231 A2 N_A_31_47#_c_776_n 0.0332055f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_232 N_A2_c_216_n N_A_31_47#_c_776_n 0.0020061f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A2_M1016_g N_A_31_47#_c_780_n 5.19281e-19 $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A2_M1021_g N_A_31_47#_c_780_n 0.00620543f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_235 N_A2_M1023_g N_A_31_47#_c_780_n 0.00620543f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_236 N_A2_M1029_g N_A_31_47#_c_780_n 5.19281e-19 $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A2_M1023_g N_A_31_47#_c_784_n 0.00844123f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A2_M1029_g N_A_31_47#_c_784_n 0.00844123f $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_239 A2 N_A_31_47#_c_784_n 0.0332055f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_240 N_A2_c_216_n N_A_31_47#_c_784_n 0.0020061f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A2_M1023_g N_A_31_47#_c_788_n 5.19281e-19 $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_242 N_A2_M1029_g N_A_31_47#_c_788_n 0.00620543f $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_243 N_A2_M1016_g N_A_31_47#_c_747_n 8.68782e-19 $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_244 A2 N_A_31_47#_c_747_n 0.0124322f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_245 N_A2_M1021_g N_A_31_47#_c_748_n 8.68782e-19 $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A2_M1023_g N_A_31_47#_c_748_n 8.68782e-19 $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_247 A2 N_A_31_47#_c_748_n 0.0219994f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_248 N_A2_c_216_n N_A_31_47#_c_748_n 0.00208088f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A2_M1029_g N_A_31_47#_c_749_n 8.68782e-19 $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_250 A2 N_A_31_47#_c_749_n 0.00852101f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_251 N_A2_M1016_g N_VGND_c_884_n 0.00146448f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A2_M1021_g N_VGND_c_884_n 0.00146448f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A2_M1023_g N_VGND_c_885_n 0.00146448f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A2_M1029_g N_VGND_c_885_n 0.00268723f $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A2_M1016_g N_VGND_c_889_n 0.00422241f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A2_M1021_g N_VGND_c_891_n 0.00422241f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_257 N_A2_M1023_g N_VGND_c_891_n 0.00422241f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A2_M1016_g N_VGND_c_895_n 0.00572376f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A2_M1021_g N_VGND_c_895_n 0.00569656f $X=2.59 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A2_M1023_g N_VGND_c_895_n 0.00569656f $X=3.01 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A2_M1029_g N_VGND_c_895_n 0.00572376f $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A2_M1029_g N_VGND_c_897_n 0.00422241f $X=3.43 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A3_M1024_g N_B1_M1003_g 0.0178641f $X=5.645 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A3_M1030_g N_B1_M1000_g 0.0178641f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_265 A3 N_B1_c_384_n 0.00213713f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_266 N_A3_c_310_n N_B1_c_384_n 0.0178641f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A3_M1004_g N_A_27_297#_c_451_n 0.00124004f $X=4.385 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A3_M1030_g N_VPWR_c_525_n 0.00126924f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A3_M1004_g N_VPWR_c_528_n 0.00357877f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A3_M1009_g N_VPWR_c_528_n 0.00357877f $X=4.805 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A3_M1028_g N_VPWR_c_528_n 0.00357877f $X=5.225 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A3_M1030_g N_VPWR_c_528_n 0.00539883f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A3_M1004_g N_VPWR_c_522_n 0.00660224f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A3_M1009_g N_VPWR_c_522_n 0.00522516f $X=4.805 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A3_M1028_g N_VPWR_c_522_n 0.00522516f $X=5.225 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A3_M1030_g N_VPWR_c_522_n 0.00961456f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A3_M1004_g N_A_449_297#_c_627_n 0.0240277f $X=4.385 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_A3_M1009_g N_A_449_297#_c_637_n 0.0187481f $X=4.805 $Y=1.985 $X2=0
+ $Y2=0
cc_279 N_A3_M1028_g N_A_449_297#_c_637_n 0.0187251f $X=5.225 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A3_M1030_g N_A_449_297#_c_637_n 0.00693298f $X=5.645 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A3_M1024_g Y 8.73151e-19 $X=5.645 $Y=0.56 $X2=0 $Y2=0
cc_282 A3 Y 0.0176835f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_283 N_A3_c_310_n Y 0.00102747f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A3_M1004_g N_Y_c_671_n 0.0113822f $X=4.385 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A3_M1009_g N_Y_c_671_n 0.010955f $X=4.805 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A3_M1028_g N_Y_c_671_n 0.010955f $X=5.225 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A3_M1030_g N_Y_c_671_n 0.0147921f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A3_c_307_n N_Y_c_671_n 0.0130423f $X=3.925 $Y=1.16 $X2=0 $Y2=0
cc_289 A3 N_Y_c_671_n 0.161122f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_290 N_A3_c_310_n N_Y_c_671_n 0.00689602f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A3_M1001_g N_A_31_47#_c_788_n 0.0109965f $X=3.85 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A3_M1001_g N_A_31_47#_c_799_n 0.0100251f $X=3.85 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A3_M1002_g N_A_31_47#_c_799_n 0.0128368f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_294 A3 N_A_31_47#_c_799_n 0.0652189f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_295 N_A3_c_309_n N_A_31_47#_c_799_n 0.0122875f $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A3_M1013_g N_A_31_47#_c_743_n 0.0118876f $X=5.105 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A3_M1024_g N_A_31_47#_c_743_n 0.0115218f $X=5.645 $Y=0.56 $X2=0 $Y2=0
cc_298 A3 N_A_31_47#_c_743_n 0.0618476f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_299 N_A3_c_310_n N_A_31_47#_c_743_n 0.00528149f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A3_M1001_g N_A_31_47#_c_749_n 8.68782e-19 $X=3.85 $Y=0.56 $X2=0 $Y2=0
cc_301 A3 N_A_31_47#_c_749_n 0.00227082f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_302 A3 N_A_31_47#_c_750_n 0.012692f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_303 N_A3_c_310_n N_A_31_47#_c_750_n 0.00251608f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A3_M1002_g N_VGND_c_886_n 8.82328e-19 $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A3_M1013_g N_VGND_c_886_n 0.00894326f $X=5.105 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A3_M1024_g N_VGND_c_886_n 0.0091746f $X=5.645 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A3_M1002_g N_VGND_c_893_n 0.00348405f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A3_M1013_g N_VGND_c_893_n 0.00348405f $X=5.105 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A3_M1024_g N_VGND_c_894_n 0.00348405f $X=5.645 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A3_M1001_g N_VGND_c_895_n 0.00660658f $X=3.85 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A3_M1002_g N_VGND_c_895_n 0.00412863f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_312 N_A3_M1013_g N_VGND_c_895_n 0.00414556f $X=5.105 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A3_M1024_g N_VGND_c_895_n 0.00417382f $X=5.645 $Y=0.56 $X2=0 $Y2=0
cc_314 N_A3_M1001_g N_VGND_c_897_n 0.00422241f $X=3.85 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A3_M1001_g N_VGND_c_898_n 0.00771502f $X=3.85 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A3_M1002_g N_VGND_c_898_n 0.0095917f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A3_M1013_g N_VGND_c_898_n 8.9098e-19 $X=5.105 $Y=0.56 $X2=0 $Y2=0
cc_318 N_B1_M1000_g N_VPWR_c_525_n 0.0116829f $X=6.065 $Y=1.985 $X2=0 $Y2=0
cc_319 N_B1_M1010_g N_VPWR_c_525_n 0.0104849f $X=6.485 $Y=1.985 $X2=0 $Y2=0
cc_320 N_B1_M1015_g N_VPWR_c_525_n 6.16378e-19 $X=6.905 $Y=1.985 $X2=0 $Y2=0
cc_321 N_B1_M1010_g N_VPWR_c_526_n 6.16378e-19 $X=6.485 $Y=1.985 $X2=0 $Y2=0
cc_322 N_B1_M1015_g N_VPWR_c_526_n 0.0104849f $X=6.905 $Y=1.985 $X2=0 $Y2=0
cc_323 N_B1_M1025_g N_VPWR_c_526_n 0.0123946f $X=7.325 $Y=1.985 $X2=0 $Y2=0
cc_324 N_B1_M1000_g N_VPWR_c_528_n 0.0046653f $X=6.065 $Y=1.985 $X2=0 $Y2=0
cc_325 N_B1_M1010_g N_VPWR_c_529_n 0.0046653f $X=6.485 $Y=1.985 $X2=0 $Y2=0
cc_326 N_B1_M1015_g N_VPWR_c_529_n 0.0046653f $X=6.905 $Y=1.985 $X2=0 $Y2=0
cc_327 N_B1_M1025_g N_VPWR_c_530_n 0.0046653f $X=7.325 $Y=1.985 $X2=0 $Y2=0
cc_328 N_B1_M1000_g N_VPWR_c_522_n 0.007919f $X=6.065 $Y=1.985 $X2=0 $Y2=0
cc_329 N_B1_M1010_g N_VPWR_c_522_n 0.00789179f $X=6.485 $Y=1.985 $X2=0 $Y2=0
cc_330 N_B1_M1015_g N_VPWR_c_522_n 0.00789179f $X=6.905 $Y=1.985 $X2=0 $Y2=0
cc_331 N_B1_M1025_g N_VPWR_c_522_n 0.00898263f $X=7.325 $Y=1.985 $X2=0 $Y2=0
cc_332 N_B1_M1003_g Y 0.0034277f $X=6.065 $Y=0.56 $X2=0 $Y2=0
cc_333 N_B1_M1000_g Y 0.00379235f $X=6.065 $Y=1.985 $X2=0 $Y2=0
cc_334 N_B1_M1006_g Y 0.00310643f $X=6.485 $Y=0.56 $X2=0 $Y2=0
cc_335 N_B1_M1010_g Y 0.00335255f $X=6.485 $Y=1.985 $X2=0 $Y2=0
cc_336 B1 Y 0.0167034f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_337 N_B1_c_384_n Y 0.014897f $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_338 N_B1_M1000_g Y 0.0184526f $X=6.065 $Y=1.985 $X2=0 $Y2=0
cc_339 N_B1_c_384_n Y 3.37401e-19 $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_340 B1 Y 0.0139517f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_341 N_B1_c_384_n Y 0.00206439f $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_342 N_B1_M1003_g N_Y_c_696_n 0.00291048f $X=6.065 $Y=0.56 $X2=0 $Y2=0
cc_343 N_B1_M1010_g N_Y_c_672_n 0.0155081f $X=6.485 $Y=1.985 $X2=0 $Y2=0
cc_344 B1 N_Y_c_672_n 0.0104851f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_345 N_B1_c_384_n N_Y_c_672_n 6.82014e-19 $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_346 N_B1_M1015_g N_Y_c_673_n 0.0148631f $X=6.905 $Y=1.985 $X2=0 $Y2=0
cc_347 N_B1_M1025_g N_Y_c_673_n 0.0154359f $X=7.325 $Y=1.985 $X2=0 $Y2=0
cc_348 B1 N_Y_c_673_n 0.0491008f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_349 N_B1_c_384_n N_Y_c_673_n 0.00311113f $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_350 B1 N_Y_c_674_n 0.0244039f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_351 N_B1_c_384_n N_Y_c_674_n 5.73441e-19 $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_352 N_B1_M1006_g N_Y_c_706_n 0.0108467f $X=6.485 $Y=0.56 $X2=0 $Y2=0
cc_353 N_B1_M1011_g N_Y_c_706_n 0.0102121f $X=6.905 $Y=0.56 $X2=0 $Y2=0
cc_354 N_B1_M1014_g N_Y_c_706_n 0.00342854f $X=7.325 $Y=0.56 $X2=0 $Y2=0
cc_355 B1 N_Y_c_706_n 0.0504243f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_356 N_B1_c_384_n N_Y_c_706_n 0.00471612f $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_357 N_B1_M1003_g N_A_31_47#_c_811_n 0.0136727f $X=6.065 $Y=0.56 $X2=0 $Y2=0
cc_358 N_B1_M1006_g N_A_31_47#_c_811_n 0.00886996f $X=6.485 $Y=0.56 $X2=0 $Y2=0
cc_359 N_B1_M1011_g N_A_31_47#_c_811_n 0.00892725f $X=6.905 $Y=0.56 $X2=0 $Y2=0
cc_360 N_B1_M1014_g N_A_31_47#_c_811_n 0.010509f $X=7.325 $Y=0.56 $X2=0 $Y2=0
cc_361 B1 N_A_31_47#_c_811_n 0.00370419f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_362 N_B1_c_384_n N_A_31_47#_c_811_n 2.51808e-19 $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_363 B1 N_A_31_47#_c_745_n 0.0234549f $X=7.505 $Y=1.105 $X2=0 $Y2=0
cc_364 N_B1_c_384_n N_A_31_47#_c_745_n 5.36066e-19 $X=7.325 $Y=1.16 $X2=0 $Y2=0
cc_365 N_B1_M1003_g N_VGND_c_886_n 0.0012797f $X=6.065 $Y=0.56 $X2=0 $Y2=0
cc_366 N_B1_M1003_g N_VGND_c_894_n 0.00357877f $X=6.065 $Y=0.56 $X2=0 $Y2=0
cc_367 N_B1_M1006_g N_VGND_c_894_n 0.00357877f $X=6.485 $Y=0.56 $X2=0 $Y2=0
cc_368 N_B1_M1011_g N_VGND_c_894_n 0.00357877f $X=6.905 $Y=0.56 $X2=0 $Y2=0
cc_369 N_B1_M1014_g N_VGND_c_894_n 0.00357877f $X=7.325 $Y=0.56 $X2=0 $Y2=0
cc_370 N_B1_M1003_g N_VGND_c_895_n 0.0052923f $X=6.065 $Y=0.56 $X2=0 $Y2=0
cc_371 N_B1_M1006_g N_VGND_c_895_n 0.00522516f $X=6.485 $Y=0.56 $X2=0 $Y2=0
cc_372 N_B1_M1011_g N_VGND_c_895_n 0.00522516f $X=6.905 $Y=0.56 $X2=0 $Y2=0
cc_373 N_B1_M1014_g N_VGND_c_895_n 0.00620254f $X=7.325 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A_27_297#_c_456_n N_VPWR_M1007_d 0.00318475f $X=0.955 $Y=1.745
+ $X2=-0.19 $Y2=1.305
cc_375 N_A_27_297#_c_464_n N_VPWR_M1026_d 0.00318475f $X=1.795 $Y=1.745 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_456_n N_VPWR_c_523_n 0.0128823f $X=0.955 $Y=1.745 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_c_464_n N_VPWR_c_524_n 0.0128823f $X=1.795 $Y=1.745 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_460_n N_VPWR_c_527_n 0.0189039f $X=1.12 $Y=2.36 $X2=0 $Y2=0
cc_379 N_A_27_297#_c_469_n N_VPWR_c_528_n 0.0190403f $X=1.96 $Y=2.205 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_c_479_n N_VPWR_c_528_n 0.0293587f $X=2.635 $Y=2.335 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_451_n N_VPWR_c_528_n 0.0544531f $X=3.64 $Y=2.36 $X2=0 $Y2=0
cc_382 N_A_27_297#_c_483_n N_VPWR_c_528_n 0.0186386f $X=2.8 $Y=2.02 $X2=0 $Y2=0
cc_383 N_A_27_297#_M1007_s N_VPWR_c_522_n 0.00225715f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_M1022_s N_VPWR_c_522_n 0.00215201f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_M1031_s N_VPWR_c_522_n 0.00215201f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_M1017_d N_VPWR_c_522_n 0.00215201f $X=2.665 $Y=1.485 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_M1027_d N_VPWR_c_522_n 0.00225742f $X=3.505 $Y=1.485 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_450_n N_VPWR_c_522_n 0.0133896f $X=0.28 $Y=2.36 $X2=0 $Y2=0
cc_389 N_A_27_297#_c_456_n N_VPWR_c_522_n 0.0111533f $X=0.955 $Y=1.745 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_460_n N_VPWR_c_522_n 0.0122217f $X=1.12 $Y=2.36 $X2=0 $Y2=0
cc_391 N_A_27_297#_c_464_n N_VPWR_c_522_n 0.0111533f $X=1.795 $Y=1.745 $X2=0
+ $Y2=0
cc_392 N_A_27_297#_c_469_n N_VPWR_c_522_n 0.0122896f $X=1.96 $Y=2.205 $X2=0
+ $Y2=0
cc_393 N_A_27_297#_c_479_n N_VPWR_c_522_n 0.0180744f $X=2.635 $Y=2.335 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_451_n N_VPWR_c_522_n 0.033284f $X=3.64 $Y=2.36 $X2=0 $Y2=0
cc_395 N_A_27_297#_c_483_n N_VPWR_c_522_n 0.0121417f $X=2.8 $Y=2.02 $X2=0 $Y2=0
cc_396 N_A_27_297#_c_450_n N_VPWR_c_532_n 0.022803f $X=0.28 $Y=2.36 $X2=0 $Y2=0
cc_397 N_A_27_297#_c_479_n N_A_449_297#_M1005_s 0.00316464f $X=2.635 $Y=2.335
+ $X2=-0.19 $Y2=1.305
cc_398 N_A_27_297#_c_451_n N_A_449_297#_M1018_s 0.00316874f $X=3.64 $Y=2.36
+ $X2=0 $Y2=0
cc_399 N_A_27_297#_c_451_n N_A_449_297#_c_627_n 0.0214559f $X=3.64 $Y=2.36 $X2=0
+ $Y2=0
cc_400 N_A_27_297#_c_479_n N_A_449_297#_c_628_n 0.0120693f $X=2.635 $Y=2.335
+ $X2=0 $Y2=0
cc_401 N_A_27_297#_M1017_d N_A_449_297#_c_630_n 0.00315327f $X=2.665 $Y=1.485
+ $X2=0 $Y2=0
cc_402 N_A_27_297#_c_479_n N_A_449_297#_c_630_n 0.00387899f $X=2.635 $Y=2.335
+ $X2=0 $Y2=0
cc_403 N_A_27_297#_c_451_n N_A_449_297#_c_630_n 0.00387899f $X=3.64 $Y=2.36
+ $X2=0 $Y2=0
cc_404 N_A_27_297#_c_483_n N_A_449_297#_c_630_n 0.016684f $X=2.8 $Y=2.02 $X2=0
+ $Y2=0
cc_405 N_A_27_297#_M1027_d N_A_449_297#_c_634_n 0.00953274f $X=3.505 $Y=1.485
+ $X2=0 $Y2=0
cc_406 N_A_27_297#_c_451_n N_A_449_297#_c_634_n 0.0464827f $X=3.64 $Y=2.36 $X2=0
+ $Y2=0
cc_407 N_A_27_297#_M1027_d N_A_449_297#_c_626_n 0.00787651f $X=3.505 $Y=1.485
+ $X2=0 $Y2=0
cc_408 N_VPWR_c_522_n N_A_449_297#_M1005_s 0.00216833f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_409 N_VPWR_c_522_n N_A_449_297#_M1018_s 0.00216833f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_522_n N_A_449_297#_M1004_s 0.00215227f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_522_n N_A_449_297#_M1028_s 0.00215227f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_528_n N_A_449_297#_c_627_n 0.0904953f $X=6.11 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_522_n N_A_449_297#_c_627_n 0.0558197f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_522_n N_A_449_297#_c_634_n 0.00676535f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_528_n N_A_449_297#_c_626_n 0.00318833f $X=6.11 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_522_n N_Y_M1004_d 0.0021699f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_522_n N_Y_M1009_d 0.00216833f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_522_n N_Y_M1030_d 0.00562358f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_419 N_VPWR_c_522_n N_Y_M1010_d 0.00562358f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_c_522_n N_Y_M1025_d 0.00387172f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_421 N_VPWR_c_528_n N_Y_c_716_n 0.0113958f $X=6.11 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_c_522_n N_Y_c_716_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_c_529_n N_Y_c_718_n 0.0113958f $X=6.95 $Y=2.72 $X2=0 $Y2=0
cc_424 N_VPWR_c_522_n N_Y_c_718_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_425 N_VPWR_M1000_s Y 0.0011179f $X=6.14 $Y=1.485 $X2=0 $Y2=0
cc_426 N_VPWR_c_525_n Y 0.0157164f $X=6.275 $Y=2.02 $X2=0 $Y2=0
cc_427 N_VPWR_c_530_n Y 0.0197934f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_522_n Y 0.0108988f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_429 N_VPWR_M1000_s N_Y_c_672_n 6.50204e-19 $X=6.14 $Y=1.485 $X2=0 $Y2=0
cc_430 N_VPWR_M1015_s N_Y_c_673_n 0.00177951f $X=6.98 $Y=1.485 $X2=0 $Y2=0
cc_431 N_VPWR_c_526_n N_Y_c_673_n 0.0157512f $X=7.115 $Y=2.02 $X2=0 $Y2=0
cc_432 N_A_449_297#_c_627_n N_Y_M1004_d 0.0111427f $X=4.68 $Y=2.165 $X2=0 $Y2=0
cc_433 N_A_449_297#_c_626_n N_Y_M1004_d 8.97565e-19 $X=4.08 $Y=2.165 $X2=0 $Y2=0
cc_434 N_A_449_297#_c_637_n N_Y_M1009_d 0.00315858f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_435 N_A_449_297#_M1004_s N_Y_c_671_n 0.00168223f $X=4.46 $Y=1.485 $X2=0 $Y2=0
cc_436 N_A_449_297#_M1028_s N_Y_c_671_n 0.00168223f $X=5.3 $Y=1.485 $X2=0 $Y2=0
cc_437 N_A_449_297#_c_634_n N_Y_c_671_n 0.00900821f $X=3.605 $Y=1.815 $X2=0
+ $Y2=0
cc_438 N_A_449_297#_c_626_n N_Y_c_671_n 0.112957f $X=4.08 $Y=2.165 $X2=0 $Y2=0
cc_439 N_Y_c_706_n N_A_31_47#_M1006_d 0.00308407f $X=7.115 $Y=0.76 $X2=0 $Y2=0
cc_440 N_Y_M1003_s N_A_31_47#_c_811_n 0.00304594f $X=6.14 $Y=0.235 $X2=0 $Y2=0
cc_441 N_Y_M1011_s N_A_31_47#_c_811_n 0.00305792f $X=6.98 $Y=0.235 $X2=0 $Y2=0
cc_442 N_Y_c_696_n N_A_31_47#_c_811_n 0.0098496f $X=6.202 $Y=0.885 $X2=0 $Y2=0
cc_443 N_Y_c_706_n N_A_31_47#_c_811_n 0.0487838f $X=7.115 $Y=0.76 $X2=0 $Y2=0
cc_444 N_Y_M1003_s N_VGND_c_895_n 0.00216833f $X=6.14 $Y=0.235 $X2=0 $Y2=0
cc_445 N_Y_M1011_s N_VGND_c_895_n 0.00216833f $X=6.98 $Y=0.235 $X2=0 $Y2=0
cc_446 N_A_31_47#_c_753_n N_VGND_M1008_d 0.00306532f $X=0.955 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_447 N_A_31_47#_c_763_n N_VGND_M1019_d 0.00306532f $X=1.795 $Y=0.8 $X2=0 $Y2=0
cc_448 N_A_31_47#_c_776_n N_VGND_M1016_s 0.00306532f $X=2.635 $Y=0.8 $X2=0 $Y2=0
cc_449 N_A_31_47#_c_784_n N_VGND_M1023_s 0.00306532f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_450 N_A_31_47#_c_799_n N_VGND_M1001_s 0.0138087f $X=4.81 $Y=0.8 $X2=0 $Y2=0
cc_451 N_A_31_47#_c_743_n N_VGND_M1013_s 0.00556882f $X=5.77 $Y=0.8 $X2=0 $Y2=0
cc_452 N_A_31_47#_c_753_n N_VGND_c_882_n 0.012179f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_453 N_A_31_47#_c_763_n N_VGND_c_883_n 0.012179f $X=1.795 $Y=0.8 $X2=0 $Y2=0
cc_454 N_A_31_47#_c_776_n N_VGND_c_884_n 0.012179f $X=2.635 $Y=0.8 $X2=0 $Y2=0
cc_455 N_A_31_47#_c_784_n N_VGND_c_885_n 0.012179f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_456 N_A_31_47#_c_743_n N_VGND_c_886_n 0.0257035f $X=5.77 $Y=0.8 $X2=0 $Y2=0
cc_457 N_A_31_47#_c_753_n N_VGND_c_887_n 0.0020257f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_458 N_A_31_47#_c_759_n N_VGND_c_887_n 0.0188215f $X=1.12 $Y=0.36 $X2=0 $Y2=0
cc_459 N_A_31_47#_c_763_n N_VGND_c_887_n 0.0020257f $X=1.795 $Y=0.8 $X2=0 $Y2=0
cc_460 N_A_31_47#_c_763_n N_VGND_c_889_n 0.0020257f $X=1.795 $Y=0.8 $X2=0 $Y2=0
cc_461 N_A_31_47#_c_767_n N_VGND_c_889_n 0.0188215f $X=1.96 $Y=0.36 $X2=0 $Y2=0
cc_462 N_A_31_47#_c_776_n N_VGND_c_889_n 0.0020257f $X=2.635 $Y=0.8 $X2=0 $Y2=0
cc_463 N_A_31_47#_c_776_n N_VGND_c_891_n 0.0020257f $X=2.635 $Y=0.8 $X2=0 $Y2=0
cc_464 N_A_31_47#_c_780_n N_VGND_c_891_n 0.0188215f $X=2.8 $Y=0.36 $X2=0 $Y2=0
cc_465 N_A_31_47#_c_784_n N_VGND_c_891_n 0.0020257f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_466 N_A_31_47#_c_799_n N_VGND_c_893_n 0.0020257f $X=4.81 $Y=0.8 $X2=0 $Y2=0
cc_467 N_A_31_47#_c_845_p N_VGND_c_893_n 0.00583301f $X=4.895 $Y=0.56 $X2=0
+ $Y2=0
cc_468 N_A_31_47#_c_743_n N_VGND_c_893_n 0.0020257f $X=5.77 $Y=0.8 $X2=0 $Y2=0
cc_469 N_A_31_47#_c_743_n N_VGND_c_894_n 0.0020257f $X=5.77 $Y=0.8 $X2=0 $Y2=0
cc_470 N_A_31_47#_c_811_n N_VGND_c_894_n 0.0832396f $X=7.45 $Y=0.365 $X2=0 $Y2=0
cc_471 N_A_31_47#_c_849_p N_VGND_c_894_n 0.0114055f $X=5.94 $Y=0.365 $X2=0 $Y2=0
cc_472 N_A_31_47#_c_744_n N_VGND_c_894_n 0.0197903f $X=7.592 $Y=0.475 $X2=0
+ $Y2=0
cc_473 N_A_31_47#_M1008_s N_VGND_c_895_n 0.00209319f $X=0.155 $Y=0.235 $X2=0
+ $Y2=0
cc_474 N_A_31_47#_M1012_s N_VGND_c_895_n 0.00215201f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_475 N_A_31_47#_M1020_s N_VGND_c_895_n 0.00215201f $X=1.825 $Y=0.235 $X2=0
+ $Y2=0
cc_476 N_A_31_47#_M1021_d N_VGND_c_895_n 0.00215201f $X=2.665 $Y=0.235 $X2=0
+ $Y2=0
cc_477 N_A_31_47#_M1029_d N_VGND_c_895_n 0.00215201f $X=3.505 $Y=0.235 $X2=0
+ $Y2=0
cc_478 N_A_31_47#_M1002_d N_VGND_c_895_n 0.00275192f $X=4.76 $Y=0.235 $X2=0
+ $Y2=0
cc_479 N_A_31_47#_M1024_d N_VGND_c_895_n 0.00240924f $X=5.72 $Y=0.235 $X2=0
+ $Y2=0
cc_480 N_A_31_47#_M1006_d N_VGND_c_895_n 0.00215227f $X=6.56 $Y=0.235 $X2=0
+ $Y2=0
cc_481 N_A_31_47#_M1014_d N_VGND_c_895_n 0.00209324f $X=7.4 $Y=0.235 $X2=0 $Y2=0
cc_482 N_A_31_47#_c_741_n N_VGND_c_895_n 0.0133626f $X=0.28 $Y=0.38 $X2=0 $Y2=0
cc_483 N_A_31_47#_c_753_n N_VGND_c_895_n 0.00841425f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_484 N_A_31_47#_c_759_n N_VGND_c_895_n 0.0121968f $X=1.12 $Y=0.36 $X2=0 $Y2=0
cc_485 N_A_31_47#_c_763_n N_VGND_c_895_n 0.00841425f $X=1.795 $Y=0.8 $X2=0 $Y2=0
cc_486 N_A_31_47#_c_767_n N_VGND_c_895_n 0.0121968f $X=1.96 $Y=0.36 $X2=0 $Y2=0
cc_487 N_A_31_47#_c_776_n N_VGND_c_895_n 0.00841425f $X=2.635 $Y=0.8 $X2=0 $Y2=0
cc_488 N_A_31_47#_c_780_n N_VGND_c_895_n 0.0121968f $X=2.8 $Y=0.36 $X2=0 $Y2=0
cc_489 N_A_31_47#_c_784_n N_VGND_c_895_n 0.00841425f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_490 N_A_31_47#_c_788_n N_VGND_c_895_n 0.0121968f $X=3.64 $Y=0.36 $X2=0 $Y2=0
cc_491 N_A_31_47#_c_799_n N_VGND_c_895_n 0.0108606f $X=4.81 $Y=0.8 $X2=0 $Y2=0
cc_492 N_A_31_47#_c_845_p N_VGND_c_895_n 0.00590828f $X=4.895 $Y=0.56 $X2=0
+ $Y2=0
cc_493 N_A_31_47#_c_743_n N_VGND_c_895_n 0.00960173f $X=5.77 $Y=0.8 $X2=0 $Y2=0
cc_494 N_A_31_47#_c_811_n N_VGND_c_895_n 0.0536017f $X=7.45 $Y=0.365 $X2=0 $Y2=0
cc_495 N_A_31_47#_c_849_p N_VGND_c_895_n 0.0065339f $X=5.94 $Y=0.365 $X2=0 $Y2=0
cc_496 N_A_31_47#_c_744_n N_VGND_c_895_n 0.010954f $X=7.592 $Y=0.475 $X2=0 $Y2=0
cc_497 N_A_31_47#_c_741_n N_VGND_c_896_n 0.0227138f $X=0.28 $Y=0.38 $X2=0 $Y2=0
cc_498 N_A_31_47#_c_753_n N_VGND_c_896_n 0.0020257f $X=0.955 $Y=0.8 $X2=0 $Y2=0
cc_499 N_A_31_47#_c_784_n N_VGND_c_897_n 0.0020257f $X=3.475 $Y=0.8 $X2=0 $Y2=0
cc_500 N_A_31_47#_c_788_n N_VGND_c_897_n 0.0188215f $X=3.64 $Y=0.36 $X2=0 $Y2=0
cc_501 N_A_31_47#_c_799_n N_VGND_c_897_n 0.00227347f $X=4.81 $Y=0.8 $X2=0 $Y2=0
cc_502 N_A_31_47#_c_788_n N_VGND_c_898_n 0.0218042f $X=3.64 $Y=0.36 $X2=0 $Y2=0
cc_503 N_A_31_47#_c_799_n N_VGND_c_898_n 0.0454767f $X=4.81 $Y=0.8 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__ha_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.055000 4.045000 1.225000 ;
        RECT 3.820000 1.225000 4.045000 1.675000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.310000 1.005000 2.615000 1.395000 ;
        RECT 2.310000 1.395000 3.595000 1.675000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 0.315000 4.965000 0.825000 ;
        RECT 4.715000 1.545000 4.965000 2.415000 ;
        RECT 4.790000 0.825000 4.965000 1.545000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.315000 0.885000 0.825000 ;
        RECT 0.555000 0.825000 0.780000 1.565000 ;
        RECT 0.555000 1.565000 0.885000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.135000  0.085000 0.375000 0.885000 ;
        RECT 1.055000  0.085000 1.250000 0.885000 ;
        RECT 2.335000  0.085000 2.665000 0.465000 ;
        RECT 4.215000  0.085000 4.465000 0.545000 ;
        RECT 5.145000  0.085000 5.385000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.135000 1.495000 0.375000 2.635000 ;
        RECT 1.055000 1.515000 1.250000 2.635000 ;
        RECT 2.850000 2.205000 3.640000 2.635000 ;
        RECT 4.215000 2.205000 4.545000 2.635000 ;
        RECT 5.145000 1.495000 5.385000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.950000 1.075000 1.590000 1.245000 ;
      RECT 1.420000 0.345000 1.745000 0.675000 ;
      RECT 1.420000 0.675000 1.590000 1.075000 ;
      RECT 1.420000 1.245000 1.590000 2.205000 ;
      RECT 1.420000 2.205000 2.220000 2.375000 ;
      RECT 1.760000 0.995000 1.930000 1.855000 ;
      RECT 1.760000 1.855000 4.465000 2.025000 ;
      RECT 1.995000 0.345000 2.165000 0.635000 ;
      RECT 1.995000 0.635000 3.005000 0.805000 ;
      RECT 2.835000 0.345000 3.005000 0.635000 ;
      RECT 3.460000 0.345000 3.630000 0.715000 ;
      RECT 3.460000 0.715000 4.465000 0.885000 ;
      RECT 3.810000 2.025000 3.980000 2.355000 ;
      RECT 4.295000 0.885000 4.465000 0.995000 ;
      RECT 4.295000 0.995000 4.620000 1.325000 ;
      RECT 4.295000 1.325000 4.465000 1.855000 ;
  END
END sky130_fd_sc_hd__ha_2
END LIBRARY

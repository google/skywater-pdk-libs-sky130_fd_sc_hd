* File: sky130_fd_sc_hd__or4b_4.spice.pex
* Created: Thu Aug 27 14:44:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4B_4%D_N 3 6 8 9 10 15 16 17
r25 15 18 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.395 $Y2=1.325
r26 15 17 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.395 $Y2=0.995
r27 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r28 9 10 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.275 $Y=1.53
+ $X2=0.275 $Y2=1.87
r29 8 9 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.275 $Y=1.19
+ $X2=0.275 $Y2=1.53
r30 8 16 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=0.275 $Y=1.19 $X2=0.275
+ $Y2=1.16
r31 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r32 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%A_109_93# 1 2 7 9 12 14 15 16 19 21 26 30
r55 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.16 $X2=1.13 $Y2=1.16
r56 26 28 14.0643 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=0.7 $Y=1.067
+ $X2=1.13 $Y2=1.067
r57 25 26 0.327078 $w=3.73e-07 $l=1e-08 $layer=LI1_cond $X=0.69 $Y=1.067 $X2=0.7
+ $Y2=1.067
r58 23 26 5.35566 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=0.7 $Y=1.325 $X2=0.7
+ $Y2=1.067
r59 23 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.7 $Y=1.325 $X2=0.7
+ $Y2=2.065
r60 19 30 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.69 $Y=2.16
+ $X2=0.69 $Y2=2.065
r61 19 21 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=0.69 $Y=2.16
+ $X2=0.69 $Y2=2.275
r62 16 25 4.6906 $w=1.9e-07 $l=2.57e-07 $layer=LI1_cond $X=0.69 $Y=0.81 $X2=0.69
+ $Y2=1.067
r63 16 18 4.49474 $w=1.9e-07 $l=7e-08 $layer=LI1_cond $X=0.69 $Y=0.81 $X2=0.69
+ $Y2=0.74
r64 14 29 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.13 $Y2=1.16
r65 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.41 $Y2=1.16
r66 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r67 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.985
r68 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r69 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
r70 2 21 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.275
r71 1 18 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%C 3 6 10 11 13 14 19 23
r48 21 23 2.24086 $w=3.58e-07 $l=7e-08 $layer=LI1_cond $X=1.975 $Y=1.8 $X2=1.975
+ $Y2=1.87
r49 13 21 0.256098 $w=3.58e-07 $l=8e-09 $layer=LI1_cond $X=1.975 $Y=1.792
+ $X2=1.975 $Y2=1.8
r50 13 29 8.73511 $w=3.58e-07 $l=1.72e-07 $layer=LI1_cond $X=1.975 $Y=1.792
+ $X2=1.975 $Y2=1.62
r51 13 14 10.6601 $w=3.58e-07 $l=3.33e-07 $layer=LI1_cond $X=1.975 $Y=1.877
+ $X2=1.975 $Y2=2.21
r52 13 23 0.224086 $w=3.58e-07 $l=7e-09 $layer=LI1_cond $X=1.975 $Y=1.877
+ $X2=1.975 $Y2=1.87
r53 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.88 $Y2=1.325
r54 11 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.88 $Y2=0.995
r55 10 29 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.88 $Y=1.16
+ $X2=1.88 $Y2=1.62
r56 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r57 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.94 $Y=1.985
+ $X2=1.94 $Y2=1.325
r58 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.94 $Y=0.56 $X2=1.94
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%B 1 3 6 10 11 14 15 31
c40 11 0 5.72837e-20 $X=2.36 $Y=1.16
c41 6 0 2.99791e-19 $X=2.36 $Y=1.985
r42 21 31 2.49696 $w=2.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.485 $Y=1.935
+ $X2=2.485 $Y2=1.87
r43 14 31 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=2.485 $Y=1.86
+ $X2=2.485 $Y2=1.87
r44 14 15 10.1799 $w=2.98e-07 $l=2.65e-07 $layer=LI1_cond $X=2.485 $Y=1.945
+ $X2=2.485 $Y2=2.21
r45 14 21 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=2.485 $Y=1.945
+ $X2=2.485 $Y2=1.935
r46 13 14 15.3247 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.43 $Y=1.45
+ $X2=2.43 $Y2=1.785
r47 10 13 12.1843 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.36 $Y=1.16
+ $X2=2.36 $Y2=1.45
r48 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r49 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.325
+ $X2=2.36 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.36 $Y=1.325 $X2=2.36
+ $Y2=1.985
r51 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=0.995
+ $X2=2.36 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.36 $Y=0.995 $X2=2.36
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%A 3 6 8 12 13 14
c41 13 0 1.24234e-19 $X=2.84 $Y=1.16
c42 8 0 1.75557e-19 $X=2.99 $Y=1.53
r43 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.16
+ $X2=2.84 $Y2=1.325
r44 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.16
+ $X2=2.84 $Y2=0.995
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.16 $X2=2.84 $Y2=1.16
r46 8 20 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.99 $Y=1.53 $X2=2.84
+ $Y2=1.53
r47 8 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=1.445
+ $X2=2.84 $Y2=1.53
r48 8 13 16.7846 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.84 $Y=1.445
+ $X2=2.84 $Y2=1.16
r49 6 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.78 $Y=1.985
+ $X2=2.78 $Y2=1.325
r50 3 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.78 $Y=0.56 $X2=2.78
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%A_215_297# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 40 43 46 48 49 52 54 57 58 63 69 74 81
c144 74 0 5.72837e-20 $X=2.57 $Y=0.74
c145 54 0 1.60701e-19 $X=3.095 $Y=0.74
r146 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.73 $Y=1.16
+ $X2=4.15 $Y2=1.16
r147 71 73 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=0.74
+ $X2=1.7 $Y2=0.74
r148 67 69 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.2 $Y=1.66
+ $X2=1.54 $Y2=1.66
r149 64 81 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.39 $Y=1.16
+ $X2=4.57 $Y2=1.16
r150 64 79 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.39 $Y=1.16
+ $X2=4.15 $Y2=1.16
r151 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.39
+ $Y=1.16 $X2=4.39 $Y2=1.16
r152 61 78 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.37 $Y=1.16
+ $X2=3.73 $Y2=1.16
r153 61 75 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.37 $Y=1.16 $X2=3.31
+ $Y2=1.16
r154 60 63 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.37 $Y=1.16
+ $X2=4.39 $Y2=1.16
r155 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.37
+ $Y=1.16 $X2=3.37 $Y2=1.16
r156 58 60 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.265 $Y=1.16
+ $X2=3.37 $Y2=1.16
r157 57 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.18 $Y=1.075
+ $X2=3.265 $Y2=1.16
r158 56 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.18 $Y=0.825
+ $X2=3.18 $Y2=1.075
r159 55 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=0.74
+ $X2=2.57 $Y2=0.74
r160 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.095 $Y=0.74
+ $X2=3.18 $Y2=0.825
r161 54 55 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.095 $Y=0.74
+ $X2=2.655 $Y2=0.74
r162 50 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0.655
+ $X2=2.57 $Y2=0.74
r163 50 52 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0.655
+ $X2=2.57 $Y2=0.49
r164 49 73 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.74
+ $X2=1.7 $Y2=0.74
r165 48 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=0.74
+ $X2=2.57 $Y2=0.74
r166 48 49 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.485 $Y=0.74
+ $X2=1.785 $Y2=0.74
r167 44 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.655
+ $X2=1.7 $Y2=0.74
r168 44 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=0.655
+ $X2=1.7 $Y2=0.49
r169 43 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.575
+ $X2=1.54 $Y2=1.66
r170 42 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.825
+ $X2=1.54 $Y2=0.74
r171 42 43 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.54 $Y=0.825
+ $X2=1.54 $Y2=1.575
r172 40 67 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.2 $Y=2.34
+ $X2=1.2 $Y2=1.745
r173 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.325
+ $X2=4.57 $Y2=1.16
r174 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.57 $Y=1.325
+ $X2=4.57 $Y2=1.985
r175 31 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=0.995
+ $X2=4.57 $Y2=1.16
r176 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.57 $Y=0.995
+ $X2=4.57 $Y2=0.56
r177 27 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.15 $Y=1.325
+ $X2=4.15 $Y2=1.16
r178 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.15 $Y=1.325
+ $X2=4.15 $Y2=1.985
r179 24 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.15 $Y=0.995
+ $X2=4.15 $Y2=1.16
r180 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.15 $Y=0.995
+ $X2=4.15 $Y2=0.56
r181 20 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.325
+ $X2=3.73 $Y2=1.16
r182 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.73 $Y=1.325
+ $X2=3.73 $Y2=1.985
r183 17 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=0.995
+ $X2=3.73 $Y2=1.16
r184 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.73 $Y=0.995
+ $X2=3.73 $Y2=0.56
r185 13 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.325
+ $X2=3.31 $Y2=1.16
r186 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.31 $Y=1.325
+ $X2=3.31 $Y2=1.985
r187 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.16
r188 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
r189 3 67 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.66
r190 3 40 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.34
r191 2 52 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.235 $X2=2.57 $Y2=0.49
r192 1 46 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.7 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%VPWR 1 2 3 4 13 15 19 23 25 27 29 31 36 41 50
+ 53 57
r65 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r66 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r68 45 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r69 45 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r71 42 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=3.94 $Y2=2.72
r72 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 41 56 3.96406 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=4.857 $Y2=2.72
r74 41 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=4.37 $Y2=2.72
r75 40 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r76 40 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r78 37 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.045 $Y2=2.72
r79 37 39 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.45 $Y2=2.72
r80 36 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.815 $Y=2.72
+ $X2=3.94 $Y2=2.72
r81 36 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.815 $Y=2.72
+ $X2=3.45 $Y2=2.72
r82 35 51 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r84 32 47 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r85 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 31 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.92 $Y=2.72
+ $X2=3.045 $Y2=2.72
r87 31 34 145.487 $w=1.68e-07 $l=2.23e-06 $layer=LI1_cond $X=2.92 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 29 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r90 25 56 3.1791 $w=2.5e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.78 $Y=2.635
+ $X2=4.857 $Y2=2.72
r91 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.78 $Y=2.635
+ $X2=4.78 $Y2=1.96
r92 21 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.94 $Y=2.635
+ $X2=3.94 $Y2=2.72
r93 21 23 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.94 $Y=2.635
+ $X2=3.94 $Y2=1.96
r94 17 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=2.635
+ $X2=3.045 $Y2=2.72
r95 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.045 $Y=2.635
+ $X2=3.045 $Y2=1.96
r96 13 47 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.182 $Y2=2.72
r97 13 15 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.225 $Y2=2.3
r98 4 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.645
+ $Y=1.485 $X2=4.78 $Y2=1.96
r99 3 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.805
+ $Y=1.485 $X2=3.94 $Y2=1.96
r100 2 19 300 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_PDIFF $count=2 $X=2.855
+ $Y=1.485 $X2=3.045 $Y2=1.96
r101 1 15 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%X 1 2 3 4 13 15 19 21 23 24 27 31 33 35 39 41
+ 43 46
r74 43 46 2.99957 $w=2.4e-07 $l=9e-08 $layer=LI1_cond $X=4.845 $Y=0.815
+ $X2=4.845 $Y2=0.905
r75 43 46 0.720277 $w=2.38e-07 $l=1.5e-08 $layer=LI1_cond $X=4.845 $Y=0.92
+ $X2=4.845 $Y2=0.905
r76 42 43 25.6899 $w=2.38e-07 $l=5.35e-07 $layer=LI1_cond $X=4.845 $Y=1.455
+ $X2=4.845 $Y2=0.92
r77 36 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=0.815
+ $X2=4.36 $Y2=0.815
r78 35 43 3.99943 $w=1.8e-07 $l=1.2e-07 $layer=LI1_cond $X=4.725 $Y=0.815
+ $X2=4.845 $Y2=0.815
r79 35 36 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=4.725 $Y=0.815
+ $X2=4.525 $Y2=0.815
r80 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.485 $Y=1.54
+ $X2=4.36 $Y2=1.54
r81 33 42 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=4.725 $Y=1.54
+ $X2=4.845 $Y2=1.455
r82 33 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.725 $Y=1.54
+ $X2=4.485 $Y2=1.54
r83 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=1.625
+ $X2=4.36 $Y2=1.54
r84 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.36 $Y=1.625
+ $X2=4.36 $Y2=2.3
r85 25 39 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.36 $Y=0.725 $X2=4.36
+ $Y2=0.815
r86 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.36 $Y=0.725
+ $X2=4.36 $Y2=0.39
r87 23 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=0.815
+ $X2=4.36 $Y2=0.815
r88 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.195 $Y=0.815
+ $X2=3.685 $Y2=0.815
r89 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.645 $Y=1.54
+ $X2=3.52 $Y2=1.54
r90 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.235 $Y=1.54
+ $X2=4.36 $Y2=1.54
r91 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.235 $Y=1.54
+ $X2=3.645 $Y2=1.54
r92 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=3.56 $Y=0.725
+ $X2=3.685 $Y2=0.815
r93 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=3.56 $Y=0.725
+ $X2=3.56 $Y2=0.485
r94 13 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=1.625
+ $X2=3.52 $Y2=1.54
r95 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.52 $Y=1.625
+ $X2=3.52 $Y2=2.3
r96 4 41 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.225
+ $Y=1.485 $X2=4.36 $Y2=1.62
r97 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.225
+ $Y=1.485 $X2=4.36 $Y2=2.3
r98 3 38 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.485 $X2=3.52 $Y2=1.62
r99 3 15 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.485 $X2=3.52 $Y2=2.3
r100 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.225
+ $Y=0.235 $X2=4.36 $Y2=0.39
r101 1 19 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.235 $X2=3.52 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_4%VGND 1 2 3 4 5 6 19 21 25 29 33 35 39 41 43
+ 45 47 52 57 62 71 74 77 80 84
c94 35 0 1.60701e-19 $X=3.855 $Y=0
r95 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r96 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r97 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r98 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r99 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r100 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r101 66 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r102 66 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r103 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r104 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=0 $X2=3.94
+ $Y2=0
r105 63 65 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=4.37
+ $Y2=0
r106 62 83 3.40825 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=4.877 $Y2=0
r107 62 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=4.37 $Y2=0
r108 61 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r109 61 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r110 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r111 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r112 58 60 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.53 $Y2=0
r113 57 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=3.065
+ $Y2=0
r114 57 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.53
+ $Y2=0
r115 56 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r116 56 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r117 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r118 53 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.16
+ $Y2=0
r119 53 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.61 $Y2=0
r120 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r121 52 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.61 $Y2=0
r122 51 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r123 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r124 48 68 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r125 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r126 47 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.16
+ $Y2=0
r127 47 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r128 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r129 45 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r130 41 83 3.40825 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=4.78 $Y=0.085
+ $X2=4.877 $Y2=0
r131 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.78 $Y=0.085
+ $X2=4.78 $Y2=0.39
r132 37 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.94 $Y=0.085
+ $X2=3.94 $Y2=0
r133 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.94 $Y=0.085
+ $X2=3.94 $Y2=0.39
r134 36 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.065
+ $Y2=0
r135 35 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.94
+ $Y2=0
r136 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.255
+ $Y2=0
r137 31 77 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0
r138 31 33 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0.4
r139 27 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r140 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.4
r141 23 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0
r142 23 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0.38
r143 19 68 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r144 19 21 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.66
r145 6 43 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.645
+ $Y=0.235 $X2=4.78 $Y2=0.39
r146 5 39 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.235 $X2=3.94 $Y2=0.39
r147 4 33 182 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.235 $X2=3.09 $Y2=0.4
r148 3 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.235 $X2=2.15 $Y2=0.4
r149 2 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
r150 1 21 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends


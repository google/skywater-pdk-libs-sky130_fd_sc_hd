* File: sky130_fd_sc_hd__dlxtn_4.spice
* Created: Thu Aug 27 14:18:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlxtn_4.pex.spice"
.subckt sky130_fd_sc_hd__dlxtn_4  VNB VPB GATE_N D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_GATE_N_M1021_g N_A_27_47#_M1021_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_193_47#_M1013_d N_A_27_47#_M1013_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g N_A_299_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 A_465_47# N_A_299_47#_M1010_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0836769 AS=0.0567 PD=0.872308 PS=0.69 NRD=41.208 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1017 N_A_561_413#_M1017_d N_A_27_47#_M1017_g A_465_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0504 AS=0.0717231 PD=0.64 PS=0.747692 NRD=0 NRS=48.072 M=1 R=2.4
+ SA=75001.1 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1008 A_659_47# N_A_193_47#_M1008_g N_A_561_413#_M1017_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0504 PD=0.687692 PS=0.64 NRD=38.076 NRS=0 M=1 R=2.4
+ SA=75001.6 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1018 N_VGND_M1018_d N_A_724_21#_M1018_g A_659_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_561_413#_M1009_g N_A_724_21#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.092625 AS=0.169 PD=0.935 PS=1.82 NRD=1.836 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1009_d N_A_724_21#_M1002_g N_Q_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.08775 PD=0.935 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_724_21#_M1012_g N_Q_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.099125 AS=0.08775 PD=0.955 PS=0.92 NRD=5.532 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1012_d N_A_724_21#_M1019_g N_Q_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.099125 AS=0.09425 PD=0.955 PS=0.94 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_A_724_21#_M1022_g N_Q_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.09425 PD=1.82 PS=0.94 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75001.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_GATE_N_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_VPWR_M1020_d N_D_M1020_g N_A_299_47#_M1020_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1015 A_465_369# N_A_299_47#_M1015_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116891 AS=0.0864 PD=1.17132 PS=0.91 NRD=39.2818 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_561_413#_M1001_d N_A_193_47#_M1001_g A_465_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09555 AS=0.0767094 PD=0.875 PS=0.768679 NRD=56.2829 NRS=59.8683
+ M=1 R=2.8 SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 A_682_413# N_A_27_47#_M1004_g N_A_561_413#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.09555 PD=0.63 PS=0.875 NRD=23.443 NRS=25.7873 M=1 R=2.8
+ SA=75001.7 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_724_21#_M1007_g A_682_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_561_413#_M1006_g N_A_724_21#_M1006_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.1425 AS=0.26 PD=1.285 PS=2.52 NRD=1.9503 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_Q_M1003_d N_A_724_21#_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1425 PD=1.27 PS=1.285 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1014 N_Q_M1003_d N_A_724_21#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1525 PD=1.27 PS=1.305 NRD=0 NRS=5.8903 M=1 R=6.66667 SA=75001
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1016 N_Q_M1016_d N_A_724_21#_M1016_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.1525 PD=1.29 PS=1.305 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1023 N_Q_M1016_d N_A_724_21#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.26 PD=1.29 PS=2.52 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=11.6844 P=17.77
c_144 VPB 0 1.57048e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dlxtn_4.pxi.spice"
*
.ends
*
*

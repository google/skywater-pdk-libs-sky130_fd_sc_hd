* File: sky130_fd_sc_hd__clkinv_16.pxi.spice
* Created: Tue Sep  1 19:01:15 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINV_16%A N_A_M1000_g N_A_M1001_g N_A_M1002_g
+ N_A_M1003_g N_A_M1004_g N_A_M1005_g N_A_M1007_g N_A_M1006_g N_A_M1008_g
+ N_A_M1009_g N_A_M1011_g N_A_M1010_g N_A_M1016_g N_A_M1012_g N_A_M1017_g
+ N_A_M1013_g N_A_M1018_g N_A_M1014_g N_A_c_159_n N_A_c_160_n N_A_M1021_g
+ N_A_M1015_g N_A_M1023_g N_A_M1019_g N_A_M1024_g N_A_M1020_g N_A_M1026_g
+ N_A_M1022_g N_A_M1032_g N_A_M1025_g N_A_M1033_g N_A_M1027_g N_A_M1035_g
+ N_A_M1028_g N_A_M1036_g N_A_M1029_g N_A_M1037_g N_A_M1030_g N_A_M1031_g
+ N_A_M1034_g N_A_M1038_g N_A_M1039_g A N_A_c_285_p N_A_c_286_p N_A_c_294_p
+ N_A_c_360_p N_A_c_371_p N_A_c_171_n N_A_c_172_n
+ PM_SKY130_FD_SC_HD__CLKINV_16%A
x_PM_SKY130_FD_SC_HD__CLKINV_16%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1010_d N_VPWR_M1013_d N_VPWR_M1015_d
+ N_VPWR_M1020_d N_VPWR_M1025_d N_VPWR_M1028_d N_VPWR_M1030_d N_VPWR_M1034_d
+ N_VPWR_M1039_d N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n
+ N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_615_p N_VPWR_c_466_n
+ N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n
+ N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n
+ N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n
+ N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n N_VPWR_c_486_n
+ N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n VPWR
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_458_n PM_SKY130_FD_SC_HD__CLKINV_16%VPWR
x_PM_SKY130_FD_SC_HD__CLKINV_16%Y N_Y_M1004_s N_Y_M1008_s N_Y_M1016_s
+ N_Y_M1018_s N_Y_M1023_s N_Y_M1026_s N_Y_M1033_s N_Y_M1036_s N_Y_M1000_s
+ N_Y_M1002_s N_Y_M1005_s N_Y_M1009_s N_Y_M1012_s N_Y_M1014_s N_Y_M1019_s
+ N_Y_M1022_s N_Y_M1027_s N_Y_M1029_s N_Y_M1031_s N_Y_M1038_s N_Y_c_638_n
+ N_Y_c_792_n N_Y_c_639_n N_Y_c_640_n N_Y_c_630_n N_Y_c_642_n N_Y_c_631_n
+ N_Y_c_644_n N_Y_c_632_n N_Y_c_646_n N_Y_c_633_n N_Y_c_634_n N_Y_c_649_n
+ N_Y_c_635_n N_Y_c_651_n N_Y_c_636_n N_Y_c_653_n N_Y_c_637_n N_Y_c_655_n
+ N_Y_c_656_n N_Y_c_657_n N_Y_c_658_n N_Y_c_818_n N_Y_c_820_n N_Y_c_659_n
+ N_Y_c_824_n N_Y_c_826_n N_Y_c_828_n N_Y_c_660_n N_Y_c_661_n N_Y_c_662_n Y Y
+ PM_SKY130_FD_SC_HD__CLKINV_16%Y
x_PM_SKY130_FD_SC_HD__CLKINV_16%VGND N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_M1011_d N_VGND_M1017_d N_VGND_M1021_d N_VGND_M1024_d N_VGND_M1032_d
+ N_VGND_M1035_d N_VGND_M1037_d N_VGND_c_862_n N_VGND_c_863_n N_VGND_c_864_n
+ N_VGND_c_865_n N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n
+ N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n
+ N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n
+ N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n N_VGND_c_883_n N_VGND_c_884_n
+ N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n VGND N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n PM_SKY130_FD_SC_HD__CLKINV_16%VGND
cc_1 VNB N_A_M1004_g 0.0383659f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=0.445
cc_2 VNB N_A_M1007_g 0.0275203f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=0.445
cc_3 VNB N_A_M1008_g 0.0275198f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=0.445
cc_4 VNB N_A_M1011_g 0.0275203f $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=0.445
cc_5 VNB N_A_M1016_g 0.0275198f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.445
cc_6 VNB N_A_M1017_g 0.028174f $X=-0.19 $Y=-0.24 $X2=4.355 $Y2=0.445
cc_7 VNB N_A_M1018_g 0.0306683f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=0.445
cc_8 VNB N_A_c_159_n 0.0217642f $X=-0.19 $Y=-0.24 $X2=5.33 $Y2=1.17
cc_9 VNB N_A_c_160_n 0.226899f $X=-0.19 $Y=-0.24 $X2=4.895 $Y2=1.17
cc_10 VNB N_A_M1021_g 0.0300266f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=0.445
cc_11 VNB N_A_M1023_g 0.0275268f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=0.445
cc_12 VNB N_A_M1024_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=6.265 $Y2=0.445
cc_13 VNB N_A_M1026_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=0.445
cc_14 VNB N_A_M1032_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=7.125 $Y2=0.445
cc_15 VNB N_A_M1033_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=7.555 $Y2=0.445
cc_16 VNB N_A_M1035_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=0.445
cc_17 VNB N_A_M1036_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=8.415 $Y2=0.445
cc_18 VNB N_A_M1037_g 0.037667f $X=-0.19 $Y=-0.24 $X2=8.845 $Y2=0.445
cc_19 VNB A 0.0767807f $X=-0.19 $Y=-0.24 $X2=1.985 $Y2=1.105
cc_20 VNB N_A_c_171_n 0.0777531f $X=-0.19 $Y=-0.24 $X2=10.46 $Y2=1.16
cc_21 VNB N_A_c_172_n 0.259413f $X=-0.19 $Y=-0.24 $X2=10.565 $Y2=1.17
cc_22 VNB N_VPWR_c_458_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_23 VNB N_Y_c_630_n 0.00675515f $X=-0.19 $Y=-0.24 $X2=5.33 $Y2=1.17
cc_24 VNB N_Y_c_631_n 0.00687652f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=1.985
cc_25 VNB N_Y_c_632_n 0.00689469f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=1.985
cc_26 VNB N_Y_c_633_n 0.00770315f $X=-0.19 $Y=-0.24 $X2=6.265 $Y2=1.985
cc_27 VNB N_Y_c_634_n 0.00700409f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=1.35
cc_28 VNB N_Y_c_635_n 0.00687169f $X=-0.19 $Y=-0.24 $X2=7.125 $Y2=1.35
cc_29 VNB N_Y_c_636_n 0.00687169f $X=-0.19 $Y=-0.24 $X2=7.555 $Y2=1.35
cc_30 VNB N_Y_c_637_n 0.00696467f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=1.35
cc_31 VNB N_VGND_c_862_n 0.01839f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=1.985
cc_32 VNB N_VGND_c_863_n 0.00402504f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=0.445
cc_33 VNB N_VGND_c_864_n 0.00405516f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=1.985
cc_34 VNB N_VGND_c_865_n 0.00466861f $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=0.445
cc_35 VNB N_VGND_c_866_n 0.00463719f $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=1.985
cc_36 VNB N_VGND_c_867_n 0.00385357f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.445
cc_37 VNB N_VGND_c_868_n 0.00407253f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=1.985
cc_38 VNB N_VGND_c_869_n 0.00402504f $X=-0.19 $Y=-0.24 $X2=4.355 $Y2=0.445
cc_39 VNB N_VGND_c_870_n 0.0165974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_871_n 0.0183325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_872_n 0.0611731f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=0.445
cc_42 VNB N_VGND_c_873_n 0.00516809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_874_n 0.0168213f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=1.985
cc_44 VNB N_VGND_c_875_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=1.985
cc_45 VNB N_VGND_c_876_n 0.0165526f $X=-0.19 $Y=-0.24 $X2=5.33 $Y2=1.17
cc_46 VNB N_VGND_c_877_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=4.895 $Y2=1.17
cc_47 VNB N_VGND_c_878_n 0.0174825f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=0.445
cc_48 VNB N_VGND_c_879_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=0.445
cc_49 VNB N_VGND_c_880_n 0.0210033f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=1.35
cc_50 VNB N_VGND_c_881_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=1.985
cc_51 VNB N_VGND_c_882_n 0.0165974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_883_n 0.00430243f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=0.99
cc_53 VNB N_VGND_c_884_n 0.0179215f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=0.445
cc_54 VNB N_VGND_c_885_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_886_n 0.0165974f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=1.35
cc_56 VNB N_VGND_c_887_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=1.985
cc_57 VNB N_VGND_c_888_n 0.0608549f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=0.445
cc_58 VNB N_VGND_c_889_n 0.649101f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=0.445
cc_59 VNB N_VGND_c_890_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=1.985
cc_60 VPB N_A_M1000_g 0.0240835f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_61 VPB N_A_M1001_g 0.0171919f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.985
cc_62 VPB N_A_M1002_g 0.0171919f $X=-0.19 $Y=1.305 $X2=1.345 $Y2=1.985
cc_63 VPB N_A_M1003_g 0.0171696f $X=-0.19 $Y=1.305 $X2=1.775 $Y2=1.985
cc_64 VPB N_A_M1005_g 0.0171412f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=1.985
cc_65 VPB N_A_M1006_g 0.0167979f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=1.985
cc_66 VPB N_A_M1009_g 0.0167978f $X=-0.19 $Y=1.305 $X2=3.065 $Y2=1.985
cc_67 VPB N_A_M1010_g 0.0167979f $X=-0.19 $Y=1.305 $X2=3.495 $Y2=1.985
cc_68 VPB N_A_M1012_g 0.0167978f $X=-0.19 $Y=1.305 $X2=3.925 $Y2=1.985
cc_69 VPB N_A_M1013_g 0.0171663f $X=-0.19 $Y=1.305 $X2=4.355 $Y2=1.985
cc_70 VPB N_A_M1014_g 0.0185867f $X=-0.19 $Y=1.305 $X2=4.82 $Y2=1.985
cc_71 VPB N_A_c_159_n 0.00935665f $X=-0.19 $Y=1.305 $X2=5.33 $Y2=1.17
cc_72 VPB N_A_c_160_n 0.049742f $X=-0.19 $Y=1.305 $X2=4.895 $Y2=1.17
cc_73 VPB N_A_M1015_g 0.0182207f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=1.985
cc_74 VPB N_A_M1019_g 0.0167992f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=1.985
cc_75 VPB N_A_M1020_g 0.016798f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=1.985
cc_76 VPB N_A_M1022_g 0.016798f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=1.985
cc_77 VPB N_A_M1025_g 0.016798f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=1.985
cc_78 VPB N_A_M1027_g 0.016798f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=1.985
cc_79 VPB N_A_M1028_g 0.016798f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=1.985
cc_80 VPB N_A_M1029_g 0.016798f $X=-0.19 $Y=1.305 $X2=8.415 $Y2=1.985
cc_81 VPB N_A_M1030_g 0.0171405f $X=-0.19 $Y=1.305 $X2=8.845 $Y2=1.985
cc_82 VPB N_A_M1031_g 0.0171685f $X=-0.19 $Y=1.305 $X2=9.275 $Y2=1.985
cc_83 VPB N_A_M1034_g 0.0171919f $X=-0.19 $Y=1.305 $X2=9.705 $Y2=1.985
cc_84 VPB N_A_M1038_g 0.0171919f $X=-0.19 $Y=1.305 $X2=10.135 $Y2=1.985
cc_85 VPB N_A_M1039_g 0.0240835f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.985
cc_86 VPB N_A_c_172_n 0.0580561f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.17
cc_87 VPB N_VPWR_c_459_n 0.0117381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_460_n 0.00465174f $X=-0.19 $Y=1.305 $X2=3.495 $Y2=0.445
cc_89 VPB N_VPWR_c_461_n 0.0040099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_462_n 0.00398868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_463_n 0.00401605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_464_n 0.0040185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_465_n 0.00461913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_466_n 0.00462176f $X=-0.19 $Y=1.305 $X2=5.33 $Y2=1.17
cc_95 VPB N_VPWR_c_467_n 0.00399476f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=0.445
cc_96 VPB N_VPWR_c_468_n 0.00399476f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=1.985
cc_97 VPB N_VPWR_c_469_n 0.00399476f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=0.445
cc_98 VPB N_VPWR_c_470_n 0.016923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_471_n 0.00399476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_472_n 0.00398868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_473_n 0.0113229f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=1.985
cc_102 VPB N_VPWR_c_474_n 0.0281366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_475_n 0.0168773f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=0.445
cc_104 VPB N_VPWR_c_476_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_477_n 0.0169317f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=1.985
cc_106 VPB N_VPWR_c_478_n 0.00497514f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=1.985
cc_107 VPB N_VPWR_c_479_n 0.0168773f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=0.99
cc_108 VPB N_VPWR_c_480_n 0.00487897f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=0.445
cc_109 VPB N_VPWR_c_481_n 0.0176508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_482_n 0.00487897f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=1.35
cc_111 VPB N_VPWR_c_483_n 0.0210316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_484_n 0.00497514f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=0.99
cc_113 VPB N_VPWR_c_485_n 0.016923f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=0.445
cc_114 VPB N_VPWR_c_486_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_487_n 0.016923f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=1.985
cc_116 VPB N_VPWR_c_488_n 0.00487897f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=1.985
cc_117 VPB N_VPWR_c_489_n 0.016923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_490_n 0.00487897f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=0.99
cc_119 VPB N_VPWR_c_491_n 0.0164391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_492_n 0.0170143f $X=-0.19 $Y=1.305 $X2=10.135 $Y2=1.985
cc_121 VPB N_VPWR_c_493_n 0.0167182f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.985
cc_122 VPB N_VPWR_c_494_n 0.00497514f $X=-0.19 $Y=1.305 $X2=9.285 $Y2=1.19
cc_123 VPB N_VPWR_c_495_n 0.00487897f $X=-0.19 $Y=1.305 $X2=9.89 $Y2=1.19
cc_124 VPB N_VPWR_c_496_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_458_n 0.0472716f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_126 VPB N_Y_c_638_n 0.00249649f $X=-0.19 $Y=1.305 $X2=4.355 $Y2=1.35
cc_127 VPB N_Y_c_639_n 0.00250643f $X=-0.19 $Y=1.305 $X2=4.82 $Y2=0.99
cc_128 VPB N_Y_c_640_n 0.00241573f $X=-0.19 $Y=1.305 $X2=4.82 $Y2=1.35
cc_129 VPB N_Y_c_630_n 0.00112034f $X=-0.19 $Y=1.305 $X2=5.33 $Y2=1.17
cc_130 VPB N_Y_c_642_n 0.00261217f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=0.445
cc_131 VPB N_Y_c_631_n 0.00104035f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=1.985
cc_132 VPB N_Y_c_644_n 0.00261217f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=0.445
cc_133 VPB N_Y_c_632_n 0.0010602f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=1.985
cc_134 VPB N_Y_c_646_n 0.00283159f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=0.445
cc_135 VPB N_Y_c_633_n 0.00109244f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=1.985
cc_136 VPB N_Y_c_634_n 0.00107025f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=1.35
cc_137 VPB N_Y_c_649_n 0.00266908f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=0.99
cc_138 VPB N_Y_c_635_n 0.00104488f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=1.35
cc_139 VPB N_Y_c_651_n 0.00266908f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=0.99
cc_140 VPB N_Y_c_636_n 0.00104488f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=1.35
cc_141 VPB N_Y_c_653_n 0.00266908f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=0.99
cc_142 VPB N_Y_c_637_n 0.00112789f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=1.35
cc_143 VPB N_Y_c_655_n 0.00218324f $X=-0.19 $Y=1.305 $X2=8.415 $Y2=0.99
cc_144 VPB N_Y_c_656_n 0.00219711f $X=-0.19 $Y=1.305 $X2=8.415 $Y2=1.35
cc_145 VPB N_Y_c_657_n 0.00173663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_Y_c_658_n 4.29584e-19 $X=-0.19 $Y=1.305 $X2=8.845 $Y2=1.985
cc_147 VPB N_Y_c_659_n 0.00306743f $X=-0.19 $Y=1.305 $X2=9.275 $Y2=1.985
cc_148 VPB N_Y_c_660_n 4.27809e-19 $X=-0.19 $Y=1.305 $X2=10.135 $Y2=1.985
cc_149 VPB N_Y_c_661_n 0.00156462f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.35
cc_150 VPB N_Y_c_662_n 0.00250177f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.985
cc_151 VPB Y 3.21417e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 N_A_M1000_g N_VPWR_c_460_n 0.00343051f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_153 A N_VPWR_c_460_n 0.00239837f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A_M1001_g N_VPWR_c_461_n 0.00160701f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_VPWR_c_461_n 0.0016204f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1003_g N_VPWR_c_462_n 0.00159632f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1005_g N_VPWR_c_462_n 0.00161113f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_M1006_g N_VPWR_c_463_n 0.00161372f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1009_g N_VPWR_c_463_n 0.0016204f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1010_g N_VPWR_c_464_n 0.00159632f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_M1012_g N_VPWR_c_464_n 0.00164413f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_M1013_g N_VPWR_c_465_n 0.0015922f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_M1014_g N_VPWR_c_465_n 0.00301162f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1015_g N_VPWR_c_466_n 0.00304967f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_M1019_g N_VPWR_c_466_n 0.0016204f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_M1020_g N_VPWR_c_467_n 0.00159632f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_M1022_g N_VPWR_c_467_n 0.00161779f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_M1025_g N_VPWR_c_468_n 0.00159632f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_M1027_g N_VPWR_c_468_n 0.00161779f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_M1028_g N_VPWR_c_469_n 0.00159632f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_M1029_g N_VPWR_c_469_n 0.00161779f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_M1029_g N_VPWR_c_470_n 0.00585385f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_M1030_g N_VPWR_c_470_n 0.00585385f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_M1030_g N_VPWR_c_471_n 0.00159632f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_M1031_g N_VPWR_c_471_n 0.00161779f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_M1034_g N_VPWR_c_472_n 0.00159632f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_M1038_g N_VPWR_c_472_n 0.00161113f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_M1039_g N_VPWR_c_474_n 0.00339991f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_c_171_n N_VPWR_c_474_n 0.00133848f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_M1002_g N_VPWR_c_475_n 0.00585385f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_M1003_g N_VPWR_c_475_n 0.00585385f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1005_g N_VPWR_c_477_n 0.00585385f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1006_g N_VPWR_c_477_n 0.00585385f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_M1009_g N_VPWR_c_479_n 0.00585385f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_M1010_g N_VPWR_c_479_n 0.00585385f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_M1012_g N_VPWR_c_481_n 0.00585385f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_M1013_g N_VPWR_c_481_n 0.00585385f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_M1014_g N_VPWR_c_483_n 0.00585385f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_M1015_g N_VPWR_c_483_n 0.00585385f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_M1019_g N_VPWR_c_485_n 0.00585385f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_M1020_g N_VPWR_c_485_n 0.00585385f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_M1022_g N_VPWR_c_487_n 0.00585385f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_M1025_g N_VPWR_c_487_n 0.00585385f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_M1027_g N_VPWR_c_489_n 0.00585385f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_M1028_g N_VPWR_c_489_n 0.00585385f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_M1000_g N_VPWR_c_491_n 0.00585385f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_M1001_g N_VPWR_c_491_n 0.00585385f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_M1031_g N_VPWR_c_492_n 0.00585385f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_M1034_g N_VPWR_c_492_n 0.00585385f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_M1038_g N_VPWR_c_493_n 0.00585385f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_M1039_g N_VPWR_c_493_n 0.00585385f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_M1000_g N_VPWR_c_458_n 0.0114189f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_M1001_g N_VPWR_c_458_n 0.0104895f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_M1002_g N_VPWR_c_458_n 0.0105203f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_M1003_g N_VPWR_c_458_n 0.0105329f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_M1005_g N_VPWR_c_458_n 0.0105203f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_M1006_g N_VPWR_c_458_n 0.0105203f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_M1009_g N_VPWR_c_458_n 0.0105203f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_M1010_g N_VPWR_c_458_n 0.0105329f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_M1012_g N_VPWR_c_458_n 0.0105203f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_M1013_g N_VPWR_c_458_n 0.0106715f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_M1014_g N_VPWR_c_458_n 0.0110562f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_M1015_g N_VPWR_c_458_n 0.010884f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_M1019_g N_VPWR_c_458_n 0.0105203f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_M1020_g N_VPWR_c_458_n 0.0105329f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_M1022_g N_VPWR_c_458_n 0.0105203f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_M1025_g N_VPWR_c_458_n 0.0105329f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_M1027_g N_VPWR_c_458_n 0.0105203f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_M1028_g N_VPWR_c_458_n 0.0105329f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A_M1029_g N_VPWR_c_458_n 0.0105203f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_M1030_g N_VPWR_c_458_n 0.0105329f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A_M1031_g N_VPWR_c_458_n 0.0105203f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_M1034_g N_VPWR_c_458_n 0.0105329f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_M1038_g N_VPWR_c_458_n 0.0105203f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_M1039_g N_VPWR_c_458_n 0.0114529f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_M1000_g N_Y_c_638_n 9.68845e-19 $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_c_160_n N_Y_c_638_n 0.00258307f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_228 A N_Y_c_638_n 0.0208016f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_229 N_A_M1001_g N_Y_c_639_n 0.0145679f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_M1002_g N_Y_c_639_n 0.0145699f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A_c_160_n N_Y_c_639_n 0.00249109f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_232 A N_Y_c_639_n 0.0435023f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A_M1003_g N_Y_c_640_n 0.0145361f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_M1005_g N_Y_c_640_n 0.0148426f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_c_160_n N_Y_c_640_n 0.00249109f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_236 A N_Y_c_640_n 0.0273253f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_237 N_A_c_285_p N_Y_c_640_n 0.0138306f $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_238 N_A_c_286_p N_Y_c_640_n 0.00428581f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_239 N_A_M1004_g N_Y_c_630_n 0.00687088f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_240 N_A_M1005_g N_Y_c_630_n 0.00163185f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A_M1007_g N_Y_c_630_n 0.00479472f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_M1006_g N_Y_c_630_n 9.05456e-19 $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_c_160_n N_Y_c_630_n 0.026551f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_244 A N_Y_c_630_n 0.0270465f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_245 N_A_c_286_p N_Y_c_630_n 0.0318015f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_246 N_A_c_294_p N_Y_c_630_n 0.00339471f $X=2.215 $Y=1.19 $X2=0 $Y2=0
cc_247 N_A_M1006_g N_Y_c_642_n 0.0164628f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_M1009_g N_Y_c_642_n 0.0165564f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_c_160_n N_Y_c_642_n 0.00443815f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_250 N_A_c_286_p N_Y_c_642_n 0.0255685f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_251 N_A_M1008_g N_Y_c_631_n 0.00483858f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_252 N_A_M1009_g N_Y_c_631_n 9.14001e-19 $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_M1011_g N_Y_c_631_n 0.00488763f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_254 N_A_M1010_g N_Y_c_631_n 9.2326e-19 $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_c_160_n N_Y_c_631_n 0.0306427f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_256 N_A_c_286_p N_Y_c_631_n 0.0373719f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_257 N_A_M1010_g N_Y_c_644_n 0.0165672f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_M1012_g N_Y_c_644_n 0.0165672f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A_c_160_n N_Y_c_644_n 0.00443815f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_260 N_A_c_286_p N_Y_c_644_n 0.0255685f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_261 N_A_M1016_g N_Y_c_632_n 0.0047937f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_M1012_g N_Y_c_632_n 9.05401e-19 $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_M1017_g N_Y_c_632_n 0.00486847f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_M1013_g N_Y_c_632_n 9.20002e-19 $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_c_160_n N_Y_c_632_n 0.0304611f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_266 N_A_c_286_p N_Y_c_632_n 0.0356193f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_267 N_A_M1013_g N_Y_c_646_n 0.0168711f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A_M1014_g N_Y_c_646_n 0.0202375f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_c_160_n N_Y_c_646_n 0.0059915f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_270 N_A_c_286_p N_Y_c_646_n 0.027541f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_271 N_A_M1018_g N_Y_c_633_n 0.00605274f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_272 N_A_M1014_g N_Y_c_633_n 0.00114052f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_c_159_n N_Y_c_633_n 0.0421728f $X=5.33 $Y=1.17 $X2=0 $Y2=0
cc_274 N_A_M1021_g N_Y_c_633_n 0.00937526f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_M1015_g N_Y_c_633_n 0.0010184f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_c_286_p N_Y_c_633_n 0.0492578f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_277 N_A_M1023_g N_Y_c_634_n 0.00507366f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_278 N_A_M1019_g N_Y_c_634_n 9.59045e-19 $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A_M1024_g N_Y_c_634_n 0.00484361f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_M1020_g N_Y_c_634_n 9.14964e-19 $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_c_286_p N_Y_c_634_n 0.0368947f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_282 N_A_c_172_n N_Y_c_634_n 0.0309751f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_283 N_A_M1020_g N_Y_c_649_n 0.0165672f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_M1022_g N_Y_c_649_n 0.0165672f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A_c_286_p N_Y_c_649_n 0.0257897f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_286 N_A_c_172_n N_Y_c_649_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_287 N_A_M1026_g N_Y_c_635_n 0.00484361f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_288 N_A_M1022_g N_Y_c_635_n 9.14964e-19 $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A_M1032_g N_Y_c_635_n 0.00484361f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_290 N_A_M1025_g N_Y_c_635_n 9.14964e-19 $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_c_286_p N_Y_c_635_n 0.0367789f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_292 N_A_c_172_n N_Y_c_635_n 0.0305483f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_293 N_A_M1025_g N_Y_c_651_n 0.0165672f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A_M1027_g N_Y_c_651_n 0.0165672f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A_c_286_p N_Y_c_651_n 0.0257897f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_296 N_A_c_172_n N_Y_c_651_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_297 N_A_M1033_g N_Y_c_636_n 0.00484361f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_M1027_g N_Y_c_636_n 9.14964e-19 $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_M1035_g N_Y_c_636_n 0.00484361f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_300 N_A_M1028_g N_Y_c_636_n 9.14964e-19 $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A_c_286_p N_Y_c_636_n 0.0367789f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_302 N_A_c_172_n N_Y_c_636_n 0.0305483f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_303 N_A_M1028_g N_Y_c_653_n 0.0165564f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A_M1029_g N_Y_c_653_n 0.0164842f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A_c_286_p N_Y_c_653_n 0.0257897f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_306 N_A_c_172_n N_Y_c_653_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_307 N_A_M1036_g N_Y_c_637_n 0.00484361f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_308 N_A_M1029_g N_Y_c_637_n 9.14964e-19 $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_M1037_g N_Y_c_637_n 0.00730344f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_310 N_A_M1030_g N_Y_c_637_n 0.00172986f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A_c_286_p N_Y_c_637_n 0.0349206f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_312 N_A_c_360_p N_Y_c_637_n 0.00117738f $X=9.4 $Y=1.19 $X2=0 $Y2=0
cc_313 N_A_c_171_n N_Y_c_637_n 0.0277667f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_c_172_n N_Y_c_637_n 0.0278283f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_315 N_A_M1030_g N_Y_c_655_n 0.0149531f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_M1031_g N_Y_c_655_n 0.0145443f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A_c_286_p N_Y_c_655_n 0.00932131f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_318 N_A_c_360_p N_Y_c_655_n 0.0019287f $X=9.4 $Y=1.19 $X2=0 $Y2=0
cc_319 N_A_c_171_n N_Y_c_655_n 0.0279415f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_c_172_n N_Y_c_655_n 0.00249109f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_321 N_A_M1034_g N_Y_c_656_n 0.0144784f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_M1038_g N_Y_c_656_n 0.0145704f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_c_371_p N_Y_c_656_n 0.0104845f $X=9.89 $Y=1.19 $X2=0 $Y2=0
cc_324 N_A_c_171_n N_Y_c_656_n 0.038728f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_c_172_n N_Y_c_656_n 0.00249109f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_326 N_A_c_160_n N_Y_c_657_n 0.00258307f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_327 A N_Y_c_657_n 0.0173133f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_328 N_A_c_285_p N_Y_c_657_n 0.00572568f $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_329 N_A_M1005_g N_Y_c_658_n 0.00128143f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A_M1015_g N_Y_c_659_n 0.0168834f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A_M1019_g N_Y_c_659_n 0.0165672f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_c_286_p N_Y_c_659_n 0.0273197f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_333 N_A_c_172_n N_Y_c_659_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_334 N_A_M1030_g N_Y_c_660_n 0.00133001f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A_c_360_p N_Y_c_661_n 0.00608613f $X=9.4 $Y=1.19 $X2=0 $Y2=0
cc_336 N_A_c_171_n N_Y_c_661_n 0.0158629f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_c_172_n N_Y_c_661_n 0.00258307f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_338 N_A_M1039_g N_Y_c_662_n 9.74928e-19 $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_c_171_n N_Y_c_662_n 0.0208016f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_c_172_n N_Y_c_662_n 0.00258307f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_341 N_A_c_286_p Y 0.00124485f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_342 N_A_M1004_g N_VGND_c_862_n 0.00372544f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_343 N_A_c_160_n N_VGND_c_862_n 0.00146648f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_344 A N_VGND_c_862_n 0.0131993f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_345 N_A_c_285_p N_VGND_c_862_n 0.00160784f $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_346 N_A_M1007_g N_VGND_c_863_n 0.00167629f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_347 N_A_M1008_g N_VGND_c_863_n 0.00169877f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_348 N_A_c_160_n N_VGND_c_863_n 0.00357354f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_349 N_A_c_286_p N_VGND_c_863_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_350 N_A_M1011_g N_VGND_c_864_n 0.00167629f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_351 N_A_M1016_g N_VGND_c_864_n 0.00173246f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_352 N_A_c_160_n N_VGND_c_864_n 0.00357354f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_353 N_A_c_286_p N_VGND_c_864_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_354 N_A_M1017_g N_VGND_c_865_n 0.00166077f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_355 N_A_M1018_g N_VGND_c_865_n 0.00315583f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_356 N_A_c_160_n N_VGND_c_865_n 0.00482428f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_357 N_A_c_286_p N_VGND_c_865_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_358 N_A_M1021_g N_VGND_c_866_n 0.00312236f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_359 N_A_M1023_g N_VGND_c_866_n 0.00169877f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_360 N_A_c_286_p N_VGND_c_866_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_361 N_A_c_172_n N_VGND_c_866_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_362 N_A_M1024_g N_VGND_c_867_n 0.00165467f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_363 N_A_M1026_g N_VGND_c_867_n 0.0015561f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_364 N_A_c_286_p N_VGND_c_867_n 0.00775425f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_365 N_A_c_172_n N_VGND_c_867_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_366 N_A_M1032_g N_VGND_c_868_n 0.00172922f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_367 N_A_M1033_g N_VGND_c_868_n 0.00169877f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_368 N_A_c_286_p N_VGND_c_868_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_369 N_A_c_172_n N_VGND_c_868_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_370 N_A_M1035_g N_VGND_c_869_n 0.00167629f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_371 N_A_M1036_g N_VGND_c_869_n 0.00169877f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_372 N_A_c_286_p N_VGND_c_869_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_373 N_A_c_172_n N_VGND_c_869_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_374 N_A_M1036_g N_VGND_c_870_n 0.00585385f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_375 N_A_M1037_g N_VGND_c_870_n 0.00585385f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_376 N_A_M1037_g N_VGND_c_871_n 0.00368624f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_377 N_A_c_286_p N_VGND_c_871_n 0.00148989f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_378 N_A_c_171_n N_VGND_c_871_n 0.0131863f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_c_172_n N_VGND_c_871_n 0.00145246f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_380 N_A_M1004_g N_VGND_c_874_n 0.00585385f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_381 N_A_M1007_g N_VGND_c_874_n 0.00585385f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_382 N_A_M1008_g N_VGND_c_876_n 0.00585385f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_383 N_A_M1011_g N_VGND_c_876_n 0.00585385f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_384 N_A_M1016_g N_VGND_c_878_n 0.00585385f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_385 N_A_M1017_g N_VGND_c_878_n 0.00585385f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_386 N_A_M1018_g N_VGND_c_880_n 0.00585385f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_387 N_A_M1021_g N_VGND_c_880_n 0.00585385f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_388 N_A_M1023_g N_VGND_c_882_n 0.00585385f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_389 N_A_M1024_g N_VGND_c_882_n 0.00585385f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_390 N_A_M1026_g N_VGND_c_884_n 0.00585385f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_391 N_A_M1032_g N_VGND_c_884_n 0.00585385f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_392 N_A_M1033_g N_VGND_c_886_n 0.00585385f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_393 N_A_M1035_g N_VGND_c_886_n 0.00585385f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_394 N_A_M1004_g N_VGND_c_889_n 0.0119802f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_395 N_A_M1007_g N_VGND_c_889_n 0.010643f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_396 N_A_M1008_g N_VGND_c_889_n 0.0106305f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_397 N_A_M1011_g N_VGND_c_889_n 0.010643f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_398 N_A_M1016_g N_VGND_c_889_n 0.0106305f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_399 N_A_M1017_g N_VGND_c_889_n 0.0107976f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_400 N_A_M1018_g N_VGND_c_889_n 0.0111111f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_401 N_A_M1021_g N_VGND_c_889_n 0.0110068f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_402 N_A_M1023_g N_VGND_c_889_n 0.0106305f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_403 N_A_M1024_g N_VGND_c_889_n 0.010643f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_404 N_A_M1026_g N_VGND_c_889_n 0.0107309f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_405 N_A_M1032_g N_VGND_c_889_n 0.010643f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_406 N_A_M1033_g N_VGND_c_889_n 0.0106305f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_407 N_A_M1035_g N_VGND_c_889_n 0.010643f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_408 N_A_M1036_g N_VGND_c_889_n 0.0106305f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_409 N_A_M1037_g N_VGND_c_889_n 0.0119927f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_410 N_VPWR_c_458_n N_Y_M1000_s 0.0031002f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_458_n N_Y_M1002_s 0.00310552f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_458_n N_Y_M1005_s 0.00414167f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_c_458_n N_Y_M1009_s 0.00310552f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_458_n N_Y_M1012_s 0.00362594f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_c_458_n N_Y_M1014_s 0.00562307f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_458_n N_Y_M1019_s 0.00327899f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_458_n N_Y_M1022_s 0.00327899f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_458_n N_Y_M1027_s 0.00327899f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_419 N_VPWR_c_458_n N_Y_M1029_s 0.00327899f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_c_458_n N_Y_M1031_s 0.00362594f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_421 N_VPWR_c_458_n N_Y_M1038_s 0.00310552f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_c_491_n N_Y_c_792_n 0.0147601f $X=1 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_c_458_n N_Y_c_792_n 0.00974347f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_424 N_VPWR_M1001_d N_Y_c_639_n 0.00177615f $X=0.99 $Y=1.485 $X2=0 $Y2=0
cc_425 N_VPWR_c_461_n N_Y_c_639_n 0.0137004f $X=1.13 $Y=2 $X2=0 $Y2=0
cc_426 N_VPWR_M1003_d N_Y_c_640_n 0.00177615f $X=1.85 $Y=1.485 $X2=0 $Y2=0
cc_427 N_VPWR_c_462_n N_Y_c_640_n 0.0132336f $X=1.99 $Y=2 $X2=0 $Y2=0
cc_428 N_VPWR_M1006_d N_Y_c_642_n 0.00178571f $X=2.71 $Y=1.485 $X2=0 $Y2=0
cc_429 N_VPWR_c_463_n N_Y_c_642_n 0.0134712f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_430 N_VPWR_M1010_d N_Y_c_644_n 0.00178571f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_431 N_VPWR_c_464_n N_Y_c_644_n 0.0134712f $X=3.71 $Y=2 $X2=0 $Y2=0
cc_432 N_VPWR_M1013_d N_Y_c_646_n 0.00216221f $X=4.43 $Y=1.485 $X2=0 $Y2=0
cc_433 N_VPWR_c_465_n N_Y_c_646_n 0.0163115f $X=4.59 $Y=2 $X2=0 $Y2=0
cc_434 N_VPWR_M1020_d N_Y_c_649_n 0.00178571f $X=6.34 $Y=1.485 $X2=0 $Y2=0
cc_435 N_VPWR_c_467_n N_Y_c_649_n 0.0134712f $X=6.48 $Y=2 $X2=0 $Y2=0
cc_436 N_VPWR_M1025_d N_Y_c_651_n 0.00178571f $X=7.2 $Y=1.485 $X2=0 $Y2=0
cc_437 N_VPWR_c_468_n N_Y_c_651_n 0.0134712f $X=7.34 $Y=2 $X2=0 $Y2=0
cc_438 N_VPWR_M1028_d N_Y_c_653_n 0.00178571f $X=8.06 $Y=1.485 $X2=0 $Y2=0
cc_439 N_VPWR_c_469_n N_Y_c_653_n 0.0134712f $X=8.2 $Y=2 $X2=0 $Y2=0
cc_440 N_VPWR_M1030_d N_Y_c_655_n 0.00177615f $X=8.92 $Y=1.485 $X2=0 $Y2=0
cc_441 N_VPWR_c_471_n N_Y_c_655_n 0.013306f $X=9.06 $Y=2 $X2=0 $Y2=0
cc_442 N_VPWR_M1034_d N_Y_c_656_n 0.00177615f $X=9.78 $Y=1.485 $X2=0 $Y2=0
cc_443 N_VPWR_c_472_n N_Y_c_656_n 0.0132336f $X=9.92 $Y=2 $X2=0 $Y2=0
cc_444 N_VPWR_c_475_n N_Y_c_657_n 0.0134834f $X=1.865 $Y=2.72 $X2=0 $Y2=0
cc_445 N_VPWR_c_458_n N_Y_c_657_n 0.00967382f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_c_477_n N_Y_c_658_n 0.0136957f $X=2.72 $Y=2.72 $X2=0 $Y2=0
cc_447 N_VPWR_c_458_n N_Y_c_658_n 0.00858812f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_448 N_VPWR_c_479_n N_Y_c_818_n 0.0134834f $X=3.585 $Y=2.72 $X2=0 $Y2=0
cc_449 N_VPWR_c_458_n N_Y_c_818_n 0.00967382f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_481_n N_Y_c_820_n 0.0129944f $X=4.465 $Y=2.72 $X2=0 $Y2=0
cc_451 N_VPWR_c_458_n N_Y_c_820_n 0.00910028f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_452 N_VPWR_M1015_d N_Y_c_659_n 0.00178571f $X=5.48 $Y=1.485 $X2=0 $Y2=0
cc_453 N_VPWR_c_615_p N_Y_c_659_n 0.0134712f $X=5.615 $Y=2 $X2=0 $Y2=0
cc_454 N_VPWR_c_485_n N_Y_c_824_n 0.0133204f $X=6.355 $Y=2.72 $X2=0 $Y2=0
cc_455 N_VPWR_c_458_n N_Y_c_824_n 0.00948264f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_456 N_VPWR_c_487_n N_Y_c_826_n 0.0133204f $X=7.215 $Y=2.72 $X2=0 $Y2=0
cc_457 N_VPWR_c_458_n N_Y_c_826_n 0.00948264f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_489_n N_Y_c_828_n 0.0133204f $X=8.075 $Y=2.72 $X2=0 $Y2=0
cc_459 N_VPWR_c_458_n N_Y_c_828_n 0.00948264f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_470_n N_Y_c_660_n 0.0133204f $X=8.935 $Y=2.72 $X2=0 $Y2=0
cc_461 N_VPWR_c_458_n N_Y_c_660_n 0.00948264f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_462 N_VPWR_c_492_n N_Y_c_661_n 0.0129944f $X=9.795 $Y=2.72 $X2=0 $Y2=0
cc_463 N_VPWR_c_458_n N_Y_c_661_n 0.00910028f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_464 N_VPWR_c_493_n N_Y_c_662_n 0.0134834f $X=10.65 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_c_458_n N_Y_c_662_n 0.00967382f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_466 N_VPWR_c_483_n Y 0.022284f $X=5.49 $Y=2.72 $X2=0 $Y2=0
cc_467 N_VPWR_c_458_n Y 0.0142622f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_468 N_Y_c_637_n N_VGND_c_870_n 0.0125932f $X=8.63 $Y=0.445 $X2=0 $Y2=0
cc_469 N_Y_c_630_n N_VGND_c_874_n 0.0118195f $X=2.42 $Y=0.445 $X2=0 $Y2=0
cc_470 N_Y_c_631_n N_VGND_c_876_n 0.012748f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_471 N_Y_c_632_n N_VGND_c_878_n 0.0122837f $X=4.14 $Y=0.445 $X2=0 $Y2=0
cc_472 N_Y_c_633_n N_VGND_c_880_n 0.0197173f $X=5.065 $Y=0.445 $X2=0 $Y2=0
cc_473 N_Y_c_634_n N_VGND_c_882_n 0.0125932f $X=6.05 $Y=0.445 $X2=0 $Y2=0
cc_474 N_Y_c_635_n N_VGND_c_884_n 0.0125932f $X=6.91 $Y=0.445 $X2=0 $Y2=0
cc_475 N_Y_c_636_n N_VGND_c_886_n 0.0125932f $X=7.77 $Y=0.445 $X2=0 $Y2=0
cc_476 N_Y_M1004_s N_VGND_c_889_n 0.00423669f $X=2.28 $Y=0.235 $X2=0 $Y2=0
cc_477 N_Y_M1008_s N_VGND_c_889_n 0.0031965f $X=3.14 $Y=0.235 $X2=0 $Y2=0
cc_478 N_Y_M1016_s N_VGND_c_889_n 0.0037166f $X=4 $Y=0.235 $X2=0 $Y2=0
cc_479 N_Y_M1018_s N_VGND_c_889_n 0.00654074f $X=4.895 $Y=0.235 $X2=0 $Y2=0
cc_480 N_Y_M1023_s N_VGND_c_889_n 0.00336987f $X=5.91 $Y=0.235 $X2=0 $Y2=0
cc_481 N_Y_M1026_s N_VGND_c_889_n 0.00336987f $X=6.77 $Y=0.235 $X2=0 $Y2=0
cc_482 N_Y_M1033_s N_VGND_c_889_n 0.00336987f $X=7.63 $Y=0.235 $X2=0 $Y2=0
cc_483 N_Y_M1036_s N_VGND_c_889_n 0.00336987f $X=8.49 $Y=0.235 $X2=0 $Y2=0
cc_484 N_Y_c_630_n N_VGND_c_889_n 0.00848423f $X=2.42 $Y=0.445 $X2=0 $Y2=0
cc_485 N_Y_c_631_n N_VGND_c_889_n 0.00962561f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_486 N_Y_c_632_n N_VGND_c_889_n 0.00905492f $X=4.14 $Y=0.445 $X2=0 $Y2=0
cc_487 N_Y_c_633_n N_VGND_c_889_n 0.01324f $X=5.065 $Y=0.445 $X2=0 $Y2=0
cc_488 N_Y_c_634_n N_VGND_c_889_n 0.00943538f $X=6.05 $Y=0.445 $X2=0 $Y2=0
cc_489 N_Y_c_635_n N_VGND_c_889_n 0.00943538f $X=6.91 $Y=0.445 $X2=0 $Y2=0
cc_490 N_Y_c_636_n N_VGND_c_889_n 0.00943538f $X=7.77 $Y=0.445 $X2=0 $Y2=0
cc_491 N_Y_c_637_n N_VGND_c_889_n 0.00943538f $X=8.63 $Y=0.445 $X2=0 $Y2=0

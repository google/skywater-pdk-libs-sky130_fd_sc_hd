* File: sky130_fd_sc_hd__a311o_4.pxi.spice
* Created: Thu Aug 27 14:04:07 2020
* 
x_PM_SKY130_FD_SC_HD__A311O_4%C1 N_C1_c_118_n N_C1_M1013_g N_C1_M1005_g
+ N_C1_c_119_n N_C1_M1027_g N_C1_M1020_g C1 C1 C1 N_C1_c_121_n
+ PM_SKY130_FD_SC_HD__A311O_4%C1
x_PM_SKY130_FD_SC_HD__A311O_4%B1 N_B1_c_161_n N_B1_M1018_g N_B1_M1001_g
+ N_B1_c_163_n N_B1_M1019_g N_B1_M1026_g B1 B1 N_B1_c_166_n N_B1_c_167_n
+ PM_SKY130_FD_SC_HD__A311O_4%B1
x_PM_SKY130_FD_SC_HD__A311O_4%A_109_47# N_A_109_47#_M1013_s N_A_109_47#_M1018_s
+ N_A_109_47#_M1004_s N_A_109_47#_M1005_s N_A_109_47#_M1009_g
+ N_A_109_47#_c_216_n N_A_109_47#_c_217_n N_A_109_47#_c_218_n
+ N_A_109_47#_M1011_g N_A_109_47#_M1007_g N_A_109_47#_c_220_n
+ N_A_109_47#_M1015_g N_A_109_47#_M1016_g N_A_109_47#_c_222_n
+ N_A_109_47#_M1025_g N_A_109_47#_c_233_n N_A_109_47#_M1017_g
+ N_A_109_47#_c_234_n N_A_109_47#_M1024_g N_A_109_47#_c_223_n
+ N_A_109_47#_c_247_n N_A_109_47#_c_261_n N_A_109_47#_c_224_n
+ N_A_109_47#_c_225_n N_A_109_47#_c_311_p N_A_109_47#_c_226_n
+ N_A_109_47#_c_227_n N_A_109_47#_c_228_n N_A_109_47#_c_238_n
+ N_A_109_47#_c_239_n N_A_109_47#_c_229_n N_A_109_47#_c_248_n
+ N_A_109_47#_c_250_n N_A_109_47#_c_265_n N_A_109_47#_c_230_n
+ N_A_109_47#_c_290_p PM_SKY130_FD_SC_HD__A311O_4%A_109_47#
x_PM_SKY130_FD_SC_HD__A311O_4%A3 N_A3_c_416_n N_A3_M1002_g N_A3_c_420_n
+ N_A3_M1008_g N_A3_c_417_n N_A3_M1010_g N_A3_c_421_n N_A3_M1012_g A3
+ N_A3_c_419_n PM_SKY130_FD_SC_HD__A311O_4%A3
x_PM_SKY130_FD_SC_HD__A311O_4%A2 N_A2_M1021_g N_A2_M1000_g N_A2_M1023_g
+ N_A2_M1003_g A2 A2 N_A2_c_471_n PM_SKY130_FD_SC_HD__A311O_4%A2
x_PM_SKY130_FD_SC_HD__A311O_4%A1 N_A1_c_513_n N_A1_M1004_g N_A1_M1014_g
+ N_A1_c_514_n N_A1_M1006_g N_A1_M1022_g A1 A1 N_A1_c_516_n
+ PM_SKY130_FD_SC_HD__A311O_4%A1
x_PM_SKY130_FD_SC_HD__A311O_4%A_27_297# N_A_27_297#_M1005_d N_A_27_297#_M1020_d
+ N_A_27_297#_M1026_s N_A_27_297#_c_563_n N_A_27_297#_c_565_n
+ N_A_27_297#_c_585_p N_A_27_297#_c_568_n N_A_27_297#_c_569_n
+ N_A_27_297#_c_574_n N_A_27_297#_c_587_p PM_SKY130_FD_SC_HD__A311O_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A311O_4%A_277_297# N_A_277_297#_M1001_d
+ N_A_277_297#_M1008_s N_A_277_297#_M1021_s N_A_277_297#_M1014_s
+ N_A_277_297#_c_636_n N_A_277_297#_c_595_n N_A_277_297#_c_596_n
+ N_A_277_297#_c_597_n N_A_277_297#_c_615_n N_A_277_297#_c_598_n
+ N_A_277_297#_c_655_p N_A_277_297#_c_624_n N_A_277_297#_c_659_p
+ N_A_277_297#_c_625_n N_A_277_297#_c_626_n N_A_277_297#_c_666_p
+ N_A_277_297#_c_627_n N_A_277_297#_c_628_n
+ PM_SKY130_FD_SC_HD__A311O_4%A_277_297#
x_PM_SKY130_FD_SC_HD__A311O_4%VPWR N_VPWR_M1007_d N_VPWR_M1016_d N_VPWR_M1024_d
+ N_VPWR_M1012_d N_VPWR_M1023_d N_VPWR_M1022_d N_VPWR_c_686_n N_VPWR_c_687_n
+ N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_690_n N_VPWR_c_691_n N_VPWR_c_692_n
+ N_VPWR_c_693_n N_VPWR_c_694_n N_VPWR_c_695_n N_VPWR_c_696_n N_VPWR_c_697_n
+ N_VPWR_c_698_n VPWR N_VPWR_c_699_n N_VPWR_c_700_n N_VPWR_c_701_n
+ N_VPWR_c_702_n N_VPWR_c_703_n N_VPWR_c_685_n PM_SKY130_FD_SC_HD__A311O_4%VPWR
x_PM_SKY130_FD_SC_HD__A311O_4%X N_X_M1009_s N_X_M1015_s N_X_M1007_s N_X_M1017_s
+ N_X_c_811_n N_X_c_816_n N_X_c_819_n N_X_c_825_n N_X_c_828_n X X N_X_c_839_n X
+ N_X_c_842_n PM_SKY130_FD_SC_HD__A311O_4%X
x_PM_SKY130_FD_SC_HD__A311O_4%VGND N_VGND_M1013_d N_VGND_M1027_d N_VGND_M1019_d
+ N_VGND_M1011_d N_VGND_M1025_d N_VGND_M1010_s N_VGND_c_867_n N_VGND_c_868_n
+ N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n
+ N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n
+ N_VGND_c_879_n VGND N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n
+ N_VGND_c_883_n N_VGND_c_884_n PM_SKY130_FD_SC_HD__A311O_4%VGND
x_PM_SKY130_FD_SC_HD__A311O_4%A_861_47# N_A_861_47#_M1002_d N_A_861_47#_M1000_s
+ N_A_861_47#_c_977_n N_A_861_47#_c_980_n N_A_861_47#_c_989_n
+ N_A_861_47#_c_978_n PM_SKY130_FD_SC_HD__A311O_4%A_861_47#
x_PM_SKY130_FD_SC_HD__A311O_4%A_1059_47# N_A_1059_47#_M1000_d
+ N_A_1059_47#_M1003_d N_A_1059_47#_M1006_d N_A_1059_47#_c_1009_n
+ N_A_1059_47#_c_1010_n N_A_1059_47#_c_1011_n N_A_1059_47#_c_1035_n
+ N_A_1059_47#_c_1015_n N_A_1059_47#_c_1012_n
+ PM_SKY130_FD_SC_HD__A311O_4%A_1059_47#
cc_1 VNB N_C1_c_118_n 0.019131f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_C1_c_119_n 0.0161198f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB C1 0.00460065f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_4 VNB N_C1_c_121_n 0.0622937f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B1_c_161_n 0.0151545f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B1_M1001_g 4.13233e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_7 VNB N_B1_c_163_n 0.0151339f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_8 VNB N_B1_M1026_g 7.19898e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_9 VNB B1 4.6614e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_10 VNB N_B1_c_166_n 0.00291062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_11 VNB N_B1_c_167_n 0.0381933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_109_47#_M1009_g 0.0179786f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_13 VNB N_A_109_47#_c_216_n 0.019268f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_14 VNB N_A_109_47#_c_217_n 0.0172086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_109_47#_c_218_n 0.0161302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_109_47#_M1007_g 7.18474e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_109_47#_c_220_n 0.0150503f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_18 VNB N_A_109_47#_M1016_g 4.12504e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_109_47#_c_222_n 0.0189164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_109_47#_c_223_n 0.0016972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_109_47#_c_224_n 0.00296614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_109_47#_c_225_n 0.00288431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_109_47#_c_226_n 0.00787824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_109_47#_c_227_n 0.0801985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_109_47#_c_228_n 5.62858e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_109_47#_c_229_n 9.9079e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_109_47#_c_230_n 0.00158557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A3_c_416_n 0.0167161f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_29 VNB N_A3_c_417_n 0.0190993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB A3 0.00347047f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_31 VNB N_A3_c_419_n 0.0445242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A2_M1021_g 4.85927e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_33 VNB N_A2_M1000_g 0.0233219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_M1023_g 5.70301e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_35 VNB N_A2_M1003_g 0.0177704f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_36 VNB N_A2_c_471_n 0.0618287f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=0.85
cc_37 VNB N_A1_c_513_n 0.0157765f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_38 VNB N_A1_c_514_n 0.0214371f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_39 VNB A1 0.00870246f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_40 VNB N_A1_c_516_n 0.0549817f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_41 VNB N_VPWR_c_685_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_811_n 0.0012044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB X 0.00235543f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.53
cc_44 VNB N_VGND_c_867_n 0.010013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_868_n 0.0177892f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_46 VNB N_VGND_c_869_n 0.00360617f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_47 VNB N_VGND_c_870_n 0.00412551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_871_n 0.00412551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_872_n 0.0190642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_873_n 0.00469317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_874_n 0.0177595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_875_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_876_n 0.0171155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_877_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_878_n 0.0182219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_879_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_880_n 0.0177913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_881_n 0.0583738f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_882_n 0.355472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_883_n 0.0158856f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_884_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_861_47#_c_977_n 0.00183208f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_63 VNB N_A_861_47#_c_978_n 0.0100526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1059_47#_c_1009_n 0.00284208f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_65 VNB N_A_1059_47#_c_1010_n 0.00248421f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_66 VNB N_A_1059_47#_c_1011_n 0.0171297f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_67 VNB N_A_1059_47#_c_1012_n 0.0104834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VPB N_C1_M1005_g 0.0218264f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_69 VPB N_C1_M1020_g 0.018742f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_70 VPB C1 0.00669483f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_71 VPB N_C1_c_121_n 0.0156439f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_72 VPB N_B1_M1001_g 0.0188487f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_73 VPB N_B1_M1026_g 0.0269411f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_74 VPB B1 0.00126587f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_75 VPB N_A_109_47#_M1007_g 0.0260026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_109_47#_M1016_g 0.0185531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_109_47#_c_233_n 0.0140178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_109_47#_c_234_n 0.0141461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_109_47#_c_223_n 0.00213728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_109_47#_c_227_n 0.0123203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_109_47#_c_228_n 0.00140742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_109_47#_c_238_n 0.0185181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_109_47#_c_239_n 3.35748e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_109_47#_c_229_n 8.75061e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A3_c_420_n 0.0135575f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_86 VPB N_A3_c_421_n 0.0142812f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_87 VPB N_A3_c_419_n 0.0122435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A2_M1021_g 0.0202785f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_89 VPB N_A2_M1023_g 0.022663f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_90 VPB N_A1_M1014_g 0.0211591f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_91 VPB N_A1_M1022_g 0.0220857f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_92 VPB A1 0.0123695f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_93 VPB N_A1_c_516_n 0.013954f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_94 VPB N_A_277_297#_c_595_n 0.0120342f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_95 VPB N_A_277_297#_c_596_n 0.00194823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_277_297#_c_597_n 0.00390423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_277_297#_c_598_n 0.00370818f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_98 VPB N_VPWR_c_686_n 0.00544578f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_99 VPB N_VPWR_c_687_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_100 VPB N_VPWR_c_688_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_689_n 0.0109642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_690_n 0.00218776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_691_n 0.0128323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_692_n 0.00273013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_693_n 0.0101444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_694_n 0.0299632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_695_n 0.011815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_696_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_697_n 0.011815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_698_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_699_n 0.0568313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_700_n 0.0231787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_701_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_702_n 0.00564807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_703_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_685_n 0.0518878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB X 0.00172967f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.53
cc_118 N_C1_c_119_n N_B1_c_161_n 0.0252415f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_119 N_C1_c_121_n N_B1_M1001_g 0.0269222f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C1_c_121_n B1 0.00279732f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C1_c_121_n N_B1_c_166_n 0.00197986f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C1_c_119_n N_B1_c_167_n 0.0220929f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_123 N_C1_c_118_n N_A_109_47#_c_223_n 8.74452e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_124 N_C1_M1005_g N_A_109_47#_c_223_n 0.00135794f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_125 N_C1_c_119_n N_A_109_47#_c_223_n 0.00259917f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_126 N_C1_M1020_g N_A_109_47#_c_223_n 0.00146782f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_127 C1 N_A_109_47#_c_223_n 0.0329105f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_128 N_C1_c_121_n N_A_109_47#_c_223_n 0.0193783f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_129 N_C1_c_119_n N_A_109_47#_c_247_n 0.0143483f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_130 N_C1_c_118_n N_A_109_47#_c_248_n 0.00339943f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_131 N_C1_c_119_n N_A_109_47#_c_248_n 0.00248939f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_132 N_C1_M1005_g N_A_109_47#_c_250_n 0.0034859f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C1_M1020_g N_A_109_47#_c_250_n 0.00338974f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_134 C1 N_A_27_297#_M1005_d 0.0104346f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_135 C1 N_A_27_297#_c_563_n 0.0145902f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_136 N_C1_c_121_n N_A_27_297#_c_563_n 6.80961e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_137 N_C1_M1005_g N_A_27_297#_c_565_n 0.0112878f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_138 N_C1_M1020_g N_A_27_297#_c_565_n 0.0112437f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_139 N_C1_M1005_g N_VPWR_c_699_n 0.00357877f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_140 N_C1_M1020_g N_VPWR_c_699_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_141 N_C1_M1005_g N_VPWR_c_685_n 0.00617937f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_142 N_C1_M1020_g N_VPWR_c_685_n 0.00525237f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_143 C1 N_VGND_M1013_d 0.00851678f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_144 N_C1_c_118_n N_VGND_c_868_n 0.00321269f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_145 C1 N_VGND_c_868_n 0.0167027f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_146 N_C1_c_121_n N_VGND_c_868_n 0.00179393f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_147 N_C1_c_119_n N_VGND_c_869_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_148 N_C1_c_118_n N_VGND_c_874_n 0.00542953f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_149 N_C1_c_119_n N_VGND_c_874_n 0.00422842f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_150 N_C1_c_118_n N_VGND_c_882_n 0.0104585f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C1_c_119_n N_VGND_c_882_n 0.00574096f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_152 C1 N_VGND_c_882_n 0.00106649f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_153 N_B1_c_163_n N_A_109_47#_M1009_g 0.0254143f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_154 N_B1_c_166_n N_A_109_47#_c_217_n 2.7761e-19 $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B1_c_167_n N_A_109_47#_c_217_n 0.0182945f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_156 B1 N_A_109_47#_c_223_n 0.0136383f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_157 N_B1_c_166_n N_A_109_47#_c_223_n 0.010735f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B1_c_167_n N_A_109_47#_c_223_n 5.8068e-19 $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_159 N_B1_c_161_n N_A_109_47#_c_247_n 0.00991871f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_160 N_B1_c_166_n N_A_109_47#_c_247_n 0.0210262f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B1_c_167_n N_A_109_47#_c_247_n 0.00132324f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_162 N_B1_c_163_n N_A_109_47#_c_261_n 0.0112845f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_163 N_B1_c_163_n N_A_109_47#_c_224_n 0.00459602f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_164 N_B1_c_166_n N_A_109_47#_c_225_n 0.00850411f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_167_n N_A_109_47#_c_225_n 0.0020541f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_166 N_B1_c_161_n N_A_109_47#_c_265_n 0.00248939f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_167 N_B1_c_163_n N_A_109_47#_c_265_n 0.00248939f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_168 N_B1_c_166_n N_A_109_47#_c_230_n 0.00479914f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B1_c_167_n N_A_109_47#_c_230_n 0.00267128f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_170 B1 N_A_27_297#_M1020_d 0.00270666f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_171 B1 N_A_27_297#_c_568_n 0.0100221f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_172 N_B1_M1001_g N_A_27_297#_c_569_n 0.0118539f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_M1026_g N_A_27_297#_c_569_n 0.00988743f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_174 B1 N_A_27_297#_c_569_n 4.22228e-19 $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_175 N_B1_M1026_g N_A_277_297#_c_595_n 0.0160452f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B1_M1001_g N_A_277_297#_c_596_n 8.20779e-19 $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_177 B1 N_A_277_297#_c_596_n 0.00694391f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_178 N_B1_c_166_n N_A_277_297#_c_596_n 0.00572021f $X=1.34 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B1_c_167_n N_A_277_297#_c_596_n 0.00244702f $X=1.73 $Y=1.135 $X2=0
+ $Y2=0
cc_180 N_B1_M1026_g N_A_277_297#_c_597_n 0.0028084f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B1_M1026_g N_VPWR_c_686_n 0.00235209f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B1_M1001_g N_VPWR_c_699_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_M1026_g N_VPWR_c_699_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1001_g N_VPWR_c_685_n 0.00525237f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1026_g N_VPWR_c_685_n 0.00655123f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_c_161_n N_VGND_c_869_n 0.00146448f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_187 N_B1_c_163_n N_VGND_c_870_n 0.00146448f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_188 N_B1_c_161_n N_VGND_c_876_n 0.00422842f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_189 N_B1_c_163_n N_VGND_c_876_n 0.00422842f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_190 N_B1_c_161_n N_VGND_c_882_n 0.00574096f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_191 N_B1_c_163_n N_VGND_c_882_n 0.00574096f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_192 N_A_109_47#_c_222_n N_A3_c_416_n 0.00648378f $X=3.43 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_193 N_A_109_47#_c_234_n N_A3_c_420_n 0.0237039f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_109_47#_c_228_n N_A3_c_420_n 0.0010783f $X=4.235 $Y=1.455 $X2=0 $Y2=0
cc_195 N_A_109_47#_c_238_n N_A3_c_420_n 0.00877405f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_196 N_A_109_47#_c_239_n N_A3_c_420_n 0.00267886f $X=4.32 $Y=1.54 $X2=0 $Y2=0
cc_197 N_A_109_47#_c_228_n N_A3_c_421_n 2.23052e-19 $X=4.235 $Y=1.455 $X2=0
+ $Y2=0
cc_198 N_A_109_47#_c_238_n N_A3_c_421_n 0.0113039f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_199 N_A_109_47#_c_226_n A3 0.0123701f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_109_47#_c_228_n A3 0.00253048f $X=4.235 $Y=1.455 $X2=0 $Y2=0
cc_201 N_A_109_47#_c_238_n A3 0.0310644f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_202 N_A_109_47#_c_226_n N_A3_c_419_n 0.0160247f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_109_47#_c_227_n N_A3_c_419_n 0.0421978f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_109_47#_c_228_n N_A3_c_419_n 0.00761155f $X=4.235 $Y=1.455 $X2=0
+ $Y2=0
cc_205 N_A_109_47#_c_238_n N_A3_c_419_n 0.00274839f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_206 N_A_109_47#_c_238_n N_A2_M1021_g 0.0121198f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_207 N_A_109_47#_c_238_n N_A2_M1023_g 0.0124755f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_208 N_A_109_47#_c_229_n N_A2_M1003_g 0.00187366f $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_209 N_A_109_47#_c_238_n A2 0.0562044f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_210 N_A_109_47#_c_229_n A2 0.00685196f $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_211 N_A_109_47#_c_238_n N_A2_c_471_n 0.0129518f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_212 N_A_109_47#_c_229_n N_A1_c_513_n 0.00335024f $X=6.6 $Y=1.455 $X2=-0.19
+ $Y2=-0.24
cc_213 N_A_109_47#_c_290_p N_A1_c_513_n 0.00240247f $X=6.68 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_109_47#_c_238_n N_A1_M1014_g 0.0149065f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_215 N_A_109_47#_c_229_n N_A1_M1014_g 0.00610341f $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_216 N_A_109_47#_c_229_n N_A1_c_514_n 0.00235578f $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_217 N_A_109_47#_c_290_p N_A1_c_514_n 0.00370555f $X=6.68 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_109_47#_c_238_n N_A1_M1022_g 0.00162687f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_219 N_A_109_47#_c_229_n N_A1_M1022_g 9.02184e-19 $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_220 N_A_109_47#_c_238_n A1 0.0095858f $X=6.515 $Y=1.54 $X2=0 $Y2=0
cc_221 N_A_109_47#_c_229_n A1 0.0197698f $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_222 N_A_109_47#_c_229_n N_A1_c_516_n 0.0201898f $X=6.6 $Y=1.455 $X2=0 $Y2=0
cc_223 N_A_109_47#_c_290_p N_A1_c_516_n 0.00178884f $X=6.68 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_109_47#_M1005_s N_A_27_297#_c_565_n 0.00312348f $X=0.545 $Y=1.485
+ $X2=0 $Y2=0
cc_225 N_A_109_47#_c_250_n N_A_27_297#_c_565_n 0.015552f $X=0.68 $Y=2.04 $X2=0
+ $Y2=0
cc_226 N_A_109_47#_M1007_g N_A_27_297#_c_574_n 0.00328747f $X=2.67 $Y=1.985
+ $X2=0 $Y2=0
cc_227 N_A_109_47#_c_238_n N_A_277_297#_M1008_s 0.00165831f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_228 N_A_109_47#_c_238_n N_A_277_297#_M1021_s 0.00165831f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_229 N_A_109_47#_c_238_n N_A_277_297#_M1014_s 0.00237967f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_230 N_A_109_47#_c_217_n N_A_277_297#_c_595_n 0.00956453f $X=2.225 $Y=1.16
+ $X2=0 $Y2=0
cc_231 N_A_109_47#_M1007_g N_A_277_297#_c_595_n 0.00384989f $X=2.67 $Y=1.985
+ $X2=0 $Y2=0
cc_232 N_A_109_47#_c_261_n N_A_277_297#_c_595_n 0.00535178f $X=1.855 $Y=0.8
+ $X2=0 $Y2=0
cc_233 N_A_109_47#_c_225_n N_A_277_297#_c_595_n 0.0120409f $X=2.025 $Y=1.16
+ $X2=0 $Y2=0
cc_234 N_A_109_47#_c_311_p N_A_277_297#_c_595_n 0.0232943f $X=2.54 $Y=1.16 $X2=0
+ $Y2=0
cc_235 N_A_109_47#_c_230_n N_A_277_297#_c_596_n 0.00364247f $X=1.52 $Y=0.72
+ $X2=0 $Y2=0
cc_236 N_A_109_47#_M1007_g N_A_277_297#_c_597_n 0.00842066f $X=2.67 $Y=1.985
+ $X2=0 $Y2=0
cc_237 N_A_109_47#_c_216_n N_A_277_297#_c_615_n 0.00355544f $X=2.515 $Y=1.16
+ $X2=0 $Y2=0
cc_238 N_A_109_47#_M1007_g N_A_277_297#_c_615_n 0.0151296f $X=2.67 $Y=1.985
+ $X2=0 $Y2=0
cc_239 N_A_109_47#_M1016_g N_A_277_297#_c_615_n 0.0116149f $X=3.09 $Y=1.985
+ $X2=0 $Y2=0
cc_240 N_A_109_47#_c_233_n N_A_277_297#_c_615_n 0.0116333f $X=3.51 $Y=1.41 $X2=0
+ $Y2=0
cc_241 N_A_109_47#_c_234_n N_A_277_297#_c_615_n 0.0131552f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_109_47#_c_311_p N_A_277_297#_c_615_n 0.00658369f $X=2.54 $Y=1.16
+ $X2=0 $Y2=0
cc_243 N_A_109_47#_c_226_n N_A_277_297#_c_615_n 0.0060034f $X=4.15 $Y=1.16 $X2=0
+ $Y2=0
cc_244 N_A_109_47#_c_238_n N_A_277_297#_c_615_n 0.00459961f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_245 N_A_109_47#_c_239_n N_A_277_297#_c_615_n 0.0058312f $X=4.32 $Y=1.54 $X2=0
+ $Y2=0
cc_246 N_A_109_47#_c_238_n N_A_277_297#_c_624_n 0.0238166f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_247 N_A_109_47#_c_238_n N_A_277_297#_c_625_n 0.0396213f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_248 N_A_109_47#_c_238_n N_A_277_297#_c_626_n 0.00747521f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_249 N_A_109_47#_c_238_n N_A_277_297#_c_627_n 0.0126766f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_250 N_A_109_47#_c_238_n N_A_277_297#_c_628_n 0.0126766f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_251 N_A_109_47#_c_239_n N_VPWR_M1024_d 0.00259754f $X=4.32 $Y=1.54 $X2=0
+ $Y2=0
cc_252 N_A_109_47#_c_238_n N_VPWR_M1012_d 0.00293855f $X=6.515 $Y=1.54 $X2=0
+ $Y2=0
cc_253 N_A_109_47#_c_238_n N_VPWR_M1023_d 0.00952312f $X=6.515 $Y=1.54 $X2=0
+ $Y2=0
cc_254 N_A_109_47#_M1007_g N_VPWR_c_686_n 0.00921014f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_A_109_47#_M1016_g N_VPWR_c_686_n 0.00110281f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_109_47#_M1007_g N_VPWR_c_687_n 0.00110281f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_A_109_47#_M1016_g N_VPWR_c_687_n 0.00810864f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A_109_47#_c_233_n N_VPWR_c_687_n 0.00810864f $X=3.51 $Y=1.41 $X2=0
+ $Y2=0
cc_259 N_A_109_47#_c_234_n N_VPWR_c_687_n 0.00110281f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_260 N_A_109_47#_c_233_n N_VPWR_c_688_n 0.00110281f $X=3.51 $Y=1.41 $X2=0
+ $Y2=0
cc_261 N_A_109_47#_c_234_n N_VPWR_c_688_n 0.00807474f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_262 N_A_109_47#_M1007_g N_VPWR_c_695_n 0.00339367f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_263 N_A_109_47#_M1016_g N_VPWR_c_695_n 0.00339367f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_264 N_A_109_47#_c_233_n N_VPWR_c_697_n 0.00339367f $X=3.51 $Y=1.41 $X2=0
+ $Y2=0
cc_265 N_A_109_47#_c_234_n N_VPWR_c_697_n 0.00339367f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_266 N_A_109_47#_M1005_s N_VPWR_c_685_n 0.00216833f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_109_47#_M1007_g N_VPWR_c_685_n 0.00398704f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A_109_47#_M1016_g N_VPWR_c_685_n 0.00398704f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A_109_47#_c_233_n N_VPWR_c_685_n 0.00398704f $X=3.51 $Y=1.41 $X2=0
+ $Y2=0
cc_270 N_A_109_47#_c_234_n N_VPWR_c_685_n 0.00398704f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_271 N_A_109_47#_c_216_n N_X_c_811_n 0.00257497f $X=2.515 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_109_47#_c_311_p N_X_c_811_n 0.0118846f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_109_47#_c_218_n N_X_c_816_n 0.00991871f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_109_47#_c_311_p N_X_c_816_n 0.0120284f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_109_47#_c_227_n N_X_c_816_n 0.00298152f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_109_47#_M1016_g N_X_c_819_n 0.00541994f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_109_47#_c_233_n N_X_c_819_n 0.00929518f $X=3.51 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_109_47#_c_234_n N_X_c_819_n 0.00374666f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_109_47#_c_226_n N_X_c_819_n 0.0231502f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_109_47#_c_227_n N_X_c_819_n 0.00460987f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_281 N_A_109_47#_c_239_n N_X_c_819_n 0.00489647f $X=4.32 $Y=1.54 $X2=0 $Y2=0
cc_282 N_A_109_47#_M1009_g N_X_c_825_n 0.00283371f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_109_47#_c_218_n N_X_c_825_n 0.00248939f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A_109_47#_c_311_p N_X_c_825_n 0.00166687f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_109_47#_c_220_n N_X_c_828_n 0.00248939f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_109_47#_c_222_n N_X_c_828_n 0.00292987f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A_109_47#_c_226_n N_X_c_828_n 0.00126101f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_109_47#_c_218_n X 0.00210489f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_109_47#_M1007_g X 0.00404077f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_290 N_A_109_47#_c_220_n X 0.00273512f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A_109_47#_M1016_g X 0.00663136f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A_109_47#_c_222_n X 0.00209246f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_109_47#_c_311_p X 0.0111129f $X=2.54 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_109_47#_c_226_n X 0.0129195f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A_109_47#_c_227_n X 0.023128f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_109_47#_M1007_g N_X_c_839_n 0.00382604f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A_109_47#_M1016_g N_X_c_839_n 0.0028141f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A_109_47#_c_227_n N_X_c_839_n 0.00208358f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_109_47#_c_220_n N_X_c_842_n 0.00822784f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_109_47#_c_226_n N_X_c_842_n 0.00169913f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A_109_47#_c_227_n N_X_c_842_n 0.00298232f $X=3.78 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_109_47#_c_247_n N_VGND_M1027_d 0.00433917f $X=1.435 $Y=0.8 $X2=0
+ $Y2=0
cc_303 N_A_109_47#_c_261_n N_VGND_M1019_d 0.00190683f $X=1.855 $Y=0.8 $X2=0
+ $Y2=0
cc_304 N_A_109_47#_c_247_n N_VGND_c_869_n 0.012179f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_305 N_A_109_47#_M1009_g N_VGND_c_870_n 0.00268723f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_306 N_A_109_47#_c_261_n N_VGND_c_870_n 0.0132198f $X=1.855 $Y=0.8 $X2=0 $Y2=0
cc_307 N_A_109_47#_c_218_n N_VGND_c_871_n 0.00268723f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_109_47#_c_220_n N_VGND_c_871_n 0.00146448f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_109_47#_c_247_n N_VGND_c_874_n 0.0020451f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_310 N_A_109_47#_c_248_n N_VGND_c_874_n 0.0148098f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_311 N_A_109_47#_c_247_n N_VGND_c_876_n 0.0020451f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_312 N_A_109_47#_c_261_n N_VGND_c_876_n 0.0020451f $X=1.855 $Y=0.8 $X2=0 $Y2=0
cc_313 N_A_109_47#_c_265_n N_VGND_c_876_n 0.0147217f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_314 N_A_109_47#_M1009_g N_VGND_c_878_n 0.00542953f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_315 N_A_109_47#_c_218_n N_VGND_c_878_n 0.00422842f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_109_47#_c_220_n N_VGND_c_880_n 0.00422842f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_109_47#_c_222_n N_VGND_c_880_n 0.00542953f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_A_109_47#_M1013_s N_VGND_c_882_n 0.00217524f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_319 N_A_109_47#_M1018_s N_VGND_c_882_n 0.00217524f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_320 N_A_109_47#_M1004_s N_VGND_c_882_n 0.00216833f $X=6.545 $Y=0.235 $X2=0
+ $Y2=0
cc_321 N_A_109_47#_M1009_g N_VGND_c_882_n 0.00958372f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_322 N_A_109_47#_c_218_n N_VGND_c_882_n 0.00576601f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_109_47#_c_220_n N_VGND_c_882_n 0.00571376f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_109_47#_c_222_n N_VGND_c_882_n 0.01021f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_109_47#_c_247_n N_VGND_c_882_n 0.00880839f $X=1.435 $Y=0.8 $X2=0
+ $Y2=0
cc_326 N_A_109_47#_c_261_n N_VGND_c_882_n 0.00477685f $X=1.855 $Y=0.8 $X2=0
+ $Y2=0
cc_327 N_A_109_47#_c_248_n N_VGND_c_882_n 0.0117588f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_328 N_A_109_47#_c_265_n N_VGND_c_882_n 0.0117318f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_329 N_A_109_47#_c_222_n N_VGND_c_883_n 0.0020985f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_330 N_A_109_47#_c_226_n N_VGND_c_883_n 0.0167914f $X=4.15 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_109_47#_c_227_n N_VGND_c_883_n 0.00836603f $X=3.78 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_109_47#_c_238_n N_A_861_47#_c_977_n 0.00505228f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_333 N_A_109_47#_c_226_n N_A_861_47#_c_980_n 9.52682e-19 $X=4.15 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_109_47#_c_238_n N_A_861_47#_c_978_n 0.00970516f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_335 N_A_109_47#_c_238_n N_A_1059_47#_c_1010_n 0.00553667f $X=6.515 $Y=1.54
+ $X2=0 $Y2=0
cc_336 N_A_109_47#_c_229_n N_A_1059_47#_c_1011_n 0.00229071f $X=6.6 $Y=1.455
+ $X2=0 $Y2=0
cc_337 N_A_109_47#_M1004_s N_A_1059_47#_c_1015_n 0.00321894f $X=6.545 $Y=0.235
+ $X2=0 $Y2=0
cc_338 N_A_109_47#_c_290_p N_A_1059_47#_c_1015_n 0.0116202f $X=6.68 $Y=0.74
+ $X2=0 $Y2=0
cc_339 N_A3_c_421_n N_A2_M1021_g 0.0248977f $X=4.77 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A3_c_419_n N_A2_M1000_g 0.00156007f $X=4.68 $Y=1.16 $X2=0 $Y2=0
cc_341 A3 A2 0.0113875f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_342 N_A3_c_419_n A2 2.03358e-19 $X=4.68 $Y=1.16 $X2=0 $Y2=0
cc_343 A3 N_A2_c_471_n 0.00189009f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A3_c_419_n N_A2_c_471_n 0.0248977f $X=4.68 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A3_c_420_n N_A_277_297#_c_615_n 0.0100732f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A3_c_421_n N_A_277_297#_c_624_n 0.0104309f $X=4.77 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A3_c_420_n N_VPWR_c_688_n 0.00661031f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A3_c_421_n N_VPWR_c_688_n 5.08801e-19 $X=4.77 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A3_c_420_n N_VPWR_c_689_n 0.00339367f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A3_c_421_n N_VPWR_c_689_n 0.00339367f $X=4.77 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A3_c_420_n N_VPWR_c_690_n 5.10594e-19 $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A3_c_421_n N_VPWR_c_690_n 0.00669517f $X=4.77 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A3_c_420_n N_VPWR_c_685_n 0.00394406f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A3_c_421_n N_VPWR_c_685_n 0.00394406f $X=4.77 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A3_c_420_n N_X_c_819_n 5.06417e-19 $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A3_c_416_n N_VGND_c_872_n 0.00542953f $X=4.23 $Y=0.96 $X2=0 $Y2=0
cc_357 N_A3_c_417_n N_VGND_c_872_n 0.00422842f $X=4.65 $Y=0.96 $X2=0 $Y2=0
cc_358 N_A3_c_417_n N_VGND_c_873_n 0.00438629f $X=4.65 $Y=0.96 $X2=0 $Y2=0
cc_359 N_A3_c_416_n N_VGND_c_882_n 0.0103104f $X=4.23 $Y=0.96 $X2=0 $Y2=0
cc_360 N_A3_c_417_n N_VGND_c_882_n 0.00703983f $X=4.65 $Y=0.96 $X2=0 $Y2=0
cc_361 N_A3_c_416_n N_VGND_c_883_n 0.00574066f $X=4.23 $Y=0.96 $X2=0 $Y2=0
cc_362 A3 N_A_861_47#_c_977_n 4.42941e-19 $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_363 N_A3_c_419_n N_A_861_47#_c_977_n 0.00331639f $X=4.68 $Y=1.16 $X2=0 $Y2=0
cc_364 N_A3_c_416_n N_A_861_47#_c_980_n 0.00310608f $X=4.23 $Y=0.96 $X2=0 $Y2=0
cc_365 N_A3_c_417_n N_A_861_47#_c_980_n 0.0025772f $X=4.65 $Y=0.96 $X2=0 $Y2=0
cc_366 N_A3_c_417_n N_A_861_47#_c_978_n 0.0120514f $X=4.65 $Y=0.96 $X2=0 $Y2=0
cc_367 A3 N_A_861_47#_c_978_n 0.0239129f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_368 N_A3_c_419_n N_A_861_47#_c_978_n 0.00340182f $X=4.68 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A2_M1003_g N_A1_c_513_n 0.0141601f $X=6.05 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_370 N_A2_M1023_g N_A1_c_516_n 0.0203125f $X=5.67 $Y=1.985 $X2=0 $Y2=0
cc_371 A2 N_A1_c_516_n 8.47849e-19 $X=5.75 $Y=1.105 $X2=0 $Y2=0
cc_372 N_A2_c_471_n N_A1_c_516_n 0.0141601f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_373 N_A2_M1021_g N_A_277_297#_c_624_n 0.0107261f $X=5.25 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A2_M1023_g N_A_277_297#_c_625_n 0.0115583f $X=5.67 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A2_M1021_g N_VPWR_c_690_n 0.00168244f $X=5.25 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A2_M1021_g N_VPWR_c_691_n 0.00424386f $X=5.25 $Y=1.985 $X2=0 $Y2=0
cc_377 N_A2_M1023_g N_VPWR_c_691_n 0.00339367f $X=5.67 $Y=1.985 $X2=0 $Y2=0
cc_378 N_A2_M1021_g N_VPWR_c_692_n 5.21357e-19 $X=5.25 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A2_M1023_g N_VPWR_c_692_n 0.00733618f $X=5.67 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A2_M1021_g N_VPWR_c_685_n 0.00570339f $X=5.25 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A2_M1023_g N_VPWR_c_685_n 0.00394406f $X=5.67 $Y=1.985 $X2=0 $Y2=0
cc_382 N_A2_M1000_g N_VGND_c_873_n 0.00182988f $X=5.63 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A2_M1000_g N_VGND_c_881_n 0.00357877f $X=5.63 $Y=0.56 $X2=0 $Y2=0
cc_384 N_A2_M1003_g N_VGND_c_881_n 0.00357877f $X=6.05 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A2_M1000_g N_VGND_c_882_n 0.00655123f $X=5.63 $Y=0.56 $X2=0 $Y2=0
cc_386 N_A2_M1003_g N_VGND_c_882_n 0.00525237f $X=6.05 $Y=0.56 $X2=0 $Y2=0
cc_387 N_A2_M1000_g N_A_861_47#_c_989_n 0.00432481f $X=5.63 $Y=0.56 $X2=0 $Y2=0
cc_388 N_A2_M1003_g N_A_861_47#_c_989_n 0.00332249f $X=6.05 $Y=0.56 $X2=0 $Y2=0
cc_389 N_A2_c_471_n N_A_861_47#_c_989_n 0.00204785f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A2_M1000_g N_A_861_47#_c_978_n 0.00963642f $X=5.63 $Y=0.56 $X2=0 $Y2=0
cc_391 A2 N_A_861_47#_c_978_n 0.0432761f $X=5.75 $Y=1.105 $X2=0 $Y2=0
cc_392 N_A2_c_471_n N_A_861_47#_c_978_n 0.0101948f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_393 N_A2_M1000_g N_A_1059_47#_c_1009_n 0.00904527f $X=5.63 $Y=0.56 $X2=0
+ $Y2=0
cc_394 N_A2_M1003_g N_A_1059_47#_c_1009_n 0.0118158f $X=6.05 $Y=0.56 $X2=0 $Y2=0
cc_395 A2 N_A_1059_47#_c_1009_n 8.50518e-19 $X=5.75 $Y=1.105 $X2=0 $Y2=0
cc_396 N_A1_M1014_g N_A_277_297#_c_625_n 0.0118343f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A1_c_516_n N_A_277_297#_c_626_n 0.00150318f $X=7.11 $Y=1.16 $X2=0 $Y2=0
cc_398 A1 N_VPWR_M1022_d 0.00277241f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_399 N_A1_M1014_g N_VPWR_c_692_n 0.0043611f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A1_M1014_g N_VPWR_c_694_n 0.0012132f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A1_M1022_g N_VPWR_c_694_n 0.0155497f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_402 A1 N_VPWR_c_694_n 0.0225966f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_403 N_A1_c_516_n N_VPWR_c_694_n 0.00112496f $X=7.11 $Y=1.16 $X2=0 $Y2=0
cc_404 N_A1_M1014_g N_VPWR_c_700_n 0.00425094f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A1_M1022_g N_VPWR_c_700_n 0.0046653f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_406 N_A1_M1014_g N_VPWR_c_685_n 0.00656687f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_407 N_A1_M1022_g N_VPWR_c_685_n 0.00789179f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A1_c_513_n N_VGND_c_881_n 0.00357877f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_409 N_A1_c_514_n N_VGND_c_881_n 0.00357877f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A1_c_513_n N_VGND_c_882_n 0.00524329f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A1_c_514_n N_VGND_c_882_n 0.00617937f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_412 N_A1_c_514_n N_A_1059_47#_c_1011_n 4.90791e-19 $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_413 A1 N_A_1059_47#_c_1011_n 0.0213585f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_414 N_A1_c_516_n N_A_1059_47#_c_1011_n 0.00602703f $X=7.11 $Y=1.16 $X2=0
+ $Y2=0
cc_415 N_A1_c_513_n N_A_1059_47#_c_1015_n 0.0113026f $X=6.47 $Y=0.995 $X2=0
+ $Y2=0
cc_416 N_A1_c_514_n N_A_1059_47#_c_1015_n 0.00925842f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_A1_c_513_n N_A_1059_47#_c_1012_n 2.24984e-19 $X=6.47 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A1_c_514_n N_A_1059_47#_c_1012_n 0.00309251f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_419 A1 N_A_1059_47#_c_1012_n 0.00131296f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_420 N_A1_c_516_n N_A_1059_47#_c_1012_n 7.35406e-19 $X=7.11 $Y=1.16 $X2=0
+ $Y2=0
cc_421 N_A_27_297#_c_569_n N_A_277_297#_M1001_d 0.00312348f $X=1.855 $Y=2.38
+ $X2=0.47 $Y2=0.995
cc_422 N_A_27_297#_c_569_n N_A_277_297#_c_636_n 0.0118729f $X=1.855 $Y=2.38
+ $X2=0.15 $Y2=0.765
cc_423 N_A_27_297#_M1026_s N_A_277_297#_c_595_n 0.00390196f $X=1.805 $Y=1.485
+ $X2=0.15 $Y2=1.445
cc_424 N_A_27_297#_c_569_n N_A_277_297#_c_595_n 0.00321995f $X=1.855 $Y=2.38
+ $X2=0.15 $Y2=1.445
cc_425 N_A_27_297#_c_574_n N_A_277_297#_c_595_n 0.0131641f $X=1.94 $Y=1.96
+ $X2=0.15 $Y2=1.445
cc_426 N_A_27_297#_c_574_n N_A_277_297#_c_597_n 0.00891455f $X=1.94 $Y=1.96
+ $X2=0 $Y2=0
cc_427 N_A_27_297#_c_574_n N_A_277_297#_c_598_n 0.0141315f $X=1.94 $Y=1.96
+ $X2=0.245 $Y2=1.16
cc_428 N_A_27_297#_c_569_n N_VPWR_c_686_n 0.010563f $X=1.855 $Y=2.38 $X2=0.245
+ $Y2=1.16
cc_429 N_A_27_297#_c_574_n N_VPWR_c_686_n 0.0022149f $X=1.94 $Y=1.96 $X2=0.245
+ $Y2=1.16
cc_430 N_A_27_297#_c_565_n N_VPWR_c_699_n 0.0358391f $X=1.015 $Y=2.38 $X2=0
+ $Y2=0
cc_431 N_A_27_297#_c_585_p N_VPWR_c_699_n 0.0116982f $X=0.345 $Y=2.38 $X2=0
+ $Y2=0
cc_432 N_A_27_297#_c_569_n N_VPWR_c_699_n 0.0475374f $X=1.855 $Y=2.38 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_c_587_p N_VPWR_c_699_n 0.0114548f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_434 N_A_27_297#_M1005_d N_VPWR_c_685_n 0.00348186f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_A_27_297#_M1020_d N_VPWR_c_685_n 0.0021521f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_436 N_A_27_297#_M1026_s N_VPWR_c_685_n 0.00348186f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_437 N_A_27_297#_c_565_n N_VPWR_c_685_n 0.0234424f $X=1.015 $Y=2.38 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_c_585_p N_VPWR_c_685_n 0.00653925f $X=0.345 $Y=2.38 $X2=0
+ $Y2=0
cc_439 N_A_27_297#_c_569_n N_VPWR_c_685_n 0.0299816f $X=1.855 $Y=2.38 $X2=0
+ $Y2=0
cc_440 N_A_27_297#_c_587_p N_VPWR_c_685_n 0.00653402f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_441 N_A_277_297#_c_595_n N_VPWR_M1007_d 0.00217528f $X=2.195 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_442 N_A_277_297#_c_597_n N_VPWR_M1007_d 0.00418328f $X=2.29 $Y=1.915
+ $X2=-0.19 $Y2=1.305
cc_443 N_A_277_297#_c_615_n N_VPWR_M1007_d 0.00458238f $X=4.475 $Y=2 $X2=-0.19
+ $Y2=1.305
cc_444 N_A_277_297#_c_598_n N_VPWR_M1007_d 0.00100151f $X=2.385 $Y=2 $X2=-0.19
+ $Y2=1.305
cc_445 N_A_277_297#_c_615_n N_VPWR_M1016_d 0.00329049f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_446 N_A_277_297#_c_615_n N_VPWR_M1024_d 0.0043761f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_447 N_A_277_297#_c_624_n N_VPWR_M1012_d 0.00514755f $X=5.375 $Y=2 $X2=0 $Y2=0
cc_448 N_A_277_297#_c_625_n N_VPWR_M1023_d 0.0171567f $X=6.595 $Y=2 $X2=0 $Y2=0
cc_449 N_A_277_297#_c_615_n N_VPWR_c_686_n 0.0136707f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_450 N_A_277_297#_c_598_n N_VPWR_c_686_n 0.00758686f $X=2.385 $Y=2 $X2=0 $Y2=0
cc_451 N_A_277_297#_c_615_n N_VPWR_c_687_n 0.0159625f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_452 N_A_277_297#_c_615_n N_VPWR_c_688_n 0.0159625f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_453 N_A_277_297#_c_615_n N_VPWR_c_689_n 0.00243651f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_454 N_A_277_297#_c_655_p N_VPWR_c_689_n 0.0113839f $X=4.56 $Y=2.3 $X2=0 $Y2=0
cc_455 N_A_277_297#_c_624_n N_VPWR_c_689_n 0.00243651f $X=5.375 $Y=2 $X2=0 $Y2=0
cc_456 N_A_277_297#_c_624_n N_VPWR_c_690_n 0.0185102f $X=5.375 $Y=2 $X2=0 $Y2=0
cc_457 N_A_277_297#_c_624_n N_VPWR_c_691_n 0.00292742f $X=5.375 $Y=2 $X2=0 $Y2=0
cc_458 N_A_277_297#_c_659_p N_VPWR_c_691_n 0.0113839f $X=5.46 $Y=2.3 $X2=0 $Y2=0
cc_459 N_A_277_297#_c_625_n N_VPWR_c_691_n 0.00243651f $X=6.595 $Y=2 $X2=0 $Y2=0
cc_460 N_A_277_297#_c_625_n N_VPWR_c_692_n 0.020494f $X=6.595 $Y=2 $X2=0 $Y2=0
cc_461 N_A_277_297#_c_615_n N_VPWR_c_695_n 0.0077537f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_462 N_A_277_297#_c_615_n N_VPWR_c_697_n 0.0077537f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_463 N_A_277_297#_c_598_n N_VPWR_c_699_n 0.00200864f $X=2.385 $Y=2 $X2=0 $Y2=0
cc_464 N_A_277_297#_c_625_n N_VPWR_c_700_n 0.00861366f $X=6.595 $Y=2 $X2=0 $Y2=0
cc_465 N_A_277_297#_c_666_p N_VPWR_c_700_n 0.0113839f $X=6.68 $Y=2.3 $X2=0 $Y2=0
cc_466 N_A_277_297#_M1001_d N_VPWR_c_685_n 0.00216833f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_A_277_297#_M1008_s N_VPWR_c_685_n 0.00249348f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_468 N_A_277_297#_M1021_s N_VPWR_c_685_n 0.00249348f $X=5.325 $Y=1.485 $X2=0
+ $Y2=0
cc_469 N_A_277_297#_M1014_s N_VPWR_c_685_n 0.00405853f $X=6.545 $Y=1.485 $X2=0
+ $Y2=0
cc_470 N_A_277_297#_c_615_n N_VPWR_c_685_n 0.034748f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_471 N_A_277_297#_c_598_n N_VPWR_c_685_n 0.00349024f $X=2.385 $Y=2 $X2=0 $Y2=0
cc_472 N_A_277_297#_c_655_p N_VPWR_c_685_n 0.00646745f $X=4.56 $Y=2.3 $X2=0
+ $Y2=0
cc_473 N_A_277_297#_c_624_n N_VPWR_c_685_n 0.0107993f $X=5.375 $Y=2 $X2=0 $Y2=0
cc_474 N_A_277_297#_c_659_p N_VPWR_c_685_n 0.00646745f $X=5.46 $Y=2.3 $X2=0
+ $Y2=0
cc_475 N_A_277_297#_c_625_n N_VPWR_c_685_n 0.0206228f $X=6.595 $Y=2 $X2=0 $Y2=0
cc_476 N_A_277_297#_c_666_p N_VPWR_c_685_n 0.00646745f $X=6.68 $Y=2.3 $X2=0
+ $Y2=0
cc_477 N_A_277_297#_c_615_n N_X_M1007_s 0.00441227f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_478 N_A_277_297#_c_615_n N_X_M1017_s 0.00438565f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_479 N_A_277_297#_c_615_n N_X_c_819_n 0.0342841f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_480 N_A_277_297#_c_595_n X 0.00326263f $X=2.195 $Y=1.54 $X2=0 $Y2=0
cc_481 N_A_277_297#_c_595_n N_X_c_839_n 0.00418573f $X=2.195 $Y=1.54 $X2=0 $Y2=0
cc_482 N_A_277_297#_c_597_n N_X_c_839_n 0.00424563f $X=2.29 $Y=1.915 $X2=0 $Y2=0
cc_483 N_A_277_297#_c_615_n N_X_c_839_n 0.0181513f $X=4.475 $Y=2 $X2=0 $Y2=0
cc_484 N_VPWR_c_685_n N_X_M1007_s 0.00315309f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_485 N_VPWR_c_685_n N_X_M1017_s 0.00315309f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_486 N_VPWR_M1016_d N_X_c_819_n 0.00394439f $X=3.165 $Y=1.485 $X2=0 $Y2=0
cc_487 N_X_c_816_n N_VGND_M1011_d 0.00415089f $X=2.91 $Y=0.8 $X2=0 $Y2=0
cc_488 N_X_c_816_n N_VGND_c_871_n 0.012179f $X=2.91 $Y=0.8 $X2=0 $Y2=0
cc_489 N_X_c_816_n N_VGND_c_878_n 0.0020451f $X=2.91 $Y=0.8 $X2=0 $Y2=0
cc_490 N_X_c_825_n N_VGND_c_878_n 0.0157702f $X=2.38 $Y=0.38 $X2=0 $Y2=0
cc_491 N_X_c_828_n N_VGND_c_880_n 0.0145181f $X=3.22 $Y=0.38 $X2=0 $Y2=0
cc_492 N_X_c_842_n N_VGND_c_880_n 0.0020451f $X=3.22 $Y=0.72 $X2=0 $Y2=0
cc_493 N_X_M1009_s N_VGND_c_882_n 0.00233757f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_494 N_X_M1015_s N_VGND_c_882_n 0.00217524f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_495 N_X_c_816_n N_VGND_c_882_n 0.00881806f $X=2.91 $Y=0.8 $X2=0 $Y2=0
cc_496 N_X_c_825_n N_VGND_c_882_n 0.0124593f $X=2.38 $Y=0.38 $X2=0 $Y2=0
cc_497 N_X_c_828_n N_VGND_c_882_n 0.0116712f $X=3.22 $Y=0.38 $X2=0 $Y2=0
cc_498 N_VGND_c_882_n N_A_861_47#_M1002_d 0.00217524f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_499 N_VGND_c_882_n N_A_861_47#_M1000_s 0.00216833f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_500 N_VGND_c_872_n N_A_861_47#_c_980_n 0.0147217f $X=4.775 $Y=0 $X2=0 $Y2=0
cc_501 N_VGND_c_882_n N_A_861_47#_c_980_n 0.0117318f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_c_883_n N_A_861_47#_c_980_n 0.0116076f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_503 N_VGND_M1010_s N_A_861_47#_c_978_n 0.00559932f $X=4.725 $Y=0.235 $X2=0
+ $Y2=0
cc_504 N_VGND_c_872_n N_A_861_47#_c_978_n 0.0020451f $X=4.775 $Y=0 $X2=0 $Y2=0
cc_505 N_VGND_c_873_n N_A_861_47#_c_978_n 0.0126475f $X=4.86 $Y=0.38 $X2=0 $Y2=0
cc_506 N_VGND_c_881_n N_A_861_47#_c_978_n 0.00477837f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_882_n N_A_861_47#_c_978_n 0.0139863f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_882_n N_A_1059_47#_M1000_d 0.00209344f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_509 N_VGND_c_882_n N_A_1059_47#_M1003_d 0.0021521f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_882_n N_A_1059_47#_M1006_d 0.00209344f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_873_n N_A_1059_47#_c_1009_n 0.0112553f $X=4.86 $Y=0.38 $X2=0
+ $Y2=0
cc_512 N_VGND_c_881_n N_A_1059_47#_c_1009_n 0.0521531f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_882_n N_A_1059_47#_c_1009_n 0.0329109f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_881_n N_A_1059_47#_c_1035_n 0.0114055f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_c_882_n N_A_1059_47#_c_1035_n 0.00653405f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_881_n N_A_1059_47#_c_1015_n 0.0522677f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_882_n N_A_1059_47#_c_1015_n 0.0330392f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_518 N_A_861_47#_c_978_n N_A_1059_47#_M1000_d 0.0049863f $X=5.675 $Y=0.765
+ $X2=-0.19 $Y2=-0.24
cc_519 N_A_861_47#_M1000_s N_A_1059_47#_c_1009_n 0.00309306f $X=5.705 $Y=0.235
+ $X2=0 $Y2=0
cc_520 N_A_861_47#_c_989_n N_A_1059_47#_c_1009_n 0.0144458f $X=5.84 $Y=0.73
+ $X2=0 $Y2=0
cc_521 N_A_861_47#_c_978_n N_A_1059_47#_c_1009_n 0.0179545f $X=5.675 $Y=0.765
+ $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_79_21# A3 a_429_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=4.3e+11p ps=2.86e+06u
M1001 a_429_297# A2 a_345_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1002 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=1.2e+12p pd=8.4e+06u as=2.7e+11p ps=2.54e+06u
M1003 VPWR B1 a_629_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.8e+11p ps=2.76e+06u
M1004 a_629_297# B2 a_79_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=8.45e+11p pd=6.5e+06u as=1.755e+11p ps=1.84e+06u
M1006 a_345_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_79_21# B2 a_345_47# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=5.655e+11p ps=5.64e+06u
M1008 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_345_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_345_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_345_47# B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_345_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

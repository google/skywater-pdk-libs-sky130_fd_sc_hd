* File: sky130_fd_sc_hd__o211a_2.pxi.spice
* Created: Tue Sep  1 19:20:35 2020
* 
x_PM_SKY130_FD_SC_HD__O211A_2%C1 N_C1_M1003_g N_C1_M1004_g C1 N_C1_c_65_n
+ N_C1_c_66_n N_C1_c_69_n C1 PM_SKY130_FD_SC_HD__O211A_2%C1
x_PM_SKY130_FD_SC_HD__O211A_2%B1 N_B1_M1000_g N_B1_M1011_g B1 N_B1_c_90_n
+ N_B1_c_91_n PM_SKY130_FD_SC_HD__O211A_2%B1
x_PM_SKY130_FD_SC_HD__O211A_2%A2 N_A2_M1002_g N_A2_M1007_g A2 N_A2_c_122_n
+ N_A2_c_123_n N_A2_c_125_n PM_SKY130_FD_SC_HD__O211A_2%A2
x_PM_SKY130_FD_SC_HD__O211A_2%A1 N_A1_M1008_g N_A1_M1006_g A1 N_A1_c_150_n
+ N_A1_c_151_n N_A1_c_152_n PM_SKY130_FD_SC_HD__O211A_2%A1
x_PM_SKY130_FD_SC_HD__O211A_2%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1004_s
+ N_A_27_47#_M1011_d N_A_27_47#_c_185_n N_A_27_47#_M1005_g N_A_27_47#_M1001_g
+ N_A_27_47#_c_186_n N_A_27_47#_M1010_g N_A_27_47#_M1009_g N_A_27_47#_c_193_n
+ N_A_27_47#_c_187_n N_A_27_47#_c_188_n N_A_27_47#_c_213_n N_A_27_47#_c_195_n
+ N_A_27_47#_c_245_p N_A_27_47#_c_218_n N_A_27_47#_c_196_n N_A_27_47#_c_189_n
+ N_A_27_47#_c_197_n N_A_27_47#_c_216_n N_A_27_47#_c_190_n
+ PM_SKY130_FD_SC_HD__O211A_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O211A_2%VPWR N_VPWR_M1004_d N_VPWR_M1008_d N_VPWR_M1009_s
+ N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n VPWR
+ N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n
+ N_VPWR_c_286_n PM_SKY130_FD_SC_HD__O211A_2%VPWR
x_PM_SKY130_FD_SC_HD__O211A_2%X N_X_M1005_d N_X_M1001_d N_X_c_346_n N_X_c_367_n
+ N_X_c_344_n N_X_c_353_n N_X_c_355_n N_X_c_347_n X N_X_c_342_n X
+ PM_SKY130_FD_SC_HD__O211A_2%X
x_PM_SKY130_FD_SC_HD__O211A_2%A_182_47# N_A_182_47#_M1000_d N_A_182_47#_M1002_d
+ N_A_182_47#_c_389_n PM_SKY130_FD_SC_HD__O211A_2%A_182_47#
x_PM_SKY130_FD_SC_HD__O211A_2%VGND N_VGND_M1002_s N_VGND_M1006_d N_VGND_M1010_s
+ N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n
+ N_VGND_c_412_n VGND N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n PM_SKY130_FD_SC_HD__O211A_2%VGND
cc_1 VNB C1 0.011737f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_2 VNB N_C1_c_65_n 0.0338286f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_3 VNB N_C1_c_66_n 0.0209404f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=0.995
cc_4 VNB B1 0.00361788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_B1_c_90_n 0.0262131f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_6 VNB N_B1_c_91_n 0.0216026f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.37
cc_7 VNB N_A2_c_122_n 0.0309573f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_8 VNB N_A2_c_123_n 0.0214255f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=0.995
cc_9 VNB N_A1_c_150_n 0.02393f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_10 VNB N_A1_c_151_n 0.00262721f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=0.995
cc_11 VNB N_A1_c_152_n 0.0170444f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.37
cc_12 VNB N_A_27_47#_c_185_n 0.0168039f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_13 VNB N_A_27_47#_c_186_n 0.0193793f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_14 VNB N_A_27_47#_c_187_n 0.0238425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_188_n 0.00279057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_189_n 0.00450395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_190_n 0.0483075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_286_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_342_n 0.00707011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.0192165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_182_47#_c_389_n 0.0129227f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_22 VNB N_VGND_c_407_n 0.00669754f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=0.995
cc_23 VNB N_VGND_c_408_n 0.00389835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_409_n 0.0126576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_410_n 0.013358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_411_n 0.0157807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_412_n 0.00448835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_413_n 0.0389455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_414_n 0.0171549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_415_n 0.00516774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_416_n 0.203591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB C1 0.00101332f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_C1_c_65_n 0.0139339f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_34 VPB N_C1_c_69_n 0.0218101f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.37
cc_35 VPB N_B1_M1011_g 0.024913f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_36 VPB B1 0.00147897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_B1_c_90_n 0.00612746f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_38 VPB N_A2_c_122_n 0.0124901f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_39 VPB N_A2_c_125_n 0.0208306f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.37
cc_40 VPB N_A1_M1008_g 0.0193896f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_41 VPB N_A1_c_150_n 0.00518771f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_42 VPB N_A1_c_151_n 9.25963e-19 $X=-0.19 $Y=1.305 $X2=0.327 $Y2=0.995
cc_43 VPB N_A_27_47#_M1001_g 0.0191803f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_44 VPB N_A_27_47#_M1009_g 0.0214522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_193_n 0.0269609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_188_n 0.00161068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_195_n 0.0111775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_196_n 0.00165093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_197_n 0.00539858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_190_n 0.0124424f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_287_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.327 $Y2=0.995
cc_52 VPB N_VPWR_c_288_n 5.66763e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_289_n 0.0128606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_290_n 0.0119106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_291_n 0.0153288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_292_n 0.034359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_293_n 0.0125091f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_294_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_295_n 0.00587791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_286_n 0.0462881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_X_c_344_n 0.00828609f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_62 VPB X 0.0236601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 N_C1_c_65_n N_B1_M1011_g 0.0272665f $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_64 N_C1_c_65_n B1 2.52061e-19 $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_65 N_C1_c_65_n N_B1_c_90_n 0.0371402f $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_66 N_C1_c_66_n N_B1_c_91_n 0.0371402f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_67 C1 N_A_27_47#_c_187_n 0.0209423f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_68 N_C1_c_65_n N_A_27_47#_c_187_n 0.00683765f $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_69 N_C1_c_66_n N_A_27_47#_c_187_n 0.0194835f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_70 C1 N_A_27_47#_c_188_n 0.023306f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_71 N_C1_c_65_n N_A_27_47#_c_188_n 0.00933493f $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C1_c_66_n N_A_27_47#_c_188_n 0.00774182f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_73 N_C1_c_69_n N_A_27_47#_c_188_n 0.00671093f $X=0.327 $Y=1.37 $X2=0 $Y2=0
cc_74 C1 N_A_27_47#_c_195_n 0.0187643f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 N_C1_c_65_n N_A_27_47#_c_195_n 0.0070044f $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_76 N_C1_c_69_n N_A_27_47#_c_195_n 0.0210839f $X=0.327 $Y=1.37 $X2=0 $Y2=0
cc_77 N_C1_c_69_n N_VPWR_c_287_n 0.0114792f $X=0.327 $Y=1.37 $X2=0 $Y2=0
cc_78 N_C1_c_69_n N_VPWR_c_291_n 0.00486043f $X=0.327 $Y=1.37 $X2=0 $Y2=0
cc_79 N_C1_c_69_n N_VPWR_c_286_n 0.00915791f $X=0.327 $Y=1.37 $X2=0 $Y2=0
cc_80 N_C1_c_66_n N_VGND_c_413_n 0.00384085f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_81 N_C1_c_66_n N_VGND_c_416_n 0.0061812f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_82 B1 A2 0.0175203f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B1_c_90_n A2 3.20197e-19 $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B1_M1011_g N_A2_c_122_n 0.00193983f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_85 B1 N_A2_c_122_n 0.00277987f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B1_c_90_n N_A2_c_122_n 0.00974493f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_c_91_n N_A_27_47#_c_187_n 8.62955e-19 $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B1_M1011_g N_A_27_47#_c_188_n 0.00411002f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_89 B1 N_A_27_47#_c_188_n 0.0250427f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B1_c_91_n N_A_27_47#_c_188_n 0.00501402f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_M1011_g N_A_27_47#_c_213_n 0.0225673f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_92 B1 N_A_27_47#_c_213_n 0.00845477f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B1_c_90_n N_A_27_47#_c_213_n 0.00190801f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_94 B1 N_A_27_47#_c_216_n 0.0167072f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B1_c_90_n N_A_27_47#_c_216_n 0.00169578f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B1_M1011_g N_VPWR_c_287_n 0.0114792f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B1_M1011_g N_VPWR_c_292_n 0.00486043f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B1_M1011_g N_VPWR_c_286_n 0.00965187f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_99 B1 N_A_182_47#_c_389_n 0.0252602f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_100 N_B1_c_90_n N_A_182_47#_c_389_n 0.00441823f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B1_c_91_n N_A_182_47#_c_389_n 0.00300687f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_91_n N_VGND_c_407_n 0.00825023f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B1_c_91_n N_VGND_c_413_n 0.00553327f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B1_c_91_n N_VGND_c_416_n 0.0110672f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A2_c_125_n N_A1_M1008_g 0.0501084f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_106 A2 N_A1_c_150_n 3.21875e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A2_c_122_n N_A1_c_150_n 0.0501084f $X=1.685 $Y=1.16 $X2=0 $Y2=0
cc_108 A2 N_A1_c_151_n 0.0260015f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_109 N_A2_c_122_n N_A1_c_151_n 0.00206466f $X=1.685 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A2_c_123_n N_A1_c_152_n 0.0248347f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_111 A2 N_A_27_47#_c_218_n 0.00792202f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_112 N_A2_c_125_n N_A_27_47#_c_218_n 0.0207361f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_113 A2 N_A_27_47#_c_216_n 0.0112033f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_114 N_A2_c_122_n N_A_27_47#_c_216_n 0.00671815f $X=1.685 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A2_c_125_n N_VPWR_c_288_n 0.00271371f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_116 N_A2_c_125_n N_VPWR_c_292_n 0.00585385f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A2_c_125_n N_VPWR_c_286_n 0.0120541f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_118 A2 N_A_182_47#_c_389_n 0.0191789f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_119 N_A2_c_122_n N_A_182_47#_c_389_n 0.00584428f $X=1.685 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A2_c_123_n N_A_182_47#_c_389_n 0.0130775f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A2_c_123_n N_VGND_c_407_n 0.00968627f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A2_c_123_n N_VGND_c_411_n 0.00339367f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A2_c_123_n N_VGND_c_416_n 0.00404074f $X=1.67 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A1_c_152_n N_A_27_47#_c_185_n 0.0232114f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A1_M1008_g N_A_27_47#_M1001_g 0.0281237f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A1_c_150_n N_A_27_47#_M1001_g 2.44719e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A1_M1008_g N_A_27_47#_c_218_n 0.018002f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A1_c_150_n N_A_27_47#_c_218_n 0.0046107f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A1_c_151_n N_A_27_47#_c_218_n 0.0197292f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_M1008_g N_A_27_47#_c_196_n 0.00353172f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_c_150_n N_A_27_47#_c_189_n 0.00229355f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A1_c_151_n N_A_27_47#_c_189_n 0.0278224f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A1_c_150_n N_A_27_47#_c_190_n 0.0201501f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A1_c_151_n N_A_27_47#_c_190_n 2.98289e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A1_M1008_g N_VPWR_c_288_n 0.0147258f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A1_M1008_g N_VPWR_c_292_n 0.00486043f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A1_M1008_g N_VPWR_c_286_n 0.00814024f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_c_152_n N_X_c_346_n 4.29205e-19 $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_c_152_n N_X_c_347_n 5.49072e-19 $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_151_n N_A_182_47#_c_389_n 0.0100609f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A1_c_152_n N_A_182_47#_c_389_n 0.00440765f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_152_n N_VGND_c_407_n 0.0011546f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_150_n N_VGND_c_408_n 0.00191959f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A1_c_152_n N_VGND_c_408_n 0.00152546f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A1_c_152_n N_VGND_c_411_n 0.0055867f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A1_c_152_n N_VGND_c_416_n 0.00996457f $X=2.23 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_188_n N_VPWR_M1004_d 5.85117e-19 $X=0.62 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_27_47#_c_213_n N_VPWR_M1004_d 0.00279092f $X=1.025 $Y=1.637 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A_27_47#_c_195_n N_VPWR_M1004_d 0.00139951f $X=0.71 $Y=1.637 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_27_47#_c_218_n N_VPWR_M1008_d 0.00887277f $X=2.495 $Y=1.637 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_c_196_n N_VPWR_M1008_d 3.00687e-19 $X=2.58 $Y=1.51 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_195_n N_VPWR_c_287_n 0.0174843f $X=0.71 $Y=1.637 $X2=0 $Y2=0
cc_153 N_A_27_47#_M1001_g N_VPWR_c_288_n 0.0177829f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_27_47#_M1009_g N_VPWR_c_288_n 6.60035e-19 $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_218_n N_VPWR_c_288_n 0.0264359f $X=2.495 $Y=1.637 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_M1001_g N_VPWR_c_290_n 5.08245e-19 $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_M1009_g N_VPWR_c_290_n 0.00749508f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_193_n N_VPWR_c_291_n 0.0182098f $X=0.26 $Y=1.82 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_245_p N_VPWR_c_292_n 0.0453367f $X=1.53 $Y=1.89 $X2=0 $Y2=0
cc_160 N_A_27_47#_M1001_g N_VPWR_c_293_n 0.00525069f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_M1009_g N_VPWR_c_293_n 0.00354752f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_M1004_s N_VPWR_c_286_n 0.00369639f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_M1011_d N_VPWR_c_286_n 0.00829096f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1001_g N_VPWR_c_286_n 0.00883958f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_M1009_g N_VPWR_c_286_n 0.00413327f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_193_n N_VPWR_c_286_n 0.0101364f $X=0.26 $Y=1.82 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_245_p N_VPWR_c_286_n 0.0257259f $X=1.53 $Y=1.89 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_218_n A_373_297# 0.00688507f $X=2.495 $Y=1.637 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_27_47#_c_185_n N_X_c_346_n 0.00462146f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_186_n N_X_c_346_n 0.00954555f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_27_47#_M1009_g N_X_c_344_n 0.0149668f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_197_n N_X_c_344_n 0.00417363f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_190_n N_X_c_344_n 0.00300016f $X=3.12 $Y=1.157 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_197_n N_X_c_353_n 0.00626655f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_190_n N_X_c_353_n 6.09191e-19 $X=3.12 $Y=1.157 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_186_n N_X_c_355_n 0.0101588f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_197_n N_X_c_355_n 0.00750973f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_190_n N_X_c_355_n 0.0052191f $X=3.12 $Y=1.157 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_185_n N_X_c_347_n 0.00352979f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_186_n N_X_c_347_n 7.52978e-19 $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_197_n N_X_c_347_n 0.0182767f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_190_n N_X_c_347_n 0.00232886f $X=3.12 $Y=1.157 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_186_n X 0.00727198f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1009_g X 0.0207007f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_197_n X 0.0251969f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_190_n X 0.0158719f $X=3.12 $Y=1.157 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_187_n A_110_47# 0.00130295f $X=0.62 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_27_47#_c_185_n N_A_182_47#_c_389_n 6.34594e-19 $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_185_n N_VGND_c_408_n 0.00160048f $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_189_n N_VGND_c_408_n 0.0021406f $X=2.665 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_186_n N_VGND_c_410_n 0.00733679f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_190_n N_VGND_c_410_n 4.52338e-19 $X=3.12 $Y=1.157 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_187_n N_VGND_c_413_n 0.0292876f $X=0.62 $Y=0.825 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_185_n N_VGND_c_414_n 0.0054895f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_186_n N_VGND_c_414_n 0.0041289f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1003_s N_VGND_c_416_n 0.00213418f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_185_n N_VGND_c_416_n 0.00984571f $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_186_n N_VGND_c_416_n 0.00666209f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_187_n N_VGND_c_416_n 0.0217454f $X=0.62 $Y=0.825 $X2=0 $Y2=0
cc_200 N_VPWR_c_286_n A_373_297# 0.00897657f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_201 N_VPWR_c_286_n N_X_M1001_d 0.00395337f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_293_n N_X_c_367_n 0.0122897f $X=3.17 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_c_286_n N_X_c_367_n 0.0072038f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_M1009_s N_X_c_344_n 0.00453229f $X=3.195 $Y=1.485 $X2=0 $Y2=0
cc_205 N_VPWR_c_289_n N_X_c_344_n 7.8746e-19 $X=3.335 $Y=2.635 $X2=0 $Y2=0
cc_206 N_VPWR_c_290_n N_X_c_344_n 0.0207804f $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_207 N_VPWR_c_293_n N_X_c_344_n 0.00241807f $X=3.17 $Y=2.72 $X2=0 $Y2=0
cc_208 N_VPWR_c_286_n N_X_c_344_n 0.00692251f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_209 N_VPWR_M1009_s X 0.00714031f $X=3.195 $Y=1.485 $X2=0 $Y2=0
cc_210 N_X_c_347_n N_A_182_47#_c_389_n 0.00462652f $X=3.05 $Y=0.7 $X2=0 $Y2=0
cc_211 N_X_c_355_n N_VGND_M1010_s 0.00247753f $X=3.345 $Y=0.7 $X2=0 $Y2=0
cc_212 N_X_c_342_n N_VGND_M1010_s 0.00360841f $X=3.442 $Y=0.785 $X2=0 $Y2=0
cc_213 X N_VGND_M1010_s 0.00144837f $X=3.455 $Y=0.85 $X2=0 $Y2=0
cc_214 N_X_c_355_n N_VGND_c_410_n 0.00853376f $X=3.345 $Y=0.7 $X2=0 $Y2=0
cc_215 N_X_c_342_n N_VGND_c_410_n 0.0163593f $X=3.442 $Y=0.785 $X2=0 $Y2=0
cc_216 N_X_c_346_n N_VGND_c_414_n 0.0186595f $X=2.885 $Y=0.36 $X2=0 $Y2=0
cc_217 N_X_c_355_n N_VGND_c_414_n 0.0025909f $X=3.345 $Y=0.7 $X2=0 $Y2=0
cc_218 N_X_M1005_d N_VGND_c_416_n 0.00223231f $X=2.745 $Y=0.235 $X2=0 $Y2=0
cc_219 N_X_c_346_n N_VGND_c_416_n 0.0121874f $X=2.885 $Y=0.36 $X2=0 $Y2=0
cc_220 N_X_c_355_n N_VGND_c_416_n 0.00482796f $X=3.345 $Y=0.7 $X2=0 $Y2=0
cc_221 N_X_c_342_n N_VGND_c_416_n 0.00101974f $X=3.442 $Y=0.785 $X2=0 $Y2=0
cc_222 A_110_47# N_VGND_c_416_n 0.00357855f $X=0.55 $Y=0.235 $X2=0.402 $Y2=0.38
cc_223 N_A_182_47#_c_389_n N_VGND_M1002_s 0.0053917f $X=1.985 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_224 N_A_182_47#_c_389_n N_VGND_c_407_n 0.0211679f $X=1.985 $Y=0.73 $X2=0
+ $Y2=0
cc_225 N_A_182_47#_c_389_n N_VGND_c_411_n 0.00640861f $X=1.985 $Y=0.73 $X2=0
+ $Y2=0
cc_226 N_A_182_47#_c_389_n N_VGND_c_413_n 0.0086677f $X=1.985 $Y=0.73 $X2=0
+ $Y2=0
cc_227 N_A_182_47#_M1000_d N_VGND_c_416_n 0.00293129f $X=0.91 $Y=0.235 $X2=0
+ $Y2=0
cc_228 N_A_182_47#_M1002_d N_VGND_c_416_n 0.00326987f $X=1.845 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_182_47#_c_389_n N_VGND_c_416_n 0.0272545f $X=1.985 $Y=0.73 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__nand3_2.spice.SKY130_FD_SC_HD__NAND3_2.pxi
* Created: Thu Aug 27 14:29:32 2020
* 
x_PM_SKY130_FD_SC_HD__NAND3_2%A N_A_c_51_n N_A_M1003_g N_A_M1001_g N_A_c_52_n
+ N_A_M1011_g N_A_M1009_g A N_A_c_54_n PM_SKY130_FD_SC_HD__NAND3_2%A
x_PM_SKY130_FD_SC_HD__NAND3_2%B N_B_M1007_g N_B_M1000_g N_B_M1008_g N_B_M1010_g
+ B B B N_B_c_96_n PM_SKY130_FD_SC_HD__NAND3_2%B
x_PM_SKY130_FD_SC_HD__NAND3_2%C N_C_M1004_g N_C_M1002_g N_C_c_145_n N_C_M1005_g
+ N_C_M1006_g C C C N_C_c_147_n PM_SKY130_FD_SC_HD__NAND3_2%C
x_PM_SKY130_FD_SC_HD__NAND3_2%VPWR N_VPWR_M1001_d N_VPWR_M1009_d N_VPWR_M1010_s
+ N_VPWR_M1002_d N_VPWR_M1006_d N_VPWR_c_185_n N_VPWR_c_186_n N_VPWR_c_187_n
+ N_VPWR_c_188_n N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n N_VPWR_c_192_n
+ VPWR N_VPWR_c_193_n N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_184_n
+ PM_SKY130_FD_SC_HD__NAND3_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND3_2%Y N_Y_M1003_s N_Y_M1001_s N_Y_M1000_d N_Y_M1002_s
+ N_Y_c_238_n N_Y_c_234_n N_Y_c_241_n N_Y_c_235_n N_Y_c_236_n N_Y_c_273_n
+ N_Y_c_237_n Y Y Y N_Y_c_244_n PM_SKY130_FD_SC_HD__NAND3_2%Y
x_PM_SKY130_FD_SC_HD__NAND3_2%A_27_47# N_A_27_47#_M1003_d N_A_27_47#_M1011_d
+ N_A_27_47#_M1008_d N_A_27_47#_c_295_n N_A_27_47#_c_296_n N_A_27_47#_c_297_n
+ PM_SKY130_FD_SC_HD__NAND3_2%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND3_2%A_277_47# N_A_277_47#_M1007_s N_A_277_47#_M1004_s
+ N_A_277_47#_c_320_n PM_SKY130_FD_SC_HD__NAND3_2%A_277_47#
x_PM_SKY130_FD_SC_HD__NAND3_2%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_c_342_n
+ N_VGND_c_343_n N_VGND_c_344_n VGND N_VGND_c_345_n N_VGND_c_346_n
+ N_VGND_c_347_n N_VGND_c_348_n PM_SKY130_FD_SC_HD__NAND3_2%VGND
cc_1 VNB N_A_c_51_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_c_52_n 0.015775f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB A 0.0134856f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_c_54_n 0.0530586f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B_M1007_g 0.0171783f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_6 VNB N_B_M1008_g 0.023095f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_7 VNB B 0.00890492f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_8 VNB N_B_c_96_n 0.0439034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_M1004_g 0.0220124f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_C_c_145_n 0.0230864f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_11 VNB C 0.0173239f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_12 VNB N_C_c_147_n 0.0492903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_184_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_295_n 0.0123949f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_15 VNB N_A_27_47#_c_296_n 0.00754845f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_16 VNB N_A_27_47#_c_297_n 0.00218948f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_17 VNB N_A_277_47#_c_320_n 0.0188238f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_18 VNB N_VGND_c_342_n 0.00552463f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_19 VNB N_VGND_c_343_n 0.0122216f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_20 VNB N_VGND_c_344_n 0.0358663f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_21 VNB N_VGND_c_345_n 0.0568341f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_22 VNB N_VGND_c_346_n 0.0158029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_347_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_348_n 0.201479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_A_M1001_g 0.025289f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_26 VPB N_A_M1009_g 0.0178886f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_27 VPB A 0.00291996f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_28 VPB N_A_c_54_n 0.0145776f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_29 VPB N_B_M1000_g 0.0194051f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_B_M1010_g 0.0266409f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_31 VPB N_B_c_96_n 0.0077444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_C_M1002_g 0.0266409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_C_M1006_g 0.0255677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_C_c_147_n 0.00875185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_185_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_186_n 0.0421978f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_37 VPB N_VPWR_c_187_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_188_n 0.0154813f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_189_n 0.0121923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_190_n 0.0528375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_191_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_192_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_193_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_194_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_195_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_184_n 0.0424721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_Y_c_234_n 0.00504979f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_48 VPB N_Y_c_235_n 0.0133774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_236_n 0.00223596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_237_n 0.00223596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 N_A_c_52_n N_B_M1007_g 0.0266303f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_52 N_A_c_54_n N_B_M1000_g 0.0297974f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_c_54_n B 0.00172151f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_54 N_A_c_54_n N_B_c_96_n 0.0201984f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_M1001_g N_VPWR_c_186_n 0.00321527f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_56 A N_VPWR_c_186_n 0.0199082f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_57 N_A_c_54_n N_VPWR_c_186_n 0.00225479f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_M1009_g N_VPWR_c_187_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_191_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_60 N_A_M1009_g N_VPWR_c_191_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_VPWR_c_184_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1009_g N_VPWR_c_184_n 0.00952874f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_M1001_g N_Y_c_238_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_64 N_A_M1009_g N_Y_c_238_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A_M1009_g N_Y_c_234_n 0.0157539f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1009_g N_Y_c_241_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1001_g Y 0.00470531f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_M1009_g Y 0.00105585f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_c_51_n N_Y_c_244_n 0.0124534f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_M1001_g N_Y_c_244_n 0.00653865f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_c_52_n N_Y_c_244_n 0.00798831f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_M1009_g N_Y_c_244_n 0.00355958f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 A N_Y_c_244_n 0.0225908f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_54_n N_Y_c_244_n 0.0229317f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 A N_A_27_47#_c_295_n 0.016487f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_54_n N_A_27_47#_c_295_n 0.00210742f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_51_n N_A_27_47#_c_297_n 0.0119513f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_c_52_n N_A_27_47#_c_297_n 0.0115553f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_c_54_n N_A_27_47#_c_297_n 2.96193e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_52_n N_A_277_47#_c_320_n 7.8374e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_51_n N_VGND_c_345_n 0.00366111f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_c_52_n N_VGND_c_345_n 0.00366111f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_c_51_n N_VGND_c_348_n 0.00626998f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_c_52_n N_VGND_c_348_n 0.00526729f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_85 B C 0.0121848f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B_c_96_n C 7.25463e-19 $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_87 B N_C_c_147_n 7.96181e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_88 N_B_c_96_n N_C_c_147_n 0.00552895f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_M1000_g N_VPWR_c_187_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_90 N_B_M1010_g N_VPWR_c_188_n 0.0033532f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_91 N_B_M1000_g N_VPWR_c_193_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B_M1010_g N_VPWR_c_193_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_93 N_B_M1000_g N_VPWR_c_184_n 0.00952874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_94 N_B_M1010_g N_VPWR_c_184_n 0.0108276f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_95 N_B_M1000_g N_Y_c_238_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_96 N_B_M1000_g N_Y_c_234_n 0.0119784f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_97 B N_Y_c_234_n 0.0209622f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B_c_96_n N_Y_c_234_n 0.00136564f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B_M1000_g N_Y_c_241_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B_M1010_g N_Y_c_241_n 0.0145598f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B_M1010_g N_Y_c_235_n 0.0147646f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_102 B N_Y_c_235_n 0.0352704f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B_c_96_n N_Y_c_235_n 0.00409692f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B_M1000_g N_Y_c_237_n 0.00149073f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B_M1010_g N_Y_c_237_n 0.00149073f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_106 B N_Y_c_237_n 0.0266429f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_107 N_B_c_96_n N_Y_c_237_n 0.00211918f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_Y_c_244_n 0.00133499f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_109 N_B_M1000_g N_Y_c_244_n 6.84328e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_110 B N_Y_c_244_n 0.0135359f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B_c_96_n N_Y_c_244_n 7.12658e-19 $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B_M1007_g N_A_27_47#_c_297_n 0.00953845f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_113 N_B_M1008_g N_A_27_47#_c_297_n 0.00789149f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_114 B N_A_27_47#_c_297_n 0.00674409f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B_c_96_n N_A_27_47#_c_297_n 8.03025e-19 $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_A_277_47#_c_320_n 0.00570702f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_117 N_B_M1008_g N_A_277_47#_c_320_n 0.0145787f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_118 B N_A_277_47#_c_320_n 0.0604314f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B_c_96_n N_A_277_47#_c_320_n 0.00640359f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_M1008_g N_VGND_c_342_n 0.00294182f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_121 N_B_M1007_g N_VGND_c_345_n 0.00366111f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_122 N_B_M1008_g N_VGND_c_345_n 0.00366111f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_123 N_B_M1007_g N_VGND_c_348_n 0.00526729f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_124 N_B_M1008_g N_VGND_c_348_n 0.00656615f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_125 N_C_M1002_g N_VPWR_c_188_n 0.0033532f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C_M1006_g N_VPWR_c_190_n 0.0041701f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_127 C N_VPWR_c_190_n 0.0317849f $X=3.385 $Y=1.105 $X2=0 $Y2=0
cc_128 N_C_c_147_n N_VPWR_c_190_n 0.00310533f $X=3.09 $Y=1.162 $X2=0 $Y2=0
cc_129 N_C_M1002_g N_VPWR_c_194_n 0.00541359f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_130 N_C_M1006_g N_VPWR_c_194_n 0.00541359f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_131 N_C_M1002_g N_VPWR_c_184_n 0.0108276f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_132 N_C_M1006_g N_VPWR_c_184_n 0.0105526f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C_M1002_g N_Y_c_235_n 0.0147646f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_134 C N_Y_c_235_n 0.0180842f $X=3.385 $Y=1.105 $X2=0 $Y2=0
cc_135 N_C_M1002_g N_Y_c_236_n 0.00149073f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_136 N_C_M1006_g N_Y_c_236_n 0.00331821f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_137 C N_Y_c_236_n 0.0266429f $X=3.385 $Y=1.105 $X2=0 $Y2=0
cc_138 N_C_c_147_n N_Y_c_236_n 0.00211918f $X=3.09 $Y=1.162 $X2=0 $Y2=0
cc_139 N_C_M1002_g N_Y_c_273_n 0.0145598f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_140 N_C_M1006_g N_Y_c_273_n 0.00902485f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_141 N_C_M1004_g N_A_277_47#_c_320_n 0.0156437f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_142 N_C_c_145_n N_A_277_47#_c_320_n 0.0049431f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_143 C N_A_277_47#_c_320_n 0.0429619f $X=3.385 $Y=1.105 $X2=0 $Y2=0
cc_144 N_C_c_147_n N_A_277_47#_c_320_n 0.00213453f $X=3.09 $Y=1.162 $X2=0 $Y2=0
cc_145 N_C_M1004_g N_VGND_c_342_n 0.00966356f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_146 N_C_c_145_n N_VGND_c_342_n 0.00115704f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_147 N_C_c_145_n N_VGND_c_344_n 0.0031688f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_148 C N_VGND_c_344_n 0.0286184f $X=3.385 $Y=1.105 $X2=0 $Y2=0
cc_149 N_C_c_147_n N_VGND_c_344_n 0.00314863f $X=3.09 $Y=1.162 $X2=0 $Y2=0
cc_150 N_C_M1004_g N_VGND_c_346_n 0.00339367f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_151 N_C_c_145_n N_VGND_c_346_n 0.00553327f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_152 N_C_M1004_g N_VGND_c_348_n 0.00398704f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_153 N_C_c_145_n N_VGND_c_348_n 0.0106771f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_154 N_VPWR_c_184_n N_Y_M1001_s 0.00215201f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_184_n N_Y_M1000_d 0.00215201f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_184_n N_Y_M1002_s 0.00215201f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_191_n N_Y_c_238_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_184_n N_Y_c_238_n 0.0122217f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_M1009_d N_Y_c_234_n 0.00167154f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_160 N_VPWR_c_187_n N_Y_c_234_n 0.0129161f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_161 N_VPWR_c_193_n N_Y_c_241_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_162 N_VPWR_c_184_n N_Y_c_241_n 0.0122217f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_M1010_s N_Y_c_235_n 0.00296777f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_164 N_VPWR_M1002_d N_Y_c_235_n 0.00296777f $X=2.335 $Y=1.485 $X2=0 $Y2=0
cc_165 N_VPWR_c_188_n N_Y_c_235_n 0.0568271f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_166 N_VPWR_c_190_n N_Y_c_236_n 0.0109319f $X=3.33 $Y=1.66 $X2=0 $Y2=0
cc_167 N_VPWR_c_194_n N_Y_c_273_n 0.0189039f $X=3.215 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_c_184_n N_Y_c_273_n 0.0122217f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_169 N_Y_M1003_s N_A_27_47#_c_297_n 0.00315577f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_170 N_Y_c_244_n N_A_27_47#_c_297_n 0.0160806f $X=0.68 $Y=0.72 $X2=0 $Y2=0
cc_171 N_Y_c_235_n N_A_277_47#_c_320_n 0.0110697f $X=2.715 $Y=1.555 $X2=0 $Y2=0
cc_172 N_Y_c_244_n N_A_277_47#_c_320_n 0.00869467f $X=0.68 $Y=0.72 $X2=0 $Y2=0
cc_173 N_Y_M1003_s N_VGND_c_348_n 0.00219239f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_297_n N_A_277_47#_M1007_s 0.00316446f $X=1.94 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_175 N_A_27_47#_M1008_d N_A_277_47#_c_320_n 0.00321334f $X=1.805 $Y=0.235
+ $X2=0 $Y2=0
cc_176 N_A_27_47#_c_297_n N_A_277_47#_c_320_n 0.0404245f $X=1.94 $Y=0.38 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_297_n N_VGND_c_342_n 0.0137364f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_296_n N_VGND_c_345_n 0.0138017f $X=0.345 $Y=0.38 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_297_n N_VGND_c_345_n 0.0780943f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1003_d N_VGND_c_348_n 0.00212393f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1011_d N_VGND_c_348_n 0.00217615f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1008_d N_VGND_c_348_n 0.00211652f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_296_n N_VGND_c_348_n 0.00953535f $X=0.345 $Y=0.38 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_297_n N_VGND_c_348_n 0.0609594f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_185 N_A_277_47#_c_320_n N_VGND_M1004_d 0.00320842f $X=2.88 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_186 N_A_277_47#_c_320_n N_VGND_c_342_n 0.0212463f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_187 N_A_277_47#_c_320_n N_VGND_c_345_n 0.00358f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_188 N_A_277_47#_c_320_n N_VGND_c_346_n 0.00643568f $X=2.88 $Y=0.72 $X2=0
+ $Y2=0
cc_189 N_A_277_47#_M1007_s N_VGND_c_348_n 0.00219239f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_190 N_A_277_47#_M1004_s N_VGND_c_348_n 0.00315309f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_191 N_A_277_47#_c_320_n N_VGND_c_348_n 0.0199318f $X=2.88 $Y=0.72 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o2bb2a_1.spice.SKY130_FD_SC_HD__O2BB2A_1.pxi
* Created: Thu Aug 27 14:38:13 2020
* 
x_PM_SKY130_FD_SC_HD__O2BB2A_1%A_76_199# N_A_76_199#_M1002_s N_A_76_199#_M1008_d
+ N_A_76_199#_M1009_g N_A_76_199#_M1003_g N_A_76_199#_c_76_n N_A_76_199#_c_77_n
+ N_A_76_199#_c_86_n N_A_76_199#_c_94_p N_A_76_199#_c_147_p N_A_76_199#_c_78_n
+ N_A_76_199#_c_88_n N_A_76_199#_c_79_n N_A_76_199#_c_80_n N_A_76_199#_c_81_n
+ N_A_76_199#_c_89_n N_A_76_199#_c_82_n PM_SKY130_FD_SC_HD__O2BB2A_1%A_76_199#
x_PM_SKY130_FD_SC_HD__O2BB2A_1%A1_N N_A1_N_M1001_g N_A1_N_M1005_g A1_N
+ N_A1_N_c_175_n A1_N PM_SKY130_FD_SC_HD__O2BB2A_1%A1_N
x_PM_SKY130_FD_SC_HD__O2BB2A_1%A2_N N_A2_N_M1010_g N_A2_N_M1011_g N_A2_N_c_213_n
+ N_A2_N_c_214_n A2_N N_A2_N_c_216_n PM_SKY130_FD_SC_HD__O2BB2A_1%A2_N
x_PM_SKY130_FD_SC_HD__O2BB2A_1%A_206_369# N_A_206_369#_M1010_d
+ N_A_206_369#_M1005_d N_A_206_369#_M1002_g N_A_206_369#_M1008_g
+ N_A_206_369#_c_262_n N_A_206_369#_c_263_n N_A_206_369#_c_264_n
+ N_A_206_369#_c_258_n N_A_206_369#_c_265_n N_A_206_369#_c_259_n
+ PM_SKY130_FD_SC_HD__O2BB2A_1%A_206_369#
x_PM_SKY130_FD_SC_HD__O2BB2A_1%B2 N_B2_M1000_g N_B2_M1004_g N_B2_c_328_n
+ N_B2_c_329_n B2 PM_SKY130_FD_SC_HD__O2BB2A_1%B2
x_PM_SKY130_FD_SC_HD__O2BB2A_1%B1 N_B1_M1007_g N_B1_M1006_g B1 B1 N_B1_c_380_n
+ PM_SKY130_FD_SC_HD__O2BB2A_1%B1
x_PM_SKY130_FD_SC_HD__O2BB2A_1%X N_X_M1009_s N_X_M1003_s N_X_c_405_n N_X_c_406_n
+ N_X_c_408_n N_X_c_407_n X N_X_c_410_n PM_SKY130_FD_SC_HD__O2BB2A_1%X
x_PM_SKY130_FD_SC_HD__O2BB2A_1%VPWR N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_M1006_d
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n VPWR N_VPWR_c_432_n
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_428_n
+ PM_SKY130_FD_SC_HD__O2BB2A_1%VPWR
x_PM_SKY130_FD_SC_HD__O2BB2A_1%VGND N_VGND_M1009_d N_VGND_M1000_d N_VGND_c_479_n
+ N_VGND_c_480_n VGND N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n
+ N_VGND_c_484_n N_VGND_c_485_n VGND PM_SKY130_FD_SC_HD__O2BB2A_1%VGND
x_PM_SKY130_FD_SC_HD__O2BB2A_1%A_489_47# N_A_489_47#_M1002_d N_A_489_47#_M1007_d
+ N_A_489_47#_c_533_n N_A_489_47#_c_534_n N_A_489_47#_c_535_n
+ N_A_489_47#_c_536_n PM_SKY130_FD_SC_HD__O2BB2A_1%A_489_47#
cc_1 VNB N_A_76_199#_c_76_n 0.00209149f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_2 VNB N_A_76_199#_c_77_n 0.0249244f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_3 VNB N_A_76_199#_c_78_n 5.22012e-19 $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.495
cc_4 VNB N_A_76_199#_c_79_n 0.00159549f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=0.485
cc_5 VNB N_A_76_199#_c_80_n 0.00320094f $X=-0.19 $Y=-0.24 $X2=2.252 $Y2=1.075
cc_6 VNB N_A_76_199#_c_81_n 0.00163916f $X=-0.19 $Y=-0.24 $X2=2.252 $Y2=1.245
cc_7 VNB N_A_76_199#_c_82_n 0.0200211f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_8 VNB N_A1_N_M1001_g 0.0304778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A1_N_c_175_n 0.0219021f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_10 VNB A1_N 0.00845745f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=1.885
cc_11 VNB N_A2_N_M1011_g 0.0133632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_N_c_213_n 0.00749846f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_A2_N_c_214_n 0.0333679f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_14 VNB A2_N 0.00142945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_N_c_216_n 0.0203025f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_16 VNB N_A_206_369#_M1002_g 0.0507849f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_17 VNB N_A_206_369#_c_258_n 0.0035652f $X=-0.19 $Y=-0.24 $X2=2.18 $Y2=1.97
cc_18 VNB N_A_206_369#_c_259_n 0.0138337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B2_M1000_g 0.0262349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B2_c_328_n 0.00540798f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_B2_c_329_n 0.0191226f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_22 VNB N_B1_M1007_g 0.0353006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB B1 0.00879609f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_24 VNB N_B1_c_380_n 0.0371837f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_25 VNB N_X_c_405_n 0.0160045f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_26 VNB N_X_c_406_n 0.00666696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_407_n 0.0218906f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_28 VNB N_VPWR_c_428_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_479_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_30 VNB N_VGND_c_480_n 0.00465965f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_31 VNB N_VGND_c_481_n 0.0573914f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=1.615
cc_32 VNB N_VGND_c_482_n 0.0176368f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.495
cc_33 VNB N_VGND_c_483_n 0.206474f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.53
cc_34 VNB N_VGND_c_484_n 0.0218339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_485_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_489_47#_c_533_n 4.75015e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_37 VNB N_A_489_47#_c_534_n 0.0165829f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_38 VNB N_A_489_47#_c_535_n 0.0032687f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_39 VNB N_A_489_47#_c_536_n 0.0164468f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_40 VPB N_A_76_199#_M1003_g 0.0234903f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_41 VPB N_A_76_199#_c_76_n 0.00141115f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_42 VPB N_A_76_199#_c_77_n 0.00487854f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_43 VPB N_A_76_199#_c_86_n 0.00184058f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.885
cc_44 VPB N_A_76_199#_c_78_n 4.42383e-19 $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.495
cc_45 VPB N_A_76_199#_c_88_n 0.00654296f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.53
cc_46 VPB N_A_76_199#_c_89_n 0.0127023f $X=-0.19 $Y=1.305 $X2=2.457 $Y2=1.97
cc_47 VPB N_A1_N_M1005_g 0.0417858f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_48 VPB N_A1_N_c_175_n 0.00437618f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_49 VPB N_A2_N_M1011_g 0.0424025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_206_369#_M1002_g 0.00287016f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_51 VPB N_A_206_369#_M1008_g 0.0209895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_206_369#_c_262_n 0.0508909f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_53 VPB N_A_206_369#_c_263_n 0.0118636f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_54 VPB N_A_206_369#_c_264_n 0.00879907f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_55 VPB N_A_206_369#_c_265_n 0.00849895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_206_369#_c_259_n 8.55232e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_B2_M1004_g 0.0343524f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_58 VPB N_B2_c_328_n 0.00147058f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_59 VPB N_B2_c_329_n 0.00515335f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_60 VPB B2 0.00697362f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_61 VPB N_B1_M1006_g 0.0465954f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_62 VPB B1 0.0162957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_63 VPB N_B1_c_380_n 0.0101292f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_64 VPB N_X_c_408_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.445
cc_65 VPB N_X_c_407_n 0.0195702f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_66 VPB N_X_c_410_n 0.0208429f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.615
cc_67 VPB N_VPWR_c_429_n 0.00763275f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_68 VPB N_VPWR_c_430_n 0.0115225f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.445
cc_69 VPB N_VPWR_c_431_n 0.0366441f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_70 VPB N_VPWR_c_432_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.885
cc_71 VPB N_VPWR_c_433_n 0.0240162f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.245
cc_72 VPB N_VPWR_c_434_n 0.0311407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_435_n 0.00507288f $X=-0.19 $Y=1.305 $X2=2.252 $Y2=1.245
cc_74 VPB N_VPWR_c_436_n 0.0153178f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=2.06
cc_75 VPB N_VPWR_c_428_n 0.0690716f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 N_A_76_199#_c_82_n N_A1_N_M1001_g 0.0187727f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_76_199#_M1003_g N_A1_N_M1005_g 0.028566f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_76_199#_c_76_n N_A1_N_M1005_g 0.00222807f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_76_199#_c_86_n N_A1_N_M1005_g 0.00415725f $X=0.74 $Y=1.885 $X2=0 $Y2=0
cc_80 N_A_76_199#_c_94_p N_A1_N_M1005_g 0.0135408f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_81 N_A_76_199#_c_88_n N_A1_N_M1005_g 0.002419f $X=0.74 $Y=1.53 $X2=0 $Y2=0
cc_82 N_A_76_199#_c_76_n N_A1_N_c_175_n 0.00102065f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_76_199#_c_77_n N_A1_N_c_175_n 0.0208346f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_76_199#_c_76_n A1_N 0.0154185f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_76_199#_c_77_n A1_N 0.00124474f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_76_199#_c_94_p A1_N 0.00353597f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_87 N_A_76_199#_c_88_n A1_N 0.00419335f $X=0.74 $Y=1.53 $X2=0 $Y2=0
cc_88 N_A_76_199#_c_94_p N_A2_N_M1011_g 0.0142668f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_89 N_A_76_199#_c_89_n N_A2_N_M1011_g 0.00433229f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_90 N_A_76_199#_c_94_p N_A_206_369#_M1005_d 0.00853544f $X=2.18 $Y=1.97 $X2=0
+ $Y2=0
cc_91 N_A_76_199#_c_78_n N_A_206_369#_M1002_g 0.0029694f $X=2.265 $Y=1.495 $X2=0
+ $Y2=0
cc_92 N_A_76_199#_c_79_n N_A_206_369#_M1002_g 0.00482007f $X=2.16 $Y=0.485 $X2=0
+ $Y2=0
cc_93 N_A_76_199#_c_80_n N_A_206_369#_M1002_g 0.0105559f $X=2.252 $Y=1.075 $X2=0
+ $Y2=0
cc_94 N_A_76_199#_c_81_n N_A_206_369#_M1002_g 0.00564727f $X=2.252 $Y=1.245
+ $X2=0 $Y2=0
cc_95 N_A_76_199#_c_89_n N_A_206_369#_M1008_g 0.0267396f $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_96 N_A_76_199#_c_94_p N_A_206_369#_c_262_n 0.00738394f $X=2.18 $Y=1.97 $X2=0
+ $Y2=0
cc_97 N_A_76_199#_c_78_n N_A_206_369#_c_262_n 0.00610077f $X=2.265 $Y=1.495
+ $X2=0 $Y2=0
cc_98 N_A_76_199#_c_79_n N_A_206_369#_c_262_n 0.00194568f $X=2.16 $Y=0.485 $X2=0
+ $Y2=0
cc_99 N_A_76_199#_c_81_n N_A_206_369#_c_262_n 7.75851e-19 $X=2.252 $Y=1.245
+ $X2=0 $Y2=0
cc_100 N_A_76_199#_c_89_n N_A_206_369#_c_262_n 0.0070745f $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_101 N_A_76_199#_c_78_n N_A_206_369#_c_263_n 0.00280991f $X=2.265 $Y=1.495
+ $X2=0 $Y2=0
cc_102 N_A_76_199#_c_89_n N_A_206_369#_c_263_n 0.0101471f $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_103 N_A_76_199#_c_86_n N_A_206_369#_c_264_n 0.00791067f $X=0.74 $Y=1.885
+ $X2=0 $Y2=0
cc_104 N_A_76_199#_c_94_p N_A_206_369#_c_264_n 0.0481175f $X=2.18 $Y=1.97 $X2=0
+ $Y2=0
cc_105 N_A_76_199#_c_88_n N_A_206_369#_c_264_n 0.0100855f $X=0.74 $Y=1.53 $X2=0
+ $Y2=0
cc_106 N_A_76_199#_c_79_n N_A_206_369#_c_258_n 0.0140162f $X=2.16 $Y=0.485 $X2=0
+ $Y2=0
cc_107 N_A_76_199#_c_94_p N_A_206_369#_c_265_n 0.0222516f $X=2.18 $Y=1.97 $X2=0
+ $Y2=0
cc_108 N_A_76_199#_c_78_n N_A_206_369#_c_265_n 0.00981918f $X=2.265 $Y=1.495
+ $X2=0 $Y2=0
cc_109 N_A_76_199#_c_89_n N_A_206_369#_c_265_n 0.0173032f $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_110 N_A_76_199#_c_78_n N_A_206_369#_c_259_n 0.00587538f $X=2.265 $Y=1.495
+ $X2=0 $Y2=0
cc_111 N_A_76_199#_c_79_n N_A_206_369#_c_259_n 0.00952847f $X=2.16 $Y=0.485
+ $X2=0 $Y2=0
cc_112 N_A_76_199#_c_80_n N_A_206_369#_c_259_n 0.0319876f $X=2.252 $Y=1.075
+ $X2=0 $Y2=0
cc_113 N_A_76_199#_c_79_n N_B2_M1000_g 2.89703e-19 $X=2.16 $Y=0.485 $X2=0 $Y2=0
cc_114 N_A_76_199#_c_80_n N_B2_M1000_g 4.47008e-19 $X=2.252 $Y=1.075 $X2=0 $Y2=0
cc_115 N_A_76_199#_c_78_n N_B2_M1004_g 5.4127e-19 $X=2.265 $Y=1.495 $X2=0 $Y2=0
cc_116 N_A_76_199#_c_89_n N_B2_M1004_g 0.00337876f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_117 N_A_76_199#_c_81_n N_B2_c_328_n 0.019763f $X=2.252 $Y=1.245 $X2=0 $Y2=0
cc_118 N_A_76_199#_c_89_n N_B2_c_328_n 0.018331f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_119 N_A_76_199#_c_80_n N_B2_c_329_n 4.28224e-19 $X=2.252 $Y=1.075 $X2=0 $Y2=0
cc_120 N_A_76_199#_c_81_n N_B2_c_329_n 2.07654e-19 $X=2.252 $Y=1.245 $X2=0 $Y2=0
cc_121 N_A_76_199#_c_89_n N_B2_c_329_n 0.00194254f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_122 N_A_76_199#_c_78_n B2 0.00432844f $X=2.265 $Y=1.495 $X2=0 $Y2=0
cc_123 N_A_76_199#_c_89_n B2 0.0439761f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_124 N_A_76_199#_c_82_n N_X_c_405_n 0.00467408f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_76_199#_c_82_n N_X_c_406_n 0.00396702f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_76_199#_M1003_g N_X_c_407_n 0.00931762f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_76_199#_c_76_n N_X_c_407_n 0.0322249f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_76_199#_c_77_n N_X_c_407_n 0.00753785f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_76_199#_c_86_n N_X_c_407_n 0.00701428f $X=0.74 $Y=1.885 $X2=0 $Y2=0
cc_130 N_A_76_199#_c_88_n N_X_c_407_n 0.0127214f $X=0.74 $Y=1.53 $X2=0 $Y2=0
cc_131 N_A_76_199#_c_82_n N_X_c_407_n 0.00497708f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_76_199#_c_86_n N_VPWR_M1003_d 0.00409302f $X=0.74 $Y=1.885 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_76_199#_c_147_p N_VPWR_M1003_d 0.00409058f $X=0.825 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_76_199#_c_88_n N_VPWR_M1003_d 0.00204498f $X=0.74 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_76_199#_c_94_p N_VPWR_M1011_d 0.0156704f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_136 N_A_76_199#_c_89_n N_VPWR_M1011_d 0.00205965f $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_137 N_A_76_199#_M1003_g N_VPWR_c_429_n 0.0100884f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_76_199#_c_147_p N_VPWR_c_429_n 0.0131715f $X=0.825 $Y=1.97 $X2=0
+ $Y2=0
cc_139 N_A_76_199#_c_88_n N_VPWR_c_429_n 0.00236443f $X=0.74 $Y=1.53 $X2=0 $Y2=0
cc_140 N_A_76_199#_M1003_g N_VPWR_c_432_n 0.0046653f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_76_199#_c_94_p N_VPWR_c_433_n 0.0124071f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_142 N_A_76_199#_c_94_p N_VPWR_c_434_n 0.00105858f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_143 N_A_76_199#_c_89_n N_VPWR_c_434_n 0.014428f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_144 N_A_76_199#_c_94_p N_VPWR_c_436_n 0.0291396f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_145 N_A_76_199#_c_89_n N_VPWR_c_436_n 0.00288761f $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_146 N_A_76_199#_M1003_g N_VPWR_c_428_n 0.008846f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_76_199#_c_94_p N_VPWR_c_428_n 0.0274652f $X=2.18 $Y=1.97 $X2=0 $Y2=0
cc_148 N_A_76_199#_c_147_p N_VPWR_c_428_n 7.95799e-19 $X=0.825 $Y=1.97 $X2=0
+ $Y2=0
cc_149 N_A_76_199#_c_89_n N_VPWR_c_428_n 0.017916f $X=2.457 $Y=1.97 $X2=0 $Y2=0
cc_150 N_A_76_199#_c_77_n N_VGND_c_479_n 0.00118907f $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_76_199#_c_82_n N_VGND_c_479_n 0.00505437f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_76_199#_c_79_n N_VGND_c_481_n 0.0106847f $X=2.16 $Y=0.485 $X2=0 $Y2=0
cc_153 N_A_76_199#_M1002_s N_VGND_c_483_n 0.00356607f $X=2.035 $Y=0.235 $X2=0
+ $Y2=0
cc_154 N_A_76_199#_c_79_n N_VGND_c_483_n 0.00903149f $X=2.16 $Y=0.485 $X2=0
+ $Y2=0
cc_155 N_A_76_199#_c_82_n N_VGND_c_483_n 0.0107684f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_156 N_A_76_199#_c_82_n N_VGND_c_484_n 0.00541359f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_76_199#_c_79_n N_A_489_47#_c_533_n 0.01717f $X=2.16 $Y=0.485 $X2=0
+ $Y2=0
cc_158 N_A_76_199#_c_80_n N_A_489_47#_c_535_n 0.0145208f $X=2.252 $Y=1.075 $X2=0
+ $Y2=0
cc_159 N_A_76_199#_c_89_n N_A_489_47#_c_535_n 9.70378e-19 $X=2.457 $Y=1.97 $X2=0
+ $Y2=0
cc_160 N_A1_N_M1005_g N_A2_N_M1011_g 0.0334182f $X=0.955 $Y=2.055 $X2=0 $Y2=0
cc_161 N_A1_N_c_175_n N_A2_N_M1011_g 0.00883344f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_162 A1_N N_A2_N_M1011_g 0.00174185f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_163 N_A1_N_M1001_g N_A2_N_c_213_n 0.00427236f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A1_N_c_175_n N_A2_N_c_213_n 0.00205827f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_165 A1_N N_A2_N_c_213_n 0.014196f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_166 N_A1_N_c_175_n N_A2_N_c_214_n 0.00686264f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A1_N_M1001_g A2_N 0.00205785f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A1_N_M1001_g N_A2_N_c_216_n 0.0317576f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A1_N_M1005_g N_A_206_369#_c_264_n 0.00676621f $X=0.955 $Y=2.055 $X2=0
+ $Y2=0
cc_170 N_A1_N_c_175_n N_A_206_369#_c_264_n 0.00231747f $X=0.995 $Y=1.16 $X2=0
+ $Y2=0
cc_171 A1_N N_A_206_369#_c_264_n 0.0137592f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_172 A1_N N_A_206_369#_c_259_n 0.00652704f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_173 N_A1_N_M1001_g N_X_c_405_n 3.76391e-19 $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A1_N_M1005_g N_VPWR_c_429_n 0.00383984f $X=0.955 $Y=2.055 $X2=0 $Y2=0
cc_175 N_A1_N_M1005_g N_VPWR_c_433_n 0.00399288f $X=0.955 $Y=2.055 $X2=0 $Y2=0
cc_176 N_A1_N_M1005_g N_VPWR_c_428_n 0.00515951f $X=0.955 $Y=2.055 $X2=0 $Y2=0
cc_177 N_A1_N_M1001_g N_VGND_c_479_n 0.00767959f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_178 A1_N N_VGND_c_479_n 9.9771e-19 $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_179 N_A1_N_M1001_g N_VGND_c_481_n 0.00585385f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A1_N_M1001_g N_VGND_c_483_n 0.0110899f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A2_N_M1011_g N_A_206_369#_M1002_g 0.00219371f $X=1.505 $Y=2.055 $X2=0
+ $Y2=0
cc_182 N_A2_N_c_214_n N_A_206_369#_M1002_g 0.00342924f $X=1.475 $Y=0.935 $X2=0
+ $Y2=0
cc_183 N_A2_N_M1011_g N_A_206_369#_c_262_n 0.0206112f $X=1.505 $Y=2.055 $X2=0
+ $Y2=0
cc_184 N_A2_N_M1011_g N_A_206_369#_c_264_n 0.0137222f $X=1.505 $Y=2.055 $X2=0
+ $Y2=0
cc_185 N_A2_N_c_213_n N_A_206_369#_c_264_n 0.0120011f $X=1.18 $Y=0.905 $X2=0
+ $Y2=0
cc_186 N_A2_N_c_214_n N_A_206_369#_c_264_n 0.00294298f $X=1.475 $Y=0.935 $X2=0
+ $Y2=0
cc_187 N_A2_N_c_213_n N_A_206_369#_c_258_n 0.00567122f $X=1.18 $Y=0.905 $X2=0
+ $Y2=0
cc_188 N_A2_N_c_214_n N_A_206_369#_c_258_n 0.00276509f $X=1.475 $Y=0.935 $X2=0
+ $Y2=0
cc_189 N_A2_N_c_216_n N_A_206_369#_c_258_n 0.00259127f $X=1.485 $Y=0.77 $X2=0
+ $Y2=0
cc_190 N_A2_N_M1011_g N_A_206_369#_c_265_n 3.07985e-19 $X=1.505 $Y=2.055 $X2=0
+ $Y2=0
cc_191 N_A2_N_M1011_g N_A_206_369#_c_259_n 0.00749157f $X=1.505 $Y=2.055 $X2=0
+ $Y2=0
cc_192 N_A2_N_c_213_n N_A_206_369#_c_259_n 0.0274487f $X=1.18 $Y=0.905 $X2=0
+ $Y2=0
cc_193 N_A2_N_c_214_n N_A_206_369#_c_259_n 0.00379772f $X=1.475 $Y=0.935 $X2=0
+ $Y2=0
cc_194 A2_N N_A_206_369#_c_259_n 0.00468916f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_195 N_A2_N_c_216_n N_A_206_369#_c_259_n 0.00220315f $X=1.485 $Y=0.77 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_213_n N_X_c_406_n 0.00221845f $X=1.18 $Y=0.905 $X2=0 $Y2=0
cc_197 N_A2_N_M1011_g N_VPWR_c_433_n 0.00399288f $X=1.505 $Y=2.055 $X2=0 $Y2=0
cc_198 N_A2_N_M1011_g N_VPWR_c_436_n 0.00631619f $X=1.505 $Y=2.055 $X2=0 $Y2=0
cc_199 N_A2_N_M1011_g N_VPWR_c_428_n 0.00515951f $X=1.505 $Y=2.055 $X2=0 $Y2=0
cc_200 N_A2_N_c_213_n N_VGND_c_479_n 8.48044e-19 $X=1.18 $Y=0.905 $X2=0 $Y2=0
cc_201 A2_N N_VGND_c_479_n 0.0110811f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_202 N_A2_N_c_213_n N_VGND_c_481_n 0.00237499f $X=1.18 $Y=0.905 $X2=0 $Y2=0
cc_203 A2_N N_VGND_c_481_n 0.00799532f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_204 N_A2_N_c_216_n N_VGND_c_481_n 0.0042834f $X=1.485 $Y=0.77 $X2=0 $Y2=0
cc_205 N_A2_N_c_213_n N_VGND_c_483_n 0.00411065f $X=1.18 $Y=0.905 $X2=0 $Y2=0
cc_206 A2_N N_VGND_c_483_n 0.00776053f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_207 N_A2_N_c_216_n N_VGND_c_483_n 0.0074896f $X=1.485 $Y=0.77 $X2=0 $Y2=0
cc_208 A2_N A_205_47# 0.00485199f $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_209 N_A_206_369#_M1002_g N_B2_M1000_g 0.0241959f $X=2.37 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A_206_369#_M1002_g N_B2_M1004_g 0.0082645f $X=2.37 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A_206_369#_c_263_n N_B2_M1004_g 0.015148f $X=2.295 $Y=1.355 $X2=0 $Y2=0
cc_212 N_A_206_369#_M1002_g N_B2_c_328_n 0.00164172f $X=2.37 $Y=0.445 $X2=0
+ $Y2=0
cc_213 N_A_206_369#_M1002_g N_B2_c_329_n 0.0197416f $X=2.37 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A_206_369#_M1002_g B2 6.34431e-19 $X=2.37 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A_206_369#_M1008_g B2 5.0288e-19 $X=2.38 $Y=2.055 $X2=0 $Y2=0
cc_216 N_A_206_369#_c_263_n B2 3.82539e-19 $X=2.295 $Y=1.355 $X2=0 $Y2=0
cc_217 N_A_206_369#_M1008_g N_VPWR_c_434_n 0.00391775f $X=2.38 $Y=2.055 $X2=0
+ $Y2=0
cc_218 N_A_206_369#_M1008_g N_VPWR_c_436_n 0.00504353f $X=2.38 $Y=2.055 $X2=0
+ $Y2=0
cc_219 N_A_206_369#_M1008_g N_VPWR_c_428_n 0.00515951f $X=2.38 $Y=2.055 $X2=0
+ $Y2=0
cc_220 N_A_206_369#_M1002_g N_VGND_c_481_n 0.00543919f $X=2.37 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_206_369#_c_258_n N_VGND_c_481_n 0.0147327f $X=1.735 $Y=0.48 $X2=0
+ $Y2=0
cc_222 N_A_206_369#_M1010_d N_VGND_c_483_n 0.00228543f $X=1.49 $Y=0.235 $X2=0
+ $Y2=0
cc_223 N_A_206_369#_M1002_g N_VGND_c_483_n 0.0111506f $X=2.37 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_206_369#_c_258_n N_VGND_c_483_n 0.0152259f $X=1.735 $Y=0.48 $X2=0
+ $Y2=0
cc_225 N_A_206_369#_M1002_g N_A_489_47#_c_533_n 4.96975e-19 $X=2.37 $Y=0.445
+ $X2=0 $Y2=0
cc_226 N_A_206_369#_M1002_g N_A_489_47#_c_535_n 0.00144502f $X=2.37 $Y=0.445
+ $X2=0 $Y2=0
cc_227 N_B2_M1000_g N_B1_M1007_g 0.0258694f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_228 N_B2_M1004_g N_B1_M1006_g 0.0419621f $X=2.85 $Y=2.055 $X2=0 $Y2=0
cc_229 B2 N_B1_M1006_g 0.00817501f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_230 N_B2_c_328_n B1 0.0208119f $X=2.905 $Y=1.2 $X2=0 $Y2=0
cc_231 N_B2_c_329_n B1 4.4849e-19 $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_232 B2 B1 0.0241065f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_233 N_B2_c_328_n N_B1_c_380_n 0.00195313f $X=2.905 $Y=1.2 $X2=0 $Y2=0
cc_234 N_B2_c_329_n N_B1_c_380_n 0.0419621f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B2_M1004_g N_VPWR_c_431_n 4.59283e-19 $X=2.85 $Y=2.055 $X2=0 $Y2=0
cc_236 B2 N_VPWR_c_431_n 0.0302744f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_237 N_B2_M1004_g N_VPWR_c_434_n 0.00462297f $X=2.85 $Y=2.055 $X2=0 $Y2=0
cc_238 B2 N_VPWR_c_434_n 0.00989629f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_239 N_B2_M1004_g N_VPWR_c_428_n 0.00450597f $X=2.85 $Y=2.055 $X2=0 $Y2=0
cc_240 B2 N_VPWR_c_428_n 0.00653087f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_241 N_B2_M1000_g N_VGND_c_480_n 0.00268723f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_242 N_B2_M1000_g N_VGND_c_481_n 0.00425893f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_243 N_B2_M1000_g N_VGND_c_483_n 0.00581681f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_244 N_B2_M1000_g N_A_489_47#_c_533_n 0.00631178f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_245 N_B2_M1000_g N_A_489_47#_c_534_n 0.00865686f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_246 N_B2_c_328_n N_A_489_47#_c_534_n 0.0260516f $X=2.905 $Y=1.2 $X2=0 $Y2=0
cc_247 N_B2_c_329_n N_A_489_47#_c_534_n 0.00173849f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B2_M1000_g N_A_489_47#_c_535_n 0.00249874f $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_249 N_B2_c_328_n N_A_489_47#_c_535_n 0.0187917f $X=2.905 $Y=1.2 $X2=0 $Y2=0
cc_250 N_B2_c_329_n N_A_489_47#_c_535_n 0.0015306f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B2_M1000_g N_A_489_47#_c_536_n 5.02919e-19 $X=2.79 $Y=0.445 $X2=0 $Y2=0
cc_252 N_B1_M1006_g N_VPWR_c_431_n 0.0112773f $X=3.21 $Y=2.055 $X2=0 $Y2=0
cc_253 B1 N_VPWR_c_431_n 0.0314133f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_254 N_B1_c_380_n N_VPWR_c_431_n 0.00115968f $X=3.415 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B1_M1006_g N_VPWR_c_434_n 0.00395287f $X=3.21 $Y=2.055 $X2=0 $Y2=0
cc_256 N_B1_M1006_g N_VPWR_c_428_n 0.00399002f $X=3.21 $Y=2.055 $X2=0 $Y2=0
cc_257 N_B1_M1007_g N_VGND_c_480_n 0.00268723f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_258 N_B1_M1007_g N_VGND_c_482_n 0.00425893f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_259 N_B1_M1007_g N_VGND_c_483_n 0.00677018f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_260 N_B1_M1007_g N_A_489_47#_c_533_n 5.04494e-19 $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_261 N_B1_M1007_g N_A_489_47#_c_534_n 0.0168974f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_262 B1 N_A_489_47#_c_534_n 0.0294383f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_263 N_B1_c_380_n N_A_489_47#_c_534_n 0.00739251f $X=3.415 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_M1007_g N_A_489_47#_c_536_n 0.00762625f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_265 N_X_c_410_n N_VPWR_c_432_n 0.0179951f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_266 N_X_M1003_s N_VPWR_c_428_n 0.00382897f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_267 N_X_c_410_n N_VPWR_c_428_n 0.00993477f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_268 N_X_c_405_n N_VGND_c_479_n 0.0329192f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_269 N_X_M1009_s N_VGND_c_483_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_270 N_X_c_405_n N_VGND_c_483_n 0.0127834f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_271 N_X_c_405_n N_VGND_c_484_n 0.0216607f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_272 N_VGND_c_483_n A_205_47# 0.00449915f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_273 N_VGND_c_483_n N_A_489_47#_M1002_d 0.00398008f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_274 N_VGND_c_483_n N_A_489_47#_M1007_d 0.00214228f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_481_n N_A_489_47#_c_533_n 0.0106087f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_483_n N_A_489_47#_c_533_n 0.00904216f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_480_n N_A_489_47#_c_534_n 0.0128746f $X=3 $Y=0.39 $X2=0 $Y2=0
cc_278 N_VGND_c_481_n N_A_489_47#_c_534_n 0.00236451f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_482_n N_A_489_47#_c_534_n 0.00236451f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_483_n N_A_489_47#_c_534_n 0.00835832f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_482_n N_A_489_47#_c_536_n 0.0152149f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_483_n N_A_489_47#_c_536_n 0.0123194f $X=3.45 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__sdfxtp_2.spice
* Created: Thu Aug 27 14:47:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfxtp_2.pex.spice"
.subckt sky130_fd_sc_hd__sdfxtp_2  VNB VPB CLK SCE D SCD VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SCD	SCD
* D	D
* SCE	SCE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_CLK_M1031_g N_A_27_47#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_193_47#_M1018_d N_A_27_47#_M1018_g N_VGND_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_SCE_M1032_g N_A_299_47#_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07455 AS=0.1176 PD=0.775 PS=1.4 NRD=21.42 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1021 A_486_47# N_A_299_47#_M1021_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.07455 PD=0.66 PS=0.775 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1022 N_A_559_369#_M1022_d N_D_M1022_g A_486_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0504 PD=0.75 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1026 A_660_47# N_SCE_M1026_g N_A_559_369#_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0483 AS=0.0693 PD=0.65 PS=0.75 NRD=17.136 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_SCD_M1020_g A_660_47# VNB NSHORT L=0.15 W=0.42 AD=0.1302
+ AS=0.0483 PD=1.46 PS=0.65 NRD=7.14 NRS=17.136 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1028 N_A_939_413#_M1028_d N_A_27_47#_M1028_g N_A_559_369#_M1028_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.0594 AS=0.1008 PD=0.69 PS=1.28 NRD=18.324 NRS=4.992 M=1
+ R=2.4 SA=75000.2 SB=75003.4 A=0.054 P=1.02 MULT=1
MM1001 A_1036_47# N_A_193_47#_M1001_g N_A_939_413#_M1028_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0634154 AS=0.0594 PD=0.701538 PS=0.69 NRD=40.38 NRS=0 M=1 R=2.4
+ SA=75000.7 SB=75002.9 A=0.054 P=1.02 MULT=1
MM1023 N_VGND_M1023_d N_A_1098_183#_M1023_g A_1036_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.118313 AS=0.0739846 PD=0.966792 PS=0.818462 NRD=47.136 NRS=34.608 M=1
+ R=2.8 SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_1098_183#_M1017_d N_A_939_413#_M1017_g N_VGND_M1023_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.126592 AS=0.180287 PD=1.2736 PS=1.47321 NRD=4.68 NRS=25.308
+ M=1 R=4.26667 SA=75001.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1003 N_A_1355_413#_M1003_d N_A_193_47#_M1003_g N_A_1098_183#_M1017_d VNB
+ NSHORT L=0.15 W=0.36 AD=0.0657 AS=0.071208 PD=0.725 PS=0.7164 NRD=26.664
+ NRS=16.656 M=1 R=2.4 SA=75002.4 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1004 A_1484_47# N_A_27_47#_M1004_g N_A_1355_413#_M1003_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0657 PD=0.687692 PS=0.725 NRD=38.076 NRS=1.656 M=1
+ R=2.4 SA=75002.9 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1027 N_VGND_M1027_d N_A_1526_315#_M1027_g A_1484_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_1355_413#_M1015_g N_A_1526_315#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.099125 AS=0.169 PD=0.955 PS=1.82 NRD=2.76 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1015_d N_A_1526_315#_M1011_g N_Q_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.099125 AS=0.08775 PD=0.955 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_1526_315#_M1013_g N_Q_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.08775 PD=1.85 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_27_47#_M1012_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1029 N_A_193_47#_M1029_d N_A_27_47#_M1029_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VPWR_M1024_d N_SCE_M1024_g N_A_299_47#_M1024_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.088 AS=0.1664 PD=0.915 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1014 A_467_369# N_SCE_M1014_g N_VPWR_M1024_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0992 AS=0.088 PD=0.95 PS=0.915 NRD=30.7714 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1016 N_A_559_369#_M1016_d N_D_M1016_g A_467_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.0992 PD=0.91 PS=0.95 NRD=0 NRS=30.7714 M=1 R=4.26667 SA=75001.1
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 A_643_369# N_A_299_47#_M1007_g N_A_559_369#_M1016_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1008 AS=0.0864 PD=0.955 PS=0.91 NRD=31.5397 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_SCD_M1005_g A_643_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1008 PD=1.85 PS=0.955 NRD=6.1464 NRS=31.5397 M=1 R=4.26667
+ SA=75002 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_939_413#_M1008_d N_A_193_47#_M1008_g N_A_559_369#_M1008_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06615 AS=0.1302 PD=0.735 PS=1.46 NRD=9.3772 NRS=21.0987 M=1
+ R=2.8 SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1030 A_1032_413# N_A_27_47#_M1030_g N_A_939_413#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0693 AS=0.06615 PD=0.75 PS=0.735 NRD=51.5943 NRS=7.0329 M=1 R=2.8
+ SA=75000.7 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_1098_183#_M1006_g A_1032_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.128423 AS=0.0693 PD=0.904615 PS=0.75 NRD=111.384 NRS=51.5943 M=1
+ R=2.8 SA=75001.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_1098_183#_M1025_d N_A_939_413#_M1025_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=0.75 AD=0.140385 AS=0.229327 PD=1.37821 PS=1.61538 NRD=0 NRS=0 M=1
+ R=5 SA=75001.2 SB=75001.1 A=0.1125 P=1.8 MULT=1
MM1009 N_A_1355_413#_M1009_d N_A_27_47#_M1009_g N_A_1098_183#_M1025_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0567 AS=0.0786154 PD=0.69 PS=0.771795 NRD=0
+ NRS=23.443 M=1 R=2.8 SA=75002.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 A_1439_413# N_A_193_47#_M1000_g N_A_1355_413#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09135 AS=0.0567 PD=0.855 PS=0.69 NRD=76.2193 NRS=0 M=1 R=2.8
+ SA=75002.7 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A_1526_315#_M1019_g A_1439_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1575 AS=0.09135 PD=1.59 PS=0.855 NRD=49.25 NRS=76.2193 M=1 R=2.8
+ SA=75003.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_1355_413#_M1002_g N_A_1526_315#_M1002_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.1525 AS=0.26 PD=1.305 PS=2.52 NRD=2.9353 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1010 N_Q_M1010_d N_A_1526_315#_M1010_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1525 PD=1.27 PS=1.305 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1033 N_Q_M1010_d N_A_1526_315#_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX34_noxref VNB VPB NWDIODE A=16.8525 P=24.21
c_109 VNB 0 8.70797e-20 $X=0.145 $Y=-0.085
c_213 VPB 0 1.42307e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__sdfxtp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o221a_4.spice.pex
* Created: Thu Aug 27 14:37:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O221A_4%C1 1 3 6 8 10 13 15 22 25
c43 8 0 1.3572e-19 $X=0.89 $Y=0.995
r44 21 22 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r45 18 21 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r46 15 25 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.23 $Y2=1.175
r47 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r52 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r54 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%B1 1 3 6 10 13 15 19 20 22 23 27 28 30
c84 28 0 1.90745e-19 $X=1.31 $Y=1.16
c85 20 0 1.87864e-19 $X=2.58 $Y=1.16
c86 1 0 1.52405e-19 $X=1.31 $Y=0.995
r87 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.16 $X2=1.31 $Y2=1.16
r88 22 23 8.21549 $w=4.93e-07 $l=3.4e-07 $layer=LI1_cond $X=1.272 $Y=1.19
+ $X2=1.272 $Y2=1.53
r89 22 28 0.724896 $w=4.93e-07 $l=3e-08 $layer=LI1_cond $X=1.272 $Y=1.19
+ $X2=1.272 $Y2=1.16
r90 20 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.16
+ $X2=2.58 $Y2=1.325
r91 20 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.16
+ $X2=2.58 $Y2=0.995
r92 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.16 $X2=2.58 $Y2=1.16
r93 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.58 $Y=1.445
+ $X2=2.58 $Y2=1.16
r94 16 23 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=1.52 $Y=1.53
+ $X2=1.272 $Y2=1.53
r95 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=1.53
+ $X2=2.58 $Y2=1.445
r96 15 16 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.415 $Y=1.53
+ $X2=1.52 $Y2=1.53
r97 13 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.985
+ $X2=2.57 $Y2=1.325
r98 10 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.56
+ $X2=2.57 $Y2=0.995
r99 4 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r100 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r101 1 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%B2 1 3 6 8 10 13 15 22
c41 6 0 1.90745e-19 $X=1.73 $Y=1.985
r42 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.94 $Y=1.16
+ $X2=2.15 $Y2=1.16
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=1.16 $X2=1.94 $Y2=1.16
r44 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.94 $Y2=1.16
r45 15 21 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=1.94 $Y2=1.175
r46 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r47 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r48 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r49 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
r50 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r51 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325 $X2=1.73
+ $Y2=1.985
r52 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995 $X2=1.73
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A1 3 6 8 10 13 15 18 19 23 24 28 31
c89 31 0 5.02546e-19 $X=4.77 $Y=1.16
c90 18 0 1.18146e-19 $X=3.44 $Y=1.16
c91 15 0 1.53436e-19 $X=4.525 $Y=1.53
r92 24 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.16 $X2=4.77 $Y2=1.16
r93 23 24 7.44331 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=4.65 $Y=1.445
+ $X2=4.65 $Y2=1.275
r94 19 29 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.445 $Y=1.16
+ $X2=3.445 $Y2=1.325
r95 19 28 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.445 $Y=1.16
+ $X2=3.445 $Y2=0.995
r96 18 21 7.37582 $w=5.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.305 $Y=1.16
+ $X2=3.305 $Y2=1.53
r97 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r98 16 21 8.31678 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=3.605 $Y=1.53 $X2=3.305
+ $Y2=1.53
r99 15 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.525 $Y=1.53
+ $X2=4.65 $Y2=1.445
r100 15 16 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.525 $Y=1.53
+ $X2=3.605 $Y2=1.53
r101 11 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.16
r102 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.985
r103 8 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.16
r104 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r105 6 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.985
+ $X2=3.51 $Y2=1.325
r106 3 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.56
+ $X2=3.51 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A2 1 3 6 8 10 13 15 21 22
c47 21 0 1.77674e-19 $X=4.14 $Y=1.16
c48 8 0 2.9244e-20 $X=4.35 $Y=0.995
c49 6 0 1.18146e-19 $X=3.93 $Y=1.985
r50 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.14 $Y=1.16
+ $X2=4.35 $Y2=1.16
r51 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.16 $X2=4.14 $Y2=1.16
r52 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.14 $Y2=1.16
r53 15 21 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=3.925 $Y=1.175
+ $X2=4.14 $Y2=1.175
r54 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.16
r55 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.985
r56 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.16
r57 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
r58 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=1.325
+ $X2=3.93 $Y2=1.16
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.93 $Y=1.325 $X2=3.93
+ $Y2=1.985
r60 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.16
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995 $X2=3.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A_109_47# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 44 47 51 53 55 58 60 61 66 70 73 74 75 80 87 95
c168 61 0 1.66254e-19 $X=5.375 $Y=1.175
c169 60 0 1.58618e-19 $X=5.29 $Y=1.445
c170 53 0 1.87864e-19 $X=4.015 $Y=1.87
c171 18 0 1.53436e-19 $X=5.19 $Y=1.985
r172 92 93 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=6.03 $Y2=1.16
r173 85 87 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.06 $Y=1.53
+ $X2=5.29 $Y2=1.53
r174 80 83 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.14 $Y=1.87 $X2=4.14
+ $Y2=1.96
r175 75 78 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.95 $Y=1.87 $X2=1.95
+ $Y2=1.96
r176 72 73 28.4433 $w=2.33e-07 $l=5.8e-07 $layer=LI1_cond $X=0.727 $Y=0.865
+ $X2=0.727 $Y2=1.445
r177 70 72 5.6861 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.68 $Y=0.73
+ $X2=0.68 $Y2=0.865
r178 67 95 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=6.45 $Y2=1.16
r179 67 93 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=6.03 $Y2=1.16
r180 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.24
+ $Y=1.16 $X2=6.24 $Y2=1.16
r181 64 92 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.4 $Y=1.16
+ $X2=5.61 $Y2=1.16
r182 64 89 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.4 $Y=1.16
+ $X2=5.19 $Y2=1.16
r183 63 66 46.5818 $w=1.98e-07 $l=8.4e-07 $layer=LI1_cond $X=5.4 $Y=1.175
+ $X2=6.24 $Y2=1.175
r184 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.4
+ $Y=1.16 $X2=5.4 $Y2=1.16
r185 61 63 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.375 $Y=1.175
+ $X2=5.4 $Y2=1.175
r186 60 87 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=1.445
+ $X2=5.29 $Y2=1.53
r187 59 61 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.29 $Y=1.275
+ $X2=5.375 $Y2=1.175
r188 59 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.29 $Y=1.275
+ $X2=5.29 $Y2=1.445
r189 57 85 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=1.615
+ $X2=5.06 $Y2=1.53
r190 57 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.06 $Y=1.615
+ $X2=5.06 $Y2=1.785
r191 56 80 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.265 $Y=1.87
+ $X2=4.14 $Y2=1.87
r192 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=1.87
+ $X2=5.06 $Y2=1.785
r193 55 56 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.975 $Y=1.87
+ $X2=4.265 $Y2=1.87
r194 54 75 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=1.87
+ $X2=1.95 $Y2=1.87
r195 53 80 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.015 $Y=1.87
+ $X2=4.14 $Y2=1.87
r196 53 54 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=4.015 $Y=1.87
+ $X2=2.075 $Y2=1.87
r197 52 74 2.98021 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.845 $Y=1.87
+ $X2=0.705 $Y2=1.87
r198 51 75 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=1.87
+ $X2=1.95 $Y2=1.87
r199 51 52 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.825 $Y=1.87
+ $X2=0.845 $Y2=1.87
r200 45 74 3.52026 $w=2.65e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.69 $Y=1.955
+ $X2=0.705 $Y2=1.87
r201 45 47 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.69 $Y=1.955
+ $X2=0.69 $Y2=2.3
r202 42 74 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.785
+ $X2=0.705 $Y2=1.87
r203 42 44 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=1.785
+ $X2=0.705 $Y2=1.62
r204 41 73 6.09362 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.705 $Y=1.585
+ $X2=0.705 $Y2=1.445
r205 41 44 1.44055 $w=2.78e-07 $l=3.5e-08 $layer=LI1_cond $X=0.705 $Y=1.585
+ $X2=0.705 $Y2=1.62
r206 37 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r207 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r208 34 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r209 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r210 30 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r211 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r212 27 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r213 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
r214 23 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.16
r215 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.985
r216 20 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r217 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r218 16 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.16
r219 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.985
r220 13 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r221 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r222 4 83 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=1.96
r223 3 78 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r224 2 47 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.3
r225 2 44 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.62
r226 1 70 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%VPWR 1 2 3 4 5 6 19 21 27 31 33 37 41 43 44
+ 45 47 67 74 75 81 86 89 91 94
r108 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r109 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 88 89 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=3.3 $Y=2.465
+ $X2=3.425 $Y2=2.465
r111 84 88 5.45271 $w=6.78e-07 $l=3.1e-07 $layer=LI1_cond $X=2.99 $Y=2.465
+ $X2=3.3 $Y2=2.465
r112 84 86 13.4907 $w=6.78e-07 $l=3.25e-07 $layer=LI1_cond $X=2.99 $Y=2.465
+ $X2=2.665 $Y2=2.465
r113 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r114 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r115 75 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r116 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r117 72 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=2.72
+ $X2=6.66 $Y2=2.72
r118 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.785 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 71 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r120 71 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r121 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r122 68 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.82 $Y2=2.72
r123 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=6.21 $Y2=2.72
r124 67 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.66 $Y2=2.72
r125 67 70 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.21 $Y2=2.72
r126 66 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r127 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 63 66 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r129 63 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r130 62 65 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r131 62 89 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.425 $Y2=2.72
r132 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 59 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r134 58 86 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.665 $Y2=2.72
r135 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r137 56 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r138 55 58 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 53 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.11 $Y2=2.72
r141 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.61 $Y2=2.72
r142 51 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r144 48 78 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r145 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 47 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=1.11 $Y2=2.72
r147 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r149 45 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r150 43 65 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.83 $Y2=2.72
r151 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.98 $Y2=2.72
r152 39 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2.72
r153 39 41 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=1.96
r154 35 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r155 35 37 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.3
r156 34 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=4.98 $Y2=2.72
r157 33 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.82 $Y2=2.72
r158 33 34 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.105 $Y2=2.72
r159 29 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r160 29 31 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.3
r161 25 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=2.635
+ $X2=1.11 $Y2=2.72
r162 25 27 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.11 $Y=2.635
+ $X2=1.11 $Y2=2.3
r163 21 24 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.27 $Y=1.65
+ $X2=0.27 $Y2=2.33
r164 19 78 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.197 $Y2=2.72
r165 19 24 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=2.33
r166 6 41 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=1.96
r167 5 37 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2.3
r168 4 31 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2.3
r169 3 88 300 $w=1.7e-07 $l=1.09455e-06 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=3.3 $Y2=2.3
r170 2 27 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.3
r171 1 24 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.33
r172 1 21 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A_277_297# 1 2 7 10 15
r21 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.37 $Y=2.3 $X2=2.37
+ $Y2=2.38
r22 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.53 $Y=2.3 $X2=1.53
+ $Y2=2.38
r23 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.655 $Y=2.38
+ $X2=1.53 $Y2=2.38
r24 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=2.38
+ $X2=2.37 $Y2=2.38
r25 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.245 $Y=2.38 $X2=1.655
+ $Y2=2.38
r26 2 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.3
r27 1 10 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A_717_297# 1 2 7 10 15
r20 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.56 $Y=2.3 $X2=4.56
+ $Y2=2.38
r21 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.72 $Y=2.3 $X2=3.72
+ $Y2=2.38
r22 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=2.38
+ $X2=3.72 $Y2=2.38
r23 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=2.38
+ $X2=4.56 $Y2=2.38
r24 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.435 $Y=2.38 $X2=3.845
+ $Y2=2.38
r25 2 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.3
r26 1 10 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%X 1 2 3 4 15 19 21 22 23 24 27 28 29 31 35
+ 39 44 45
r75 43 45 13.5704 $w=5.13e-07 $l=5.4e-07 $layer=LI1_cond $X=6.747 $Y=0.905
+ $X2=6.747 $Y2=1.445
r76 40 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.365 $Y=1.53
+ $X2=6.24 $Y2=1.53
r77 39 45 5.28309 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.575 $Y=1.53
+ $X2=6.747 $Y2=1.53
r78 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.575 $Y=1.53
+ $X2=6.365 $Y2=1.53
r79 35 37 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=6.24 $Y=1.62
+ $X2=6.24 $Y2=2.3
r80 33 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=1.615
+ $X2=6.24 $Y2=1.53
r81 33 35 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.24 $Y=1.615
+ $X2=6.24 $Y2=1.62
r82 29 43 35.7538 $w=1.73e-07 $l=5.07e-07 $layer=LI1_cond $X=6.24 $Y=0.815
+ $X2=6.747 $Y2=0.815
r83 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.24 $Y2=0.39
r84 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.115 $Y=1.53
+ $X2=6.24 $Y2=1.53
r85 27 28 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.115 $Y=1.53
+ $X2=5.9 $Y2=1.53
r86 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.815 $Y=1.615
+ $X2=5.9 $Y2=1.53
r87 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.815 $Y=1.615
+ $X2=5.815 $Y2=1.785
r88 23 29 11.1833 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=6.24 $Y2=0.815
r89 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=5.565 $Y2=0.815
r90 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.73 $Y=1.87
+ $X2=5.815 $Y2=1.785
r91 21 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.73 $Y=1.87
+ $X2=5.525 $Y2=1.87
r92 17 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.42 $Y=1.955
+ $X2=5.525 $Y2=1.87
r93 17 19 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=5.42 $Y=1.955
+ $X2=5.42 $Y2=1.96
r94 13 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.4 $Y=0.725
+ $X2=5.565 $Y2=0.815
r95 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.4 $Y=0.725 $X2=5.4
+ $Y2=0.39
r96 4 37 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=2.3
r97 4 35 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.62
r98 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.96
r99 2 31 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.39
r100 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A_27_47# 1 2 3 4 13 15 17 21 27 32
c42 21 0 2.88125e-19 $X=1.1 $Y=0.73
r43 25 27 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=1.94 $Y=0.365
+ $X2=2.78 $Y2=0.365
r44 23 32 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.365
+ $X2=1.1 $Y2=0.365
r45 23 25 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=1.185 $Y=0.365
+ $X2=1.94 $Y2=0.365
r46 19 32 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.1 $Y=0.475 $X2=1.1
+ $Y2=0.365
r47 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.1 $Y=0.475
+ $X2=1.1 $Y2=0.73
r48 18 30 3.72571 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=0.365
+ $X2=0.215 $Y2=0.365
r49 17 32 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.365
+ $X2=1.1 $Y2=0.365
r50 17 18 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.365
+ $X2=0.345 $Y2=0.365
r51 13 30 3.15253 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=0.215 $Y=0.475
+ $X2=0.215 $Y2=0.365
r52 13 15 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=0.475
+ $X2=0.215 $Y2=0.73
r53 4 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.38
r54 3 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r55 2 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r56 2 21 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.73
r57 1 30 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
r58 1 15 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%A_277_47# 1 2 3 4 13 19 23 25 29 31 32
c66 32 0 2.9244e-20 $X=3.72 $Y=0.81
r67 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.725
+ $X2=4.56 $Y2=0.39
r68 26 32 8.10876 $w=1.85e-07 $l=1.67481e-07 $layer=LI1_cond $X=3.885 $Y=0.815
+ $X2=3.72 $Y2=0.81
r69 25 27 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.395 $Y=0.815
+ $X2=4.56 $Y2=0.725
r70 25 26 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.395 $Y=0.815
+ $X2=3.885 $Y2=0.815
r71 21 32 0.63164 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.72 $Y=0.715
+ $X2=3.72 $Y2=0.81
r72 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.72 $Y=0.715
+ $X2=3.72 $Y2=0.42
r73 19 32 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0.81
+ $X2=3.72 $Y2=0.81
r74 19 31 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=3.555 $Y=0.81
+ $X2=2.535 $Y2=0.81
r75 15 18 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=1.52 $Y=0.775
+ $X2=2.36 $Y2=0.775
r76 13 31 6.61899 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.405 $Y=0.775
+ $X2=2.535 $Y2=0.775
r77 13 18 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=2.405 $Y=0.775
+ $X2=2.36 $Y2=0.775
r78 4 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.39
r79 3 23 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.42
r80 2 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.73
r81 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_4%VGND 1 2 3 4 5 18 22 26 28 32 36 39 40 42 43
+ 44 45 46 61 68 69 72 75
r107 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r108 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r109 69 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=6.67
+ $Y2=0
r110 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r111 66 75 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=6.702
+ $Y2=0
r112 66 68 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=7.13
+ $Y2=0
r113 65 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r114 65 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r115 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r116 62 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0 $X2=5.82
+ $Y2=0
r117 62 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.21 $Y2=0
r118 61 75 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.702 $Y2=0
r119 61 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.21 $Y2=0
r120 60 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r121 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r122 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r123 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r124 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r125 53 54 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r126 49 53 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.99
+ $Y2=0
r127 46 54 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=2.99 $Y2=0
r128 46 49 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r129 44 59 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.83
+ $Y2=0
r130 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r131 42 56 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=0
+ $X2=3.91 $Y2=0
r132 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0 $X2=4.14
+ $Y2=0
r133 41 59 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.83 $Y2=0
r134 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.14
+ $Y2=0
r135 39 53 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.145 $Y=0
+ $X2=2.99 $Y2=0
r136 39 40 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.265
+ $Y2=0
r137 38 56 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=3.91 $Y2=0
r138 38 40 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.265
+ $Y2=0
r139 34 75 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=6.702 $Y=0.085
+ $X2=6.702 $Y2=0
r140 34 36 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=6.702 $Y=0.085
+ $X2=6.702 $Y2=0.39
r141 30 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r142 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.39
r143 29 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r144 28 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.82
+ $Y2=0
r145 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.065 $Y2=0
r146 24 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r147 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r148 20 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r149 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.39
r150 16 40 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0.085
+ $X2=3.265 $Y2=0
r151 16 18 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.265 $Y=0.085
+ $X2=3.265 $Y2=0.38
r152 5 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.39
r153 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.39
r154 3 26 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.39
r155 2 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.39
r156 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.3 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a41o_2.pxi.spice
* Created: Thu Aug 27 14:06:08 2020
* 
x_PM_SKY130_FD_SC_HD__A41O_2%A_79_21# N_A_79_21#_M1002_s N_A_79_21#_M1006_d
+ N_A_79_21#_M1012_s N_A_79_21#_c_70_n N_A_79_21#_M1007_g N_A_79_21#_M1004_g
+ N_A_79_21#_c_71_n N_A_79_21#_M1013_g N_A_79_21#_M1010_g N_A_79_21#_c_72_n
+ N_A_79_21#_c_73_n N_A_79_21#_c_74_n N_A_79_21#_c_138_p N_A_79_21#_c_80_n
+ N_A_79_21#_c_115_p N_A_79_21#_c_81_n N_A_79_21#_c_147_p N_A_79_21#_c_83_p
+ N_A_79_21#_c_155_p N_A_79_21#_c_75_n N_A_79_21#_c_91_p
+ PM_SKY130_FD_SC_HD__A41O_2%A_79_21#
x_PM_SKY130_FD_SC_HD__A41O_2%B1 N_B1_c_171_n N_B1_M1002_g N_B1_M1012_g B1
+ N_B1_c_173_n PM_SKY130_FD_SC_HD__A41O_2%B1
x_PM_SKY130_FD_SC_HD__A41O_2%A4 N_A4_c_203_n N_A4_M1005_g N_A4_M1011_g A4 A4
+ N_A4_c_204_n N_A4_c_205_n PM_SKY130_FD_SC_HD__A41O_2%A4
x_PM_SKY130_FD_SC_HD__A41O_2%A3 N_A3_M1008_g N_A3_M1009_g N_A3_c_240_n
+ N_A3_c_241_n A3 N_A3_c_242_n PM_SKY130_FD_SC_HD__A41O_2%A3
x_PM_SKY130_FD_SC_HD__A41O_2%A2 N_A2_c_281_n N_A2_M1003_g N_A2_M1001_g A2 A2 A2
+ N_A2_c_284_n PM_SKY130_FD_SC_HD__A41O_2%A2
x_PM_SKY130_FD_SC_HD__A41O_2%A1 N_A1_c_322_n N_A1_M1006_g N_A1_M1000_g A1 A1 A1
+ N_A1_c_324_n PM_SKY130_FD_SC_HD__A41O_2%A1
x_PM_SKY130_FD_SC_HD__A41O_2%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1011_d
+ N_VPWR_M1001_d N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n
+ N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n VPWR N_VPWR_c_357_n
+ N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_349_n N_VPWR_c_361_n N_VPWR_c_362_n
+ PM_SKY130_FD_SC_HD__A41O_2%VPWR
x_PM_SKY130_FD_SC_HD__A41O_2%X N_X_M1007_s N_X_M1004_s N_X_c_428_p X X X X X X
+ PM_SKY130_FD_SC_HD__A41O_2%X
x_PM_SKY130_FD_SC_HD__A41O_2%A_381_297# N_A_381_297#_M1012_d
+ N_A_381_297#_M1009_d N_A_381_297#_M1000_d N_A_381_297#_c_433_n
+ N_A_381_297#_c_440_n N_A_381_297#_c_436_n N_A_381_297#_c_441_n
+ N_A_381_297#_c_448_n PM_SKY130_FD_SC_HD__A41O_2%A_381_297#
x_PM_SKY130_FD_SC_HD__A41O_2%VGND N_VGND_M1007_d N_VGND_M1013_d N_VGND_M1002_d
+ N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n VGND
+ N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n
+ N_VGND_c_478_n PM_SKY130_FD_SC_HD__A41O_2%VGND
cc_1 VNB N_A_79_21#_c_70_n 0.0210549f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_71_n 0.0182277f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_72_n 0.00220089f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.16
cc_4 VNB N_A_79_21#_c_73_n 0.0582519f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.16
cc_5 VNB N_A_79_21#_c_74_n 0.0117345f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.72
cc_6 VNB N_A_79_21#_c_75_n 0.00877038f $X=-0.19 $Y=-0.24 $X2=3.88 $Y2=0.38
cc_7 VNB N_B1_c_171_n 0.0201215f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_8 VNB B1 0.00214266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_173_n 0.0328006f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_10 VNB N_A4_c_203_n 0.0162214f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_11 VNB N_A4_c_204_n 0.0203911f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_12 VNB N_A4_c_205_n 0.00420204f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_13 VNB N_A3_c_240_n 0.00165924f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A3_c_241_n 0.0251692f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB N_A3_c_242_n 0.017822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_281_n 0.0177942f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_17 VNB A2 0.00269554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB A2 0.00492685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_284_n 0.0196965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A1_c_322_n 0.0193697f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_21 VNB A1 0.0046014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_324_n 0.0422983f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_23 VNB N_VPWR_c_349_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_24 VNB X 0.00165916f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_25 VNB N_VGND_c_469_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_26 VNB N_VGND_c_470_n 0.0262563f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_27 VNB N_VGND_c_471_n 0.00469218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_472_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_29 VNB N_VGND_c_473_n 0.012531f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=0.805
cc_30 VNB N_VGND_c_474_n 0.0145503f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.72
cc_31 VNB N_VGND_c_475_n 0.0474174f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=0.42
cc_32 VNB N_VGND_c_476_n 0.221296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_477_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=3.88 $Y2=0.38
cc_34 VNB N_VGND_c_478_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=0.72
cc_35 VPB N_A_79_21#_M1004_g 0.025043f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB N_A_79_21#_M1010_g 0.0218133f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_37 VPB N_A_79_21#_c_72_n 0.00320403f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.16
cc_38 VPB N_A_79_21#_c_73_n 0.0125744f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.16
cc_39 VPB N_A_79_21#_c_80_n 0.015238f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.58
cc_40 VPB N_A_79_21#_c_81_n 0.00786871f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=2
cc_41 VPB N_B1_M1012_g 0.0235946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B1_c_173_n 0.00954548f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_43 VPB N_A4_M1011_g 0.0172558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A4_c_204_n 0.00460828f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_45 VPB N_A4_c_205_n 0.00309295f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_46 VPB N_A3_M1009_g 0.0197723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A3_c_240_n 0.00135347f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_48 VPB N_A3_c_241_n 0.00563612f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_49 VPB A3 0.00742947f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_50 VPB N_A2_M1001_g 0.0206293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB A2 0.00238272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A2_c_284_n 0.00463524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A1_M1000_g 0.0221492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB A1 0.00669587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A1_c_324_n 0.00970694f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_56 VPB N_VPWR_c_350_n 0.0103102f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_57 VPB N_VPWR_c_351_n 0.0425289f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_58 VPB N_VPWR_c_352_n 0.0110503f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_59 VPB N_VPWR_c_353_n 0.00516508f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.495
cc_60 VPB N_VPWR_c_354_n 0.00516508f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.72
cc_61 VPB N_VPWR_c_355_n 0.0288082f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.58
cc_62 VPB N_VPWR_c_356_n 0.00478085f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.665
cc_63 VPB N_VPWR_c_357_n 0.0158959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_358_n 0.0201757f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=0.38
cc_65 VPB N_VPWR_c_359_n 0.0174804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_349_n 0.0533468f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_67 VPB N_VPWR_c_361_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_362_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB X 0.00242024f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_70 N_A_79_21#_c_72_n N_B1_c_171_n 0.00412051f $X=1.065 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_71 N_A_79_21#_c_83_p N_B1_c_171_n 0.0180917f $X=2.375 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_79_21#_c_72_n N_B1_M1012_g 0.00368448f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_80_n N_B1_M1012_g 0.0079637f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_81_n N_B1_M1012_g 0.0120362f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_72_n B1 0.0124033f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_73_n B1 0.00157011f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_74_n B1 0.00499907f $X=1.495 $Y=0.72 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_80_n B1 0.0219172f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_91_p B1 0.0114015f $X=1.6 $Y=0.72 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_72_n N_B1_c_173_n 9.79693e-19 $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_73_n N_B1_c_173_n 0.0205554f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_74_n N_B1_c_173_n 0.00149223f $X=1.495 $Y=0.72 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_80_n N_B1_c_173_n 0.00750174f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_91_p N_B1_c_173_n 0.00501508f $X=1.6 $Y=0.72 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_83_p N_A4_c_203_n 0.0110469f $X=2.375 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_79_21#_c_80_n N_A4_M1011_g 3.02206e-19 $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_81_n N_A4_M1011_g 5.75749e-19 $X=1.62 $Y=2 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_83_p N_A4_c_204_n 5.4424e-19 $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_80_n N_A4_c_205_n 0.00894055f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_83_p N_A4_c_205_n 0.0217942f $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_75_n N_A3_c_240_n 0.00420507f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_75_n N_A3_c_241_n 0.00171533f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_75_n N_A3_c_242_n 0.0136285f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_75_n N_A2_c_281_n 0.0126588f $X=3.88 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_79_21#_c_75_n A2 0.00743184f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_75_n A2 0.00530414f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_75_n N_A2_c_284_n 9.55082e-19 $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_75_n N_A1_c_322_n 0.012398f $X=3.88 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_79_21#_M1006_d A1 0.00970914f $X=3.745 $Y=0.235 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_75_n A1 0.0106245f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_75_n N_A1_c_324_n 8.1644e-19 $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_80_n N_VPWR_M1010_d 0.00296009f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_115_p N_VPWR_M1010_d 0.00253899f $X=1.15 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A_79_21#_M1004_g N_VPWR_c_351_n 0.0169088f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_79_21#_M1010_g N_VPWR_c_351_n 7.65745e-19 $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_M1010_g N_VPWR_c_352_n 0.00311793f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_107 N_A_79_21#_c_73_n N_VPWR_c_352_n 6.01176e-19 $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_80_n N_VPWR_c_352_n 0.00935937f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_115_p N_VPWR_c_352_n 0.0114956f $X=1.15 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_81_n N_VPWR_c_352_n 0.0444962f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_81_n N_VPWR_c_355_n 0.016757f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_112 N_A_79_21#_M1004_g N_VPWR_c_357_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_79_21#_M1010_g N_VPWR_c_357_n 0.00585385f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_79_21#_M1012_s N_VPWR_c_349_n 0.00211564f $X=1.495 $Y=1.485 $X2=0
+ $Y2=0
cc_115 N_A_79_21#_M1004_g N_VPWR_c_349_n 0.00789179f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_79_21#_M1010_g N_VPWR_c_349_n 0.0118632f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_81_n N_VPWR_c_349_n 0.0121755f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_70_n X 0.00360646f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_79_21#_M1004_g X 0.00503223f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_71_n X 0.00139758f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_79_21#_M1010_g X 0.00242672f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_72_n X 0.0386771f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_73_n X 0.0279635f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_72_n N_VGND_M1013_d 0.00139313f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_74_n N_VGND_M1013_d 0.00297499f $X=1.495 $Y=0.72 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_138_p N_VGND_M1013_d 0.00249951f $X=1.15 $Y=0.72 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_83_p N_VGND_M1002_d 0.00435389f $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_70_n N_VGND_c_470_n 0.012622f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_71_n N_VGND_c_470_n 6.89759e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_70_n N_VGND_c_471_n 5.8955e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_71_n N_VGND_c_471_n 0.00904117f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_73_n N_VGND_c_471_n 6.40396e-19 $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_74_n N_VGND_c_471_n 0.00877789f $X=1.495 $Y=0.72 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_138_p N_VGND_c_471_n 0.010787f $X=1.15 $Y=0.72 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_147_p N_VGND_c_471_n 0.0133761f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_83_p N_VGND_c_472_n 0.0159625f $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_70_n N_VGND_c_473_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_71_n N_VGND_c_473_n 0.0046653f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_74_n N_VGND_c_474_n 0.00418519f $X=1.495 $Y=0.72 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_147_p N_VGND_c_474_n 0.0141996f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_83_p N_VGND_c_474_n 0.00244309f $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_83_p N_VGND_c_475_n 0.00244309f $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_155_p N_VGND_c_475_n 0.00894629f $X=2.545 $Y=0.38 $X2=0
+ $Y2=0
cc_144 N_A_79_21#_c_75_n N_VGND_c_475_n 0.0677453f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_145 N_A_79_21#_M1002_s N_VGND_c_476_n 0.00225589f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_146 N_A_79_21#_M1006_d N_VGND_c_476_n 0.0021084f $X=3.745 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_79_21#_c_70_n N_VGND_c_476_n 0.00796766f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_71_n N_VGND_c_476_n 0.00796766f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_74_n N_VGND_c_476_n 0.00705575f $X=1.495 $Y=0.72 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_138_p N_VGND_c_476_n 8.57032e-19 $X=1.15 $Y=0.72 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_147_p N_VGND_c_476_n 0.0079665f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_83_p N_VGND_c_476_n 0.00988417f $X=2.375 $Y=0.72 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_155_p N_VGND_c_476_n 0.00636368f $X=2.545 $Y=0.38 $X2=0
+ $Y2=0
cc_154 N_A_79_21#_c_75_n N_VGND_c_476_n 0.0523446f $X=3.88 $Y=0.38 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_83_p A_465_47# 0.00696224f $X=2.375 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_79_21#_c_155_p A_465_47# 0.00192457f $X=2.545 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A_79_21#_c_75_n A_549_47# 0.0129829f $X=3.88 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_79_21#_c_75_n A_665_47# 0.00363803f $X=3.88 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_159 N_B1_c_171_n N_A4_c_203_n 0.0266891f $X=1.83 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_160 N_B1_M1012_g N_A4_M1011_g 0.0260247f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B1_c_173_n N_A4_c_204_n 0.0209651f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_162 B1 N_A4_c_205_n 0.012274f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_163 N_B1_c_173_n N_A4_c_205_n 0.0100722f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B1_M1012_g N_VPWR_c_352_n 0.00283988f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B1_M1012_g N_VPWR_c_355_n 0.00542953f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_166 N_B1_M1012_g N_VPWR_c_349_n 0.0109803f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_167 N_B1_c_171_n N_VGND_c_471_n 0.00180458f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B1_c_171_n N_VGND_c_472_n 0.00699641f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B1_c_171_n N_VGND_c_474_n 0.00339367f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B1_c_171_n N_VGND_c_476_n 0.00527013f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A4_M1011_g N_A3_M1009_g 0.0445693f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A4_c_205_n N_A3_M1009_g 0.00148463f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A4_c_204_n N_A3_c_240_n 0.00100444f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A4_c_205_n N_A3_c_240_n 0.0180705f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A4_c_204_n N_A3_c_241_n 0.0202199f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A4_c_205_n N_A3_c_241_n 0.00111877f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A4_M1011_g A3 2.0959e-19 $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A4_c_205_n A3 0.00530702f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A4_c_203_n N_A3_c_242_n 0.0401184f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A4_M1011_g N_VPWR_c_353_n 0.00302074f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A4_M1011_g N_VPWR_c_355_n 0.00441875f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A4_M1011_g N_VPWR_c_349_n 0.00591459f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A4_c_205_n N_A_381_297#_M1012_d 0.00260187f $X=2.25 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_184 N_A4_M1011_g N_A_381_297#_c_433_n 0.0101783f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A4_c_204_n N_A_381_297#_c_433_n 7.90399e-19 $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A4_c_205_n N_A_381_297#_c_433_n 0.0113192f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A4_c_205_n N_A_381_297#_c_436_n 0.0104779f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A4_c_203_n N_VGND_c_472_n 0.00811949f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A4_c_203_n N_VGND_c_475_n 0.00339367f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A4_c_203_n N_VGND_c_476_n 0.00401529f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A3_c_242_n N_A2_c_281_n 0.0257323f $X=2.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_192 N_A3_M1009_g N_A2_M1001_g 0.0231944f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A3_c_240_n N_A2_M1001_g 8.58478e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_194 A3 N_A2_M1001_g 0.00191002f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_195 N_A3_c_240_n A2 0.00237303f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A3_c_241_n A2 2.04198e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A3_c_240_n A2 0.0169297f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A3_c_241_n A2 0.00130496f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_199 A3 A2 0.00784382f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_200 N_A3_c_240_n N_A2_c_284_n 7.74181e-19 $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A3_c_241_n N_A2_c_284_n 0.0206301f $X=2.77 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A3_M1009_g N_VPWR_c_353_n 0.00302074f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A3_M1009_g N_VPWR_c_358_n 0.00441875f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A3_M1009_g N_VPWR_c_349_n 0.00625799f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_205 A3 N_A_381_297#_M1009_d 0.00552876f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_206 N_A3_M1009_g N_A_381_297#_c_433_n 0.0129195f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_207 A3 N_A_381_297#_c_433_n 0.00403356f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_208 A3 N_A_381_297#_c_440_n 0.00911921f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_209 A3 N_A_381_297#_c_441_n 0.0133455f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_210 N_A3_c_242_n N_VGND_c_472_n 0.00146555f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A3_c_242_n N_VGND_c_475_n 0.00366111f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A3_c_242_n N_VGND_c_476_n 0.00569218f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A2_c_281_n N_A1_c_322_n 0.0417537f $X=3.25 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_214 A2 N_A1_c_322_n 0.00212896f $X=3.36 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_215 N_A2_M1001_g N_A1_M1000_g 0.0428204f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_216 A2 A1 0.0114509f $X=3.36 $Y=0.765 $X2=0 $Y2=0
cc_217 A2 A1 0.025042f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_218 N_A2_c_284_n A1 2.42069e-19 $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_219 A2 N_A1_c_324_n 0.00404544f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_220 N_A2_c_284_n N_A1_c_324_n 0.0206846f $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_221 A2 N_VPWR_M1001_d 0.00265857f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A2_M1001_g N_VPWR_c_354_n 0.00302074f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A2_M1001_g N_VPWR_c_358_n 0.00441875f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A2_M1001_g N_VPWR_c_349_n 0.00631719f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A2_M1001_g N_A_381_297#_c_440_n 0.0147927f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_226 A2 N_A_381_297#_c_440_n 0.0177664f $X=3.36 $Y=1.105 $X2=0 $Y2=0
cc_227 N_A2_c_284_n N_A_381_297#_c_440_n 0.00101759f $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A2_M1001_g N_A_381_297#_c_441_n 0.00690125f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A2_c_281_n N_VGND_c_475_n 0.00366111f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A2_c_281_n N_VGND_c_476_n 0.00569218f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_231 A2 A_665_47# 0.00266747f $X=3.36 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_232 N_A1_M1000_g N_VPWR_c_354_n 0.00302074f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_M1000_g N_VPWR_c_359_n 0.00441875f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_M1000_g N_VPWR_c_349_n 0.00684159f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_235 A1 N_A_381_297#_M1000_d 0.0103551f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_236 N_A1_M1000_g N_A_381_297#_c_440_n 0.0147351f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_237 A1 N_A_381_297#_c_448_n 0.0146803f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A1_c_324_n N_A_381_297#_c_448_n 6.87511e-19 $X=3.87 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A1_c_322_n N_VGND_c_475_n 0.00366111f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A1_c_322_n N_VGND_c_476_n 0.00622254f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_241 N_VPWR_c_349_n N_X_M1004_s 0.00492927f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_242 N_VPWR_c_357_n X 0.0121054f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_243 N_VPWR_c_349_n X 0.00724021f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_349_n N_A_381_297#_M1012_d 0.00414531f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_245 N_VPWR_c_349_n N_A_381_297#_M1009_d 0.00484415f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_349_n N_A_381_297#_M1000_d 0.00377405f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_247 N_VPWR_M1011_d N_A_381_297#_c_433_n 0.00761236f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_353_n N_A_381_297#_c_433_n 0.0102407f $X=2.46 $Y=2.34 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_355_n N_A_381_297#_c_433_n 0.0023033f $X=2.335 $Y=2.72 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_358_n N_A_381_297#_c_433_n 0.0023033f $X=3.335 $Y=2.72 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_349_n N_A_381_297#_c_433_n 0.010153f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_252 N_VPWR_M1001_d N_A_381_297#_c_440_n 0.00340098f $X=3.325 $Y=1.485 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_354_n N_A_381_297#_c_440_n 0.0102407f $X=3.46 $Y=2.34 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_358_n N_A_381_297#_c_440_n 0.00443964f $X=3.335 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_359_n N_A_381_297#_c_440_n 0.0023033f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_349_n N_A_381_297#_c_440_n 0.0143308f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_355_n N_A_381_297#_c_436_n 0.0113839f $X=2.335 $Y=2.72 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_349_n N_A_381_297#_c_436_n 0.00646745f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_358_n N_A_381_297#_c_441_n 0.0115924f $X=3.335 $Y=2.72 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_349_n N_A_381_297#_c_441_n 0.00646745f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_359_n N_A_381_297#_c_448_n 0.0115924f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_349_n N_A_381_297#_c_448_n 0.00646745f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_263 N_X_c_428_p N_VGND_c_473_n 0.00906544f $X=0.68 $Y=0.46 $X2=0 $Y2=0
cc_264 N_X_M1007_s N_VGND_c_476_n 0.00512397f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_265 N_X_c_428_p N_VGND_c_476_n 0.00634211f $X=0.68 $Y=0.46 $X2=0 $Y2=0
cc_266 X N_VGND_c_476_n 5.23187e-19 $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_267 N_VGND_c_476_n A_465_47# 0.00236972f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_268 N_VGND_c_476_n A_549_47# 0.00350336f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_269 N_VGND_c_476_n A_665_47# 0.00219239f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a21bo_1.spice.pex
* Created: Thu Aug 27 14:00:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BO_1%B1_N 1 2 3 5 6 8 13 15 16 17 18 24
r38 17 18 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.16
+ $X2=0.22 $Y2=1.53
r39 17 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r40 16 17 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.22 $Y=0.85
+ $X2=0.22 $Y2=1.16
r41 15 16 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=0.51
+ $X2=0.22 $Y2=0.85
r42 11 24 145.524 $w=2.7e-07 $l=6.55e-07 $layer=POLY_cond $X=0.24 $Y=1.815
+ $X2=0.24 $Y2=1.16
r43 11 13 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.89
+ $X2=0.47 $Y2=1.89
r44 9 24 56.6543 $w=2.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=0.905
+ $X2=0.24 $Y2=1.16
r45 6 8 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.815 $Y=0.755
+ $X2=0.815 $Y2=0.445
r46 3 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.965
+ $X2=0.47 $Y2=1.89
r47 3 5 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.47 $Y=1.965 $X2=0.47
+ $Y2=2.275
r48 2 9 29.8935 $w=1.5e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.375 $Y=0.83
+ $X2=0.24 $Y2=0.905
r49 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.74 $Y=0.83
+ $X2=0.815 $Y2=0.755
r50 1 2 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.74 $Y=0.83 $X2=0.375
+ $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%A_27_413# 1 2 7 11 13 15 16 19 23 25 26 28
+ 35
c65 25 0 1.83237e-19 $X=0.685 $Y=1.335
r66 29 35 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=0.72 $Y=1.44
+ $X2=0.72 $Y2=1.285
r67 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.44 $X2=0.72 $Y2=1.44
r68 26 28 13.7276 $w=3.38e-07 $l=4.05e-07 $layer=LI1_cond $X=0.685 $Y=1.845
+ $X2=0.685 $Y2=1.44
r69 25 34 6.97447 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.685 $Y=1.335
+ $X2=0.685 $Y2=1.165
r70 25 28 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=0.685 $Y=1.335
+ $X2=0.685 $Y2=1.44
r71 23 34 35.8259 $w=2.28e-07 $l=7.15e-07 $layer=LI1_cond $X=0.63 $Y=0.45
+ $X2=0.63 $Y2=1.165
r72 17 26 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.225 $Y=1.945
+ $X2=0.685 $Y2=1.945
r73 17 19 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=2.27
r74 13 16 25.7466 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.415 $Y=1.385
+ $X2=1.415 $Y2=1.285
r75 13 15 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.415 $Y=1.385 $X2=1.415
+ $Y2=1.985
r76 9 16 25.7466 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.415 $Y=1.185
+ $X2=1.415 $Y2=1.285
r77 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.415 $Y=1.185
+ $X2=1.415 $Y2=0.56
r78 8 35 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.855 $Y=1.285
+ $X2=0.72 $Y2=1.285
r79 7 16 1.30468 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.34 $Y=1.285 $X2=1.415
+ $Y2=1.285
r80 7 8 160.815 $w=2e-07 $l=4.85e-07 $layer=POLY_cond $X=1.34 $Y=1.285 $X2=0.855
+ $Y2=1.285
r81 2 19 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.27
r82 1 23 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.475
+ $Y=0.235 $X2=0.6 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%A1 3 6 8 9 13 14 15
c37 13 0 1.88495e-19 $X=1.845 $Y=1.16
c38 6 0 6.97181e-20 $X=1.835 $Y=1.985
r39 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.16
+ $X2=1.845 $Y2=1.325
r40 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.16
+ $X2=1.845 $Y2=0.995
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.16 $X2=1.845 $Y2=1.16
r42 8 9 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.962 $Y=1.19
+ $X2=1.962 $Y2=1.53
r43 8 14 0.813489 $w=4.23e-07 $l=3e-08 $layer=LI1_cond $X=1.962 $Y=1.19
+ $X2=1.962 $Y2=1.16
r44 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.835 $Y=1.985
+ $X2=1.835 $Y2=1.325
r45 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.835 $Y=0.56
+ $X2=1.835 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%A2 1 3 6 8 9 15
r35 12 15 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.265 $Y=1.16
+ $X2=2.475 $Y2=1.16
r36 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.5 $Y=1.16 $X2=2.5
+ $Y2=1.53
r37 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.475
+ $Y=1.16 $X2=2.475 $Y2=1.16
r38 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.325
+ $X2=2.265 $Y2=1.16
r39 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.265 $Y=1.325
+ $X2=2.265 $Y2=1.985
r40 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=0.995
+ $X2=2.265 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.265 $Y=0.995
+ $X2=2.265 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%A_215_297# 1 2 7 9 12 16 21 22 26 31 34 40
c76 31 0 6.97181e-20 $X=1.47 $Y=1.195
r77 36 37 5.28703 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.575 $Y=0.72
+ $X2=1.575 $Y2=0.815
r78 34 36 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.575 $Y=0.38
+ $X2=1.575 $Y2=0.72
r79 29 31 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=1.2 $Y=1.195 $X2=1.47
+ $Y2=1.195
r80 27 40 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.005 $Y=1.16
+ $X2=3.21 $Y2=1.16
r81 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.005
+ $Y=1.16 $X2=3.005 $Y2=1.16
r82 24 26 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=2.97 $Y=0.815
+ $X2=2.97 $Y2=1.16
r83 23 36 5.54258 $w=1.9e-07 $l=2.15e-07 $layer=LI1_cond $X=1.79 $Y=0.72
+ $X2=1.575 $Y2=0.72
r84 22 24 7.03324 $w=1.9e-07 $l=1.71026e-07 $layer=LI1_cond $X=2.84 $Y=0.72
+ $X2=2.97 $Y2=0.815
r85 22 23 61.2919 $w=1.88e-07 $l=1.05e-06 $layer=LI1_cond $X=2.84 $Y=0.72
+ $X2=1.79 $Y2=0.72
r86 21 31 2.55512 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=1.47 $Y=1.045
+ $X2=1.47 $Y2=1.195
r87 21 37 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=1.47 $Y=1.045
+ $X2=1.47 $Y2=0.815
r88 16 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.63 $X2=1.2
+ $Y2=2.31
r89 14 29 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.2 $Y=1.345 $X2=1.2
+ $Y2=1.195
r90 14 16 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.2 $Y=1.345
+ $X2=1.2 $Y2=1.63
r91 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r92 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.985
r93 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r94 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995 $X2=3.21
+ $Y2=0.56
r95 2 18 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.31
r96 2 16 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.63
r97 1 34 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.49
+ $Y=0.235 $X2=1.625 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%VPWR 1 2 3 12 16 20 24 26 31 36 43 44 47 50
+ 53
r59 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 44 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r63 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 41 53 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.11 $Y=2.72
+ $X2=2.967 $Y2=2.72
r65 41 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.11 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 40 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 40 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.05 $Y2=2.72
r70 37 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 36 53 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.967 $Y2=2.72
r72 36 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.53 $Y2=2.72
r73 35 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 35 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 32 47 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 32 34 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=1.61 $Y2=2.72
r78 31 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=2.05 $Y2=2.72
r79 31 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=1.61 $Y2=2.72
r80 26 47 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r82 24 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r84 20 23 27.4969 $w=2.83e-07 $l=6.8e-07 $layer=LI1_cond $X=2.967 $Y=1.66
+ $X2=2.967 $Y2=2.34
r85 18 53 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.967 $Y=2.635
+ $X2=2.967 $Y2=2.72
r86 18 23 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=2.967 $Y=2.635
+ $X2=2.967 $Y2=2.34
r87 14 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.635
+ $X2=2.05 $Y2=2.72
r88 14 16 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.05 $Y=2.635
+ $X2=2.05 $Y2=2.24
r89 10 47 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=2.72
r90 10 12 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=2.34
r91 3 23 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.485 $X2=3 $Y2=2.34
r92 3 20 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.485 $X2=3 $Y2=1.66
r93 2 16 600 $w=1.7e-07 $l=8.22025e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.485 $X2=2.05 $Y2=2.24
r94 1 12 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%A_298_297# 1 2 9 14 16
c19 9 0 1.88495e-19 $X=2.39 $Y=1.885
r20 10 14 3.24051 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=1.715 $Y=1.885 $X2=1.625
+ $Y2=1.885
r21 9 16 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=1.885 $X2=2.475
+ $Y2=1.885
r22 9 10 37.4318 $w=1.98e-07 $l=6.75e-07 $layer=LI1_cond $X=2.39 $Y=1.885
+ $X2=1.715 $Y2=1.885
r23 2 16 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=2.34
+ $Y=1.485 $X2=2.475 $Y2=1.95
r24 1 14 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=1.485 $X2=1.625 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%X 1 2 7 8 9 10 11 12
r11 11 12 16.8751 $w=2.78e-07 $l=4.1e-07 $layer=LI1_cond $X=3.44 $Y=1.8 $X2=3.44
+ $Y2=2.21
r12 10 11 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.44 $Y=1.53
+ $X2=3.44 $Y2=1.8
r13 9 10 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.44 $Y=1.19 $X2=3.44
+ $Y2=1.53
r14 8 9 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.44 $Y=0.85 $X2=3.44
+ $Y2=1.19
r15 7 8 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.44 $Y=0.51 $X2=3.44
+ $Y2=0.85
r16 2 11 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.8
r17 1 7 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_1%VGND 1 2 9 13 15 27 28 31 36 42
r46 40 42 8.54973 $w=5.38e-07 $l=1.1e-07 $layer=LI1_cond $X=2.99 $Y=0.185
+ $X2=3.1 $Y2=0.185
r47 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r48 38 40 1.77197 $w=5.38e-07 $l=8e-08 $layer=LI1_cond $X=2.91 $Y=0.185 $X2=2.99
+ $Y2=0.185
r49 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r50 34 38 8.41685 $w=5.38e-07 $l=3.8e-07 $layer=LI1_cond $X=2.53 $Y=0.185
+ $X2=2.91 $Y2=0.185
r51 34 36 9.65721 $w=5.38e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=0.185
+ $X2=2.37 $Y2=0.185
r52 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r53 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 28 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r55 27 42 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.1
+ $Y2=0
r56 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r58 24 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r59 23 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.37
+ $Y2=0
r60 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r61 21 31 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=1.067
+ $Y2=0
r62 21 23 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=2.07
+ $Y2=0
r63 18 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r64 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r65 15 31 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.067
+ $Y2=0
r66 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.69
+ $Y2=0
r67 13 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r68 9 11 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.067 $Y=0.36
+ $X2=1.067 $Y2=0.7
r69 7 31 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.067 $Y=0.085
+ $X2=1.067 $Y2=0
r70 7 9 12.9356 $w=2.43e-07 $l=2.75e-07 $layer=LI1_cond $X=1.067 $Y=0.085
+ $X2=1.067 $Y2=0.36
r71 2 38 91 $w=1.7e-07 $l=6.29404e-07 $layer=licon1_NDIFF $count=2 $X=2.34
+ $Y=0.235 $X2=2.91 $Y2=0.36
r72 1 11 182 $w=1.7e-07 $l=5.62317e-07 $layer=licon1_NDIFF $count=1 $X=0.89
+ $Y=0.235 $X2=1.105 $Y2=0.7
r73 1 9 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.89
+ $Y=0.235 $X2=1.105 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__clkdlybuf4s50_2.pxi.spice
* Created: Thu Aug 27 14:12:09 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A N_A_M1003_g N_A_M1006_g A N_A_c_69_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_27_47# N_A_27_47#_M1003_s
+ N_A_27_47#_M1006_s N_A_27_47#_M1002_g N_A_27_47#_M1008_g N_A_27_47#_c_99_n
+ N_A_27_47#_c_105_n N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_106_n
+ N_A_27_47#_c_107_n N_A_27_47#_c_102_n N_A_27_47#_c_103_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_283_47# N_A_283_47#_M1002_d
+ N_A_283_47#_M1008_d N_A_283_47#_M1000_g N_A_283_47#_M1007_g
+ N_A_283_47#_c_164_n N_A_283_47#_c_165_n N_A_283_47#_c_166_n
+ N_A_283_47#_c_167_n N_A_283_47#_c_173_n N_A_283_47#_c_168_n
+ N_A_283_47#_c_169_n N_A_283_47#_c_170_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_283_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_390_47# N_A_390_47#_M1000_s
+ N_A_390_47#_M1007_s N_A_390_47#_M1001_g N_A_390_47#_M1004_g
+ N_A_390_47#_c_230_n N_A_390_47#_c_231_n N_A_390_47#_M1005_g
+ N_A_390_47#_M1009_g N_A_390_47#_c_234_n N_A_390_47#_c_246_n
+ N_A_390_47#_c_240_n N_A_390_47#_c_250_n N_A_390_47#_c_235_n
+ N_A_390_47#_c_256_n N_A_390_47#_c_241_n N_A_390_47#_c_236_n
+ N_A_390_47#_c_265_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_390_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%VPWR N_VPWR_M1006_d N_VPWR_M1007_d
+ N_VPWR_M1009_d N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_319_n VPWR N_VPWR_c_320_n N_VPWR_c_321_n
+ N_VPWR_c_322_n N_VPWR_c_313_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%X N_X_M1001_d N_X_M1004_s X X X X X X X
+ N_X_c_361_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%VGND N_VGND_M1003_d N_VGND_M1000_d
+ N_VGND_M1005_s N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n
+ N_VGND_c_388_n N_VGND_c_389_n VGND N_VGND_c_390_n N_VGND_c_391_n
+ N_VGND_c_392_n N_VGND_c_393_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%VGND
cc_1 VNB N_A_M1003_g 0.0386035f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.445
cc_2 VNB A 0.00912554f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_69_n 0.0335458f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_4 VNB N_A_27_47#_M1002_g 0.0436537f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_M1008_g 8.77414e-19 $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_6 VNB N_A_27_47#_c_99_n 0.0187625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_100_n 0.00427248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_101_n 0.00988546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_102_n 0.00409488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_103_n 0.0382272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_283_47#_M1000_g 0.043309f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_A_283_47#_c_164_n 0.00600833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_283_47#_c_165_n 0.00431044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_283_47#_c_166_n 0.0122986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_283_47#_c_167_n 0.0381658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_283_47#_c_168_n 0.00139809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_283_47#_c_169_n 0.00961938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_283_47#_c_170_n 0.0021445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_390_47#_M1001_g 0.0291724f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A_390_47#_c_230_n 0.0129031f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_21 VNB N_A_390_47#_c_231_n 0.0167616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_390_47#_M1005_g 0.0344922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_390_47#_M1009_g 5.18715e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_390_47#_c_234_n 0.0120043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_390_47#_c_235_n 0.0015085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_390_47#_c_236_n 0.00286356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_313_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB X 0.0273854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_384_n 0.00557217f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_30 VNB N_VGND_c_385_n 0.00278429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_386_n 0.00988902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_387_n 0.0223464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_388_n 0.0469211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_389_n 0.0051069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_390_n 0.0171347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_391_n 0.0207419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_392_n 0.00632006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_393_n 0.22551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_A_M1006_g 0.0281332f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_40 VPB N_A_c_69_n 0.0060125f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_41 VPB N_A_27_47#_M1008_g 0.064802f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_42 VPB N_A_27_47#_c_105_n 0.0331199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_106_n 0.00361619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_107_n 0.00966686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_102_n 0.00238782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_283_47#_M1007_g 0.0671574f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_47 VPB N_A_283_47#_c_167_n 0.00582278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_283_47#_c_173_n 0.00858648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_283_47#_c_168_n 0.00978399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_390_47#_M1004_g 0.0194939f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_51 VPB N_A_390_47#_c_231_n 0.00525792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_390_47#_M1009_g 0.0235992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_390_47#_c_240_n 3.17803e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_390_47#_c_241_n 0.00307087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_390_47#_c_236_n 0.00300682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_314_n 0.00284395f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_57 VPB N_VPWR_c_315_n 0.0027881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_316_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_317_n 0.0331646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_318_n 0.047311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_319_n 0.00510509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_320_n 0.0178855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_321_n 0.0203644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_322_n 0.00516427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_313_n 0.0506567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB X 0.00827921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_A_27_47#_M1002_g 0.0185276f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_69_n N_A_27_47#_M1008_g 0.0292706f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_A_27_47#_c_99_n 0.00760017f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_M1006_g N_A_27_47#_c_105_n 0.013155f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_M1003_g N_A_27_47#_c_100_n 0.0109242f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_100_n 0.0044446f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_A_27_47#_c_101_n 0.00376303f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_101_n 0.0270462f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_69_n N_A_27_47#_c_101_n 0.00620362f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_A_27_47#_c_106_n 0.0125565f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_77 A N_A_27_47#_c_106_n 0.00341853f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A_M1006_g N_A_27_47#_c_107_n 0.00434938f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_79 A N_A_27_47#_c_107_n 0.0283632f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_c_69_n N_A_27_47#_c_107_n 0.00593193f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_M1003_g N_A_27_47#_c_102_n 0.00264753f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_82 A N_A_27_47#_c_102_n 0.0106709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_c_69_n N_A_27_47#_c_102_n 0.00467276f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_84 A N_A_27_47#_c_103_n 3.33924e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A_c_69_n N_A_27_47#_c_103_n 0.018018f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_VPWR_c_314_n 0.00669214f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1006_g N_VPWR_c_320_n 0.0054895f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1006_g N_VPWR_c_313_n 0.0109548f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VGND_c_384_n 0.00312855f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_M1003_g N_VGND_c_390_n 0.00435476f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VGND_c_393_n 0.00707288f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_M1002_g N_A_283_47#_c_165_n 0.0030022f $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_c_102_n N_A_283_47#_c_165_n 0.00768466f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_103_n N_A_283_47#_c_165_n 5.95992e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_103_n N_A_283_47#_c_167_n 0.00458499f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_M1008_g N_A_283_47#_c_173_n 0.0193272f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_102_n N_A_283_47#_c_173_n 9.56133e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_M1008_g N_A_283_47#_c_168_n 0.0138427f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_102_n N_A_283_47#_c_168_n 0.0172793f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_103_n N_A_283_47#_c_168_n 5.95992e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_M1002_g N_A_283_47#_c_169_n 0.0070844f $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_102_n N_A_283_47#_c_169_n 0.00754188f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_102_n N_A_283_47#_c_170_n 0.0139147f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_103_n N_A_283_47#_c_170_n 8.02526e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_106_n N_VPWR_M1006_d 0.00205346f $X=0.85 $Y=1.542 $X2=-0.19
+ $Y2=-0.24
cc_106 N_A_27_47#_M1008_g N_VPWR_c_314_n 0.0230203f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_106_n N_VPWR_c_314_n 0.0194235f $X=0.85 $Y=1.542 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_102_n N_VPWR_c_314_n 0.00454861f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_27_47#_M1008_g N_VPWR_c_318_n 0.0185453f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_c_105_n N_VPWR_c_320_n 0.0221174f $X=0.265 $Y=1.965 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1006_s N_VPWR_c_313_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_M1008_g N_VPWR_c_313_n 0.0308452f $X=1.165 $Y=2.075 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_105_n N_VPWR_c_313_n 0.0130273f $X=0.265 $Y=1.965 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_100_n N_VGND_M1003_d 0.00191084f $X=0.85 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_27_47#_M1002_g N_VGND_c_384_n 0.00338626f $X=1.165 $Y=0.56 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_100_n N_VGND_c_384_n 0.0196209f $X=0.85 $Y=0.82 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_102_n N_VGND_c_384_n 6.93596e-19 $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_27_47#_M1002_g N_VGND_c_388_n 0.016042f $X=1.165 $Y=0.56 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_102_n N_VGND_c_388_n 0.00512243f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_99_n N_VGND_c_390_n 0.0192004f $X=0.265 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_100_n N_VGND_c_390_n 0.0022703f $X=0.85 $Y=0.82 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1003_s N_VGND_c_393_n 0.00218887f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_M1002_g N_VGND_c_393_n 0.0225454f $X=1.165 $Y=0.56 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_99_n N_VGND_c_393_n 0.0124763f $X=0.265 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_100_n N_VGND_c_393_n 0.00470124f $X=0.85 $Y=0.82 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_102_n N_VGND_c_393_n 0.00837329f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_283_47#_M1000_g N_A_390_47#_M1001_g 0.0209755f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_128 N_A_283_47#_M1007_g N_A_390_47#_M1004_g 0.022375f $X=2.46 $Y=2.075 $X2=0
+ $Y2=0
cc_129 N_A_283_47#_M1000_g N_A_390_47#_c_231_n 0.0215083f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_130 N_A_283_47#_M1000_g N_A_390_47#_c_246_n 0.0169818f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_131 N_A_283_47#_c_164_n N_A_390_47#_c_246_n 0.0345007f $X=1.555 $Y=0.435
+ $X2=0 $Y2=0
cc_132 N_A_283_47#_M1007_g N_A_390_47#_c_240_n 0.0276946f $X=2.46 $Y=2.075 $X2=0
+ $Y2=0
cc_133 N_A_283_47#_c_168_n N_A_390_47#_c_240_n 0.0619222f $X=1.592 $Y=1.785
+ $X2=0 $Y2=0
cc_134 N_A_283_47#_M1000_g N_A_390_47#_c_250_n 0.0161808f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_135 N_A_283_47#_c_166_n N_A_390_47#_c_250_n 0.00471073f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_283_47#_M1000_g N_A_390_47#_c_235_n 0.00395261f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_137 N_A_283_47#_c_166_n N_A_390_47#_c_235_n 0.0199392f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_283_47#_c_167_n N_A_390_47#_c_235_n 0.00547388f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_283_47#_c_169_n N_A_390_47#_c_235_n 0.0133135f $X=1.617 $Y=0.9 $X2=0
+ $Y2=0
cc_140 N_A_283_47#_M1007_g N_A_390_47#_c_256_n 0.0207576f $X=2.46 $Y=2.075 $X2=0
+ $Y2=0
cc_141 N_A_283_47#_c_166_n N_A_390_47#_c_256_n 0.00390417f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_283_47#_M1007_g N_A_390_47#_c_241_n 0.00401616f $X=2.46 $Y=2.075
+ $X2=0 $Y2=0
cc_143 N_A_283_47#_c_166_n N_A_390_47#_c_241_n 0.0168098f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_283_47#_c_167_n N_A_390_47#_c_241_n 0.00537291f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_283_47#_c_168_n N_A_390_47#_c_241_n 0.0129229f $X=1.592 $Y=1.785
+ $X2=0 $Y2=0
cc_146 N_A_283_47#_M1000_g N_A_390_47#_c_236_n 0.00290526f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_147 N_A_283_47#_M1007_g N_A_390_47#_c_236_n 0.00293731f $X=2.46 $Y=2.075
+ $X2=0 $Y2=0
cc_148 N_A_283_47#_c_167_n N_A_390_47#_c_236_n 0.00571204f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_283_47#_M1000_g N_A_390_47#_c_265_n 0.0173815f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_150 N_A_283_47#_M1007_g N_A_390_47#_c_265_n 0.0249116f $X=2.46 $Y=2.075 $X2=0
+ $Y2=0
cc_151 N_A_283_47#_c_166_n N_A_390_47#_c_265_n 0.0127974f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_283_47#_c_167_n N_A_390_47#_c_265_n 0.0128312f $X=2.14 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A_283_47#_c_173_n N_VPWR_c_314_n 0.0225936f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_154 N_A_283_47#_M1007_g N_VPWR_c_315_n 0.0240668f $X=2.46 $Y=2.075 $X2=0
+ $Y2=0
cc_155 N_A_283_47#_M1007_g N_VPWR_c_318_n 0.0181551f $X=2.46 $Y=2.075 $X2=0
+ $Y2=0
cc_156 N_A_283_47#_c_173_n N_VPWR_c_318_n 0.026426f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_157 N_A_283_47#_M1008_d N_VPWR_c_313_n 0.00213418f $X=1.415 $Y=1.665 $X2=0
+ $Y2=0
cc_158 N_A_283_47#_M1007_g N_VPWR_c_313_n 0.030231f $X=2.46 $Y=2.075 $X2=0 $Y2=0
cc_159 N_A_283_47#_c_173_n N_VPWR_c_313_n 0.015338f $X=1.555 $Y=1.965 $X2=0
+ $Y2=0
cc_160 N_A_283_47#_M1007_g X 0.00116786f $X=2.46 $Y=2.075 $X2=0 $Y2=0
cc_161 N_A_283_47#_M1000_g N_X_c_361_n 3.0423e-19 $X=2.46 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_283_47#_M1000_g N_VGND_c_385_n 0.0150249f $X=2.46 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A_283_47#_M1000_g N_VGND_c_388_n 0.0141825f $X=2.46 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A_283_47#_c_164_n N_VGND_c_388_n 0.0217634f $X=1.555 $Y=0.435 $X2=0
+ $Y2=0
cc_165 N_A_283_47#_M1002_d N_VGND_c_393_n 0.00300709f $X=1.415 $Y=0.235 $X2=0
+ $Y2=0
cc_166 N_A_283_47#_M1000_g N_VGND_c_393_n 0.0174764f $X=2.46 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_283_47#_c_164_n N_VGND_c_393_n 0.0134826f $X=1.555 $Y=0.435 $X2=0
+ $Y2=0
cc_168 N_A_390_47#_M1004_g N_VPWR_c_315_n 0.00311401f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_390_47#_c_231_n N_VPWR_c_315_n 0.00165851f $X=3.19 $Y=1.16 $X2=0
+ $Y2=0
cc_170 N_A_390_47#_c_240_n N_VPWR_c_315_n 0.0222064f $X=2.075 $Y=1.96 $X2=0
+ $Y2=0
cc_171 N_A_390_47#_c_236_n N_VPWR_c_315_n 0.0111699f $X=3.055 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_390_47#_M1009_g N_VPWR_c_317_n 0.00899682f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_390_47#_c_240_n N_VPWR_c_318_n 0.0153696f $X=2.075 $Y=1.96 $X2=0
+ $Y2=0
cc_174 N_A_390_47#_M1004_g N_VPWR_c_321_n 0.00579312f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_390_47#_M1009_g N_VPWR_c_321_n 0.00357668f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_390_47#_M1007_s N_VPWR_c_313_n 0.00334295f $X=1.95 $Y=1.665 $X2=0
+ $Y2=0
cc_177 N_A_390_47#_M1004_g N_VPWR_c_313_n 0.0105173f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_390_47#_M1009_g N_VPWR_c_313_n 0.00633656f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_390_47#_c_240_n N_VPWR_c_313_n 0.00936871f $X=2.075 $Y=1.96 $X2=0
+ $Y2=0
cc_180 N_A_390_47#_M1001_g X 0.00837437f $X=3.115 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A_390_47#_c_230_n X 0.0079865f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_390_47#_c_231_n X 0.00493234f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_390_47#_M1005_g X 0.0140958f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_390_47#_M1009_g X 0.00806081f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_390_47#_c_234_n X 0.00758359f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_390_47#_c_236_n X 0.025593f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_390_47#_M1004_g X 0.00637177f $X=3.115 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_390_47#_c_230_n X 0.00263886f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_390_47#_M1009_g X 0.00876628f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_390_47#_c_265_n X 0.00283299f $X=2.56 $Y=0.82 $X2=0 $Y2=0
cc_191 N_A_390_47#_M1004_g X 0.00690713f $X=3.115 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_390_47#_M1009_g X 0.0214295f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_390_47#_M1001_g N_X_c_361_n 0.00399649f $X=3.115 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_390_47#_c_230_n N_X_c_361_n 0.00218757f $X=3.465 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_390_47#_M1005_g N_X_c_361_n 0.0121195f $X=3.54 $Y=0.445 $X2=0 $Y2=0
cc_196 N_A_390_47#_M1001_g N_VGND_c_385_n 0.00311401f $X=3.115 $Y=0.445 $X2=0
+ $Y2=0
cc_197 N_A_390_47#_c_231_n N_VGND_c_385_n 0.00171461f $X=3.19 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_390_47#_c_246_n N_VGND_c_385_n 0.00985096f $X=2.075 $Y=0.47 $X2=0
+ $Y2=0
cc_199 N_A_390_47#_c_236_n N_VGND_c_385_n 0.0120075f $X=3.055 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_390_47#_M1005_g N_VGND_c_387_n 0.00740335f $X=3.54 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_390_47#_c_246_n N_VGND_c_388_n 0.0139983f $X=2.075 $Y=0.47 $X2=0
+ $Y2=0
cc_202 N_A_390_47#_c_250_n N_VGND_c_388_n 0.00313989f $X=2.475 $Y=0.82 $X2=0
+ $Y2=0
cc_203 N_A_390_47#_c_265_n N_VGND_c_388_n 0.00242772f $X=2.56 $Y=0.82 $X2=0
+ $Y2=0
cc_204 N_A_390_47#_M1001_g N_VGND_c_391_n 0.00577905f $X=3.115 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_390_47#_M1005_g N_VGND_c_391_n 0.00361001f $X=3.54 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_390_47#_M1000_s N_VGND_c_393_n 0.00335569f $X=1.95 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_A_390_47#_M1001_g N_VGND_c_393_n 0.010547f $X=3.115 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_390_47#_M1005_g N_VGND_c_393_n 0.00637982f $X=3.54 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_390_47#_c_246_n N_VGND_c_393_n 0.00935388f $X=2.075 $Y=0.47 $X2=0
+ $Y2=0
cc_210 N_A_390_47#_c_250_n N_VGND_c_393_n 0.00509412f $X=2.475 $Y=0.82 $X2=0
+ $Y2=0
cc_211 N_A_390_47#_c_265_n N_VGND_c_393_n 0.00383132f $X=2.56 $Y=0.82 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_313_n N_X_M1004_s 0.00219216f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_321_n X 0.0261201f $X=3.795 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_313_n X 0.016019f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_215 N_X_c_361_n N_VGND_c_391_n 0.0230043f $X=3.485 $Y=0.455 $X2=0 $Y2=0
cc_216 N_X_M1001_d N_VGND_c_393_n 0.00221452f $X=3.19 $Y=0.235 $X2=0 $Y2=0
cc_217 N_X_c_361_n N_VGND_c_393_n 0.0158294f $X=3.485 $Y=0.455 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nand4b_1.pxi.spice
* Created: Tue Sep  1 19:16:57 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4B_1%A_N N_A_N_M1009_g N_A_N_M1003_g A_N N_A_N_c_57_n
+ N_A_N_c_58_n PM_SKY130_FD_SC_HD__NAND4B_1%A_N
x_PM_SKY130_FD_SC_HD__NAND4B_1%D N_D_M1002_g N_D_M1008_g D N_D_c_88_n N_D_c_89_n
+ PM_SKY130_FD_SC_HD__NAND4B_1%D
x_PM_SKY130_FD_SC_HD__NAND4B_1%C N_C_M1000_g N_C_M1001_g C C N_C_c_123_n
+ N_C_c_124_n PM_SKY130_FD_SC_HD__NAND4B_1%C
x_PM_SKY130_FD_SC_HD__NAND4B_1%B N_B_M1007_g N_B_M1006_g B B N_B_c_161_n
+ N_B_c_162_n PM_SKY130_FD_SC_HD__NAND4B_1%B
x_PM_SKY130_FD_SC_HD__NAND4B_1%A_41_93# N_A_41_93#_M1009_s N_A_41_93#_M1003_s
+ N_A_41_93#_M1004_g N_A_41_93#_M1005_g N_A_41_93#_c_199_n N_A_41_93#_c_214_n
+ N_A_41_93#_c_228_n N_A_41_93#_c_200_n N_A_41_93#_c_201_n N_A_41_93#_c_207_n
+ N_A_41_93#_c_221_n N_A_41_93#_c_202_n N_A_41_93#_c_203_n N_A_41_93#_c_204_n
+ PM_SKY130_FD_SC_HD__NAND4B_1%A_41_93#
x_PM_SKY130_FD_SC_HD__NAND4B_1%VPWR N_VPWR_M1003_d N_VPWR_M1001_d N_VPWR_M1005_d
+ N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n
+ N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n VPWR
+ N_VPWR_c_293_n N_VPWR_c_283_n PM_SKY130_FD_SC_HD__NAND4B_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND4B_1%Y N_Y_M1004_d N_Y_M1008_d N_Y_M1006_d N_Y_c_329_n
+ N_Y_c_331_n N_Y_c_334_n N_Y_c_337_n N_Y_c_327_n N_Y_c_325_n N_Y_c_342_n Y
+ N_Y_c_326_n PM_SKY130_FD_SC_HD__NAND4B_1%Y
x_PM_SKY130_FD_SC_HD__NAND4B_1%VGND N_VGND_M1009_d N_VGND_c_371_n VGND
+ N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n PM_SKY130_FD_SC_HD__NAND4B_1%VGND
cc_1 VNB A_N 0.00282198f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_2 VNB N_A_N_c_57_n 0.0256803f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_A_N_c_58_n 0.0216082f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_4 VNB D 0.00238161f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_5 VNB N_D_c_88_n 0.0234624f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_6 VNB N_D_c_89_n 0.0195981f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_7 VNB C 6.78145e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_8 VNB N_C_c_123_n 0.0262217f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_9 VNB N_C_c_124_n 0.0168332f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_10 VNB B 0.00332104f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_11 VNB N_B_c_161_n 0.0212752f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_12 VNB N_B_c_162_n 0.0172109f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_13 VNB N_A_41_93#_c_199_n 0.0224415f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_14 VNB N_A_41_93#_c_200_n 0.00110967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_41_93#_c_201_n 0.0207556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_41_93#_c_202_n 0.00226835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_41_93#_c_203_n 0.0275164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_41_93#_c_204_n 0.0200719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_283_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_325_n 0.0230125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_326_n 0.0256632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_371_n 0.0107612f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_23 VNB N_VGND_c_372_n 0.0591634f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_24 VNB N_VGND_c_373_n 0.186431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_374_n 0.0260149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_N_M1003_g 0.0253918f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_27 VPB A_N 0.0020516f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_28 VPB N_A_N_c_57_n 0.00653301f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_29 VPB N_D_M1008_g 0.0221988f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_30 VPB D 3.20519e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_31 VPB N_D_c_88_n 0.00692673f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_32 VPB N_C_M1001_g 0.0203709f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_33 VPB C 0.00162853f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_34 VPB N_C_c_123_n 0.00642581f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_35 VPB N_B_M1006_g 0.0216215f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_36 VPB B 0.00113058f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_37 VPB N_B_c_161_n 0.00433855f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_38 VPB N_A_41_93#_M1005_g 0.023865f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_39 VPB N_A_41_93#_c_199_n 0.0149536f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_40 VPB N_A_41_93#_c_207_n 0.0236179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_41_93#_c_202_n 0.00150608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_41_93#_c_203_n 0.00576159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_284_n 0.022704f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_44 VPB N_VPWR_c_285_n 0.00474998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_286_n 0.00498362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_287_n 0.0247369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_288_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_289_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_290_n 0.00544936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_291_n 0.0218642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_292_n 0.00410958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_293_n 0.0116899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_283_n 0.0611597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_Y_c_327_n 0.016286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_Y_c_325_n 0.00987107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 N_A_N_M1003_g N_D_M1008_g 0.0143222f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_57 A_N D 0.0238604f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_N_c_57_n D 3.00886e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_59 A_N N_D_c_88_n 0.00219735f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_60 N_A_N_c_57_n N_D_c_88_n 0.0204854f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_N_c_58_n N_D_c_89_n 0.0163053f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A_N_M1003_g N_A_41_93#_c_199_n 0.0067114f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_63 A_N N_A_41_93#_c_199_n 0.0248817f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_N_c_57_n N_A_41_93#_c_199_n 0.00816168f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_N_c_58_n N_A_41_93#_c_199_n 0.00552893f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_66 N_A_N_c_58_n N_A_41_93#_c_214_n 0.00979936f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_67 A_N N_A_41_93#_c_201_n 0.022175f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_N_c_57_n N_A_41_93#_c_201_n 0.00394703f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_N_c_58_n N_A_41_93#_c_201_n 0.00455452f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_N_M1003_g N_A_41_93#_c_207_n 4.58643e-19 $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_71 A_N N_A_41_93#_c_207_n 0.00343051f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_72 N_A_N_c_57_n N_A_41_93#_c_207_n 0.00472985f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_N_c_58_n N_A_41_93#_c_221_n 8.58928e-19 $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A_N_M1003_g N_VPWR_c_284_n 0.0052717f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_75 A_N N_VPWR_c_284_n 0.00460569f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_N_M1003_g N_VPWR_c_287_n 0.00327927f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_77 N_A_N_M1003_g N_VPWR_c_283_n 0.00417489f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_78 N_A_N_c_58_n N_VGND_c_371_n 0.00353636f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_N_c_58_n N_VGND_c_373_n 0.00512902f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_N_c_58_n N_VGND_c_374_n 0.00392672f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_81 N_D_M1008_g N_C_M1001_g 0.0151563f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_82 D C 0.0178021f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_83 N_D_c_88_n C 3.5587e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_84 N_D_c_89_n C 9.66904e-19 $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_85 D N_C_c_123_n 0.00214521f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_86 N_D_c_88_n N_C_c_123_n 0.0207134f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_87 N_D_c_89_n N_C_c_124_n 0.0415308f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_88 D N_A_41_93#_c_214_n 0.0120433f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_89 N_D_c_88_n N_A_41_93#_c_214_n 0.00301183f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_90 N_D_c_89_n N_A_41_93#_c_214_n 0.010702f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_91 N_D_c_89_n N_A_41_93#_c_201_n 5.59292e-19 $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_92 D N_A_41_93#_c_221_n 0.00396267f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_93 N_D_c_89_n N_A_41_93#_c_221_n 0.00716949f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_94 N_D_M1008_g N_VPWR_c_284_n 0.00321269f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_95 N_D_c_88_n N_VPWR_c_284_n 0.00217348f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_96 N_D_M1008_g N_VPWR_c_289_n 0.00541359f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_97 N_D_M1008_g N_VPWR_c_283_n 0.0108548f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_98 N_D_M1008_g N_Y_c_329_n 0.00216132f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_99 D N_Y_c_329_n 0.0060702f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_100 N_D_M1008_g N_Y_c_331_n 0.00885586f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_101 N_D_c_89_n N_VGND_c_371_n 0.00478313f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_102 N_D_c_89_n N_VGND_c_372_n 0.00428075f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_103 N_D_c_89_n N_VGND_c_373_n 0.0069836f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_104 N_C_M1001_g N_B_M1006_g 0.0198628f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_105 C B 0.0384972f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_106 N_C_c_123_n B 0.0018146f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_107 N_C_c_124_n B 3.52085e-19 $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_108 C N_B_c_161_n 3.82942e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_109 N_C_c_123_n N_B_c_161_n 0.0206074f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_110 C N_B_c_162_n 7.6277e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_111 N_C_c_124_n N_B_c_162_n 0.0292182f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_112 C N_A_41_93#_c_228_n 0.0143973f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_113 N_C_c_123_n N_A_41_93#_c_228_n 6.42489e-19 $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_114 N_C_c_124_n N_A_41_93#_c_228_n 0.0125738f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_115 C N_A_41_93#_c_221_n 0.00435518f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_116 N_C_c_124_n N_A_41_93#_c_221_n 0.00451965f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C_M1001_g N_VPWR_c_285_n 0.0016963f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_118 N_C_M1001_g N_VPWR_c_289_n 0.00541359f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_119 N_C_M1001_g N_VPWR_c_283_n 0.00981263f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_120 N_C_M1001_g N_Y_c_329_n 0.00196977f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_121 N_C_M1001_g N_Y_c_331_n 0.010277f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_122 N_C_M1001_g N_Y_c_334_n 0.0126503f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_123 C N_Y_c_334_n 0.01693f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_124 N_C_c_123_n N_Y_c_334_n 0.00110224f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_125 N_C_M1001_g N_Y_c_337_n 5.96051e-19 $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C_c_124_n N_VGND_c_372_n 0.00390868f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_127 N_C_c_124_n N_VGND_c_373_n 0.00575332f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_128 C A_316_47# 0.00229559f $X=1.525 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_129 N_B_M1006_g N_A_41_93#_M1005_g 0.0220159f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_130 B N_A_41_93#_c_228_n 0.0117784f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_131 N_B_c_161_n N_A_41_93#_c_228_n 0.00170799f $X=2.1 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B_c_162_n N_A_41_93#_c_228_n 0.0118148f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_133 B N_A_41_93#_c_200_n 0.0175596f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_134 N_B_c_162_n N_A_41_93#_c_200_n 0.00405271f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_135 B N_A_41_93#_c_202_n 0.026043f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_136 N_B_c_161_n N_A_41_93#_c_202_n 0.00230841f $X=2.1 $Y=1.16 $X2=0 $Y2=0
cc_137 B N_A_41_93#_c_203_n 2.98157e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_138 N_B_c_161_n N_A_41_93#_c_203_n 0.0145996f $X=2.1 $Y=1.16 $X2=0 $Y2=0
cc_139 B N_A_41_93#_c_204_n 5.94804e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_140 N_B_c_162_n N_A_41_93#_c_204_n 0.026699f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B_M1006_g N_VPWR_c_285_n 0.00299999f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B_M1006_g N_VPWR_c_291_n 0.00541359f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B_M1006_g N_VPWR_c_283_n 0.0100793f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B_M1006_g N_Y_c_331_n 5.96051e-19 $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B_M1006_g N_Y_c_334_n 0.0112741f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_146 B N_Y_c_334_n 0.0107269f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_147 N_B_M1006_g N_Y_c_337_n 0.010277f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B_M1006_g N_Y_c_342_n 8.8334e-19 $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_149 B N_Y_c_342_n 0.00583661f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_150 N_B_c_161_n N_Y_c_342_n 0.00263989f $X=2.1 $Y=1.16 $X2=0 $Y2=0
cc_151 N_B_c_162_n N_VGND_c_372_n 0.00390868f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B_c_162_n N_VGND_c_373_n 0.00603026f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_153 B A_423_47# 0.00120781f $X=1.985 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_154 N_A_41_93#_c_214_n N_VPWR_c_284_n 0.00511975f $X=1.155 $Y=0.74 $X2=0
+ $Y2=0
cc_155 N_A_41_93#_c_207_n N_VPWR_c_284_n 0.00133957f $X=0.39 $Y=1.76 $X2=0 $Y2=0
cc_156 N_A_41_93#_M1005_g N_VPWR_c_286_n 0.00445216f $X=2.58 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_41_93#_M1005_g N_VPWR_c_291_n 0.00585385f $X=2.58 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_41_93#_M1005_g N_VPWR_c_283_n 0.0120002f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_41_93#_c_207_n N_VPWR_c_283_n 0.0161088f $X=0.39 $Y=1.76 $X2=0 $Y2=0
cc_160 N_A_41_93#_c_221_n N_Y_c_329_n 0.00303746f $X=1.245 $Y=0.51 $X2=0 $Y2=0
cc_161 N_A_41_93#_M1005_g N_Y_c_337_n 0.010959f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_41_93#_M1005_g N_Y_c_327_n 0.0173403f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_41_93#_c_202_n N_Y_c_327_n 0.020935f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_41_93#_c_203_n N_Y_c_327_n 0.00430395f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_41_93#_M1005_g N_Y_c_325_n 0.00532965f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_41_93#_c_200_n N_Y_c_325_n 0.00641422f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_41_93#_c_202_n N_Y_c_325_n 0.0255425f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_41_93#_c_203_n N_Y_c_325_n 0.00820562f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_41_93#_c_204_n N_Y_c_325_n 0.00325724f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_41_93#_c_202_n N_Y_c_342_n 0.00520145f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_41_93#_c_202_n N_Y_c_326_n 0.00410432f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_41_93#_c_203_n N_Y_c_326_n 0.00369177f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_41_93#_c_214_n N_VGND_M1009_d 0.00746632f $X=1.155 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_41_93#_c_214_n N_VGND_c_371_n 0.0211878f $X=1.155 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_41_93#_c_201_n N_VGND_c_371_n 0.00216362f $X=0.475 $Y=0.635 $X2=0
+ $Y2=0
cc_176 N_A_41_93#_c_214_n N_VGND_c_372_n 0.00248883f $X=1.155 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_41_93#_c_228_n N_VGND_c_372_n 0.032231f $X=2.355 $Y=0.51 $X2=0 $Y2=0
cc_178 N_A_41_93#_c_221_n N_VGND_c_372_n 0.00488204f $X=1.245 $Y=0.51 $X2=0
+ $Y2=0
cc_179 N_A_41_93#_c_204_n N_VGND_c_372_n 0.00559425f $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_41_93#_c_214_n N_VGND_c_373_n 0.0102792f $X=1.155 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_41_93#_c_228_n N_VGND_c_373_n 0.0382125f $X=2.355 $Y=0.51 $X2=0 $Y2=0
cc_182 N_A_41_93#_c_201_n N_VGND_c_373_n 0.0131201f $X=0.475 $Y=0.635 $X2=0
+ $Y2=0
cc_183 N_A_41_93#_c_221_n N_VGND_c_373_n 0.0060711f $X=1.245 $Y=0.51 $X2=0 $Y2=0
cc_184 N_A_41_93#_c_204_n N_VGND_c_373_n 0.0115227f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_41_93#_c_214_n N_VGND_c_374_n 0.00257535f $X=1.155 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_41_93#_c_201_n N_VGND_c_374_n 0.0120273f $X=0.475 $Y=0.635 $X2=0
+ $Y2=0
cc_187 N_A_41_93#_c_228_n A_232_47# 0.00235031f $X=2.355 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_41_93#_c_221_n A_232_47# 0.00671709f $X=1.245 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_41_93#_c_228_n A_316_47# 0.010698f $X=2.355 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_41_93#_c_228_n A_423_47# 0.00925372f $X=2.355 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_41_93#_c_200_n A_423_47# 0.00309549f $X=2.44 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_192 N_VPWR_c_283_n N_Y_M1008_d 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_283_n N_Y_M1006_d 0.00628276f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_c_289_n N_Y_c_331_n 0.0189039f $X=1.63 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_283_n N_Y_c_331_n 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_M1001_d N_Y_c_334_n 0.00995379f $X=1.58 $Y=1.485 $X2=0 $Y2=0
cc_197 N_VPWR_c_285_n N_Y_c_334_n 0.0220482f $X=1.775 $Y=2 $X2=0 $Y2=0
cc_198 N_VPWR_c_291_n N_Y_c_337_n 0.0209845f $X=2.705 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_283_n N_Y_c_337_n 0.0124268f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_M1005_d N_Y_c_327_n 0.00693734f $X=2.655 $Y=1.485 $X2=0 $Y2=0
cc_201 N_VPWR_c_286_n N_Y_c_327_n 0.0168412f $X=2.79 $Y=2 $X2=0 $Y2=0
cc_202 N_Y_c_326_n N_VGND_c_372_n 0.0302286f $X=2.86 $Y=0.38 $X2=0 $Y2=0
cc_203 N_Y_M1004_d N_VGND_c_373_n 0.00426238f $X=2.655 $Y=0.235 $X2=0 $Y2=0
cc_204 N_Y_c_326_n N_VGND_c_373_n 0.0168278f $X=2.86 $Y=0.38 $X2=0 $Y2=0
cc_205 N_VGND_c_373_n A_232_47# 0.00242407f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_206 N_VGND_c_373_n A_316_47# 0.00347185f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_207 N_VGND_c_373_n A_423_47# 0.00351546f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__dlrtn_2.pxi.spice
* Created: Tue Sep  1 19:05:19 2020
* 
x_PM_SKY130_FD_SC_HD__DLRTN_2%GATE_N N_GATE_N_c_146_n N_GATE_N_c_141_n
+ N_GATE_N_M1018_g N_GATE_N_c_147_n N_GATE_N_M1008_g N_GATE_N_c_142_n
+ N_GATE_N_c_148_n GATE_N GATE_N N_GATE_N_c_144_n N_GATE_N_c_145_n
+ PM_SKY130_FD_SC_HD__DLRTN_2%GATE_N
x_PM_SKY130_FD_SC_HD__DLRTN_2%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1008_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_M1017_g N_A_27_47#_M1020_g
+ N_A_27_47#_c_337_p N_A_27_47#_c_186_n N_A_27_47#_c_187_n N_A_27_47#_c_196_n
+ N_A_27_47#_c_197_n N_A_27_47#_c_198_n N_A_27_47#_c_199_n N_A_27_47#_c_188_n
+ N_A_27_47#_c_189_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n N_A_27_47#_c_201_n
+ N_A_27_47#_c_202_n N_A_27_47#_c_203_n N_A_27_47#_c_204_n N_A_27_47#_c_205_n
+ N_A_27_47#_c_192_n N_A_27_47#_c_193_n PM_SKY130_FD_SC_HD__DLRTN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRTN_2%D N_D_M1002_g N_D_M1016_g D N_D_c_352_n
+ N_D_c_353_n PM_SKY130_FD_SC_HD__DLRTN_2%D
x_PM_SKY130_FD_SC_HD__DLRTN_2%A_299_47# N_A_299_47#_M1002_s N_A_299_47#_M1016_s
+ N_A_299_47#_c_390_n N_A_299_47#_M1004_g N_A_299_47#_M1012_g
+ N_A_299_47#_c_398_n N_A_299_47#_c_392_n N_A_299_47#_c_399_n
+ N_A_299_47#_c_400_n N_A_299_47#_c_393_n N_A_299_47#_c_394_n
+ N_A_299_47#_c_395_n N_A_299_47#_c_396_n PM_SKY130_FD_SC_HD__DLRTN_2%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRTN_2%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1001_g N_A_193_47#_c_472_n N_A_193_47#_c_473_n
+ N_A_193_47#_M1011_g N_A_193_47#_c_479_n N_A_193_47#_c_475_n
+ N_A_193_47#_c_481_n N_A_193_47#_c_482_n N_A_193_47#_c_483_n
+ N_A_193_47#_c_484_n N_A_193_47#_c_485_n N_A_193_47#_c_486_n
+ N_A_193_47#_c_487_n PM_SKY130_FD_SC_HD__DLRTN_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRTN_2%A_711_307# N_A_711_307#_M1015_s
+ N_A_711_307#_M1013_d N_A_711_307#_M1009_g N_A_711_307#_M1021_g
+ N_A_711_307#_M1006_g N_A_711_307#_c_586_n N_A_711_307#_M1003_g
+ N_A_711_307#_c_587_n N_A_711_307#_M1005_g N_A_711_307#_M1014_g
+ N_A_711_307#_c_597_n N_A_711_307#_c_598_n N_A_711_307#_c_588_n
+ N_A_711_307#_c_611_p N_A_711_307#_c_589_n N_A_711_307#_c_657_p
+ N_A_711_307#_c_629_p N_A_711_307#_c_599_n N_A_711_307#_c_643_p
+ N_A_711_307#_c_590_n N_A_711_307#_c_591_n N_A_711_307#_c_592_n
+ PM_SKY130_FD_SC_HD__DLRTN_2%A_711_307#
x_PM_SKY130_FD_SC_HD__DLRTN_2%A_560_47# N_A_560_47#_M1017_d N_A_560_47#_M1001_d
+ N_A_560_47#_M1013_g N_A_560_47#_M1015_g N_A_560_47#_c_721_n
+ N_A_560_47#_c_722_n N_A_560_47#_c_729_n N_A_560_47#_c_733_n
+ N_A_560_47#_c_723_n N_A_560_47#_c_727_n N_A_560_47#_c_724_n
+ N_A_560_47#_c_725_n PM_SKY130_FD_SC_HD__DLRTN_2%A_560_47#
x_PM_SKY130_FD_SC_HD__DLRTN_2%RESET_B N_RESET_B_M1019_g N_RESET_B_c_806_n
+ N_RESET_B_M1007_g RESET_B N_RESET_B_c_807_n N_RESET_B_c_808_n
+ PM_SKY130_FD_SC_HD__DLRTN_2%RESET_B
x_PM_SKY130_FD_SC_HD__DLRTN_2%VPWR N_VPWR_M1008_d N_VPWR_M1016_d N_VPWR_M1009_d
+ N_VPWR_M1013_s N_VPWR_M1019_d N_VPWR_M1014_s N_VPWR_c_847_n N_VPWR_c_848_n
+ N_VPWR_c_849_n N_VPWR_c_850_n N_VPWR_c_851_n N_VPWR_c_852_n N_VPWR_c_853_n
+ VPWR N_VPWR_c_854_n N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n
+ N_VPWR_c_858_n N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n
+ N_VPWR_c_846_n PM_SKY130_FD_SC_HD__DLRTN_2%VPWR
x_PM_SKY130_FD_SC_HD__DLRTN_2%Q N_Q_M1003_d N_Q_M1006_d N_Q_c_962_n N_Q_c_965_n
+ N_Q_c_969_n N_Q_c_972_n N_Q_c_960_n Q Q Q N_Q_c_959_n Q
+ PM_SKY130_FD_SC_HD__DLRTN_2%Q
x_PM_SKY130_FD_SC_HD__DLRTN_2%VGND N_VGND_M1018_d N_VGND_M1002_d N_VGND_M1021_d
+ N_VGND_M1007_d N_VGND_M1005_s N_VGND_c_1006_n N_VGND_c_1007_n N_VGND_c_1008_n
+ N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n VGND N_VGND_c_1012_n
+ N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n
+ N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n
+ N_VGND_c_1021_n PM_SKY130_FD_SC_HD__DLRTN_2%VGND
cc_1 VNB N_GATE_N_c_141_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_142_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_144_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_145_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0397896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_M1017_g 0.0207626f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_8 VNB N_A_27_47#_c_186_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_187_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_188_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_189_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_190_n 0.0265912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_191_n 0.00779739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_192_n 0.0230671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_193_n 0.00251875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1002_g 0.0258823f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_M1016_g 0.00623887f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_352_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_353_n 0.0421319f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_20 VNB N_A_299_47#_c_390_n 0.0166762f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_21 VNB N_A_299_47#_M1012_g 0.0126741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_392_n 0.00251174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_393_n 0.00494173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_299_47#_c_394_n 0.00328354f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_25 VNB N_A_299_47#_c_395_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_26 VNB N_A_299_47#_c_396_n 0.026293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_472_n 0.0131123f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_28 VNB N_A_193_47#_c_473_n 0.0048068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_M1011_g 0.0472201f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_30 VNB N_A_193_47#_c_475_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_711_307#_M1021_g 0.0520206f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_32 VNB N_A_711_307#_c_586_n 0.0162836f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_33 VNB N_A_711_307#_c_587_n 0.019249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_711_307#_c_588_n 0.00485875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_711_307#_c_589_n 0.00322373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_711_307#_c_590_n 0.00231489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_711_307#_c_591_n 0.00115194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_711_307#_c_592_n 0.0381104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_560_47#_M1015_g 0.0239034f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_40 VNB N_A_560_47#_c_721_n 0.0514663f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_41 VNB N_A_560_47#_c_722_n 0.00860675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_560_47#_c_723_n 0.00802419f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_43 VNB N_A_560_47#_c_724_n 0.00353042f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_44 VNB N_A_560_47#_c_725_n 0.0108934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_806_n 0.016907f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_46 VNB N_RESET_B_c_807_n 0.0200615f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_47 VNB N_RESET_B_c_808_n 0.0039239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_846_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB Q 0.0191391f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_50 VNB N_Q_c_959_n 0.00583005f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_51 VNB N_VGND_c_1006_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1007_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1008_n 0.00605666f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_54 VNB N_VGND_c_1009_n 0.00222645f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1010_n 0.00988417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1011_n 0.0186875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1012_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1013_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1014_n 0.0407825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1015_n 0.0259377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1016_n 0.0172773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1017_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1018_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1019_n 0.00517156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1020_n 0.00506955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1021_n 0.333506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VPB N_GATE_N_c_146_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_68 VPB N_GATE_N_c_147_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_69 VPB N_GATE_N_c_148_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_70 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_71 VPB N_GATE_N_c_144_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_72 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_73 VPB N_A_27_47#_M1020_g 0.0200937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_196_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_75 VPB N_A_27_47#_c_197_n 0.0048535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_198_n 0.0270819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_199_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_188_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_201_n 0.027681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_202_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_203_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_204_n 0.00270156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_205_n 0.00363453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_192_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_193_n 2.87635e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_D_M1016_g 0.0462839f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_87 VPB N_D_c_352_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_88 VPB N_A_299_47#_M1012_g 0.0366887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_299_47#_c_398_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_299_47#_c_399_n 0.00403449f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_91 VPB N_A_299_47#_c_400_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_299_47#_c_394_n 0.00362722f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_93 VPB N_A_193_47#_M1001_g 0.0297186f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_94 VPB N_A_193_47#_c_472_n 0.0171022f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_95 VPB N_A_193_47#_c_473_n 0.00604992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_193_47#_c_479_n 0.0117991f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_97 VPB N_A_193_47#_c_475_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_193_47#_c_481_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_99 VPB N_A_193_47#_c_482_n 0.00515531f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_100 VPB N_A_193_47#_c_483_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_101 VPB N_A_193_47#_c_484_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_193_47#_c_485_n 0.00114133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_193_47#_c_486_n 0.0104341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_47#_c_487_n 0.0110271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_711_307#_M1009_g 0.0291236f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_106 VPB N_A_711_307#_M1021_g 0.01873f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_107 VPB N_A_711_307#_M1006_g 0.0187064f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_108 VPB N_A_711_307#_M1014_g 0.0226986f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_109 VPB N_A_711_307#_c_597_n 0.00572936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_711_307#_c_598_n 0.0478629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_711_307#_c_599_n 0.00169248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_711_307#_c_590_n 5.87434e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_711_307#_c_592_n 0.00710672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_560_47#_M1013_g 0.0267095f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_115 VPB N_A_560_47#_c_727_n 0.00679787f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_116 VPB N_A_560_47#_c_724_n 0.00488257f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_117 VPB N_RESET_B_M1019_g 0.0195761f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_118 VPB N_RESET_B_c_807_n 0.00411246f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_119 VPB N_RESET_B_c_808_n 0.00302832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_847_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_848_n 0.00342009f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_122 VPB N_VPWR_c_849_n 0.00803208f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_850_n 0.00107106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_851_n 3.26211e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_852_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_853_n 0.0359479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_854_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_855_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_856_n 0.0392932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_857_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_858_n 0.0154541f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_859_n 0.0164495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_860_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_861_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_862_n 0.00490136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_846_n 0.0571775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_Q_c_960_n 0.00642382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB Q 0.00390984f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_139 N_GATE_N_c_141_n N_A_27_47#_M1010_g 0.0187834f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_140 N_GATE_N_c_145_n N_A_27_47#_M1010_g 0.0041981f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_141 N_GATE_N_c_148_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_142 N_GATE_N_c_144_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_143 N_GATE_N_c_141_n N_A_27_47#_c_186_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_144 N_GATE_N_c_142_n N_A_27_47#_c_186_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_145 N_GATE_N_c_142_n N_A_27_47#_c_187_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_146 GATE_N N_A_27_47#_c_187_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_147 N_GATE_N_c_144_n N_A_27_47#_c_187_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_148 N_GATE_N_c_147_n N_A_27_47#_c_196_n 0.0135489f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_149 N_GATE_N_c_148_n N_A_27_47#_c_196_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_150 N_GATE_N_c_147_n N_A_27_47#_c_199_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_151 N_GATE_N_c_148_n N_A_27_47#_c_199_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_152 GATE_N N_A_27_47#_c_199_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_153 N_GATE_N_c_144_n N_A_27_47#_c_199_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_154 N_GATE_N_c_144_n N_A_27_47#_c_188_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_155 N_GATE_N_c_142_n N_A_27_47#_c_189_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_156 GATE_N N_A_27_47#_c_189_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_157 N_GATE_N_c_145_n N_A_27_47#_c_189_n 0.0015185f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_158 N_GATE_N_c_146_n N_A_27_47#_c_202_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_159 N_GATE_N_c_148_n N_A_27_47#_c_202_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_160 GATE_N N_A_27_47#_c_202_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_161 N_GATE_N_c_146_n N_A_27_47#_c_203_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_162 N_GATE_N_c_148_n N_A_27_47#_c_203_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_163 GATE_N N_A_27_47#_c_192_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_164 N_GATE_N_c_144_n N_A_27_47#_c_192_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_165 N_GATE_N_c_147_n N_VPWR_c_847_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_166 N_GATE_N_c_147_n N_VPWR_c_854_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_167 N_GATE_N_c_147_n N_VPWR_c_846_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_168 N_GATE_N_c_141_n N_VGND_c_1006_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_169 N_GATE_N_c_141_n N_VGND_c_1012_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_170 N_GATE_N_c_142_n N_VGND_c_1012_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_171 N_GATE_N_c_141_n N_VGND_c_1021_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_201_n N_D_M1016_g 0.00583826f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_201_n N_D_c_352_n 0.0087134f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1010_g N_D_c_353_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1017_g N_A_299_47#_c_390_n 0.0260428f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_191_n N_A_299_47#_c_390_n 2.11196e-19 $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_191_n N_A_299_47#_M1012_g 9.31407e-19 $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_201_n N_A_299_47#_M1012_g 0.00493352f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_193_n N_A_299_47#_M1012_g 0.00261248f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_180 N_A_27_47#_c_201_n N_A_299_47#_c_399_n 0.0114299f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_201_n N_A_299_47#_c_400_n 0.0115067f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_190_n N_A_299_47#_c_393_n 9.2948e-19 $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_191_n N_A_299_47#_c_393_n 0.0172223f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_201_n N_A_299_47#_c_393_n 0.00675641f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_191_n N_A_299_47#_c_394_n 0.0017693f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_201_n N_A_299_47#_c_394_n 0.0112945f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_190_n N_A_299_47#_c_396_n 0.0165895f $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_191_n N_A_299_47#_c_396_n 0.00208631f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_201_n N_A_299_47#_c_396_n 9.68438e-19 $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1020_g N_A_193_47#_M1001_g 0.0192024f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_197_n N_A_193_47#_M1001_g 0.00212148f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_198_n N_A_193_47#_c_472_n 0.0179236f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_191_n N_A_193_47#_c_472_n 0.00109701f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_201_n N_A_193_47#_c_472_n 0.00144279f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_204_n N_A_193_47#_c_472_n 0.00140497f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_205_n N_A_193_47#_c_472_n 0.00494665f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_193_n N_A_193_47#_c_472_n 0.0123877f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_190_n N_A_193_47#_c_473_n 0.0196536f $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_191_n N_A_193_47#_c_473_n 0.00521073f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_M1017_g N_A_193_47#_M1011_g 0.0121054f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_190_n N_A_193_47#_M1011_g 0.0157721f $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_191_n N_A_193_47#_M1011_g 0.00535958f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_193_n N_A_193_47#_M1011_g 0.00229612f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_204 N_A_27_47#_c_198_n N_A_193_47#_c_479_n 0.016035f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_201_n N_A_193_47#_c_479_n 0.00274258f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_204_n N_A_193_47#_c_479_n 7.88621e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_205_n N_A_193_47#_c_479_n 0.00212148f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_M1010_g N_A_193_47#_c_475_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_186_n N_A_193_47#_c_475_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_188_n N_A_193_47#_c_475_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_189_n N_A_193_47#_c_475_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_201_n N_A_193_47#_c_475_n 0.0184539f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_202_n N_A_193_47#_c_475_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_203_n N_A_193_47#_c_475_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_196_n N_A_193_47#_c_481_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_201_n N_A_193_47#_c_481_n 0.00195186f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_192_n N_A_193_47#_c_481_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_201_n N_A_193_47#_c_482_n 0.0871075f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_M1000_g N_A_193_47#_c_483_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_196_n N_A_193_47#_c_483_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_201_n N_A_193_47#_c_483_n 0.0259095f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_203_n N_A_193_47#_c_483_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_M1000_g N_A_193_47#_c_484_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_197_n N_A_193_47#_c_485_n 0.00155445f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_201_n N_A_193_47#_c_485_n 0.0255946f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_201_n N_A_193_47#_c_486_n 0.00162915f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_204_n N_A_193_47#_c_486_n 0.00124306f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_193_n N_A_193_47#_c_486_n 0.00212148f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_229 N_A_27_47#_c_198_n N_A_193_47#_c_487_n 2.60298e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_190_n N_A_193_47#_c_487_n 5.77836e-19 $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_191_n N_A_193_47#_c_487_n 0.00519043f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_201_n N_A_193_47#_c_487_n 0.0220946f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_204_n N_A_193_47#_c_487_n 0.00272314f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_193_n N_A_193_47#_c_487_n 0.0454941f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_M1020_g N_A_711_307#_M1009_g 0.0268652f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_197_n N_A_711_307#_M1009_g 3.32912e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_197_n N_A_711_307#_c_598_n 2.34066e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_198_n N_A_711_307#_c_598_n 0.0167148f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_205_n N_A_711_307#_c_598_n 3.81333e-19 $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_240 N_A_27_47#_M1020_g N_A_560_47#_c_729_n 0.00869479f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_197_n N_A_560_47#_c_729_n 0.0143694f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_198_n N_A_560_47#_c_729_n 0.00230542f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_204_n N_A_560_47#_c_729_n 0.00263773f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_190_n N_A_560_47#_c_733_n 6.30778e-19 $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_191_n N_A_560_47#_c_733_n 0.0196066f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_191_n N_A_560_47#_c_723_n 0.0205767f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_M1020_g N_A_560_47#_c_727_n 0.00558999f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_198_n N_A_560_47#_c_727_n 0.00167434f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_204_n N_A_560_47#_c_727_n 0.00129859f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_205_n N_A_560_47#_c_727_n 0.0436531f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_193_n N_A_560_47#_c_727_n 0.00387374f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_252 N_A_27_47#_c_198_n N_A_560_47#_c_725_n 5.33621e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_191_n N_A_560_47#_c_725_n 0.00854989f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_193_n N_A_560_47#_c_725_n 0.0105774f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_196_n N_VPWR_M1008_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A_27_47#_M1000_g N_VPWR_c_847_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_196_n N_VPWR_c_847_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_199_n N_VPWR_c_847_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_202_n N_VPWR_c_847_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_201_n N_VPWR_c_848_n 0.00195141f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_196_n N_VPWR_c_854_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_199_n N_VPWR_c_854_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_263 N_A_27_47#_M1000_g N_VPWR_c_855_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1020_g N_VPWR_c_856_n 0.00366111f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1000_g N_VPWR_c_846_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1020_g N_VPWR_c_846_n 0.00544154f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_196_n N_VPWR_c_846_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_199_n N_VPWR_c_846_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_186_n N_VGND_M1018_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_270 N_A_27_47#_M1010_g N_VGND_c_1006_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_186_n N_VGND_c_1006_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_188_n N_VGND_c_1006_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_192_n N_VGND_c_1006_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1017_g N_VGND_c_1007_n 0.00184233f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_337_p N_VGND_c_1012_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_186_n N_VGND_c_1012_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_M1010_g N_VGND_c_1013_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1017_g N_VGND_c_1014_n 0.00460154f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_190_n N_VGND_c_1014_n 0.00105849f $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_191_n N_VGND_c_1014_n 0.00203207f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_M1018_s N_VGND_c_1021_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1010_g N_VGND_c_1021_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1017_g N_VGND_c_1021_n 0.00720224f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_337_p N_VGND_c_1021_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_186_n N_VGND_c_1021_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_190_n N_VGND_c_1021_n 0.00125829f $X=2.765 $Y=0.9 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_191_n N_VGND_c_1021_n 0.00373364f $X=3.01 $Y=0.925 $X2=0
+ $Y2=0
cc_288 N_D_M1002_g N_A_299_47#_c_390_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_289 N_D_c_353_n N_A_299_47#_M1012_g 0.0381981f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_290 N_D_M1016_g N_A_299_47#_c_398_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_291 N_D_M1002_g N_A_299_47#_c_392_n 0.0144458f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_292 N_D_c_352_n N_A_299_47#_c_392_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_293 N_D_c_353_n N_A_299_47#_c_392_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_294 N_D_M1016_g N_A_299_47#_c_399_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_295 N_D_M1016_g N_A_299_47#_c_400_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_296 N_D_c_352_n N_A_299_47#_c_400_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_297 N_D_c_353_n N_A_299_47#_c_400_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_298 N_D_M1002_g N_A_299_47#_c_393_n 0.00569145f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_299 N_D_c_352_n N_A_299_47#_c_393_n 0.0112581f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_300 N_D_c_352_n N_A_299_47#_c_394_n 0.0172838f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_301 N_D_c_353_n N_A_299_47#_c_394_n 0.00562919f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_302 N_D_M1002_g N_A_299_47#_c_395_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_303 N_D_c_352_n N_A_299_47#_c_395_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_304 N_D_c_353_n N_A_299_47#_c_395_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_305 N_D_M1002_g N_A_299_47#_c_396_n 0.0203127f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_306 N_D_M1002_g N_A_193_47#_c_475_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_307 N_D_M1016_g N_A_193_47#_c_475_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_308 N_D_c_352_n N_A_193_47#_c_475_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_309 N_D_c_353_n N_A_193_47#_c_475_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_310 N_D_M1016_g N_A_193_47#_c_481_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_311 N_D_M1016_g N_A_193_47#_c_482_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_312 N_D_M1016_g N_VPWR_c_848_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_313 N_D_M1016_g N_VPWR_c_855_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_314 N_D_M1016_g N_VPWR_c_846_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_315 N_D_M1002_g N_VGND_c_1007_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_316 N_D_M1002_g N_VGND_c_1013_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_317 N_D_M1002_g N_VGND_c_1021_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_318 N_D_c_353_n N_VGND_c_1021_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_319 N_A_299_47#_M1012_g N_A_193_47#_M1001_g 0.0340556f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_320 N_A_299_47#_M1012_g N_A_193_47#_c_473_n 0.024821f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_321 N_A_299_47#_c_398_n N_A_193_47#_c_475_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_322 N_A_299_47#_c_400_n N_A_193_47#_c_475_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_323 N_A_299_47#_c_395_n N_A_193_47#_c_475_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_324 N_A_299_47#_c_398_n N_A_193_47#_c_481_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_325 N_A_299_47#_M1012_g N_A_193_47#_c_482_n 0.00365242f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_326 N_A_299_47#_c_398_n N_A_193_47#_c_482_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_327 N_A_299_47#_c_399_n N_A_193_47#_c_482_n 0.00558649f $X=1.96 $Y=1.58 $X2=0
+ $Y2=0
cc_328 N_A_299_47#_c_398_n N_A_193_47#_c_483_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_299_47#_M1012_g N_A_193_47#_c_485_n 0.00149195f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_330 N_A_299_47#_M1012_g N_A_193_47#_c_487_n 0.00673436f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_331 N_A_299_47#_c_399_n N_A_193_47#_c_487_n 0.00754519f $X=1.96 $Y=1.58 $X2=0
+ $Y2=0
cc_332 N_A_299_47#_c_394_n N_A_193_47#_c_487_n 0.00647732f $X=2.05 $Y=1.495
+ $X2=0 $Y2=0
cc_333 N_A_299_47#_M1012_g N_A_560_47#_c_729_n 5.00797e-19 $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_334 N_A_299_47#_M1012_g N_VPWR_c_848_n 0.0220604f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_398_n N_VPWR_c_848_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_336 N_A_299_47#_c_399_n N_VPWR_c_848_n 0.0133983f $X=1.96 $Y=1.58 $X2=0 $Y2=0
cc_337 N_A_299_47#_c_398_n N_VPWR_c_855_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_338 N_A_299_47#_M1012_g N_VPWR_c_856_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_339 N_A_299_47#_M1016_s N_VPWR_c_846_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_M1012_g N_VPWR_c_846_n 0.00262666f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_341 N_A_299_47#_c_398_n N_VPWR_c_846_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_342 N_A_299_47#_c_393_n N_VGND_M1002_d 0.00165422f $X=2.05 $Y=1.095 $X2=0
+ $Y2=0
cc_343 N_A_299_47#_c_390_n N_VGND_c_1007_n 0.00946131f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_344 N_A_299_47#_c_392_n N_VGND_c_1007_n 0.0020169f $X=1.96 $Y=0.7 $X2=0 $Y2=0
cc_345 N_A_299_47#_c_393_n N_VGND_c_1007_n 0.0148674f $X=2.05 $Y=1.095 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_c_392_n N_VGND_c_1013_n 0.00255672f $X=1.96 $Y=0.7 $X2=0
+ $Y2=0
cc_347 N_A_299_47#_c_395_n N_VGND_c_1013_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_348 N_A_299_47#_c_390_n N_VGND_c_1014_n 0.0046653f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_349 N_A_299_47#_c_396_n N_VGND_c_1014_n 8.97291e-19 $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_350 N_A_299_47#_M1002_s N_VGND_c_1021_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_351 N_A_299_47#_c_390_n N_VGND_c_1021_n 0.00440683f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_352 N_A_299_47#_c_392_n N_VGND_c_1021_n 0.00468534f $X=1.96 $Y=0.7 $X2=0
+ $Y2=0
cc_353 N_A_299_47#_c_393_n N_VGND_c_1021_n 0.00557078f $X=2.05 $Y=1.095 $X2=0
+ $Y2=0
cc_354 N_A_299_47#_c_395_n N_VGND_c_1021_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_355 N_A_299_47#_c_396_n N_VGND_c_1021_n 0.0010595f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_356 N_A_193_47#_M1011_g N_A_711_307#_M1021_g 0.0424218f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_357 N_A_193_47#_M1001_g N_A_560_47#_c_729_n 0.00454949f $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_358 N_A_193_47#_M1011_g N_A_560_47#_c_733_n 0.0125446f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_359 N_A_193_47#_M1011_g N_A_560_47#_c_723_n 0.00583764f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_360 N_A_193_47#_M1001_g N_A_560_47#_c_727_n 4.33428e-19 $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_361 N_A_193_47#_c_472_n N_A_560_47#_c_727_n 6.91978e-19 $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_362 N_A_193_47#_c_472_n N_A_560_47#_c_725_n 9.24158e-19 $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_M1011_g N_A_560_47#_c_725_n 0.00228104f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_364 N_A_193_47#_c_482_n N_VPWR_M1016_d 6.81311e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_365 N_A_193_47#_c_484_n N_VPWR_c_847_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_193_47#_M1001_g N_VPWR_c_848_n 0.00354746f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_367 N_A_193_47#_c_482_n N_VPWR_c_848_n 0.0171704f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_368 N_A_193_47#_c_485_n N_VPWR_c_848_n 0.0013481f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_193_47#_c_487_n N_VPWR_c_848_n 0.00972665f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_484_n N_VPWR_c_855_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_371 N_A_193_47#_M1001_g N_VPWR_c_856_n 0.00443167f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_487_n N_VPWR_c_856_n 0.00456724f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_373 N_A_193_47#_M1001_g N_VPWR_c_846_n 0.00660849f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_482_n N_VPWR_c_846_n 0.0516753f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_375 N_A_193_47#_c_483_n N_VPWR_c_846_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_376 N_A_193_47#_c_484_n N_VPWR_c_846_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_485_n N_VPWR_c_846_n 0.0151013f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_c_487_n N_VPWR_c_846_n 0.00403974f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_482_n A_465_369# 0.00119229f $X=2.41 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_380 N_A_193_47#_c_485_n A_465_369# 0.00120144f $X=2.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_381 N_A_193_47#_c_487_n A_465_369# 0.0030615f $X=2.67 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_193_47#_M1011_g N_VGND_c_1008_n 0.00172953f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_c_475_n N_VGND_c_1013_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_M1011_g N_VGND_c_1014_n 0.0037981f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_385 N_A_193_47#_M1010_d N_VGND_c_1021_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_386 N_A_193_47#_M1011_g N_VGND_c_1021_n 0.00570274f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_387 N_A_193_47#_c_475_n N_VGND_c_1021_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_388 N_A_711_307#_c_597_n N_A_560_47#_M1013_g 0.0166405f $X=4.73 $Y=1.7 $X2=0
+ $Y2=0
cc_389 N_A_711_307#_c_598_n N_A_560_47#_M1013_g 0.00687993f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_390 N_A_711_307#_c_588_n N_A_560_47#_M1015_g 0.00755158f $X=4.42 $Y=0.4 $X2=0
+ $Y2=0
cc_391 N_A_711_307#_c_611_p N_A_560_47#_M1015_g 0.00793834f $X=5.415 $Y=0.74
+ $X2=0 $Y2=0
cc_392 N_A_711_307#_c_589_n N_A_560_47#_M1015_g 0.00101901f $X=4.59 $Y=0.74
+ $X2=0 $Y2=0
cc_393 N_A_711_307#_M1021_g N_A_560_47#_c_721_n 0.0170245f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_394 N_A_711_307#_c_597_n N_A_560_47#_c_721_n 0.00823747f $X=4.73 $Y=1.7 $X2=0
+ $Y2=0
cc_395 N_A_711_307#_c_598_n N_A_560_47#_c_721_n 0.00424117f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_396 N_A_711_307#_c_589_n N_A_560_47#_c_721_n 0.00886838f $X=4.59 $Y=0.74
+ $X2=0 $Y2=0
cc_397 N_A_711_307#_M1009_g N_A_560_47#_c_729_n 0.00500469f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_398 N_A_711_307#_M1021_g N_A_560_47#_c_733_n 0.00159883f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_399 N_A_711_307#_M1021_g N_A_560_47#_c_723_n 0.0110627f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_400 N_A_711_307#_M1009_g N_A_560_47#_c_727_n 0.0159393f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_401 N_A_711_307#_M1021_g N_A_560_47#_c_727_n 0.00748409f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_711_307#_c_597_n N_A_560_47#_c_727_n 0.0206864f $X=4.73 $Y=1.7 $X2=0
+ $Y2=0
cc_403 N_A_711_307#_c_598_n N_A_560_47#_c_727_n 0.0101307f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_404 N_A_711_307#_M1021_g N_A_560_47#_c_724_n 0.0238827f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_405 N_A_711_307#_c_597_n N_A_560_47#_c_724_n 0.0338662f $X=4.73 $Y=1.7 $X2=0
+ $Y2=0
cc_406 N_A_711_307#_c_598_n N_A_560_47#_c_724_n 0.00653921f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_407 N_A_711_307#_c_589_n N_A_560_47#_c_724_n 0.0050906f $X=4.59 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_711_307#_M1006_g N_RESET_B_M1019_g 0.0221506f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_711_307#_c_629_p N_RESET_B_M1019_g 0.0131717f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_410 N_A_711_307#_c_599_n N_RESET_B_M1019_g 0.00299828f $X=5.5 $Y=1.535 $X2=0
+ $Y2=0
cc_411 N_A_711_307#_c_586_n N_RESET_B_c_806_n 0.0240078f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_412 N_A_711_307#_c_588_n N_RESET_B_c_806_n 0.00152503f $X=4.42 $Y=0.4 $X2=0
+ $Y2=0
cc_413 N_A_711_307#_c_611_p N_RESET_B_c_806_n 0.0118724f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_414 N_A_711_307#_c_591_n N_RESET_B_c_806_n 0.00311071f $X=5.482 $Y=0.995
+ $X2=0 $Y2=0
cc_415 N_A_711_307#_c_611_p N_RESET_B_c_807_n 0.0025449f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_711_307#_c_629_p N_RESET_B_c_807_n 0.00176617f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_417 N_A_711_307#_c_590_n N_RESET_B_c_807_n 0.00186324f $X=5.53 $Y=1.16 $X2=0
+ $Y2=0
cc_418 N_A_711_307#_c_592_n N_RESET_B_c_807_n 0.0203929f $X=5.97 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_711_307#_c_597_n N_RESET_B_c_808_n 0.0131995f $X=4.73 $Y=1.7 $X2=0
+ $Y2=0
cc_420 N_A_711_307#_c_611_p N_RESET_B_c_808_n 0.037239f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_421 N_A_711_307#_c_589_n N_RESET_B_c_808_n 0.00663756f $X=4.59 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A_711_307#_c_629_p N_RESET_B_c_808_n 0.0123079f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_423 N_A_711_307#_c_643_p N_RESET_B_c_808_n 0.0128063f $X=4.825 $Y=1.755 $X2=0
+ $Y2=0
cc_424 N_A_711_307#_c_590_n N_RESET_B_c_808_n 0.0259555f $X=5.53 $Y=1.16 $X2=0
+ $Y2=0
cc_425 N_A_711_307#_c_592_n N_RESET_B_c_808_n 3.60538e-19 $X=5.97 $Y=1.16 $X2=0
+ $Y2=0
cc_426 N_A_711_307#_c_597_n N_VPWR_M1013_s 0.00664759f $X=4.73 $Y=1.7 $X2=0
+ $Y2=0
cc_427 N_A_711_307#_c_629_p N_VPWR_M1019_d 0.00911213f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_428 N_A_711_307#_M1009_g N_VPWR_c_849_n 0.0065946f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_429 N_A_711_307#_c_597_n N_VPWR_c_849_n 0.015605f $X=4.73 $Y=1.7 $X2=0 $Y2=0
cc_430 N_A_711_307#_c_598_n N_VPWR_c_849_n 0.00593927f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_431 N_A_711_307#_c_597_n N_VPWR_c_850_n 0.0120619f $X=4.73 $Y=1.7 $X2=0 $Y2=0
cc_432 N_A_711_307#_M1006_g N_VPWR_c_851_n 0.0106598f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_433 N_A_711_307#_M1014_g N_VPWR_c_851_n 7.49e-19 $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_434 N_A_711_307#_c_629_p N_VPWR_c_851_n 0.0205447f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_435 N_A_711_307#_M1014_g N_VPWR_c_853_n 0.00442893f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_436 N_A_711_307#_M1009_g N_VPWR_c_856_n 0.00512226f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_437 N_A_711_307#_c_657_p N_VPWR_c_857_n 0.0121054f $X=4.825 $Y=2.27 $X2=0
+ $Y2=0
cc_438 N_A_711_307#_M1006_g N_VPWR_c_859_n 0.00505556f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_439 N_A_711_307#_M1014_g N_VPWR_c_859_n 0.00541359f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_440 N_A_711_307#_M1013_d N_VPWR_c_846_n 0.00385995f $X=4.69 $Y=1.485 $X2=0
+ $Y2=0
cc_441 N_A_711_307#_M1009_g N_VPWR_c_846_n 0.0103819f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_442 N_A_711_307#_M1006_g N_VPWR_c_846_n 0.00859622f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_443 N_A_711_307#_M1014_g N_VPWR_c_846_n 0.0105459f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_711_307#_c_597_n N_VPWR_c_846_n 0.0135362f $X=4.73 $Y=1.7 $X2=0 $Y2=0
cc_445 N_A_711_307#_c_598_n N_VPWR_c_846_n 0.00230567f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_446 N_A_711_307#_c_657_p N_VPWR_c_846_n 0.00724021f $X=4.825 $Y=2.27 $X2=0
+ $Y2=0
cc_447 N_A_711_307#_c_586_n N_Q_c_962_n 0.00407088f $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A_711_307#_c_587_n N_Q_c_962_n 0.00971895f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_449 N_A_711_307#_c_611_p N_Q_c_962_n 0.00860939f $X=5.415 $Y=0.74 $X2=0 $Y2=0
cc_450 N_A_711_307#_c_586_n N_Q_c_965_n 0.00360736f $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_451 N_A_711_307#_c_587_n N_Q_c_965_n 0.00285458f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_452 N_A_711_307#_c_590_n N_Q_c_965_n 5.67058e-19 $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_453 N_A_711_307#_c_592_n N_Q_c_965_n 0.00115756f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_454 N_A_711_307#_M1006_g N_Q_c_969_n 0.00304202f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_711_307#_M1014_g N_Q_c_969_n 0.00283598f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_456 N_A_711_307#_c_592_n N_Q_c_969_n 0.00228063f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_711_307#_M1006_g N_Q_c_972_n 0.00476088f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_A_711_307#_M1014_g N_Q_c_972_n 0.0120309f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_459 N_A_711_307#_c_629_p N_Q_c_972_n 0.0133619f $X=5.415 $Y=1.62 $X2=0 $Y2=0
cc_460 N_A_711_307#_c_599_n N_Q_c_972_n 0.00238698f $X=5.5 $Y=1.535 $X2=0 $Y2=0
cc_461 N_A_711_307#_M1006_g N_Q_c_960_n 7.59735e-19 $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_462 N_A_711_307#_M1014_g N_Q_c_960_n 0.0110611f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_463 N_A_711_307#_c_599_n N_Q_c_960_n 0.00895287f $X=5.5 $Y=1.535 $X2=0 $Y2=0
cc_464 N_A_711_307#_c_592_n N_Q_c_960_n 9.62648e-19 $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_465 N_A_711_307#_M1014_g Q 0.00617274f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_466 N_A_711_307#_M1006_g Q 3.91463e-19 $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_467 N_A_711_307#_c_586_n Q 6.9963e-19 $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_468 N_A_711_307#_c_587_n Q 0.00417216f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_469 N_A_711_307#_M1014_g Q 0.00239602f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_470 N_A_711_307#_c_599_n Q 0.00413456f $X=5.5 $Y=1.535 $X2=0 $Y2=0
cc_471 N_A_711_307#_c_590_n Q 0.0254346f $X=5.53 $Y=1.16 $X2=0 $Y2=0
cc_472 N_A_711_307#_c_591_n Q 0.00728749f $X=5.482 $Y=0.995 $X2=0 $Y2=0
cc_473 N_A_711_307#_c_592_n Q 0.0202106f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_474 N_A_711_307#_c_586_n N_Q_c_959_n 8.34038e-19 $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_475 N_A_711_307#_c_587_n N_Q_c_959_n 0.00811298f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_476 N_A_711_307#_c_611_p N_Q_c_959_n 0.00519448f $X=5.415 $Y=0.74 $X2=0 $Y2=0
cc_477 N_A_711_307#_c_591_n N_Q_c_959_n 0.00492401f $X=5.482 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_711_307#_c_592_n N_Q_c_959_n 8.81346e-19 $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_711_307#_c_611_p N_VGND_M1007_d 0.00920577f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_480 N_A_711_307#_c_591_n N_VGND_M1007_d 7.52091e-19 $X=5.482 $Y=0.995 $X2=0
+ $Y2=0
cc_481 N_A_711_307#_M1021_g N_VGND_c_1008_n 0.0115353f $X=3.69 $Y=0.445 $X2=0
+ $Y2=0
cc_482 N_A_711_307#_c_588_n N_VGND_c_1008_n 0.0230272f $X=4.42 $Y=0.4 $X2=0
+ $Y2=0
cc_483 N_A_711_307#_c_586_n N_VGND_c_1009_n 0.00295374f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_A_711_307#_c_588_n N_VGND_c_1009_n 0.00712945f $X=4.42 $Y=0.4 $X2=0
+ $Y2=0
cc_485 N_A_711_307#_c_611_p N_VGND_c_1009_n 0.020151f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_711_307#_c_587_n N_VGND_c_1011_n 0.00360303f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_A_711_307#_M1021_g N_VGND_c_1014_n 0.0046653f $X=3.69 $Y=0.445 $X2=0
+ $Y2=0
cc_488 N_A_711_307#_c_588_n N_VGND_c_1015_n 0.022192f $X=4.42 $Y=0.4 $X2=0 $Y2=0
cc_489 N_A_711_307#_c_611_p N_VGND_c_1015_n 0.00732922f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_490 N_A_711_307#_c_586_n N_VGND_c_1016_n 0.00424377f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_491 N_A_711_307#_c_587_n N_VGND_c_1016_n 0.00539883f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_492 N_A_711_307#_c_611_p N_VGND_c_1016_n 0.00234481f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_A_711_307#_M1015_s N_VGND_c_1021_n 0.00209319f $X=4.295 $Y=0.235 $X2=0
+ $Y2=0
cc_494 N_A_711_307#_M1021_g N_VGND_c_1021_n 0.00813035f $X=3.69 $Y=0.445 $X2=0
+ $Y2=0
cc_495 N_A_711_307#_c_586_n N_VGND_c_1021_n 0.00617479f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_496 N_A_711_307#_c_587_n N_VGND_c_1021_n 0.00674774f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_A_711_307#_c_588_n N_VGND_c_1021_n 0.0131132f $X=4.42 $Y=0.4 $X2=0
+ $Y2=0
cc_498 N_A_711_307#_c_611_p N_VGND_c_1021_n 0.0185208f $X=5.415 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_711_307#_c_611_p A_941_47# 0.00441372f $X=5.415 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_500 N_A_560_47#_M1013_g N_RESET_B_M1019_g 0.0244798f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_501 N_A_560_47#_M1015_g N_RESET_B_c_806_n 0.0424066f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_502 N_A_560_47#_M1013_g N_RESET_B_c_807_n 0.00145765f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_503 N_A_560_47#_M1015_g N_RESET_B_c_807_n 0.0198038f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_504 N_A_560_47#_M1013_g N_RESET_B_c_808_n 0.00315875f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_505 N_A_560_47#_M1015_g N_RESET_B_c_808_n 0.00319632f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_506 N_A_560_47#_c_721_n N_RESET_B_c_808_n 0.00709983f $X=4.54 $Y=1.16 $X2=0
+ $Y2=0
cc_507 N_A_560_47#_c_722_n N_RESET_B_c_808_n 0.00730491f $X=4.622 $Y=1.162 $X2=0
+ $Y2=0
cc_508 N_A_560_47#_c_724_n N_RESET_B_c_808_n 0.0255162f $X=4.145 $Y=1.16 $X2=0
+ $Y2=0
cc_509 N_A_560_47#_c_729_n N_VPWR_c_848_n 0.00547986f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_510 N_A_560_47#_M1013_g N_VPWR_c_849_n 0.00103168f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_A_560_47#_c_729_n N_VPWR_c_849_n 0.0125356f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_512 N_A_560_47#_c_727_n N_VPWR_c_849_n 0.00791951f $X=3.52 $Y=2.255 $X2=0
+ $Y2=0
cc_513 N_A_560_47#_M1013_g N_VPWR_c_850_n 0.00851573f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_514 N_A_560_47#_M1013_g N_VPWR_c_851_n 6.54137e-19 $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_515 N_A_560_47#_c_729_n N_VPWR_c_856_n 0.0370561f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_516 N_A_560_47#_M1013_g N_VPWR_c_858_n 0.00535584f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_517 N_A_560_47#_M1001_d N_VPWR_c_846_n 0.00217615f $X=2.805 $Y=2.065 $X2=0
+ $Y2=0
cc_518 N_A_560_47#_M1013_g N_VPWR_c_846_n 0.00478989f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_519 N_A_560_47#_c_729_n N_VPWR_c_846_n 0.029179f $X=3.435 $Y=2.34 $X2=0 $Y2=0
cc_520 N_A_560_47#_c_729_n A_645_413# 0.00648275f $X=3.435 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_521 N_A_560_47#_c_727_n A_645_413# 0.00225548f $X=3.52 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_522 N_A_560_47#_M1015_g N_VGND_c_1008_n 0.0023728f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_523 N_A_560_47#_c_721_n N_VGND_c_1008_n 0.00160278f $X=4.54 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_A_560_47#_c_733_n N_VGND_c_1008_n 0.0106425f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_525 N_A_560_47#_c_724_n N_VGND_c_1008_n 0.0115522f $X=4.145 $Y=1.16 $X2=0
+ $Y2=0
cc_526 N_A_560_47#_M1015_g N_VGND_c_1009_n 0.00181288f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_527 N_A_560_47#_c_733_n N_VGND_c_1014_n 0.0235028f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_528 N_A_560_47#_M1015_g N_VGND_c_1015_n 0.00413124f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_529 N_A_560_47#_M1017_d N_VGND_c_1021_n 0.0029318f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_530 N_A_560_47#_M1015_g N_VGND_c_1021_n 0.00707749f $X=4.63 $Y=0.56 $X2=0
+ $Y2=0
cc_531 N_A_560_47#_c_733_n N_VGND_c_1021_n 0.0234633f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_532 N_A_560_47#_c_733_n A_658_47# 0.0037502f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_533 N_A_560_47#_c_723_n A_658_47# 0.00152789f $X=3.415 $Y=1.025 $X2=-0.19
+ $Y2=-0.24
cc_534 N_RESET_B_M1019_g N_VPWR_c_850_n 5.74285e-19 $X=5.035 $Y=1.985 $X2=0
+ $Y2=0
cc_535 N_RESET_B_M1019_g N_VPWR_c_851_n 0.0100483f $X=5.035 $Y=1.985 $X2=0 $Y2=0
cc_536 N_RESET_B_M1019_g N_VPWR_c_857_n 0.00505556f $X=5.035 $Y=1.985 $X2=0
+ $Y2=0
cc_537 N_RESET_B_M1019_g N_VPWR_c_846_n 0.00861019f $X=5.035 $Y=1.985 $X2=0
+ $Y2=0
cc_538 N_RESET_B_c_806_n N_VGND_c_1009_n 0.00968908f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_539 N_RESET_B_c_806_n N_VGND_c_1015_n 0.00341689f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_RESET_B_c_806_n N_VGND_c_1021_n 0.00405445f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_846_n A_465_369# 0.00373974f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_542 N_VPWR_c_846_n A_645_413# 0.00267918f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_543 N_VPWR_c_846_n N_Q_M1006_d 0.00468958f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_544 N_VPWR_c_851_n N_Q_c_969_n 0.0408895f $X=5.275 $Y=2.02 $X2=0 $Y2=0
cc_545 N_VPWR_M1014_s N_Q_c_960_n 0.00231287f $X=6.045 $Y=1.485 $X2=0 $Y2=0
cc_546 N_VPWR_c_853_n N_Q_c_960_n 0.022894f $X=6.18 $Y=1.835 $X2=0 $Y2=0
cc_547 N_VPWR_c_859_n Q 0.0166934f $X=6.095 $Y=2.72 $X2=0 $Y2=0
cc_548 N_VPWR_c_846_n Q 0.010102f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_549 N_Q_c_959_n N_VGND_M1005_s 0.00273341f $X=6.07 $Y=0.89 $X2=0 $Y2=0
cc_550 N_Q_c_959_n N_VGND_c_1011_n 0.0221752f $X=6.07 $Y=0.89 $X2=0 $Y2=0
cc_551 N_Q_c_965_n N_VGND_c_1016_n 0.0178243f $X=5.84 $Y=0.37 $X2=0 $Y2=0
cc_552 N_Q_M1003_d N_VGND_c_1021_n 0.00215227f $X=5.625 $Y=0.235 $X2=0 $Y2=0
cc_553 N_Q_c_965_n N_VGND_c_1021_n 0.0119575f $X=5.84 $Y=0.37 $X2=0 $Y2=0
cc_554 N_Q_c_959_n N_VGND_c_1021_n 0.00719248f $X=6.07 $Y=0.89 $X2=0 $Y2=0
cc_555 N_VGND_c_1021_n A_465_47# 0.0111582f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_556 N_VGND_c_1021_n A_658_47# 0.00669936f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_557 N_VGND_c_1021_n A_941_47# 0.00323135f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24

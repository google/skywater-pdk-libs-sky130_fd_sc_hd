* File: sky130_fd_sc_hd__o311ai_2.pex.spice
* Created: Tue Sep  1 19:24:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311AI_2%A1 3 7 11 15 17 18 26 28
c40 26 0 6.18781e-20 $X=0.94 $Y=1.16
c41 11 0 7.11327e-20 $X=1.01 $Y=1.985
r42 27 28 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=1.01 $Y=1.16 $X2=1.03
+ $Y2=1.16
r43 25 27 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=0.94 $Y=1.16 $X2=1.01
+ $Y2=1.16
r44 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r45 23 25 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=0.61 $Y=1.16
+ $X2=0.94 $Y2=1.16
r46 21 23 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=0.59 $Y=1.16 $X2=0.61
+ $Y2=1.16
r47 18 26 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=1.185
+ $X2=0.94 $Y2=1.185
r48 17 18 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=0.23 $Y=1.185
+ $X2=0.69 $Y2=1.185
r49 13 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.03 $Y=1.025
+ $X2=1.03 $Y2=1.16
r50 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.03 $Y=1.025
+ $X2=1.03 $Y2=0.56
r51 9 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.01 $Y=1.295
+ $X2=1.01 $Y2=1.16
r52 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.01 $Y=1.295
+ $X2=1.01 $Y2=1.985
r53 5 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.61 $Y=1.025
+ $X2=0.61 $Y2=1.16
r54 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.61 $Y=1.025
+ $X2=0.61 $Y2=0.56
r55 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.59 $Y=1.295
+ $X2=0.59 $Y2=1.16
r56 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.59 $Y=1.295 $X2=0.59
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%A2 3 7 11 15 17 18 28
c50 28 0 1.83965e-19 $X=1.87 $Y=1.16
c51 18 0 1.37236e-19 $X=2.07 $Y=1.19
c52 11 0 8.77293e-20 $X=1.85 $Y=1.985
c53 3 0 6.18781e-20 $X=1.43 $Y=1.985
r54 27 28 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=1.85 $Y=1.16 $X2=1.87
+ $Y2=1.16
r55 25 27 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=1.82 $Y=1.16 $X2=1.85
+ $Y2=1.16
r56 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.16 $X2=1.82 $Y2=1.16
r57 23 25 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=1.45 $Y=1.16
+ $X2=1.82 $Y2=1.16
r58 21 23 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=1.43 $Y=1.16 $X2=1.45
+ $Y2=1.16
r59 18 26 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=2.07 $Y=1.185
+ $X2=1.82 $Y2=1.185
r60 17 26 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.61 $Y=1.185
+ $X2=1.82 $Y2=1.185
r61 13 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.87 $Y=1.025
+ $X2=1.87 $Y2=1.16
r62 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.87 $Y=1.025
+ $X2=1.87 $Y2=0.56
r63 9 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.85 $Y=1.295
+ $X2=1.85 $Y2=1.16
r64 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.85 $Y=1.295
+ $X2=1.85 $Y2=1.985
r65 5 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.45 $Y=1.025
+ $X2=1.45 $Y2=1.16
r66 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.45 $Y=1.025
+ $X2=1.45 $Y2=0.56
r67 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.43 $Y=1.295
+ $X2=1.43 $Y2=1.16
r68 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.43 $Y=1.295 $X2=1.43
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%A3 3 7 11 15 17 18 19 22 31
c48 19 0 5.92676e-19 $X=2.99 $Y=1.19
c49 7 0 6.61036e-20 $X=2.79 $Y=1.985
r50 30 31 13.3304 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=3.15 $Y=1.16 $X2=3.21
+ $Y2=1.16
r51 28 30 71.0956 $w=2.7e-07 $l=3.2e-07 $layer=POLY_cond $X=2.83 $Y=1.16
+ $X2=3.15 $Y2=1.16
r52 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.16 $X2=2.83 $Y2=1.16
r53 26 28 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=2.79 $Y=1.16 $X2=2.83
+ $Y2=1.16
r54 22 26 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.715 $Y=1.16
+ $X2=2.79 $Y2=1.16
r55 22 24 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=2.715 $Y=1.16
+ $X2=2.49 $Y2=1.16
r56 19 29 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=2.99 $Y=1.185
+ $X2=2.83 $Y2=1.185
r57 18 29 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.49 $Y=1.185
+ $X2=2.83 $Y2=1.185
r58 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.16 $X2=2.49 $Y2=1.16
r59 17 24 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.365 $Y=1.16
+ $X2=2.49 $Y2=1.16
r60 13 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.21 $Y=1.295
+ $X2=3.21 $Y2=1.16
r61 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.21 $Y=1.295
+ $X2=3.21 $Y2=1.985
r62 9 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.15 $Y=1.025
+ $X2=3.15 $Y2=1.16
r63 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.15 $Y=1.025
+ $X2=3.15 $Y2=0.56
r64 5 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.79 $Y=1.295
+ $X2=2.79 $Y2=1.16
r65 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.79 $Y=1.295 $X2=2.79
+ $Y2=1.985
r66 1 17 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.29 $Y=1.025
+ $X2=2.365 $Y2=1.16
r67 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.29 $Y=1.025
+ $X2=2.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%B1 3 7 11 15 17 18 27 28
c44 28 0 2.34477e-19 $X=4.39 $Y=1.16
c45 27 0 1.85039e-19 $X=4 $Y=1.16
r46 26 28 86.6477 $w=2.7e-07 $l=3.9e-07 $layer=POLY_cond $X=4 $Y=1.16 $X2=4.39
+ $Y2=1.16
r47 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4 $Y=1.16
+ $X2=4 $Y2=1.16
r48 24 26 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=3.99 $Y=1.16 $X2=4
+ $Y2=1.16
r49 23 24 79.9825 $w=2.7e-07 $l=3.6e-07 $layer=POLY_cond $X=3.63 $Y=1.16
+ $X2=3.99 $Y2=1.16
r50 21 23 13.3304 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=3.57 $Y=1.16 $X2=3.63
+ $Y2=1.16
r51 18 27 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=3.91 $Y=1.185 $X2=4
+ $Y2=1.185
r52 17 18 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=3.45 $Y=1.185
+ $X2=3.91 $Y2=1.185
r53 13 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.39 $Y=1.295
+ $X2=4.39 $Y2=1.16
r54 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.39 $Y=1.295
+ $X2=4.39 $Y2=1.985
r55 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.99 $Y=1.025
+ $X2=3.99 $Y2=1.16
r56 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.99 $Y=1.025
+ $X2=3.99 $Y2=0.56
r57 5 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.63 $Y=1.295
+ $X2=3.63 $Y2=1.16
r58 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.63 $Y=1.295 $X2=3.63
+ $Y2=1.985
r59 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.57 $Y=1.025
+ $X2=3.57 $Y2=1.16
r60 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.57 $Y=1.025
+ $X2=3.57 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%C1 3 7 11 15 17 18 21 23
c43 21 0 1.85039e-19 $X=5.465 $Y=1.16
r44 32 33 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=5.37 $Y=1.16 $X2=5.39
+ $Y2=1.16
r45 30 32 26.6608 $w=2.7e-07 $l=1.2e-07 $layer=POLY_cond $X=5.25 $Y=1.16
+ $X2=5.37 $Y2=1.16
r46 28 30 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=4.97 $Y=1.16
+ $X2=5.25 $Y2=1.16
r47 26 28 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=4.95 $Y=1.16 $X2=4.97
+ $Y2=1.16
r48 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.16 $X2=5.59 $Y2=1.16
r49 21 33 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.465 $Y=1.16
+ $X2=5.39 $Y2=1.16
r50 21 23 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=5.465 $Y=1.16
+ $X2=5.59 $Y2=1.16
r51 18 24 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=5.75 $Y=1.185
+ $X2=5.59 $Y2=1.185
r52 17 24 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=5.25 $Y=1.185
+ $X2=5.59 $Y2=1.185
r53 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.16 $X2=5.25 $Y2=1.16
r54 13 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.39 $Y=1.025
+ $X2=5.39 $Y2=1.16
r55 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.39 $Y=1.025
+ $X2=5.39 $Y2=0.56
r56 9 32 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.37 $Y=1.295
+ $X2=5.37 $Y2=1.16
r57 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.37 $Y=1.295
+ $X2=5.37 $Y2=1.985
r58 5 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.97 $Y=1.025
+ $X2=4.97 $Y2=1.16
r59 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.97 $Y=1.025
+ $X2=4.97 $Y2=0.56
r60 1 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.95 $Y=1.295
+ $X2=4.95 $Y2=1.16
r61 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.95 $Y=1.295 $X2=4.95
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%A_51_297# 1 2 3 12 14 15 18 20 22 25
r37 22 24 4.392 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.1 $Y=1.725 $X2=2.1
+ $Y2=1.815
r38 21 25 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=1.605
+ $X2=1.22 $Y2=1.605
r39 20 22 6.82018 $w=2.4e-07 $l=1.75e-07 $layer=LI1_cond $X=1.975 $Y=1.605
+ $X2=2.1 $Y2=1.725
r40 20 21 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=1.605
+ $X2=1.305 $Y2=1.605
r41 16 25 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.22 $Y=1.725
+ $X2=1.22 $Y2=1.605
r42 16 18 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.22 $Y=1.725 $X2=1.22
+ $Y2=1.815
r43 14 25 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.605
+ $X2=1.22 $Y2=1.605
r44 14 15 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=1.135 $Y=1.605
+ $X2=0.465 $Y2=1.605
r45 10 15 7.27854 $w=2.4e-07 $l=2.42693e-07 $layer=LI1_cond $X=0.275 $Y=1.725
+ $X2=0.465 $Y2=1.605
r46 10 12 2.72947 $w=3.78e-07 $l=9e-08 $layer=LI1_cond $X=0.275 $Y=1.725
+ $X2=0.275 $Y2=1.815
r47 3 24 600 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=1.485 $X2=2.06 $Y2=1.815
r48 2 18 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.485 $X2=1.22 $Y2=1.815
r49 1 12 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.255
+ $Y=1.485 $X2=0.38 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%VPWR 1 2 3 14 18 22 25 26 27 29 42 43 46 49
r70 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r73 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r74 40 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 37 49 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.345 $Y=2.72
+ $X2=4.01 $Y2=2.72
r77 37 39 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.345 $Y=2.72
+ $X2=4.83 $Y2=2.72
r78 36 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r80 33 36 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 32 35 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=2.72
+ $X2=0.8 $Y2=2.72
r85 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.965 $Y=2.72
+ $X2=1.15 $Y2=2.72
r86 29 49 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=4.01 $Y2=2.72
r87 29 35 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.45 $Y2=2.72
r88 27 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 25 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=2.72
+ $X2=4.83 $Y2=2.72
r90 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=2.72
+ $X2=5.16 $Y2=2.72
r91 24 42 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.75 $Y2=2.72
r92 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.16 $Y2=2.72
r93 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=2.635
+ $X2=5.16 $Y2=2.72
r94 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=5.16 $Y=2.635
+ $X2=5.16 $Y2=2.02
r95 16 49 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.01 $Y=2.635
+ $X2=4.01 $Y2=2.72
r96 16 18 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.01 $Y=2.635
+ $X2=4.01 $Y2=2.02
r97 12 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=2.635 $X2=0.8
+ $Y2=2.72
r98 12 14 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.8 $Y=2.635
+ $X2=0.8 $Y2=2.02
r99 3 22 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.025
+ $Y=1.485 $X2=5.16 $Y2=2.02
r100 2 18 150 $w=1.7e-07 $l=7.35085e-07 $layer=licon1_PDIFF $count=4 $X=3.705
+ $Y=1.485 $X2=4.18 $Y2=2.02
r101 1 14 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=0.665
+ $Y=1.485 $X2=0.8 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%A_301_297# 1 2 9 11 12 15
r26 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3 $Y=2.295 $X2=3
+ $Y2=2.02
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.835 $Y=2.38
+ $X2=3 $Y2=2.295
r28 11 12 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.835 $Y=2.38
+ $X2=1.805 $Y2=2.38
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=2.295
+ $X2=1.805 $Y2=2.38
r30 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.64 $Y=2.295
+ $X2=1.64 $Y2=2.02
r31 2 15 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.865
+ $Y=1.485 $X2=3 $Y2=2.02
r32 1 9 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.505
+ $Y=1.485 $X2=1.64 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%Y 1 2 3 4 5 6 19 20 23 25 29 32 33 35 37 38
+ 39 40 41 42 43 59 71
c79 32 0 5.36204e-20 $X=3.42 $Y=1.605
r80 42 43 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=5.695 $Y=1.87
+ $X2=5.695 $Y2=2.21
r81 42 71 1.58461 $w=3.98e-07 $l=5.5e-08 $layer=LI1_cond $X=5.695 $Y=1.87
+ $X2=5.695 $Y2=1.815
r82 41 69 1.51637 $w=3.78e-07 $l=5e-08 $layer=LI1_cond $X=5.705 $Y=0.51
+ $X2=5.705 $Y2=0.56
r83 40 60 2.09911 $w=3.6e-07 $l=1.29615e-07 $layer=LI1_cond $X=4.715 $Y=1.605
+ $X2=4.735 $Y2=1.485
r84 40 60 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=4.735 $Y=1.465
+ $X2=4.735 $Y2=1.485
r85 39 40 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=4.735 $Y=1.19
+ $X2=4.735 $Y2=1.465
r86 38 59 2.8286 $w=3.6e-07 $l=1.15e-07 $layer=LI1_cond $X=4.735 $Y=0.77
+ $X2=4.735 $Y2=0.885
r87 38 39 8.96345 $w=3.58e-07 $l=2.8e-07 $layer=LI1_cond $X=4.735 $Y=0.91
+ $X2=4.735 $Y2=1.19
r88 38 59 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=4.735 $Y=0.91
+ $X2=4.735 $Y2=0.885
r89 36 69 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=5.705 $Y=0.655
+ $X2=5.705 $Y2=0.56
r90 35 38 21.0068 $w=3.48e-07 $l=6e-07 $layer=LI1_cond $X=5.515 $Y=0.77
+ $X2=4.915 $Y2=0.77
r91 35 36 7.36673 $w=2.3e-07 $l=2.40728e-07 $layer=LI1_cond $X=5.515 $Y=0.77
+ $X2=5.705 $Y2=0.655
r92 34 71 2.593 $w=3.98e-07 $l=9e-08 $layer=LI1_cond $X=5.695 $Y=1.725 $X2=5.695
+ $Y2=1.815
r93 33 40 19.2962 $w=3.68e-07 $l=5.8e-07 $layer=LI1_cond $X=5.495 $Y=1.605
+ $X2=4.915 $Y2=1.605
r94 33 34 7.38573 $w=2.4e-07 $l=2.52982e-07 $layer=LI1_cond $X=5.495 $Y=1.605
+ $X2=5.695 $Y2=1.725
r95 31 37 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.54 $Y=1.725 $X2=2.54
+ $Y2=1.815
r96 27 40 2.09911 $w=3.1e-07 $l=1.40712e-07 $layer=LI1_cond $X=4.67 $Y=1.725
+ $X2=4.715 $Y2=1.605
r97 27 29 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=4.67 $Y=1.725 $X2=4.67
+ $Y2=1.815
r98 26 32 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=1.605
+ $X2=3.42 $Y2=1.605
r99 25 40 4.12331 $w=2.4e-07 $l=2e-07 $layer=LI1_cond $X=4.515 $Y=1.605
+ $X2=4.715 $Y2=1.605
r100 25 26 48.4986 $w=2.38e-07 $l=1.01e-06 $layer=LI1_cond $X=4.515 $Y=1.605
+ $X2=3.505 $Y2=1.605
r101 21 32 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.42 $Y=1.725
+ $X2=3.42 $Y2=1.605
r102 21 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.42 $Y=1.725
+ $X2=3.42 $Y2=1.815
r103 20 31 6.82018 $w=2.4e-07 $l=1.75e-07 $layer=LI1_cond $X=2.665 $Y=1.605
+ $X2=2.54 $Y2=1.725
r104 19 32 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.605
+ $X2=3.42 $Y2=1.605
r105 19 20 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=3.335 $Y=1.605
+ $X2=2.665 $Y2=1.605
r106 6 71 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=5.445
+ $Y=1.485 $X2=5.58 $Y2=1.815
r107 5 29 300 $w=1.7e-07 $l=4.20179e-07 $layer=licon1_PDIFF $count=2 $X=4.465
+ $Y=1.485 $X2=4.67 $Y2=1.815
r108 4 23 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.815
r109 3 37 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.485 $X2=2.58 $Y2=1.815
r110 2 69 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=5.465
+ $Y=0.235 $X2=5.6 $Y2=0.56
r111 1 38 182 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.235 $X2=4.76 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%A_55_47# 1 2 3 4 5 16 18 21 23 26 28 33 36
+ 40 41 42
r68 36 38 6.05033 $w=3.98e-07 $l=2.1e-07 $layer=LI1_cond $X=0.285 $Y=0.56
+ $X2=0.285 $Y2=0.77
r69 31 42 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=0.77
+ $X2=3.36 $Y2=0.77
r70 31 33 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=3.445 $Y=0.77
+ $X2=4.2 $Y2=0.77
r71 28 42 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.36 $Y=0.655
+ $X2=3.36 $Y2=0.77
r72 28 30 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.36 $Y=0.655
+ $X2=3.36 $Y2=0.56
r73 27 41 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.77
+ $X2=2.08 $Y2=0.77
r74 26 42 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0.77
+ $X2=3.36 $Y2=0.77
r75 26 27 55.6179 $w=2.28e-07 $l=1.11e-06 $layer=LI1_cond $X=3.275 $Y=0.77
+ $X2=2.165 $Y2=0.77
r76 23 41 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.08 $Y=0.655
+ $X2=2.08 $Y2=0.77
r77 23 25 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.08 $Y=0.655
+ $X2=2.08 $Y2=0.56
r78 22 40 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=0.77
+ $X2=1.24 $Y2=0.77
r79 21 41 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0.77
+ $X2=2.08 $Y2=0.77
r80 21 22 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.995 $Y=0.77
+ $X2=1.325 $Y2=0.77
r81 18 40 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.24 $Y=0.655
+ $X2=1.24 $Y2=0.77
r82 18 20 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.24 $Y=0.655
+ $X2=1.24 $Y2=0.56
r83 17 38 3.97524 $w=2.3e-07 $l=2e-07 $layer=LI1_cond $X=0.485 $Y=0.77 $X2=0.285
+ $Y2=0.77
r84 16 40 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.77
+ $X2=1.24 $Y2=0.77
r85 16 17 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.155 $Y=0.77
+ $X2=0.485 $Y2=0.77
r86 5 33 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.235 $X2=4.2 $Y2=0.76
r87 4 30 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.36 $Y2=0.56
r88 3 25 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.235 $X2=2.08 $Y2=0.56
r89 2 20 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.235 $X2=1.24 $Y2=0.56
r90 1 36 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.235 $X2=0.4 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%VGND 1 2 3 14 18 20 22 37 38 41 44 49 55
r80 53 55 8.91182 $w=5.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=0.2
+ $X2=3.105 $Y2=0.2
r81 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r82 51 53 2.09838 $w=5.68e-07 $l=1e-07 $layer=LI1_cond $X=2.89 $Y=0.2 $X2=2.99
+ $Y2=0.2
r83 48 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r84 47 51 7.55418 $w=5.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.53 $Y=0.2 $X2=2.89
+ $Y2=0.2
r85 47 49 10.5905 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.53 $Y=0.2
+ $X2=2.335 $Y2=0.2
r86 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r87 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r88 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r89 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r90 35 38 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=5.75
+ $Y2=0
r91 35 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r92 34 37 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=5.75
+ $Y2=0
r93 34 55 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.105
+ $Y2=0
r94 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r95 31 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r96 31 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r97 30 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.335
+ $Y2=0
r98 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r99 28 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.66
+ $Y2=0
r100 28 30 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=2.07
+ $Y2=0
r101 26 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r102 26 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r103 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r104 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.82
+ $Y2=0
r105 23 25 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=1.15 $Y2=0
r106 22 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.66
+ $Y2=0
r107 22 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.15
+ $Y2=0
r108 20 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r109 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0
r110 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0.36
r111 12 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0
r112 12 14 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0.36
r113 3 51 91 $w=1.7e-07 $l=5.84166e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.235 $X2=2.89 $Y2=0.36
r114 2 18 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.525
+ $Y=0.235 $X2=1.66 $Y2=0.36
r115 1 14 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.235 $X2=0.82 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_2%A_729_47# 1 2 11
r17 8 11 70.1487 $w=2.28e-07 $l=1.4e-06 $layer=LI1_cond $X=3.78 $Y=0.37 $X2=5.18
+ $Y2=0.37
r18 2 11 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.18 $Y2=0.36
r19 1 8 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.235 $X2=3.78 $Y2=0.36
.ends


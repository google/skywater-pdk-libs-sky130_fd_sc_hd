* File: sky130_fd_sc_hd__a22o_2.spice.SKY130_FD_SC_HD__A22O_2.pxi
* Created: Thu Aug 27 14:02:34 2020
* 
x_PM_SKY130_FD_SC_HD__A22O_2%B2 N_B2_M1011_g N_B2_M1008_g B2 N_B2_c_62_n
+ N_B2_c_63_n N_B2_c_64_n PM_SKY130_FD_SC_HD__A22O_2%B2
x_PM_SKY130_FD_SC_HD__A22O_2%B1 N_B1_M1000_g N_B1_M1002_g B1 B1 N_B1_c_91_n
+ N_B1_c_92_n PM_SKY130_FD_SC_HD__A22O_2%B1
x_PM_SKY130_FD_SC_HD__A22O_2%A1 N_A1_M1001_g N_A1_M1010_g A1 A1 N_A1_c_131_n
+ N_A1_c_132_n PM_SKY130_FD_SC_HD__A22O_2%A1
x_PM_SKY130_FD_SC_HD__A22O_2%A2 N_A2_M1006_g N_A2_M1005_g A2 N_A2_c_167_n
+ N_A2_c_168_n N_A2_c_169_n PM_SKY130_FD_SC_HD__A22O_2%A2
x_PM_SKY130_FD_SC_HD__A22O_2%A_27_297# N_A_27_297#_M1000_d N_A_27_297#_M1001_s
+ N_A_27_297#_M1008_s N_A_27_297#_M1002_d N_A_27_297#_c_204_n
+ N_A_27_297#_M1007_g N_A_27_297#_M1003_g N_A_27_297#_c_205_n
+ N_A_27_297#_M1009_g N_A_27_297#_M1004_g N_A_27_297#_c_213_n
+ N_A_27_297#_c_214_n N_A_27_297#_c_215_n N_A_27_297#_c_216_n
+ N_A_27_297#_c_206_n N_A_27_297#_c_248_n N_A_27_297#_c_207_n
+ N_A_27_297#_c_208_n N_A_27_297#_c_209_n N_A_27_297#_c_218_n
+ N_A_27_297#_c_228_n N_A_27_297#_c_210_n PM_SKY130_FD_SC_HD__A22O_2%A_27_297#
x_PM_SKY130_FD_SC_HD__A22O_2%A_109_297# N_A_109_297#_M1008_d
+ N_A_109_297#_M1010_d N_A_109_297#_c_327_n N_A_109_297#_c_337_n
+ N_A_109_297#_c_342_p N_A_109_297#_c_329_n
+ PM_SKY130_FD_SC_HD__A22O_2%A_109_297#
x_PM_SKY130_FD_SC_HD__A22O_2%VPWR N_VPWR_M1010_s N_VPWR_M1005_d N_VPWR_M1004_d
+ N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n VPWR
+ N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n
+ N_VPWR_c_350_n PM_SKY130_FD_SC_HD__A22O_2%VPWR
x_PM_SKY130_FD_SC_HD__A22O_2%X N_X_M1007_d N_X_M1003_s N_X_c_407_n X X X
+ PM_SKY130_FD_SC_HD__A22O_2%X
x_PM_SKY130_FD_SC_HD__A22O_2%VGND N_VGND_M1011_s N_VGND_M1006_d N_VGND_M1009_s
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n
+ VGND N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n
+ PM_SKY130_FD_SC_HD__A22O_2%VGND
cc_1 VNB N_B2_c_62_n 0.0271486f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_2 VNB N_B2_c_63_n 0.0142681f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_3 VNB N_B2_c_64_n 0.0202523f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_4 VNB B1 0.00559744f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB B1 0.00553086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_B1_c_91_n 0.0241176f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_7 VNB N_B1_c_92_n 0.0190454f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_8 VNB A1 0.00265473f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_9 VNB A1 0.00206851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A1_c_131_n 0.0295813f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_11 VNB N_A1_c_132_n 0.0199376f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_12 VNB N_A2_c_167_n 0.0194031f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_13 VNB N_A2_c_168_n 0.00501659f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_14 VNB N_A2_c_169_n 0.0168697f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_15 VNB N_A_27_297#_c_204_n 0.0159674f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_16 VNB N_A_27_297#_c_205_n 0.0189287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_206_n 0.01475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_207_n 0.00359049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_208_n 0.00180044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_209_n 9.16142e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_297#_c_210_n 0.0497764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_350_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB X 6.52027e-19 $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_24 VNB N_VGND_c_426_n 0.0119341f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_25 VNB N_VGND_c_427_n 0.027794f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_26 VNB N_VGND_c_428_n 0.00224727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_429_n 0.0112093f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.175
cc_28 VNB N_VGND_c_430_n 0.0111495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_431_n 0.0419729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_432_n 0.0174317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_433_n 0.00507731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_434_n 0.203659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_B2_M1008_g 0.0255346f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_34 VPB N_B2_c_62_n 0.00476167f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_35 VPB N_B1_M1002_g 0.0255531f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB N_B1_c_91_n 0.00488357f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_37 VPB N_A1_M1010_g 0.0251751f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_38 VPB N_A1_c_131_n 0.00672831f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_39 VPB N_A2_M1005_g 0.0198907f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_40 VPB N_A2_c_167_n 0.00407683f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_41 VPB N_A_27_297#_M1003_g 0.0180715f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.175
cc_42 VPB N_A_27_297#_M1004_g 0.0242693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_297#_c_213_n 0.00746643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_297#_c_214_n 0.025859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_297#_c_215_n 0.0320347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_297#_c_216_n 0.00971545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_297#_c_209_n 0.00132789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_297#_c_218_n 0.00256417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_297#_c_210_n 0.00820056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_109_297#_c_327_n 0.00819467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_351_n 0.0059122f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_52 VPB N_VPWR_c_352_n 0.00210405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_353_n 0.0111834f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.175
cc_54 VPB N_VPWR_c_354_n 0.00833811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_355_n 0.0364036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_356_n 0.0146389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_357_n 0.0154264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_358_n 0.0054066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_359_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_350_n 0.0483412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 9.51109e-19 $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_62 N_B2_M1008_g N_B1_M1002_g 0.0437171f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_63 N_B2_c_62_n B1 3.38478e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B2_c_62_n B1 9.18012e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_65 N_B2_c_63_n B1 0.0162583f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_66 N_B2_c_62_n N_B1_c_91_n 0.0338406f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B2_c_63_n N_B1_c_91_n 7.15179e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B2_c_64_n N_B1_c_92_n 0.0338406f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B2_M1008_g N_A_27_297#_c_213_n 7.12665e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_70 N_B2_M1008_g N_A_27_297#_c_214_n 0.00966083f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_71 N_B2_M1008_g N_A_27_297#_c_215_n 0.0088291f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_72 N_B2_c_63_n N_A_27_297#_c_215_n 0.0100322f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B2_M1008_g N_A_27_297#_c_216_n 0.00149869f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_74 N_B2_c_62_n N_A_27_297#_c_216_n 0.00295538f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B2_c_63_n N_A_27_297#_c_216_n 0.0263428f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B2_c_64_n N_A_27_297#_c_206_n 7.24737e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_77 N_B2_M1008_g N_A_27_297#_c_228_n 0.00819053f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B2_M1008_g N_VPWR_c_355_n 0.00357835f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B2_M1008_g N_VPWR_c_350_n 0.00620759f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_80 N_B2_c_62_n N_VGND_c_427_n 0.00275758f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B2_c_63_n N_VGND_c_427_n 0.0270634f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B2_c_64_n N_VGND_c_427_n 0.0264669f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B2_c_64_n N_VGND_c_434_n 7.20442e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_84 B1 A1 0.0223083f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_85 N_B1_c_91_n A1 2.2062e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_86 B1 A1 0.0129839f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B1_c_91_n A1 6.20311e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_88 B1 N_A1_c_131_n 2.97885e-19 $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_89 B1 N_A1_c_131_n 8.83743e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B1_c_91_n N_A1_c_131_n 0.00758269f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_91 B1 N_A_27_297#_M1000_d 0.00558122f $X=1.07 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_92 N_B1_M1002_g N_A_27_297#_c_214_n 0.00147562f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 N_B1_M1002_g N_A_27_297#_c_215_n 0.0124265f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_94 B1 N_A_27_297#_c_215_n 0.0346626f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B1_c_91_n N_A_27_297#_c_215_n 0.00345472f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_96 B1 N_A_27_297#_c_206_n 0.0168276f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_97 B1 N_A_27_297#_c_206_n 0.00462247f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B1_c_91_n N_A_27_297#_c_206_n 0.0018138f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B1_c_92_n N_A_27_297#_c_206_n 0.00810253f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_A_27_297#_c_218_n 0.00185095f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B1_M1002_g N_A_27_297#_c_228_n 0.00681763f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_M1002_g N_A_109_297#_c_327_n 0.0131306f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_M1002_g N_A_109_297#_c_329_n 0.00406201f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_B1_M1002_g N_VPWR_c_351_n 0.00237859f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B1_M1002_g N_VPWR_c_355_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B1_M1002_g N_VPWR_c_350_n 0.00657948f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_107 B1 N_VGND_c_427_n 0.00606397f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_108 N_B1_c_92_n N_VGND_c_427_n 0.00412676f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B1_c_92_n N_VGND_c_431_n 0.0042613f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B1_c_92_n N_VGND_c_434_n 0.0081372f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A1_M1010_g N_A2_M1005_g 0.0229849f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_112 A1 N_A2_c_167_n 3.78337e-19 $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_113 A1 N_A2_c_167_n 2.41928e-19 $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_114 N_A1_c_131_n N_A2_c_167_n 0.0216734f $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_115 A1 N_A2_c_168_n 0.016083f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A1_c_131_n N_A2_c_168_n 0.00131294f $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A1_c_132_n N_A2_c_169_n 0.0295033f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_118 A1 N_A_27_297#_M1001_s 0.00586103f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_119 N_A1_M1010_g N_A_27_297#_c_215_n 0.0147495f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_120 A1 N_A_27_297#_c_215_n 0.02377f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A1_c_131_n N_A_27_297#_c_215_n 0.00505271f $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_122 A1 N_A_27_297#_c_206_n 0.0143007f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_123 A1 N_A_27_297#_c_206_n 0.00271225f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A1_c_131_n N_A_27_297#_c_206_n 6.23547e-19 $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A1_c_132_n N_A_27_297#_c_206_n 0.01264f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A1_c_132_n N_A_27_297#_c_248_n 0.0045799f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_127 A1 N_A_27_297#_c_208_n 0.00624318f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_128 N_A1_c_132_n N_A_27_297#_c_208_n 0.00172045f $X=1.722 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_A1_M1010_g N_A_109_297#_c_327_n 0.0141907f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A1_M1010_g N_VPWR_c_351_n 0.00990552f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_M1010_g N_VPWR_c_356_n 0.00273041f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A1_M1010_g N_VPWR_c_350_n 0.00348631f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A1_c_132_n N_VGND_c_428_n 0.00127092f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A1_c_132_n N_VGND_c_431_n 0.00357877f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A1_c_132_n N_VGND_c_434_n 0.00672549f $X=1.722 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A2_c_169_n N_A_27_297#_c_204_n 0.0203582f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A2_M1005_g N_A_27_297#_M1003_g 0.0223671f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A2_M1005_g N_A_27_297#_c_215_n 0.015518f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A2_c_167_n N_A_27_297#_c_215_n 0.0028355f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A2_c_168_n N_A_27_297#_c_215_n 0.0280408f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_c_169_n N_A_27_297#_c_206_n 0.00222116f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_169_n N_A_27_297#_c_248_n 0.00442179f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A2_c_167_n N_A_27_297#_c_207_n 0.00221567f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_c_168_n N_A_27_297#_c_207_n 0.0190591f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A2_c_169_n N_A_27_297#_c_207_n 0.0118724f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A2_c_167_n N_A_27_297#_c_208_n 7.67796e-19 $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_c_168_n N_A_27_297#_c_208_n 0.0113712f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_M1005_g N_A_27_297#_c_209_n 0.00243411f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A2_c_167_n N_A_27_297#_c_209_n 0.0010489f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_168_n N_A_27_297#_c_209_n 0.0121929f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_c_169_n N_A_27_297#_c_209_n 0.00167934f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_167_n N_A_27_297#_c_210_n 0.0225009f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A2_c_168_n N_A_27_297#_c_210_n 0.0013901f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_M1005_g N_VPWR_c_351_n 5.43585e-19 $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A2_M1005_g N_VPWR_c_352_n 0.00166715f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A2_M1005_g N_VPWR_c_356_n 0.00585385f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A2_M1005_g N_VPWR_c_350_n 0.0107512f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A2_c_169_n N_VGND_c_428_n 0.0091562f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_169_n N_VGND_c_431_n 0.00350562f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_169_n N_VGND_c_434_n 0.00436f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_27_297#_c_215_n N_A_109_297#_M1008_d 0.00166235f $X=2.645 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_162 N_A_27_297#_c_228_n N_A_109_297#_M1008_d 0.00312752f $X=0.935 $Y=2.36
+ $X2=-0.19 $Y2=-0.24
cc_163 N_A_27_297#_c_215_n N_A_109_297#_M1010_d 0.00229659f $X=2.645 $Y=1.54
+ $X2=0 $Y2=0
cc_164 N_A_27_297#_M1002_d N_A_109_297#_c_327_n 0.00554761f $X=0.965 $Y=1.485
+ $X2=0 $Y2=0
cc_165 N_A_27_297#_c_218_n N_A_109_297#_c_327_n 0.0157397f $X=1.1 $Y=2.34 $X2=0
+ $Y2=0
cc_166 N_A_27_297#_c_228_n N_A_109_297#_c_327_n 0.0048504f $X=0.935 $Y=2.36
+ $X2=0 $Y2=0
cc_167 N_A_27_297#_c_215_n N_A_109_297#_c_337_n 0.0160896f $X=2.645 $Y=1.54
+ $X2=0 $Y2=0
cc_168 N_A_27_297#_c_215_n N_A_109_297#_c_329_n 0.0851707f $X=2.645 $Y=1.54
+ $X2=0 $Y2=0
cc_169 N_A_27_297#_c_228_n N_A_109_297#_c_329_n 0.0118327f $X=0.935 $Y=2.36
+ $X2=0 $Y2=0
cc_170 N_A_27_297#_c_215_n N_VPWR_M1010_s 0.00277869f $X=2.645 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_27_297#_c_215_n N_VPWR_M1005_d 0.00253908f $X=2.645 $Y=1.54 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_c_218_n N_VPWR_c_351_n 0.0169231f $X=1.1 $Y=2.34 $X2=0 $Y2=0
cc_173 N_A_27_297#_M1003_g N_VPWR_c_352_n 0.0108609f $X=2.775 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_M1004_g N_VPWR_c_352_n 4.83856e-19 $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_c_215_n N_VPWR_c_352_n 0.0140564f $X=2.645 $Y=1.54 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_M1004_g N_VPWR_c_354_n 0.00673095f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_c_213_n N_VPWR_c_355_n 0.021178f $X=0.26 $Y=2.295 $X2=0 $Y2=0
cc_178 N_A_27_297#_c_228_n N_VPWR_c_355_n 0.0481435f $X=0.935 $Y=2.36 $X2=0
+ $Y2=0
cc_179 N_A_27_297#_M1003_g N_VPWR_c_357_n 0.0046653f $X=2.775 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_27_297#_M1004_g N_VPWR_c_357_n 0.00526178f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_27_297#_M1008_s N_VPWR_c_350_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_A_27_297#_M1002_d N_VPWR_c_350_n 0.00209344f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_M1003_g N_VPWR_c_350_n 0.00789179f $X=2.775 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_27_297#_M1004_g N_VPWR_c_350_n 0.0101251f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_27_297#_c_213_n N_VPWR_c_350_n 0.0124992f $X=0.26 $Y=2.295 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_c_228_n N_VPWR_c_350_n 0.030037f $X=0.935 $Y=2.36 $X2=0 $Y2=0
cc_187 N_A_27_297#_c_205_n N_X_c_407_n 0.0042988f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_27_297#_c_210_n N_X_c_407_n 0.00170475f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_204_n X 0.00460679f $X=2.775 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_27_297#_M1003_g X 0.00506951f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_27_297#_c_205_n X 0.0078344f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_27_297#_M1004_g X 0.020111f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_27_297#_c_215_n X 0.0131028f $X=2.645 $Y=1.54 $X2=0 $Y2=0
cc_194 N_A_27_297#_c_207_n X 0.0130895f $X=2.645 $Y=0.82 $X2=0 $Y2=0
cc_195 N_A_27_297#_c_209_n X 0.0371162f $X=2.73 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_210_n X 0.0255973f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_207_n N_VGND_M1006_d 0.00208738f $X=2.645 $Y=0.82 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_206_n N_VGND_c_427_n 0.0137634f $X=1.975 $Y=0.38 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_204_n N_VGND_c_428_n 0.00174093f $X=2.775 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_c_206_n N_VGND_c_428_n 0.0175383f $X=1.975 $Y=0.38 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_c_248_n N_VGND_c_428_n 0.00373345f $X=2.06 $Y=0.735 $X2=0
+ $Y2=0
cc_202 N_A_27_297#_c_207_n N_VGND_c_428_n 0.0178614f $X=2.645 $Y=0.82 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_205_n N_VGND_c_430_n 0.00715217f $X=3.195 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_206_n N_VGND_c_431_n 0.0817349f $X=1.975 $Y=0.38 $X2=0
+ $Y2=0
cc_205 N_A_27_297#_c_207_n N_VGND_c_431_n 0.00245781f $X=2.645 $Y=0.82 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_204_n N_VGND_c_432_n 0.00473211f $X=2.775 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_27_297#_c_205_n N_VGND_c_432_n 0.00524716f $X=3.195 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_27_297#_c_207_n N_VGND_c_432_n 0.00176795f $X=2.645 $Y=0.82 $X2=0
+ $Y2=0
cc_209 N_A_27_297#_M1000_d N_VGND_c_434_n 0.00209344f $X=0.925 $Y=0.235 $X2=0
+ $Y2=0
cc_210 N_A_27_297#_M1001_s N_VGND_c_434_n 0.00209344f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_211 N_A_27_297#_c_204_n N_VGND_c_434_n 0.00701835f $X=2.775 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_27_297#_c_205_n N_VGND_c_434_n 0.0100791f $X=3.195 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_206_n N_VGND_c_434_n 0.048613f $X=1.975 $Y=0.38 $X2=0 $Y2=0
cc_214 N_A_27_297#_c_207_n N_VGND_c_434_n 0.00917387f $X=2.645 $Y=0.82 $X2=0
+ $Y2=0
cc_215 N_A_27_297#_c_206_n A_381_47# 0.00539739f $X=1.975 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_216 N_A_27_297#_c_248_n A_381_47# 0.00521283f $X=2.06 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_27_297#_c_207_n A_381_47# 6.20362e-19 $X=2.645 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_27_297#_c_208_n A_381_47# 0.00216212f $X=2.145 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_109_297#_c_327_n N_VPWR_M1010_s 0.00520183f $X=1.98 $Y=1.915
+ $X2=-0.19 $Y2=1.305
cc_220 N_A_109_297#_c_327_n N_VPWR_c_351_n 0.0221078f $X=1.98 $Y=1.915 $X2=0
+ $Y2=0
cc_221 N_A_109_297#_c_342_p N_VPWR_c_351_n 0.0191044f $X=2.065 $Y=2.3 $X2=0
+ $Y2=0
cc_222 N_A_109_297#_c_327_n N_VPWR_c_355_n 0.00320421f $X=1.98 $Y=1.915 $X2=0
+ $Y2=0
cc_223 N_A_109_297#_c_327_n N_VPWR_c_356_n 0.00217595f $X=1.98 $Y=1.915 $X2=0
+ $Y2=0
cc_224 N_A_109_297#_c_342_p N_VPWR_c_356_n 0.0156476f $X=2.065 $Y=2.3 $X2=0
+ $Y2=0
cc_225 N_A_109_297#_M1008_d N_VPWR_c_350_n 0.00216833f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_226 N_A_109_297#_M1010_d N_VPWR_c_350_n 0.00314787f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_227 N_A_109_297#_c_327_n N_VPWR_c_350_n 0.0120275f $X=1.98 $Y=1.915 $X2=0
+ $Y2=0
cc_228 N_A_109_297#_c_342_p N_VPWR_c_350_n 0.00954719f $X=2.065 $Y=2.3 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_350_n N_X_M1003_s 0.0038878f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_354_n X 0.0731451f $X=3.415 $Y=1.63 $X2=0 $Y2=0
cc_231 N_VPWR_c_357_n X 0.0158317f $X=3.33 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_350_n X 0.00968523f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_c_354_n N_VGND_c_430_n 0.00786978f $X=3.415 $Y=1.63 $X2=0 $Y2=0
cc_234 N_X_c_407_n N_VGND_c_430_n 0.0238996f $X=3.075 $Y=0.42 $X2=0 $Y2=0
cc_235 X N_VGND_c_430_n 0.0282127f $X=2.93 $Y=1.785 $X2=0 $Y2=0
cc_236 N_X_c_407_n N_VGND_c_432_n 0.0151483f $X=3.075 $Y=0.42 $X2=0 $Y2=0
cc_237 N_X_M1007_d N_VGND_c_434_n 0.00385329f $X=2.85 $Y=0.235 $X2=0 $Y2=0
cc_238 N_X_c_407_n N_VGND_c_434_n 0.00957453f $X=3.075 $Y=0.42 $X2=0 $Y2=0
cc_239 N_VGND_c_434_n A_109_47# 0.00978874f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_240 N_VGND_c_434_n A_381_47# 0.00311078f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

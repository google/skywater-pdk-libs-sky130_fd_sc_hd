* File: sky130_fd_sc_hd__a21boi_4.spice.SKY130_FD_SC_HD__A21BOI_4.pxi
* Created: Thu Aug 27 14:00:47 2020
* 
x_PM_SKY130_FD_SC_HD__A21BOI_4%B1_N N_B1_N_M1025_g N_B1_N_M1016_g B1_N
+ N_B1_N_c_102_n N_B1_N_c_103_n PM_SKY130_FD_SC_HD__A21BOI_4%B1_N
x_PM_SKY130_FD_SC_HD__A21BOI_4%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1025_s
+ N_A_27_47#_c_135_n N_A_27_47#_M1001_g N_A_27_47#_M1000_g N_A_27_47#_c_136_n
+ N_A_27_47#_M1009_g N_A_27_47#_M1005_g N_A_27_47#_c_137_n N_A_27_47#_M1018_g
+ N_A_27_47#_M1010_g N_A_27_47#_c_138_n N_A_27_47#_M1019_g N_A_27_47#_M1020_g
+ N_A_27_47#_c_139_n N_A_27_47#_c_140_n N_A_27_47#_c_159_n N_A_27_47#_c_148_n
+ N_A_27_47#_c_141_n N_A_27_47#_c_149_n N_A_27_47#_c_150_n N_A_27_47#_c_151_n
+ N_A_27_47#_c_142_n N_A_27_47#_c_143_n PM_SKY130_FD_SC_HD__A21BOI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__A21BOI_4%A2 N_A2_M1002_g N_A2_M1007_g N_A2_c_252_n
+ N_A2_M1014_g N_A2_M1004_g N_A2_c_253_n N_A2_M1015_g N_A2_M1013_g N_A2_c_254_n
+ N_A2_M1024_g N_A2_M1017_g N_A2_c_255_n N_A2_c_256_n N_A2_c_275_n N_A2_c_257_n
+ N_A2_c_268_n A2 N_A2_c_258_n N_A2_c_259_n N_A2_c_260_n
+ PM_SKY130_FD_SC_HD__A21BOI_4%A2
x_PM_SKY130_FD_SC_HD__A21BOI_4%A1 N_A1_c_378_n N_A1_M1006_g N_A1_M1003_g
+ N_A1_c_380_n N_A1_M1011_g N_A1_M1008_g N_A1_c_382_n N_A1_M1021_g N_A1_M1012_g
+ N_A1_c_384_n N_A1_M1022_g N_A1_M1023_g A1 PM_SKY130_FD_SC_HD__A21BOI_4%A1
x_PM_SKY130_FD_SC_HD__A21BOI_4%VPWR N_VPWR_M1025_d N_VPWR_M1002_d N_VPWR_M1008_d
+ N_VPWR_M1023_d N_VPWR_M1013_d N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n
+ N_VPWR_c_459_n VPWR N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n
+ N_VPWR_c_450_n N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_466_n
+ PM_SKY130_FD_SC_HD__A21BOI_4%VPWR
x_PM_SKY130_FD_SC_HD__A21BOI_4%A_223_297# N_A_223_297#_M1000_d
+ N_A_223_297#_M1005_d N_A_223_297#_M1020_d N_A_223_297#_M1003_s
+ N_A_223_297#_M1012_s N_A_223_297#_M1004_s N_A_223_297#_M1017_s
+ N_A_223_297#_c_610_n N_A_223_297#_c_569_n N_A_223_297#_c_573_n
+ N_A_223_297#_c_584_n N_A_223_297#_c_575_n N_A_223_297#_c_626_n
+ N_A_223_297#_c_588_n N_A_223_297#_c_633_n N_A_223_297#_c_590_n
+ N_A_223_297#_c_567_n N_A_223_297#_c_568_n N_A_223_297#_c_596_n
+ N_A_223_297#_c_597_n PM_SKY130_FD_SC_HD__A21BOI_4%A_223_297#
x_PM_SKY130_FD_SC_HD__A21BOI_4%Y N_Y_M1001_s N_Y_M1018_s N_Y_M1006_s N_Y_M1021_s
+ N_Y_M1000_s N_Y_M1010_s N_Y_c_653_n N_Y_c_709_p N_Y_c_657_n N_Y_c_648_n
+ N_Y_c_649_n N_Y_c_650_n N_Y_c_664_n N_Y_c_666_n N_Y_c_668_n N_Y_c_651_n Y
+ N_Y_c_669_n Y PM_SKY130_FD_SC_HD__A21BOI_4%Y
x_PM_SKY130_FD_SC_HD__A21BOI_4%VGND N_VGND_M1016_d N_VGND_M1009_d N_VGND_M1019_d
+ N_VGND_M1014_d N_VGND_M1024_d N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n
+ N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n N_VGND_c_734_n
+ N_VGND_c_735_n N_VGND_c_736_n VGND N_VGND_c_737_n N_VGND_c_738_n
+ N_VGND_c_739_n N_VGND_c_740_n PM_SKY130_FD_SC_HD__A21BOI_4%VGND
x_PM_SKY130_FD_SC_HD__A21BOI_4%A_658_47# N_A_658_47#_M1007_s N_A_658_47#_M1011_d
+ N_A_658_47#_M1022_d N_A_658_47#_M1015_s N_A_658_47#_c_830_n
+ N_A_658_47#_c_831_n N_A_658_47#_c_832_n N_A_658_47#_c_828_n
+ N_A_658_47#_c_829_n N_A_658_47#_c_843_n PM_SKY130_FD_SC_HD__A21BOI_4%A_658_47#
cc_1 VNB B1_N 0.013842f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_2 VNB N_B1_N_c_102_n 0.0297894f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.16
cc_3 VNB N_B1_N_c_103_n 0.0231202f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=0.995
cc_4 VNB N_A_27_47#_c_135_n 0.0164085f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=0.56
cc_5 VNB N_A_27_47#_c_136_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.325
cc_6 VNB N_A_27_47#_c_137_n 0.0160015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_138_n 0.0183771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_139_n 0.00937296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_140_n 0.0144029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_141_n 0.00154426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_142_n 0.0023212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_143_n 0.0814771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_252_n 0.016129f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_14 VNB N_A2_c_253_n 0.0159999f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.16
cc_15 VNB N_A2_c_254_n 0.0219817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_255_n 0.00159939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A2_c_256_n 0.0238251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_257_n 0.00237446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_258_n 0.0187412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_259_n 0.0615981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_260_n 0.00961897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_378_n 0.0160486f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.325
cc_23 VNB N_A1_M1003_g 3.5465e-19 $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=0.56
cc_24 VNB N_A1_c_380_n 0.0158334f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_25 VNB N_A1_M1008_g 3.82449e-19 $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=0.995
cc_26 VNB N_A1_c_382_n 0.0158329f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.16
cc_27 VNB N_A1_M1012_g 3.82449e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A1_c_384_n 0.0879521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A1_M1023_g 4.33197e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB A1 0.00170867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_450_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_648_n 0.00423887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_649_n 4.56702e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_650_n 0.00972875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_651_n 0.00656144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_727_n 3.08929e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_728_n 0.00421457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_729_n 0.0359713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_730_n 0.0297204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_731_n 0.0125281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_732_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_733_n 0.0550106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_734_n 0.00362081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_735_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_736_n 0.00499771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_737_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_738_n 0.341178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_739_n 0.0114607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_740_n 0.0143321f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_658_47#_c_828_n 0.00452179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_658_47#_c_829_n 0.003364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VPB N_B1_N_M1025_g 0.0275226f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_53 VPB B1_N 0.0146528f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_54 VPB N_B1_N_c_102_n 0.0052048f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_55 VPB N_A_27_47#_M1000_g 0.0227058f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_56 VPB N_A_27_47#_M1005_g 0.0185953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_M1010_g 0.0185649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_M1020_g 0.0177211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_148_n 0.00461041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_149_n 0.00762873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_150_n 0.0126004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_151_n 0.0282991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_142_n 0.00503429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_143_n 0.0211271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A2_M1002_g 0.0176318f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_66 VPB N_A2_M1004_g 0.0171445f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=0.995
cc_67 VPB N_A2_M1013_g 0.017124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A2_M1017_g 0.0222503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A2_c_255_n 0.00276621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A2_c_256_n 0.00631169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A2_c_257_n 0.00197902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A2_c_268_n 0.0136346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A2_c_259_n 0.0123305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A2_c_260_n 0.00733094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A1_M1003_g 0.0196283f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=0.56
cc_76 VPB N_A1_M1008_g 0.0193016f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=0.995
cc_77 VPB N_A1_M1012_g 0.0193016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A1_M1023_g 0.0196386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB A1 0.00799673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_451_n 0.00871222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_452_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_453_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_454_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_455_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_456_n 0.0113516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_457_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_458_n 0.0113994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_459_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_460_n 0.0546787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_461_n 0.0122674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_462_n 0.0209462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_450_n 0.0607309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_464_n 0.023139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_465_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_466_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_223_297#_c_567_n 0.0112688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_223_297#_c_568_n 0.0137952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_648_n 0.00268101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 B1_N N_A_27_47#_M1025_s 0.00289727f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_100 N_B1_N_c_103_n N_A_27_47#_c_135_n 0.0148378f $X=0.565 $Y=0.995 $X2=0
+ $Y2=0
cc_101 B1_N N_A_27_47#_c_139_n 0.0185209f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_102 N_B1_N_c_102_n N_A_27_47#_c_139_n 4.15056e-19 $X=0.565 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_B1_N_c_103_n N_A_27_47#_c_140_n 0.0111225f $X=0.565 $Y=0.995 $X2=0
+ $Y2=0
cc_104 B1_N N_A_27_47#_c_159_n 0.0114513f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_105 N_B1_N_c_102_n N_A_27_47#_c_159_n 0.00126544f $X=0.565 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_B1_N_c_103_n N_A_27_47#_c_159_n 0.0160313f $X=0.565 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_B1_N_M1025_g N_A_27_47#_c_148_n 0.0120787f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_108 B1_N N_A_27_47#_c_148_n 0.0106319f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_109 N_B1_N_c_102_n N_A_27_47#_c_148_n 0.00175404f $X=0.565 $Y=1.16 $X2=0
+ $Y2=0
cc_110 B1_N N_A_27_47#_c_141_n 0.00295838f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_111 N_B1_N_c_103_n N_A_27_47#_c_141_n 0.00538638f $X=0.565 $Y=0.995 $X2=0
+ $Y2=0
cc_112 N_B1_N_M1025_g N_A_27_47#_c_149_n 0.00697957f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_113 B1_N N_A_27_47#_c_149_n 0.0218242f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_114 N_B1_N_M1025_g N_A_27_47#_c_151_n 0.0118608f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_115 B1_N N_A_27_47#_c_151_n 0.0223603f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_116 B1_N N_A_27_47#_c_142_n 0.0268954f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_117 N_B1_N_c_102_n N_A_27_47#_c_142_n 0.00257049f $X=0.565 $Y=1.16 $X2=0
+ $Y2=0
cc_118 B1_N N_A_27_47#_c_143_n 2.67713e-19 $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_119 N_B1_N_c_102_n N_A_27_47#_c_143_n 0.0148378f $X=0.565 $Y=1.16 $X2=0 $Y2=0
cc_120 B1_N N_VPWR_M1025_d 0.00157293f $X=0.145 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_121 N_B1_N_M1025_g N_VPWR_c_451_n 0.00454665f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_N_M1025_g N_VPWR_c_450_n 0.00802324f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_N_M1025_g N_VPWR_c_464_n 0.00424868f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_N_M1025_g N_A_223_297#_c_569_n 0.00425622f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_B1_N_c_103_n N_VGND_c_730_n 0.00872204f $X=0.565 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_N_c_103_n N_VGND_c_738_n 0.00702962f $X=0.565 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1020_g N_A2_M1002_g 0.0357673f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1020_g N_A2_c_255_n 5.08272e-19 $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_143_n N_A2_c_255_n 2.96609e-19 $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_143_n N_A2_c_256_n 0.0207157f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_27_47#_M1020_g N_A2_c_275_n 8.40721e-19 $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_138_n N_A2_c_258_n 0.00899944f $X=2.445 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_148_n N_VPWR_M1025_d 0.00874894f $X=0.82 $Y=1.895 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_27_47#_c_149_n N_VPWR_M1025_d 0.00356612f $X=0.905 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_27_47#_M1000_g N_VPWR_c_451_n 0.00228791f $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_148_n N_VPWR_c_451_n 0.0201051f $X=0.82 $Y=1.895 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1020_g N_VPWR_c_452_n 0.00101195f $X=2.745 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_M1000_g N_VPWR_c_460_n 0.00357877f $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_M1005_g N_VPWR_c_460_n 0.00357842f $X=1.885 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1010_g N_VPWR_c_460_n 0.00357668f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_M1020_g N_VPWR_c_460_n 0.00357668f $X=2.745 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_148_n N_VPWR_c_460_n 0.0018132f $X=0.82 $Y=1.895 $X2=0 $Y2=0
cc_143 N_A_27_47#_M1025_s N_VPWR_c_450_n 0.00213418f $X=0.165 $Y=1.485 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_M1000_g N_VPWR_c_450_n 0.00657863f $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_M1005_g N_VPWR_c_450_n 0.00527891f $X=1.885 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_M1010_g N_VPWR_c_450_n 0.00527877f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_M1020_g N_VPWR_c_450_n 0.00537502f $X=2.745 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_148_n N_VPWR_c_450_n 0.00796907f $X=0.82 $Y=1.895 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_151_n N_VPWR_c_450_n 0.0124497f $X=0.29 $Y=2 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_148_n N_VPWR_c_464_n 0.00208303f $X=0.82 $Y=1.895 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_c_151_n N_VPWR_c_464_n 0.0210489f $X=0.29 $Y=2 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_148_n N_A_223_297#_c_569_n 0.0176158f $X=0.82 $Y=1.895 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_150_n N_A_223_297#_c_569_n 0.00759562f $X=2.235 $Y=1.16
+ $X2=0 $Y2=0
cc_154 N_A_27_47#_c_143_n N_A_223_297#_c_569_n 0.00113237f $X=2.745 $Y=1.16
+ $X2=0 $Y2=0
cc_155 N_A_27_47#_M1000_g N_A_223_297#_c_573_n 0.0146159f $X=1.455 $Y=1.985
+ $X2=0 $Y2=0
cc_156 N_A_27_47#_M1005_g N_A_223_297#_c_573_n 0.00863478f $X=1.885 $Y=1.985
+ $X2=0 $Y2=0
cc_157 N_A_27_47#_M1005_g N_A_223_297#_c_575_n 0.00128732f $X=1.885 $Y=1.985
+ $X2=0 $Y2=0
cc_158 N_A_27_47#_M1010_g N_A_223_297#_c_575_n 0.0100298f $X=2.315 $Y=1.985
+ $X2=0 $Y2=0
cc_159 N_A_27_47#_M1020_g N_A_223_297#_c_575_n 0.0166494f $X=2.745 $Y=1.985
+ $X2=0 $Y2=0
cc_160 N_A_27_47#_c_136_n N_Y_c_653_n 0.0122034f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_137_n N_Y_c_653_n 0.0115395f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_150_n N_Y_c_653_n 0.0420392f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_143_n N_Y_c_653_n 0.00278364f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_138_n N_Y_c_657_n 0.0146315f $X=2.445 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_150_n N_Y_c_657_n 0.00377018f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_27_47#_M1010_g N_Y_c_648_n 0.00550767f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_138_n N_Y_c_648_n 0.00302208f $X=2.445 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_27_47#_M1020_g N_Y_c_648_n 0.0190837f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_150_n N_Y_c_648_n 0.0245207f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_143_n N_Y_c_648_n 0.0197399f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_150_n N_Y_c_664_n 0.0141276f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_143_n N_Y_c_664_n 0.0025826f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_150_n N_Y_c_666_n 0.0144259f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_143_n N_Y_c_666_n 0.00284454f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_138_n N_Y_c_668_n 4.93918e-19 $X=2.445 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1005_g N_Y_c_669_n 0.0170373f $X=1.885 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1010_g N_Y_c_669_n 0.0174728f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_150_n N_Y_c_669_n 0.0457478f $X=2.235 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_143_n N_Y_c_669_n 0.00491429f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_159_n N_VGND_M1016_d 0.00536666f $X=0.82 $Y=0.705 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_27_47#_c_141_n N_VGND_M1016_d 0.00116546f $X=0.962 $Y=1.035 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_27_47#_c_135_n N_VGND_c_727_n 7.79461e-19 $X=1.155 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_136_n N_VGND_c_727_n 0.00709932f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_137_n N_VGND_c_727_n 0.0062525f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_138_n N_VGND_c_727_n 4.98169e-19 $X=2.445 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_135_n N_VGND_c_730_n 0.00728604f $X=1.155 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_136_n N_VGND_c_730_n 7.82447e-19 $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_140_n N_VGND_c_730_n 0.0244675f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_159_n N_VGND_c_730_n 0.0278519f $X=0.82 $Y=0.705 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_135_n N_VGND_c_731_n 0.00487821f $X=1.155 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_136_n N_VGND_c_731_n 0.00351072f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1016_s N_VGND_c_738_n 0.00371687f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_135_n N_VGND_c_738_n 0.00830224f $X=1.155 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_136_n N_VGND_c_738_n 0.00411677f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_137_n N_VGND_c_738_n 0.0040731f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_138_n N_VGND_c_738_n 0.00421891f $X=2.445 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_140_n N_VGND_c_738_n 0.0135138f $X=0.28 $Y=0.36 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_159_n N_VGND_c_738_n 0.00910161f $X=0.82 $Y=0.705 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_137_n N_VGND_c_739_n 0.00351072f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_138_n N_VGND_c_739_n 0.00360664f $X=2.445 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_137_n N_VGND_c_740_n 5.33636e-19 $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_138_n N_VGND_c_740_n 0.00802208f $X=2.445 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_143_n N_VGND_c_740_n 9.94449e-19 $X=2.745 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_A2_c_258_n N_A1_c_378_n 0.0245688f $X=3.195 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_205 N_A2_M1002_g N_A1_M1003_g 0.0422562f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A2_c_255_n N_A1_M1003_g 0.00392475f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A2_c_268_n N_A1_M1003_g 0.0125777f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_208 N_A2_c_268_n N_A1_M1008_g 0.0125621f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_209 N_A2_c_268_n N_A1_M1012_g 0.0125621f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_210 N_A2_c_252_n N_A1_c_384_n 0.0240407f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A2_c_255_n N_A1_c_384_n 7.52702e-19 $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_c_256_n N_A1_c_384_n 0.0223423f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A2_c_257_n N_A1_c_384_n 0.0065184f $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_214 N_A2_c_268_n N_A1_c_384_n 0.00207346f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_215 N_A2_c_259_n N_A1_c_384_n 0.0240407f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_M1004_g N_A1_M1023_g 0.0240407f $X=5.365 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A2_c_268_n N_A1_M1023_g 0.0137744f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_218 N_A2_c_255_n A1 0.0215566f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A2_c_256_n A1 8.88438e-19 $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A2_c_257_n A1 0.0162397f $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_221 N_A2_c_268_n A1 0.108295f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_222 N_A2_c_259_n A1 3.07858e-19 $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A2_c_275_n N_VPWR_M1002_d 4.097e-19 $X=3.375 $Y=1.592 $X2=0 $Y2=0
cc_224 N_A2_c_268_n N_VPWR_M1002_d 0.00147256f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_225 N_A2_c_268_n N_VPWR_M1008_d 0.00178427f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_226 N_A2_c_257_n N_VPWR_M1023_d 3.10624e-19 $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_227 N_A2_c_268_n N_VPWR_M1023_d 0.00147256f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_228 N_A2_c_260_n N_VPWR_M1013_d 0.00184156f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A2_M1002_g N_VPWR_c_452_n 0.00685925f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A2_M1004_g N_VPWR_c_454_n 0.00621909f $X=5.365 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A2_M1013_g N_VPWR_c_454_n 4.98572e-19 $X=5.795 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A2_M1004_g N_VPWR_c_455_n 5.01519e-19 $X=5.365 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A2_M1013_g N_VPWR_c_455_n 0.0062985f $X=5.795 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A2_M1017_g N_VPWR_c_455_n 0.00788945f $X=6.225 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A2_M1004_g N_VPWR_c_458_n 0.00351072f $X=5.365 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A2_M1013_g N_VPWR_c_458_n 0.00351072f $X=5.795 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A2_M1002_g N_VPWR_c_460_n 0.00379212f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A2_M1017_g N_VPWR_c_462_n 0.00351072f $X=6.225 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A2_M1002_g N_VPWR_c_450_n 0.00445145f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A2_M1004_g N_VPWR_c_450_n 0.0040731f $X=5.365 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A2_M1013_g N_VPWR_c_450_n 0.0040731f $X=5.795 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A2_M1017_g N_VPWR_c_450_n 0.00514785f $X=6.225 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A2_c_275_n N_A_223_297#_M1020_d 0.00239676f $X=3.375 $Y=1.592 $X2=0
+ $Y2=0
cc_244 N_A2_c_268_n N_A_223_297#_M1003_s 0.00178427f $X=5.205 $Y=1.39 $X2=0
+ $Y2=0
cc_245 N_A2_c_268_n N_A_223_297#_M1012_s 0.00177993f $X=5.205 $Y=1.39 $X2=0
+ $Y2=0
cc_246 N_A2_c_257_n N_A_223_297#_M1004_s 2.54531e-19 $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_247 N_A2_c_260_n N_A_223_297#_M1004_s 0.00157145f $X=6.285 $Y=1.16 $X2=0
+ $Y2=0
cc_248 N_A2_c_260_n N_A_223_297#_M1017_s 0.0109084f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A2_M1002_g N_A_223_297#_c_584_n 0.0135032f $X=3.205 $Y=1.985 $X2=0
+ $Y2=0
cc_250 N_A2_c_275_n N_A_223_297#_c_584_n 0.0147522f $X=3.375 $Y=1.592 $X2=0
+ $Y2=0
cc_251 N_A2_c_268_n N_A_223_297#_c_584_n 0.0674146f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_252 N_A2_c_275_n N_A_223_297#_c_575_n 0.00381962f $X=3.375 $Y=1.592 $X2=0
+ $Y2=0
cc_253 N_A2_M1004_g N_A_223_297#_c_588_n 0.0137977f $X=5.365 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_A2_c_268_n N_A_223_297#_c_588_n 0.0348689f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_255 N_A2_M1013_g N_A_223_297#_c_590_n 0.0138609f $X=5.795 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A2_M1017_g N_A_223_297#_c_590_n 0.01108f $X=6.225 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A2_c_259_n N_A_223_297#_c_590_n 3.267e-19 $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A2_c_260_n N_A_223_297#_c_590_n 0.03668f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A2_c_259_n N_A_223_297#_c_567_n 2.48761e-19 $X=6.285 $Y=1.16 $X2=0
+ $Y2=0
cc_260 N_A2_c_260_n N_A_223_297#_c_567_n 0.00821211f $X=6.285 $Y=1.16 $X2=0
+ $Y2=0
cc_261 N_A2_c_268_n N_A_223_297#_c_596_n 0.01361f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_262 N_A2_c_257_n N_A_223_297#_c_597_n 0.0146138f $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_263 N_A2_c_259_n N_A_223_297#_c_597_n 3.5494e-19 $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A2_M1002_g N_Y_c_648_n 0.0015018f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A2_c_255_n N_Y_c_648_n 0.0332134f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A2_c_256_n N_Y_c_648_n 0.0030338f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A2_c_275_n N_Y_c_648_n 0.00488521f $X=3.375 $Y=1.592 $X2=0 $Y2=0
cc_268 N_A2_c_258_n N_Y_c_648_n 0.0022552f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A2_c_256_n N_Y_c_649_n 0.00171462f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A2_c_258_n N_Y_c_649_n 0.00517698f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A2_c_268_n N_Y_c_650_n 0.00563538f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_272 N_A2_c_255_n N_Y_c_651_n 0.0270822f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A2_c_256_n N_Y_c_651_n 0.00274735f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A2_c_258_n N_Y_c_651_n 0.01036f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_252_n N_VGND_c_728_n 0.00275982f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A2_c_253_n N_VGND_c_728_n 0.00151324f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A2_c_254_n N_VGND_c_729_n 0.00325061f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A2_c_259_n N_VGND_c_729_n 0.00183945f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A2_c_260_n N_VGND_c_729_n 0.00793512f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A2_c_252_n N_VGND_c_733_n 0.00425616f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_c_258_n N_VGND_c_733_n 0.00420889f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A2_c_253_n N_VGND_c_735_n 0.00427134f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A2_c_254_n N_VGND_c_735_n 0.0054895f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A2_c_252_n N_VGND_c_738_n 0.00583934f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A2_c_253_n N_VGND_c_738_n 0.00580493f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A2_c_254_n N_VGND_c_738_n 0.0108014f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A2_c_258_n N_VGND_c_738_n 0.00641769f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A2_c_258_n N_VGND_c_740_n 0.00348622f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A2_c_258_n N_A_658_47#_c_830_n 0.0032509f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A2_c_252_n N_A_658_47#_c_831_n 0.00274319f $X=5.365 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A2_c_252_n N_A_658_47#_c_832_n 0.00354489f $X=5.365 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A2_c_253_n N_A_658_47#_c_832_n 4.5244e-19 $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A2_c_252_n N_A_658_47#_c_828_n 0.00883987f $X=5.365 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A2_c_253_n N_A_658_47#_c_828_n 0.00975354f $X=5.795 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A2_c_254_n N_A_658_47#_c_828_n 0.00312188f $X=6.225 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A2_c_257_n N_A_658_47#_c_828_n 0.040856f $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_297 N_A2_c_259_n N_A_658_47#_c_828_n 0.00502404f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A2_c_260_n N_A_658_47#_c_828_n 0.0287976f $X=6.285 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A2_c_252_n N_A_658_47#_c_829_n 9.23859e-19 $X=5.365 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_A2_c_257_n N_A_658_47#_c_829_n 0.00994332f $X=5.52 $Y=1.39 $X2=0 $Y2=0
cc_301 N_A2_c_268_n N_A_658_47#_c_829_n 0.00548957f $X=5.205 $Y=1.39 $X2=0 $Y2=0
cc_302 N_A2_c_252_n N_A_658_47#_c_843_n 5.22552e-19 $X=5.365 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A2_c_253_n N_A_658_47#_c_843_n 0.00627823f $X=5.795 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A2_c_254_n N_A_658_47#_c_843_n 0.00529965f $X=6.225 $Y=0.995 $X2=0
+ $Y2=0
cc_305 N_A1_M1003_g N_VPWR_c_452_n 0.00765922f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A1_M1008_g N_VPWR_c_452_n 0.00104385f $X=4.075 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A1_M1003_g N_VPWR_c_453_n 0.00104385f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A1_M1008_g N_VPWR_c_453_n 0.00765006f $X=4.075 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A1_M1012_g N_VPWR_c_453_n 0.00625485f $X=4.505 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A1_M1023_g N_VPWR_c_453_n 4.98572e-19 $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A1_M1012_g N_VPWR_c_454_n 4.98572e-19 $X=4.505 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A1_M1023_g N_VPWR_c_454_n 0.00621909f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A1_M1012_g N_VPWR_c_456_n 0.00351072f $X=4.505 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A1_M1023_g N_VPWR_c_456_n 0.00351072f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A1_M1003_g N_VPWR_c_461_n 0.00351072f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A1_M1008_g N_VPWR_c_461_n 0.00351072f $X=4.075 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A1_M1003_g N_VPWR_c_450_n 0.00411677f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A1_M1008_g N_VPWR_c_450_n 0.00411677f $X=4.075 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A1_M1012_g N_VPWR_c_450_n 0.0040731f $X=4.505 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A1_M1023_g N_VPWR_c_450_n 0.0040731f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A1_M1003_g N_A_223_297#_c_584_n 0.0110962f $X=3.645 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A1_M1008_g N_A_223_297#_c_584_n 0.01108f $X=4.075 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A1_M1012_g N_A_223_297#_c_584_n 0.01108f $X=4.505 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A1_M1023_g N_A_223_297#_c_588_n 0.0110168f $X=4.935 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A1_c_378_n N_Y_c_650_n 0.00981933f $X=3.645 $Y=0.99 $X2=0 $Y2=0
cc_326 N_A1_c_380_n N_Y_c_650_n 0.00987975f $X=4.075 $Y=0.99 $X2=0 $Y2=0
cc_327 N_A1_c_382_n N_Y_c_650_n 0.00987975f $X=4.505 $Y=0.99 $X2=0 $Y2=0
cc_328 N_A1_c_384_n N_Y_c_650_n 0.0102606f $X=4.935 $Y=0.99 $X2=0 $Y2=0
cc_329 A1 N_Y_c_650_n 0.0987456f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_330 N_A1_c_378_n N_VGND_c_733_n 0.00357877f $X=3.645 $Y=0.99 $X2=0 $Y2=0
cc_331 N_A1_c_380_n N_VGND_c_733_n 0.00357877f $X=4.075 $Y=0.99 $X2=0 $Y2=0
cc_332 N_A1_c_382_n N_VGND_c_733_n 0.00357877f $X=4.505 $Y=0.99 $X2=0 $Y2=0
cc_333 N_A1_c_384_n N_VGND_c_733_n 0.00357877f $X=4.935 $Y=0.99 $X2=0 $Y2=0
cc_334 N_A1_c_378_n N_VGND_c_738_n 0.00530427f $X=3.645 $Y=0.99 $X2=0 $Y2=0
cc_335 N_A1_c_380_n N_VGND_c_738_n 0.00527894f $X=4.075 $Y=0.99 $X2=0 $Y2=0
cc_336 N_A1_c_382_n N_VGND_c_738_n 0.00527894f $X=4.505 $Y=0.99 $X2=0 $Y2=0
cc_337 N_A1_c_384_n N_VGND_c_738_n 0.00530427f $X=4.935 $Y=0.99 $X2=0 $Y2=0
cc_338 N_A1_c_378_n N_A_658_47#_c_830_n 0.00979905f $X=3.645 $Y=0.99 $X2=0 $Y2=0
cc_339 N_A1_c_380_n N_A_658_47#_c_830_n 0.00979905f $X=4.075 $Y=0.99 $X2=0 $Y2=0
cc_340 N_A1_c_382_n N_A_658_47#_c_830_n 0.00979905f $X=4.505 $Y=0.99 $X2=0 $Y2=0
cc_341 N_A1_c_384_n N_A_658_47#_c_830_n 0.012154f $X=4.935 $Y=0.99 $X2=0 $Y2=0
cc_342 A1 N_A_658_47#_c_830_n 0.00229035f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_343 N_A1_c_384_n N_A_658_47#_c_829_n 4.2252e-19 $X=4.935 $Y=0.99 $X2=0 $Y2=0
cc_344 N_VPWR_c_450_n N_A_223_297#_M1000_d 0.00369641f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_345 N_VPWR_c_450_n N_A_223_297#_M1005_d 0.00223231f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_450_n N_A_223_297#_M1020_d 0.00258751f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_450_n N_A_223_297#_M1003_s 0.00318969f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_450_n N_A_223_297#_M1012_s 0.00251209f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_450_n N_A_223_297#_M1004_s 0.00254571f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_450_n N_A_223_297#_M1017_s 0.00227407f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_451_n N_A_223_297#_c_610_n 0.0150673f $X=0.72 $Y=2.34 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_460_n N_A_223_297#_c_610_n 0.0125853f $X=3.265 $Y=2.72 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_450_n N_A_223_297#_c_610_n 0.00750689f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_451_n N_A_223_297#_c_569_n 0.00216477f $X=0.72 $Y=2.34 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_460_n N_A_223_297#_c_573_n 0.0330048f $X=3.265 $Y=2.72 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_450_n N_A_223_297#_c_573_n 0.0204525f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_M1002_d N_A_223_297#_c_584_n 0.00367764f $X=3.28 $Y=1.485 $X2=0
+ $Y2=0
cc_358 N_VPWR_M1008_d N_A_223_297#_c_584_n 0.00339518f $X=4.15 $Y=1.485 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_452_n N_A_223_297#_c_584_n 0.0162775f $X=3.43 $Y=2.36 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_453_n N_A_223_297#_c_584_n 0.0162283f $X=4.29 $Y=2.36 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_456_n N_A_223_297#_c_584_n 0.00263122f $X=4.985 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_460_n N_A_223_297#_c_584_n 0.00270999f $X=3.265 $Y=2.72 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_461_n N_A_223_297#_c_584_n 0.00860985f $X=4.125 $Y=2.72 $X2=0
+ $Y2=0
cc_364 N_VPWR_c_450_n N_A_223_297#_c_584_n 0.02585f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_c_460_n N_A_223_297#_c_575_n 0.0668997f $X=3.265 $Y=2.72 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_450_n N_A_223_297#_c_575_n 0.0420965f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_456_n N_A_223_297#_c_626_n 0.0123333f $X=4.985 $Y=2.72 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_450_n N_A_223_297#_c_626_n 0.00721345f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_M1023_d N_A_223_297#_c_588_n 0.00349236f $X=5.01 $Y=1.485 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_454_n N_A_223_297#_c_588_n 0.0162283f $X=5.15 $Y=2.36 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_456_n N_A_223_297#_c_588_n 0.00263122f $X=4.985 $Y=2.72 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_458_n N_A_223_297#_c_588_n 0.00263838f $X=5.845 $Y=2.72 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_450_n N_A_223_297#_c_588_n 0.0101396f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_458_n N_A_223_297#_c_633_n 0.0119785f $X=5.845 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_450_n N_A_223_297#_c_633_n 0.00682467f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_376 N_VPWR_M1013_d N_A_223_297#_c_590_n 0.00338714f $X=5.87 $Y=1.485 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_455_n N_A_223_297#_c_590_n 0.0162283f $X=6.01 $Y=2.36 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_458_n N_A_223_297#_c_590_n 0.00274153f $X=5.845 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_462_n N_A_223_297#_c_590_n 0.00263122f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_450_n N_A_223_297#_c_590_n 0.0104307f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_462_n N_A_223_297#_c_568_n 0.0176323f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_450_n N_A_223_297#_c_568_n 0.00989931f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_450_n N_Y_M1000_s 0.00224864f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_450_n N_Y_M1010_s 0.00224837f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_385 N_A_223_297#_c_573_n N_Y_M1000_s 0.00341119f $X=1.935 $Y=2.34 $X2=0 $Y2=0
cc_386 N_A_223_297#_c_575_n N_Y_M1010_s 0.00335287f $X=3.095 $Y=1.99 $X2=0 $Y2=0
cc_387 N_A_223_297#_c_575_n N_Y_c_648_n 0.0245809f $X=3.095 $Y=1.99 $X2=0 $Y2=0
cc_388 N_A_223_297#_M1005_d N_Y_c_669_n 0.00363318f $X=1.96 $Y=1.485 $X2=0 $Y2=0
cc_389 N_A_223_297#_c_573_n N_Y_c_669_n 0.0206064f $X=1.935 $Y=2.34 $X2=0 $Y2=0
cc_390 N_A_223_297#_c_575_n N_Y_c_669_n 0.0349576f $X=3.095 $Y=1.99 $X2=0 $Y2=0
cc_391 N_Y_c_653_n N_VGND_M1009_d 0.00325948f $X=2.135 $Y=0.74 $X2=0 $Y2=0
cc_392 N_Y_c_668_n N_VGND_M1019_d 0.00411293f $X=2.715 $Y=0.795 $X2=0 $Y2=0
cc_393 N_Y_c_651_n N_VGND_M1019_d 0.00296219f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_394 N_Y_c_653_n N_VGND_c_727_n 0.0163189f $X=2.135 $Y=0.74 $X2=0 $Y2=0
cc_395 N_Y_c_653_n N_VGND_c_731_n 0.00264265f $X=2.135 $Y=0.74 $X2=0 $Y2=0
cc_396 N_Y_c_664_n N_VGND_c_731_n 0.00699602f $X=1.37 $Y=0.535 $X2=0 $Y2=0
cc_397 N_Y_c_651_n N_VGND_c_733_n 0.00210662f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_398 N_Y_M1001_s N_VGND_c_738_n 0.00408233f $X=1.23 $Y=0.235 $X2=0 $Y2=0
cc_399 N_Y_M1018_s N_VGND_c_738_n 0.00256331f $X=2.09 $Y=0.235 $X2=0 $Y2=0
cc_400 N_Y_M1006_s N_VGND_c_738_n 0.00224864f $X=3.72 $Y=0.235 $X2=0 $Y2=0
cc_401 N_Y_M1021_s N_VGND_c_738_n 0.00224864f $X=4.58 $Y=0.235 $X2=0 $Y2=0
cc_402 N_Y_c_653_n N_VGND_c_738_n 0.0102198f $X=2.135 $Y=0.74 $X2=0 $Y2=0
cc_403 N_Y_c_709_p N_VGND_c_738_n 0.00721967f $X=2.23 $Y=0.42 $X2=0 $Y2=0
cc_404 N_Y_c_657_n N_VGND_c_738_n 0.00420955f $X=2.57 $Y=0.78 $X2=0 $Y2=0
cc_405 N_Y_c_649_n N_VGND_c_738_n 0.00313233f $X=3.365 $Y=0.785 $X2=0 $Y2=0
cc_406 N_Y_c_664_n N_VGND_c_738_n 0.00672198f $X=1.37 $Y=0.535 $X2=0 $Y2=0
cc_407 N_Y_c_668_n N_VGND_c_738_n 0.00132048f $X=2.715 $Y=0.795 $X2=0 $Y2=0
cc_408 N_Y_c_651_n N_VGND_c_738_n 0.00489978f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_409 N_Y_c_653_n N_VGND_c_739_n 0.00264265f $X=2.135 $Y=0.74 $X2=0 $Y2=0
cc_410 N_Y_c_709_p N_VGND_c_739_n 0.0123614f $X=2.23 $Y=0.42 $X2=0 $Y2=0
cc_411 N_Y_c_657_n N_VGND_c_739_n 0.0021487f $X=2.57 $Y=0.78 $X2=0 $Y2=0
cc_412 N_Y_c_657_n N_VGND_c_740_n 0.00176606f $X=2.57 $Y=0.78 $X2=0 $Y2=0
cc_413 N_Y_c_668_n N_VGND_c_740_n 0.0241502f $X=2.715 $Y=0.795 $X2=0 $Y2=0
cc_414 N_Y_c_651_n N_VGND_c_740_n 0.0173755f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_415 N_Y_c_650_n N_A_658_47#_M1007_s 0.00152947f $X=4.72 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_416 N_Y_c_650_n N_A_658_47#_M1011_d 0.00172716f $X=4.72 $Y=0.76 $X2=0 $Y2=0
cc_417 N_Y_M1006_s N_A_658_47#_c_830_n 0.00324321f $X=3.72 $Y=0.235 $X2=0 $Y2=0
cc_418 N_Y_M1021_s N_A_658_47#_c_830_n 0.00324321f $X=4.58 $Y=0.235 $X2=0 $Y2=0
cc_419 N_Y_c_649_n N_A_658_47#_c_830_n 0.0821126f $X=3.365 $Y=0.785 $X2=0 $Y2=0
cc_420 N_Y_c_650_n N_A_658_47#_c_829_n 0.00710427f $X=4.72 $Y=0.76 $X2=0 $Y2=0
cc_421 N_VGND_c_738_n N_A_658_47#_M1007_s 0.00223258f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_422 N_VGND_c_738_n N_A_658_47#_M1011_d 0.00223258f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_738_n N_A_658_47#_M1022_d 0.00223235f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_738_n N_A_658_47#_M1015_s 0.00223231f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_733_n N_A_658_47#_c_830_n 0.100183f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_738_n N_A_658_47#_c_830_n 0.064026f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_733_n N_A_658_47#_c_831_n 0.0157493f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_738_n N_A_658_47#_c_831_n 0.00981451f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_M1014_d N_A_658_47#_c_828_n 0.00172391f $X=5.44 $Y=0.235 $X2=0
+ $Y2=0
cc_430 N_VGND_c_728_n N_A_658_47#_c_828_n 0.0130261f $X=5.58 $Y=0.4 $X2=0 $Y2=0
cc_431 N_VGND_c_733_n N_A_658_47#_c_828_n 0.00196536f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_735_n N_A_658_47#_c_828_n 0.00196536f $X=6.345 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_c_738_n N_A_658_47#_c_828_n 0.00828266f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_735_n N_A_658_47#_c_843_n 0.0188765f $X=6.345 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_738_n N_A_658_47#_c_843_n 0.0122527f $X=6.67 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__a211oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__a211oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 1.035000 3.080000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.740000 1.035000 4.500000 1.285000 ;
        RECT 4.175000 1.285000 4.500000 1.655000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.035000 1.785000 1.285000 ;
        RECT 1.035000 1.285000 1.255000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.405000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.826000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.255000 0.835000 0.655000 ;
        RECT 0.575000 0.655000 3.145000 0.855000 ;
        RECT 0.575000 0.855000 0.855000 1.785000 ;
        RECT 0.575000 1.785000 0.905000 2.105000 ;
        RECT 1.505000 0.285000 1.695000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.145000  0.085000 0.395000 0.815000 ;
      RECT 0.145000  1.785000 0.405000 2.285000 ;
      RECT 0.145000  2.285000 2.215000 2.455000 ;
      RECT 1.005000  0.085000 1.335000 0.475000 ;
      RECT 1.075000  1.785000 1.265000 2.255000 ;
      RECT 1.075000  2.255000 2.215000 2.285000 ;
      RECT 1.435000  1.455000 3.975000 1.655000 ;
      RECT 1.435000  1.655000 1.765000 2.075000 ;
      RECT 1.865000  0.085000 2.195000 0.475000 ;
      RECT 1.935000  1.835000 2.215000 2.255000 ;
      RECT 2.385000  0.265000 3.495000 0.475000 ;
      RECT 2.435000  1.835000 2.665000 2.635000 ;
      RECT 2.845000  1.655000 3.115000 2.465000 ;
      RECT 3.295000  1.835000 3.525000 2.635000 ;
      RECT 3.325000  0.475000 3.495000 0.635000 ;
      RECT 3.325000  0.635000 4.435000 0.855000 ;
      RECT 3.675000  0.085000 4.005000 0.455000 ;
      RECT 3.705000  1.655000 3.975000 2.465000 ;
      RECT 4.155000  1.835000 4.385000 2.635000 ;
      RECT 4.185000  0.265000 4.435000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_2

* File: sky130_fd_sc_hd__o21ba_2.pxi.spice
* Created: Thu Aug 27 14:36:06 2020
* 
x_PM_SKY130_FD_SC_HD__O21BA_2%B1_N N_B1_N_M1010_g N_B1_N_M1006_g B1_N B1_N
+ N_B1_N_c_75_n N_B1_N_c_76_n PM_SKY130_FD_SC_HD__O21BA_2%B1_N
x_PM_SKY130_FD_SC_HD__O21BA_2%A_174_21# N_A_174_21#_M1003_s N_A_174_21#_M1004_d
+ N_A_174_21#_c_110_n N_A_174_21#_M1002_g N_A_174_21#_M1007_g
+ N_A_174_21#_c_111_n N_A_174_21#_M1011_g N_A_174_21#_M1009_g
+ N_A_174_21#_c_112_n N_A_174_21#_c_113_n N_A_174_21#_c_114_n
+ N_A_174_21#_c_115_n N_A_174_21#_c_116_n N_A_174_21#_c_152_p
+ N_A_174_21#_c_121_n N_A_174_21#_c_117_n PM_SKY130_FD_SC_HD__O21BA_2%A_174_21#
x_PM_SKY130_FD_SC_HD__O21BA_2%A_27_93# N_A_27_93#_M1010_s N_A_27_93#_M1006_s
+ N_A_27_93#_c_211_n N_A_27_93#_M1003_g N_A_27_93#_M1004_g N_A_27_93#_c_212_n
+ N_A_27_93#_c_213_n N_A_27_93#_c_220_n N_A_27_93#_c_221_n N_A_27_93#_c_222_n
+ N_A_27_93#_c_223_n N_A_27_93#_c_214_n N_A_27_93#_c_215_n N_A_27_93#_c_216_n
+ PM_SKY130_FD_SC_HD__O21BA_2%A_27_93#
x_PM_SKY130_FD_SC_HD__O21BA_2%A2 N_A2_M1005_g N_A2_M1000_g A2 N_A2_c_287_n
+ N_A2_c_288_n N_A2_c_289_n PM_SKY130_FD_SC_HD__O21BA_2%A2
x_PM_SKY130_FD_SC_HD__O21BA_2%A1 N_A1_M1001_g N_A1_M1008_g A1 A1 N_A1_c_324_n
+ N_A1_c_325_n N_A1_c_326_n PM_SKY130_FD_SC_HD__O21BA_2%A1
x_PM_SKY130_FD_SC_HD__O21BA_2%VPWR N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_M1001_d
+ N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n VPWR N_VPWR_c_357_n
+ N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_353_n
+ PM_SKY130_FD_SC_HD__O21BA_2%VPWR
x_PM_SKY130_FD_SC_HD__O21BA_2%X N_X_M1002_s N_X_M1007_s N_X_c_408_n N_X_c_414_n
+ X N_X_c_425_n PM_SKY130_FD_SC_HD__O21BA_2%X
x_PM_SKY130_FD_SC_HD__O21BA_2%VGND N_VGND_M1010_d N_VGND_M1011_d N_VGND_M1005_d
+ N_VGND_c_438_n N_VGND_c_439_n N_VGND_c_440_n VGND N_VGND_c_441_n
+ N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n
+ N_VGND_c_447_n N_VGND_c_448_n PM_SKY130_FD_SC_HD__O21BA_2%VGND
x_PM_SKY130_FD_SC_HD__O21BA_2%A_478_47# N_A_478_47#_M1003_d N_A_478_47#_M1008_d
+ N_A_478_47#_c_505_n N_A_478_47#_c_500_n N_A_478_47#_c_501_n
+ N_A_478_47#_c_502_n PM_SKY130_FD_SC_HD__O21BA_2%A_478_47#
cc_1 VNB B1_N 0.00302066f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_2 VNB N_B1_N_c_75_n 0.0242164f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_B1_N_c_76_n 0.02048f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_4 VNB N_A_174_21#_c_110_n 0.0185884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_174_21#_c_111_n 0.0186092f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_6 VNB N_A_174_21#_c_112_n 0.00626998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_174_21#_c_113_n 0.00488265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_174_21#_c_114_n 0.0011214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_174_21#_c_115_n 0.00579898f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_174_21#_c_116_n 6.70754e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_174_21#_c_117_n 0.0354183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_93#_c_211_n 0.0206731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_93#_c_212_n 0.0364621f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_14 VNB N_A_27_93#_c_213_n 0.0101833f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_15 VNB N_A_27_93#_c_214_n 0.0015776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_93#_c_215_n 0.0181192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_93#_c_216_n 0.0220555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_287_n 0.0193059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_288_n 0.0080067f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_20 VNB N_A2_c_289_n 0.0167156f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_21 VNB N_A1_c_324_n 0.0321205f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_22 VNB N_A1_c_325_n 0.0105018f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_23 VNB N_A1_c_326_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_24 VNB N_VPWR_c_353_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_408_n 6.67958e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_26 VNB N_VGND_c_438_n 0.0088337f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_27 VNB N_VGND_c_439_n 0.00597916f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.325
cc_28 VNB N_VGND_c_440_n 0.00465817f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_29 VNB N_VGND_c_441_n 0.0193449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_442_n 0.0161981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_443_n 0.0294862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_444_n 0.0174072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_445_n 0.210401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_446_n 0.00345893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_447_n 0.00564938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_448_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_478_47#_c_500_n 0.0156944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_478_47#_c_501_n 0.00226847f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_39 VNB N_A_478_47#_c_502_n 0.0184083f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_40 VPB N_B1_N_M1006_g 0.0220679f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_41 VPB B1_N 4.80488e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_42 VPB B1_N 0.00247149f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_43 VPB N_B1_N_c_75_n 0.0047062f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_44 VPB N_A_174_21#_M1007_g 0.0202136f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_45 VPB N_A_174_21#_M1009_g 0.0214596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_174_21#_c_114_n 0.00137925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_174_21#_c_121_n 0.00485734f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_174_21#_c_117_n 0.00627021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_93#_M1004_g 0.0237823f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_50 VPB N_A_27_93#_c_212_n 0.0204081f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_51 VPB N_A_27_93#_c_213_n 6.59856e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_52 VPB N_A_27_93#_c_220_n 0.00601347f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.53
cc_53 VPB N_A_27_93#_c_221_n 0.00826367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_93#_c_222_n 6.28953e-19 $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_55 VPB N_A_27_93#_c_223_n 0.0119472f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_56 VPB N_A_27_93#_c_214_n 0.00272957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_93#_c_216_n 0.00888141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A2_M1000_g 0.0188676f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_59 VPB N_A2_c_287_n 0.00408489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A1_M1001_g 0.021722f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.675
cc_61 VPB N_A1_c_324_n 0.00736483f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_62 VPB N_A1_c_325_n 0.0156899f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_63 VPB N_VPWR_c_354_n 0.0154239f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_64 VPB N_VPWR_c_355_n 0.0120646f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_65 VPB N_VPWR_c_356_n 0.0260645f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.325
cc_66 VPB N_VPWR_c_357_n 0.016934f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_67 VPB N_VPWR_c_358_n 0.0258873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_359_n 0.00622792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_360_n 0.011884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_361_n 0.0197769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_353_n 0.0502642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_408_n 0.00157803f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_73 N_B1_N_c_76_n N_A_174_21#_c_110_n 0.00850967f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B1_N_M1006_g N_A_174_21#_M1007_g 0.022536f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_75 B1_N N_A_174_21#_M1007_g 0.00260914f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_76 B1_N N_A_174_21#_c_117_n 0.00244321f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_77 N_B1_N_c_75_n N_A_174_21#_c_117_n 0.0196228f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_N_M1006_g N_A_27_93#_c_222_n 0.0109407f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_79 B1_N N_A_27_93#_c_222_n 0.00409821f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_80 B1_N N_A_27_93#_c_222_n 0.0133274f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_81 N_B1_N_M1006_g N_A_27_93#_c_223_n 0.00340695f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_82 N_B1_N_c_76_n N_A_27_93#_c_215_n 8.00287e-19 $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B1_N_M1006_g N_A_27_93#_c_216_n 0.00350801f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_84 B1_N N_A_27_93#_c_216_n 0.0248826f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_85 B1_N N_A_27_93#_c_216_n 0.00763889f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_86 N_B1_N_c_75_n N_A_27_93#_c_216_n 0.00755993f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_N_c_76_n N_A_27_93#_c_216_n 0.00547137f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_88 B1_N N_VPWR_M1006_d 0.0052227f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_89 N_B1_N_M1006_g N_VPWR_c_354_n 6.50777e-19 $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_90 N_B1_N_M1006_g N_VPWR_c_357_n 0.00215805f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_91 N_B1_N_M1006_g N_VPWR_c_353_n 0.00350691f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_92 B1_N N_X_c_408_n 0.025008f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_93 B1_N N_X_c_408_n 0.0121667f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_94 N_B1_N_c_75_n N_X_c_408_n 2.89837e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B1_N_c_76_n N_X_c_408_n 8.85159e-19 $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_96 B1_N N_X_c_414_n 0.0149922f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_97 B1_N N_VGND_c_438_n 0.0149603f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B1_N_c_75_n N_VGND_c_438_n 0.0011232f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B1_N_c_76_n N_VGND_c_438_n 0.00268459f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B1_N_c_76_n N_VGND_c_441_n 0.00510437f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_N_c_76_n N_VGND_c_445_n 0.00512902f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_174_21#_c_113_n N_A_27_93#_c_211_n 0.0056297f $X=2.105 $Y=0.38 $X2=0
+ $Y2=0
cc_103 N_A_174_21#_c_114_n N_A_27_93#_c_211_n 0.00434463f $X=2.19 $Y=1.455 $X2=0
+ $Y2=0
cc_104 N_A_174_21#_c_115_n N_A_27_93#_c_211_n 6.74391e-19 $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_105 N_A_174_21#_c_116_n N_A_27_93#_c_211_n 0.001852f $X=2.107 $Y=0.74 $X2=0
+ $Y2=0
cc_106 N_A_174_21#_c_114_n N_A_27_93#_M1004_g 0.00470087f $X=2.19 $Y=1.455 $X2=0
+ $Y2=0
cc_107 N_A_174_21#_c_121_n N_A_27_93#_M1004_g 0.0279709f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_108 N_A_174_21#_c_112_n N_A_27_93#_c_212_n 0.00330825f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_109 N_A_174_21#_c_114_n N_A_27_93#_c_212_n 0.0140274f $X=2.19 $Y=1.455 $X2=0
+ $Y2=0
cc_110 N_A_174_21#_c_115_n N_A_27_93#_c_212_n 0.00145398f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_111 N_A_174_21#_c_116_n N_A_27_93#_c_212_n 0.0071269f $X=2.107 $Y=0.74 $X2=0
+ $Y2=0
cc_112 N_A_174_21#_c_121_n N_A_27_93#_c_212_n 7.55821e-19 $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_113 N_A_174_21#_c_117_n N_A_27_93#_c_212_n 0.0225029f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_A_174_21#_c_114_n N_A_27_93#_c_213_n 0.00430976f $X=2.19 $Y=1.455 $X2=0
+ $Y2=0
cc_115 N_A_174_21#_M1007_g N_A_27_93#_c_222_n 0.0139133f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_174_21#_M1009_g N_A_27_93#_c_222_n 0.0146102f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_174_21#_c_115_n N_A_27_93#_c_222_n 0.00294414f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_118 N_A_174_21#_c_121_n N_A_27_93#_c_222_n 0.0151336f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_119 N_A_174_21#_M1009_g N_A_27_93#_c_214_n 0.0119886f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_174_21#_c_112_n N_A_27_93#_c_214_n 0.0134259f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_174_21#_c_114_n N_A_27_93#_c_214_n 0.0321559f $X=2.19 $Y=1.455 $X2=0
+ $Y2=0
cc_122 N_A_174_21#_c_115_n N_A_27_93#_c_214_n 0.016052f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_123 N_A_174_21#_c_121_n N_A_27_93#_c_214_n 0.0330781f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_124 N_A_174_21#_c_117_n N_A_27_93#_c_214_n 0.00106127f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_125 N_A_174_21#_c_114_n N_A2_M1000_g 6.31887e-19 $X=2.19 $Y=1.455 $X2=0 $Y2=0
cc_126 N_A_174_21#_c_152_p N_A2_M1000_g 0.00636844f $X=2.562 $Y=1.745 $X2=0
+ $Y2=0
cc_127 N_A_174_21#_c_121_n N_A2_M1000_g 0.00927355f $X=2.585 $Y=1.62 $X2=0 $Y2=0
cc_128 N_A_174_21#_c_114_n N_A2_c_287_n 8.29066e-19 $X=2.19 $Y=1.455 $X2=0 $Y2=0
cc_129 N_A_174_21#_c_121_n N_A2_c_287_n 0.0029336f $X=2.585 $Y=1.62 $X2=0 $Y2=0
cc_130 N_A_174_21#_c_114_n N_A2_c_288_n 0.0162992f $X=2.19 $Y=1.455 $X2=0 $Y2=0
cc_131 N_A_174_21#_c_121_n N_A2_c_288_n 0.0230718f $X=2.585 $Y=1.62 $X2=0 $Y2=0
cc_132 N_A_174_21#_c_113_n N_A2_c_289_n 4.31957e-19 $X=2.105 $Y=0.38 $X2=0 $Y2=0
cc_133 N_A_174_21#_c_114_n N_A2_c_289_n 4.95557e-19 $X=2.19 $Y=1.455 $X2=0 $Y2=0
cc_134 N_A_174_21#_c_152_p N_A1_M1001_g 0.00113093f $X=2.562 $Y=1.745 $X2=0
+ $Y2=0
cc_135 N_A_174_21#_c_121_n N_A1_M1001_g 0.00202926f $X=2.585 $Y=1.62 $X2=0 $Y2=0
cc_136 N_A_174_21#_c_121_n N_A1_c_325_n 0.0072862f $X=2.585 $Y=1.62 $X2=0 $Y2=0
cc_137 N_A_174_21#_c_121_n N_VPWR_M1009_d 0.00644856f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_138 N_A_174_21#_M1007_g N_VPWR_c_354_n 0.0101377f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_174_21#_M1009_g N_VPWR_c_354_n 0.00124983f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_174_21#_c_152_p N_VPWR_c_356_n 0.0139781f $X=2.562 $Y=1.745 $X2=0
+ $Y2=0
cc_141 N_A_174_21#_c_121_n N_VPWR_c_356_n 0.00544786f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_142 N_A_174_21#_c_152_p N_VPWR_c_358_n 0.0185827f $X=2.562 $Y=1.745 $X2=0
+ $Y2=0
cc_143 N_A_174_21#_c_121_n N_VPWR_c_358_n 0.00255839f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_144 N_A_174_21#_M1007_g N_VPWR_c_360_n 0.00345093f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_174_21#_M1009_g N_VPWR_c_360_n 0.00330683f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_174_21#_M1007_g N_VPWR_c_361_n 0.00127272f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_174_21#_M1009_g N_VPWR_c_361_n 0.0109001f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_174_21#_c_121_n N_VPWR_c_361_n 0.0065293f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_149 N_A_174_21#_M1004_d N_VPWR_c_353_n 0.00267758f $X=2.39 $Y=1.485 $X2=0
+ $Y2=0
cc_150 N_A_174_21#_M1007_g N_VPWR_c_353_n 0.0040856f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_174_21#_M1009_g N_VPWR_c_353_n 0.00392244f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_174_21#_c_152_p N_VPWR_c_353_n 0.0122055f $X=2.562 $Y=1.745 $X2=0
+ $Y2=0
cc_153 N_A_174_21#_c_121_n N_VPWR_c_353_n 0.00463302f $X=2.585 $Y=1.62 $X2=0
+ $Y2=0
cc_154 N_A_174_21#_c_110_n N_X_c_408_n 0.00935263f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_174_21#_M1007_g N_X_c_408_n 0.00353062f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_174_21#_c_111_n N_X_c_408_n 0.00311425f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_174_21#_M1009_g N_X_c_408_n 0.00164983f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_174_21#_c_115_n N_X_c_408_n 0.0423187f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_174_21#_c_117_n N_X_c_408_n 0.0117034f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_174_21#_M1007_g N_X_c_414_n 0.00422686f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_174_21#_M1009_g N_X_c_414_n 0.00503697f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_174_21#_c_115_n N_X_c_414_n 0.00426886f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_174_21#_c_117_n N_X_c_414_n 0.00347997f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_174_21#_c_110_n N_X_c_425_n 0.00549377f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_174_21#_c_117_n N_X_c_425_n 0.00275312f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_174_21#_c_112_n N_VGND_M1011_d 0.00573967f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_174_21#_c_115_n N_VGND_M1011_d 0.00192584f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_174_21#_c_110_n N_VGND_c_438_n 0.00688572f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_174_21#_c_110_n N_VGND_c_439_n 5.00906e-19 $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_174_21#_c_111_n N_VGND_c_439_n 0.00842215f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_174_21#_c_112_n N_VGND_c_439_n 0.0135256f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_174_21#_c_113_n N_VGND_c_439_n 0.0193004f $X=2.105 $Y=0.38 $X2=0
+ $Y2=0
cc_173 N_A_174_21#_c_115_n N_VGND_c_439_n 0.00972384f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_174_21#_c_110_n N_VGND_c_442_n 0.00471631f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A_174_21#_c_111_n N_VGND_c_442_n 0.0046653f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_174_21#_c_112_n N_VGND_c_443_n 0.00296166f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_174_21#_c_113_n N_VGND_c_443_n 0.0212296f $X=2.105 $Y=0.38 $X2=0
+ $Y2=0
cc_178 N_A_174_21#_M1003_s N_VGND_c_445_n 0.00209319f $X=1.98 $Y=0.235 $X2=0
+ $Y2=0
cc_179 N_A_174_21#_c_110_n N_VGND_c_445_n 0.00935686f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_174_21#_c_111_n N_VGND_c_445_n 0.00789179f $X=1.365 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_174_21#_c_112_n N_VGND_c_445_n 0.00552058f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_182 N_A_174_21#_c_113_n N_VGND_c_445_n 0.0125676f $X=2.105 $Y=0.38 $X2=0
+ $Y2=0
cc_183 N_A_174_21#_c_115_n N_VGND_c_445_n 7.8771e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_174_21#_c_114_n N_A_478_47#_c_501_n 0.00357582f $X=2.19 $Y=1.455
+ $X2=0 $Y2=0
cc_185 N_A_27_93#_M1004_g N_A2_M1000_g 0.0115077f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_93#_c_213_n N_A2_c_287_n 0.0223337f $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_93#_c_213_n N_A2_c_288_n 0.00168903f $X=2.315 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_27_93#_c_211_n N_A2_c_289_n 0.0185121f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_27_93#_c_222_n N_VPWR_M1006_d 0.00570778f $X=1.765 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_27_93#_c_222_n N_VPWR_M1009_d 0.0175753f $X=1.765 $Y=1.95 $X2=0 $Y2=0
cc_191 N_A_27_93#_c_214_n N_VPWR_M1009_d 0.0115999f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_93#_c_222_n N_VPWR_c_354_n 0.0256561f $X=1.765 $Y=1.95 $X2=0 $Y2=0
cc_193 N_A_27_93#_c_222_n N_VPWR_c_357_n 0.00181145f $X=1.765 $Y=1.95 $X2=0
+ $Y2=0
cc_194 N_A_27_93#_c_223_n N_VPWR_c_357_n 0.00563795f $X=0.395 $Y=1.95 $X2=0
+ $Y2=0
cc_195 N_A_27_93#_M1004_g N_VPWR_c_358_n 0.00432313f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_27_93#_c_222_n N_VPWR_c_360_n 0.00684751f $X=1.765 $Y=1.95 $X2=0
+ $Y2=0
cc_197 N_A_27_93#_M1004_g N_VPWR_c_361_n 0.00518337f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_27_93#_c_222_n N_VPWR_c_361_n 0.0367075f $X=1.765 $Y=1.95 $X2=0 $Y2=0
cc_199 N_A_27_93#_M1004_g N_VPWR_c_353_n 0.00717985f $X=2.315 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_27_93#_c_222_n N_VPWR_c_353_n 0.0196784f $X=1.765 $Y=1.95 $X2=0 $Y2=0
cc_201 N_A_27_93#_c_223_n N_VPWR_c_353_n 0.00893864f $X=0.395 $Y=1.95 $X2=0
+ $Y2=0
cc_202 N_A_27_93#_c_222_n N_X_M1007_s 0.00444151f $X=1.765 $Y=1.95 $X2=0 $Y2=0
cc_203 N_A_27_93#_c_214_n N_X_c_408_n 0.00493741f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_27_93#_c_222_n N_X_c_414_n 0.0206325f $X=1.765 $Y=1.95 $X2=0 $Y2=0
cc_205 N_A_27_93#_c_214_n N_X_c_414_n 0.00747202f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_27_93#_c_215_n N_VGND_c_438_n 0.00197424f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_207 N_A_27_93#_c_211_n N_VGND_c_439_n 0.00244811f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_27_93#_c_215_n N_VGND_c_441_n 0.00842023f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_209 N_A_27_93#_c_211_n N_VGND_c_443_n 0.00533769f $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_27_93#_c_211_n N_VGND_c_445_n 0.011004f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_27_93#_c_215_n N_VGND_c_445_n 0.00885431f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_212 N_A_27_93#_c_211_n N_A_478_47#_c_501_n 6.9769e-19 $X=2.315 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A2_M1000_g N_A1_M1001_g 0.0490473f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A2_c_287_n N_A1_c_324_n 0.0490473f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A2_c_288_n N_A1_c_324_n 0.00127973f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_c_287_n N_A1_c_325_n 0.00186401f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A2_c_288_n N_A1_c_325_n 0.0175619f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A2_c_289_n N_A1_c_326_n 0.0258192f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A2_M1000_g N_VPWR_c_356_n 0.00286602f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A2_M1000_g N_VPWR_c_358_n 0.00578292f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A2_M1000_g N_VPWR_c_353_n 0.0105848f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A2_c_289_n N_VGND_c_440_n 0.00268723f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_289_n N_VGND_c_443_n 0.0042866f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_289_n N_VGND_c_445_n 0.0059799f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A2_c_289_n N_A_478_47#_c_505_n 0.00570335f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A2_c_288_n N_A_478_47#_c_500_n 0.0131891f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A2_c_289_n N_A_478_47#_c_500_n 0.00845772f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A2_c_287_n N_A_478_47#_c_501_n 0.00292653f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A2_c_288_n N_A_478_47#_c_501_n 0.024539f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A2_c_289_n N_A_478_47#_c_501_n 0.00231212f $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A2_c_289_n N_A_478_47#_c_502_n 5.47074e-19 $X=2.735 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A1_c_325_n N_VPWR_M1001_d 0.00358226f $X=3.265 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A1_M1001_g N_VPWR_c_356_n 0.0165737f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_c_324_n N_VPWR_c_356_n 7.27962e-19 $X=3.265 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A1_c_325_n N_VPWR_c_356_n 0.0179278f $X=3.265 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A1_M1001_g N_VPWR_c_358_n 0.0046653f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A1_M1001_g N_VPWR_c_353_n 0.00783311f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A1_c_326_n N_VGND_c_440_n 0.00268723f $X=3.255 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A1_c_326_n N_VGND_c_444_n 0.00425021f $X=3.255 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A1_c_326_n N_VGND_c_445_n 0.00671814f $X=3.255 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A1_c_326_n N_A_478_47#_c_505_n 5.19634e-19 $X=3.255 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A1_c_324_n N_A_478_47#_c_500_n 0.0056401f $X=3.265 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A1_c_325_n N_A_478_47#_c_500_n 0.0414457f $X=3.265 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A1_c_326_n N_A_478_47#_c_500_n 0.00972067f $X=3.255 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A1_c_326_n N_A_478_47#_c_502_n 0.00634641f $X=3.255 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_353_n N_X_M1007_s 0.00335014f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_247 N_VPWR_c_353_n A_574_297# 0.00897657f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_248 N_X_c_408_n N_VGND_c_438_n 0.0162189f $X=1.03 $Y=1.495 $X2=0 $Y2=0
cc_249 N_X_c_425_n N_VGND_c_438_n 0.0249733f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_250 N_X_c_425_n N_VGND_c_442_n 0.0174312f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_251 N_X_M1002_s N_VGND_c_445_n 0.00385329f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_252 N_X_c_425_n N_VGND_c_445_n 0.0107455f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_253 N_VGND_c_445_n N_A_478_47#_M1003_d 0.00467811f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_254 N_VGND_c_445_n N_A_478_47#_M1008_d 0.00209863f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_443_n N_A_478_47#_c_505_n 0.0108847f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_445_n N_A_478_47#_c_505_n 0.0105737f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_M1005_d N_A_478_47#_c_500_n 0.00165819f $X=2.865 $Y=0.235 $X2=0
+ $Y2=0
cc_258 N_VGND_c_440_n N_A_478_47#_c_500_n 0.0116529f $X=3 $Y=0.39 $X2=0 $Y2=0
cc_259 N_VGND_c_443_n N_A_478_47#_c_500_n 0.00193763f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_444_n N_A_478_47#_c_500_n 0.00193763f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_445_n N_A_478_47#_c_500_n 0.00827287f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_444_n N_A_478_47#_c_502_n 0.0194423f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_445_n N_A_478_47#_c_502_n 0.012503f $X=3.45 $Y=0 $X2=0 $Y2=0

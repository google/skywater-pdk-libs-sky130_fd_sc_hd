* File: sky130_fd_sc_hd__a2111o_2.spice.SKY130_FD_SC_HD__A2111O_2.pxi
* Created: Thu Aug 27 13:58:37 2020
* 
x_PM_SKY130_FD_SC_HD__A2111O_2%A_86_235# N_A_86_235#_M1008_d N_A_86_235#_M1001_d
+ N_A_86_235#_M1002_s N_A_86_235#_M1005_g N_A_86_235#_c_74_n N_A_86_235#_M1004_g
+ N_A_86_235#_M1012_g N_A_86_235#_c_75_n N_A_86_235#_M1009_g N_A_86_235#_c_76_n
+ N_A_86_235#_c_77_n N_A_86_235#_c_83_n N_A_86_235#_c_84_n N_A_86_235#_c_92_p
+ N_A_86_235#_c_138_p N_A_86_235#_c_105_p N_A_86_235#_c_102_p
+ N_A_86_235#_c_113_p N_A_86_235#_c_78_n N_A_86_235#_c_85_n N_A_86_235#_c_98_p
+ N_A_86_235#_c_79_n PM_SKY130_FD_SC_HD__A2111O_2%A_86_235#
x_PM_SKY130_FD_SC_HD__A2111O_2%D1 N_D1_M1008_g N_D1_M1002_g D1 D1 D1 D1
+ N_D1_c_169_n N_D1_c_170_n N_D1_c_171_n PM_SKY130_FD_SC_HD__A2111O_2%D1
x_PM_SKY130_FD_SC_HD__A2111O_2%C1 N_C1_M1006_g N_C1_M1011_g C1 C1 C1 C1
+ N_C1_c_209_n N_C1_c_210_n PM_SKY130_FD_SC_HD__A2111O_2%C1
x_PM_SKY130_FD_SC_HD__A2111O_2%B1 N_B1_M1010_g N_B1_M1001_g B1 B1 N_B1_c_244_n
+ N_B1_c_245_n PM_SKY130_FD_SC_HD__A2111O_2%B1
x_PM_SKY130_FD_SC_HD__A2111O_2%A1 N_A1_M1013_g N_A1_M1000_g A1 A1 A1
+ N_A1_c_279_n N_A1_c_280_n N_A1_c_281_n A1 A1 PM_SKY130_FD_SC_HD__A2111O_2%A1
x_PM_SKY130_FD_SC_HD__A2111O_2%A2 N_A2_M1003_g N_A2_M1007_g A2 A2 N_A2_c_323_n
+ N_A2_c_324_n N_A2_c_325_n PM_SKY130_FD_SC_HD__A2111O_2%A2
x_PM_SKY130_FD_SC_HD__A2111O_2%VPWR N_VPWR_M1005_d N_VPWR_M1012_d N_VPWR_M1000_d
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_357_n VPWR N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_351_n
+ N_VPWR_c_361_n PM_SKY130_FD_SC_HD__A2111O_2%VPWR
x_PM_SKY130_FD_SC_HD__A2111O_2%X N_X_M1004_d N_X_M1005_s X X X X X X N_X_c_407_n
+ PM_SKY130_FD_SC_HD__A2111O_2%X
x_PM_SKY130_FD_SC_HD__A2111O_2%A_607_297# N_A_607_297#_M1010_d
+ N_A_607_297#_M1007_d N_A_607_297#_c_430_n N_A_607_297#_c_442_n
+ N_A_607_297#_c_428_n PM_SKY130_FD_SC_HD__A2111O_2%A_607_297#
x_PM_SKY130_FD_SC_HD__A2111O_2%VGND N_VGND_M1004_s N_VGND_M1009_s N_VGND_M1011_d
+ N_VGND_M1003_d N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_467_n N_VGND_c_451_n
+ N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n
+ N_VGND_c_457_n VGND N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n
+ N_VGND_c_461_n PM_SKY130_FD_SC_HD__A2111O_2%VGND
cc_1 VNB N_A_86_235#_c_74_n 0.0216065f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.995
cc_2 VNB N_A_86_235#_c_75_n 0.0189482f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=0.995
cc_3 VNB N_A_86_235#_c_76_n 0.00129763f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=1.2
cc_4 VNB N_A_86_235#_c_77_n 0.00439183f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.075
cc_5 VNB N_A_86_235#_c_78_n 0.00232761f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.2
cc_6 VNB N_A_86_235#_c_79_n 0.0694993f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=1.16
cc_7 VNB N_D1_c_169_n 0.0259755f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.325
cc_8 VNB N_D1_c_170_n 0.00402909f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.985
cc_9 VNB N_D1_c_171_n 0.0189641f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.985
cc_10 VNB C1 0.00357663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_C1_c_209_n 0.0241582f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.325
cc_12 VNB N_C1_c_210_n 0.0175047f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.985
cc_13 VNB B1 0.0013952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B1_c_244_n 0.026154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_245_n 0.0179785f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_16 VNB N_A1_c_279_n 0.0232f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_17 VNB N_A1_c_280_n 0.0060727f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.325
cc_18 VNB N_A1_c_281_n 0.0165041f $X=-0.19 $Y=-0.24 $X2=0.935 $Y2=1.985
cc_19 VNB A1 0.0017574f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=0.56
cc_20 VNB N_A2_c_323_n 0.0280197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_324_n 0.0203618f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.995
cc_22 VNB N_A2_c_325_n 0.0231176f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_23 VNB N_VPWR_c_351_n 0.193827f $X=-0.19 $Y=-0.24 $X2=3.09 $Y2=0.7
cc_24 VNB N_X_c_407_n 0.00100421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_449_n 0.0116412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_450_n 0.0469232f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_27 VNB N_VGND_c_451_n 0.00493598f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=0.56
cc_28 VNB N_VGND_c_452_n 0.0116445f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.2
cc_29 VNB N_VGND_c_453_n 0.0287931f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.16
cc_30 VNB N_VGND_c_454_n 0.0103329f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.075
cc_31 VNB N_VGND_c_455_n 0.0043718f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=1.64
cc_32 VNB N_VGND_c_456_n 0.0133821f $X=-0.19 $Y=-0.24 $X2=1.7 $Y2=1.66
cc_33 VNB N_VGND_c_457_n 0.00630985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_458_n 0.016088f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=0.615
cc_35 VNB N_VGND_c_459_n 0.0321696f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=0.7
cc_36 VNB N_VGND_c_460_n 0.00427278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_461_n 0.236287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_86_235#_M1005_g 0.0251848f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_39 VPB N_A_86_235#_M1012_g 0.0223785f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.985
cc_40 VPB N_A_86_235#_c_76_n 0.0028457f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.2
cc_41 VPB N_A_86_235#_c_83_n 0.00145687f $X=-0.19 $Y=1.305 $X2=1.64 $Y2=1.64
cc_42 VPB N_A_86_235#_c_84_n 0.00900369f $X=-0.19 $Y=1.305 $X2=1.7 $Y2=1.66
cc_43 VPB N_A_86_235#_c_85_n 0.00373334f $X=-0.19 $Y=1.305 $X2=1.64 $Y2=1.495
cc_44 VPB N_A_86_235#_c_79_n 0.0206662f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.16
cc_45 VPB N_D1_M1002_g 0.0216253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB D1 0.00263934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_D1_c_169_n 0.00832809f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.325
cc_48 VPB N_D1_c_170_n 0.00287817f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.985
cc_49 VPB N_C1_M1006_g 0.018719f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.485
cc_50 VPB C1 0.00108331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_C1_c_209_n 0.00637716f $X=-0.19 $Y=1.305 $X2=0.935 $Y2=1.325
cc_52 VPB N_B1_M1010_g 0.0206266f $X=-0.19 $Y=1.305 $X2=1.575 $Y2=1.485
cc_53 VPB B1 9.99185e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_B1_c_244_n 0.00658824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A1_M1000_g 0.0197733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A1_c_279_n 0.00625292f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=0.56
cc_57 VPB A1 0.0022916f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=0.56
cc_58 VPB N_A2_M1007_g 0.023648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A2_c_323_n 0.00662171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A2_c_324_n 0.0212638f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=0.995
cc_61 VPB N_VPWR_c_352_n 0.0105238f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.325
cc_62 VPB N_VPWR_c_353_n 0.0404788f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_63 VPB N_VPWR_c_354_n 0.0142037f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=0.56
cc_64 VPB N_VPWR_c_355_n 0.0055721f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=0.56
cc_65 VPB N_VPWR_c_356_n 0.0611249f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.2
cc_66 VPB N_VPWR_c_357_n 0.0063111f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.16
cc_67 VPB N_VPWR_c_358_n 0.0165977f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=0.785
cc_68 VPB N_VPWR_c_359_n 0.018915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_351_n 0.0522391f $X=-0.19 $Y=1.305 $X2=3.09 $Y2=0.7
cc_70 VPB N_VPWR_c_361_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.2
cc_71 VPB N_X_c_407_n 0.00153327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_607_297#_c_428_n 0.0261041f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_73 N_A_86_235#_c_83_n N_D1_M1002_g 0.00593816f $X=1.64 $Y=1.64 $X2=0 $Y2=0
cc_74 N_A_86_235#_c_84_n N_D1_M1002_g 0.00388782f $X=1.7 $Y=1.66 $X2=0 $Y2=0
cc_75 N_A_86_235#_c_85_n N_D1_M1002_g 0.00106688f $X=1.64 $Y=1.495 $X2=0 $Y2=0
cc_76 N_A_86_235#_c_85_n D1 0.0097859f $X=1.64 $Y=1.495 $X2=0 $Y2=0
cc_77 N_A_86_235#_c_77_n N_D1_c_169_n 7.10858e-19 $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_78 N_A_86_235#_c_92_p N_D1_c_169_n 0.00344203f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_79 N_A_86_235#_c_78_n N_D1_c_169_n 0.00243509f $X=1.6 $Y=1.2 $X2=0 $Y2=0
cc_80 N_A_86_235#_c_79_n N_D1_c_169_n 0.00875872f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_86_235#_c_77_n N_D1_c_170_n 0.00586608f $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_82 N_A_86_235#_c_92_p N_D1_c_170_n 0.0160027f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_83 N_A_86_235#_c_78_n N_D1_c_170_n 0.0202508f $X=1.6 $Y=1.2 $X2=0 $Y2=0
cc_84 N_A_86_235#_c_98_p N_D1_c_170_n 0.00528418f $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_85 N_A_86_235#_c_79_n N_D1_c_170_n 2.09472e-19 $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_86_235#_c_77_n N_D1_c_171_n 0.00652155f $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_87 N_A_86_235#_c_92_p N_D1_c_171_n 0.0135133f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_88 N_A_86_235#_c_102_p C1 0.0187053f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_89 N_A_86_235#_c_102_p N_C1_c_209_n 6.01575e-19 $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_90 N_A_86_235#_c_98_p N_C1_c_209_n 0.00190299f $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_91 N_A_86_235#_c_105_p N_C1_c_210_n 0.00485598f $X=2.275 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_86_235#_c_102_p N_C1_c_210_n 0.0102875f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_93 N_A_86_235#_c_98_p N_C1_c_210_n 0.0020634f $X=2.3 $Y=0.7 $X2=0 $Y2=0
cc_94 N_A_86_235#_c_102_p B1 0.0162735f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_95 N_A_86_235#_c_102_p N_B1_c_244_n 0.00145768f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_96 N_A_86_235#_c_105_p N_B1_c_245_n 3.01204e-19 $X=2.275 $Y=0.42 $X2=0 $Y2=0
cc_97 N_A_86_235#_c_102_p N_B1_c_245_n 0.0122036f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_98 N_A_86_235#_c_102_p N_A1_c_280_n 0.0145086f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_99 N_A_86_235#_c_113_p N_A1_c_280_n 0.025507f $X=3.23 $Y=0.42 $X2=0 $Y2=0
cc_100 N_A_86_235#_c_102_p N_A1_c_281_n 0.00138694f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_101 N_A_86_235#_M1005_g N_VPWR_c_353_n 0.0153334f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_102 N_A_86_235#_M1012_g N_VPWR_c_353_n 9.85584e-19 $X=0.935 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_86_235#_M1012_g N_VPWR_c_354_n 0.00313429f $X=0.935 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_86_235#_c_76_n N_VPWR_c_354_n 0.020114f $X=1.495 $Y=1.2 $X2=0 $Y2=0
cc_105 N_A_86_235#_c_83_n N_VPWR_c_354_n 0.0751944f $X=1.64 $Y=1.64 $X2=0 $Y2=0
cc_106 N_A_86_235#_c_79_n N_VPWR_c_354_n 0.00586894f $X=1.015 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_86_235#_c_84_n N_VPWR_c_356_n 0.0203609f $X=1.7 $Y=1.66 $X2=0 $Y2=0
cc_108 N_A_86_235#_M1005_g N_VPWR_c_358_n 0.00564095f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_86_235#_M1012_g N_VPWR_c_358_n 0.00537216f $X=0.935 $Y=1.985 $X2=0
+ $Y2=0
cc_110 N_A_86_235#_M1002_s N_VPWR_c_351_n 0.00948669f $X=1.575 $Y=1.485 $X2=0
+ $Y2=0
cc_111 N_A_86_235#_M1005_g N_VPWR_c_351_n 0.00953074f $X=0.505 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_86_235#_M1012_g N_VPWR_c_351_n 0.0107307f $X=0.935 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_86_235#_c_84_n N_VPWR_c_351_n 0.0110914f $X=1.7 $Y=1.66 $X2=0 $Y2=0
cc_114 N_A_86_235#_M1005_g N_X_c_407_n 0.00514976f $X=0.505 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_86_235#_c_74_n N_X_c_407_n 0.0143751f $X=0.585 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_86_235#_M1012_g N_X_c_407_n 0.0174543f $X=0.935 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_86_235#_c_75_n N_X_c_407_n 0.00148958f $X=1.015 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_86_235#_c_76_n N_X_c_407_n 0.0195174f $X=1.495 $Y=1.2 $X2=0 $Y2=0
cc_119 N_A_86_235#_c_77_n N_X_c_407_n 0.00618087f $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_120 N_A_86_235#_c_85_n N_X_c_407_n 0.00490303f $X=1.64 $Y=1.495 $X2=0 $Y2=0
cc_121 N_A_86_235#_c_79_n N_X_c_407_n 0.0328107f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_86_235#_c_77_n N_VGND_M1009_s 0.0034711f $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_123 N_A_86_235#_c_92_p N_VGND_M1009_s 0.00831775f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_124 N_A_86_235#_c_138_p N_VGND_M1009_s 0.00582981f $X=1.705 $Y=0.7 $X2=0
+ $Y2=0
cc_125 N_A_86_235#_c_102_p N_VGND_M1011_d 0.00965831f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_126 N_A_86_235#_c_74_n N_VGND_c_450_n 0.00519652f $X=0.585 $Y=0.995 $X2=0
+ $Y2=0
cc_127 N_A_86_235#_c_75_n N_VGND_c_467_n 0.00460671f $X=1.015 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_86_235#_c_76_n N_VGND_c_467_n 0.0154693f $X=1.495 $Y=1.2 $X2=0 $Y2=0
cc_129 N_A_86_235#_c_77_n N_VGND_c_467_n 0.00605754f $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_130 N_A_86_235#_c_138_p N_VGND_c_467_n 0.0142383f $X=1.705 $Y=0.7 $X2=0 $Y2=0
cc_131 N_A_86_235#_c_79_n N_VGND_c_467_n 0.00565812f $X=1.015 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_86_235#_c_102_p N_VGND_c_451_n 0.0197859f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_133 N_A_86_235#_c_76_n N_VGND_c_454_n 0.00507909f $X=1.495 $Y=1.2 $X2=0 $Y2=0
cc_134 N_A_86_235#_c_92_p N_VGND_c_454_n 0.0184621f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_135 N_A_86_235#_c_138_p N_VGND_c_454_n 0.0174866f $X=1.705 $Y=0.7 $X2=0 $Y2=0
cc_136 N_A_86_235#_c_79_n N_VGND_c_454_n 0.00163441f $X=1.015 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_86_235#_c_92_p N_VGND_c_456_n 0.00259773f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_138 N_A_86_235#_c_105_p N_VGND_c_456_n 0.0141125f $X=2.275 $Y=0.42 $X2=0
+ $Y2=0
cc_139 N_A_86_235#_c_102_p N_VGND_c_456_n 0.00272761f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_140 N_A_86_235#_c_74_n N_VGND_c_458_n 0.00503406f $X=0.585 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_86_235#_c_75_n N_VGND_c_458_n 0.00486043f $X=1.015 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_A_86_235#_c_102_p N_VGND_c_459_n 0.00276179f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_143 N_A_86_235#_c_113_p N_VGND_c_459_n 0.0149005f $X=3.23 $Y=0.42 $X2=0 $Y2=0
cc_144 N_A_86_235#_c_74_n N_VGND_c_460_n 5.05522e-19 $X=0.585 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_86_235#_c_75_n N_VGND_c_460_n 0.00775004f $X=1.015 $Y=0.995 $X2=0
+ $Y2=0
cc_146 N_A_86_235#_M1008_d N_VGND_c_461_n 0.0023722f $X=2.135 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_86_235#_M1001_d N_VGND_c_461_n 0.00579837f $X=3.09 $Y=0.235 $X2=0
+ $Y2=0
cc_148 N_A_86_235#_c_74_n N_VGND_c_461_n 0.00971369f $X=0.585 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_86_235#_c_75_n N_VGND_c_461_n 0.00817678f $X=1.015 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A_86_235#_c_92_p N_VGND_c_461_n 0.00561394f $X=2.18 $Y=0.7 $X2=0 $Y2=0
cc_151 N_A_86_235#_c_138_p N_VGND_c_461_n 0.00110124f $X=1.705 $Y=0.7 $X2=0
+ $Y2=0
cc_152 N_A_86_235#_c_105_p N_VGND_c_461_n 0.00901671f $X=2.275 $Y=0.42 $X2=0
+ $Y2=0
cc_153 N_A_86_235#_c_102_p N_VGND_c_461_n 0.00969987f $X=3.09 $Y=0.7 $X2=0 $Y2=0
cc_154 N_A_86_235#_c_113_p N_VGND_c_461_n 0.00929827f $X=3.23 $Y=0.42 $X2=0
+ $Y2=0
cc_155 N_D1_M1002_g N_C1_M1006_g 0.0488723f $X=2.06 $Y=1.985 $X2=0 $Y2=0
cc_156 D1 N_C1_M1006_g 0.00417035f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_157 N_D1_c_169_n C1 0.00119777f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_158 N_D1_c_170_n C1 0.105292f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_159 N_D1_c_169_n N_C1_c_209_n 0.0488723f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_160 N_D1_c_170_n N_C1_c_209_n 0.00417035f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_161 N_D1_c_171_n N_C1_c_210_n 0.0248182f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_162 N_D1_M1002_g N_VPWR_c_354_n 0.00198883f $X=2.06 $Y=1.985 $X2=0 $Y2=0
cc_163 N_D1_M1002_g N_VPWR_c_356_n 0.0037962f $X=2.06 $Y=1.985 $X2=0 $Y2=0
cc_164 D1 N_VPWR_c_356_n 0.0101792f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_165 N_D1_M1002_g N_VPWR_c_351_n 0.00658426f $X=2.06 $Y=1.985 $X2=0 $Y2=0
cc_166 D1 N_VPWR_c_351_n 0.00989771f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_167 D1 A_427_297# 0.00800054f $X=1.985 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_168 N_D1_c_171_n N_VGND_c_467_n 0.00313316f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_169 N_D1_c_171_n N_VGND_c_455_n 0.00797606f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_170 N_D1_c_171_n N_VGND_c_456_n 0.00351072f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_171 N_D1_c_171_n N_VGND_c_461_n 0.00408313f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_172 N_C1_M1006_g N_B1_M1010_g 0.0349499f $X=2.42 $Y=1.985 $X2=0 $Y2=0
cc_173 N_C1_M1006_g B1 3.6572e-19 $X=2.42 $Y=1.985 $X2=0 $Y2=0
cc_174 C1 B1 0.0577002f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_175 N_C1_c_209_n B1 3.5391e-19 $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_176 C1 N_B1_c_244_n 0.013463f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_177 N_C1_c_209_n N_B1_c_244_n 0.02057f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_178 N_C1_c_210_n N_B1_c_245_n 0.0197813f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_179 N_C1_M1006_g N_VPWR_c_356_n 0.00490733f $X=2.42 $Y=1.985 $X2=0 $Y2=0
cc_180 C1 N_VPWR_c_356_n 0.0113978f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_181 N_C1_M1006_g N_VPWR_c_351_n 0.0084661f $X=2.42 $Y=1.985 $X2=0 $Y2=0
cc_182 C1 N_VPWR_c_351_n 0.0108343f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_183 C1 A_499_297# 0.0140317f $X=2.445 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_184 N_C1_c_210_n N_VGND_c_451_n 0.00169893f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_185 N_C1_c_210_n N_VGND_c_455_n 4.84906e-19 $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_186 N_C1_c_210_n N_VGND_c_456_n 0.00421482f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_187 N_C1_c_210_n N_VGND_c_461_n 0.00582215f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_M1010_g N_A1_M1000_g 0.0267839f $X=2.96 $Y=1.985 $X2=0 $Y2=0
cc_189 B1 N_A1_M1000_g 0.00134529f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_190 B1 N_A1_c_279_n 3.55626e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_191 N_B1_c_244_n N_A1_c_279_n 0.0205668f $X=3.05 $Y=1.16 $X2=0 $Y2=0
cc_192 B1 N_A1_c_280_n 0.0132291f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_193 N_B1_c_244_n N_A1_c_280_n 9.90028e-19 $X=3.05 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B1_c_245_n N_A1_c_280_n 0.00189858f $X=3.05 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B1_c_245_n N_A1_c_281_n 0.0183423f $X=3.05 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B1_M1010_g A1 0.00113211f $X=2.96 $Y=1.985 $X2=0 $Y2=0
cc_197 B1 A1 0.0471306f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_198 N_B1_c_244_n A1 9.87238e-19 $X=3.05 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_M1010_g N_VPWR_c_356_n 0.00585385f $X=2.96 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_M1010_g N_VPWR_c_351_n 0.011422f $X=2.96 $Y=1.985 $X2=0 $Y2=0
cc_201 B1 N_A_607_297#_M1010_d 0.00336012f $X=2.905 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_202 B1 N_A_607_297#_c_430_n 0.00885845f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_203 N_B1_c_244_n N_A_607_297#_c_430_n 9.65699e-19 $X=3.05 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B1_c_245_n N_VGND_c_451_n 0.00321276f $X=3.05 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B1_c_245_n N_VGND_c_459_n 0.00422112f $X=3.05 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B1_c_245_n N_VGND_c_461_n 0.00598811f $X=3.05 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_M1000_g N_A2_M1007_g 0.0335504f $X=3.5 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A1_c_280_n N_A2_c_323_n 5.37878e-19 $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_209 A1 N_A2_c_323_n 0.00210719f $X=3.45 $Y=1.19 $X2=0 $Y2=0
cc_210 N_A1_M1000_g N_A2_c_324_n 5.93261e-19 $X=3.5 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A1_c_279_n N_A2_c_324_n 0.00114342f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A1_c_280_n N_A2_c_324_n 0.0180047f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_213 A1 N_A2_c_324_n 0.0391448f $X=3.45 $Y=1.19 $X2=0 $Y2=0
cc_214 N_A1_c_279_n N_A2_c_325_n 0.0222729f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A1_c_280_n N_A2_c_325_n 0.0194258f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A1_c_281_n N_A2_c_325_n 0.0254791f $X=3.59 $Y=0.98 $X2=0 $Y2=0
cc_217 A1 N_VPWR_M1000_d 0.00404968f $X=3.45 $Y=1.19 $X2=0 $Y2=0
cc_218 N_A1_M1000_g N_VPWR_c_355_n 0.00326685f $X=3.5 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A1_M1000_g N_VPWR_c_356_n 0.00425094f $X=3.5 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A1_M1000_g N_VPWR_c_351_n 0.00616819f $X=3.5 $Y=1.985 $X2=0 $Y2=0
cc_221 A1 N_A_607_297#_M1010_d 0.00233256f $X=3.45 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_222 N_A1_M1000_g N_A_607_297#_c_428_n 0.0110046f $X=3.5 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A1_c_279_n N_A_607_297#_c_428_n 4.81123e-19 $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_224 A1 N_A_607_297#_c_428_n 0.0224336f $X=3.45 $Y=1.19 $X2=0 $Y2=0
cc_225 N_A1_c_280_n N_VGND_c_459_n 0.0245745f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A1_c_281_n N_VGND_c_459_n 0.0048249f $X=3.59 $Y=0.98 $X2=0 $Y2=0
cc_227 N_A1_c_280_n N_VGND_c_461_n 0.0180216f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A1_c_281_n N_VGND_c_461_n 0.00863638f $X=3.59 $Y=0.98 $X2=0 $Y2=0
cc_229 N_A1_c_280_n A_715_47# 0.0103245f $X=3.59 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_230 N_A2_M1007_g N_VPWR_c_355_n 0.00438997f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A2_M1007_g N_VPWR_c_359_n 0.00415375f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A2_M1007_g N_VPWR_c_351_n 0.0069265f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A2_c_324_n N_A_607_297#_M1007_d 0.00343567f $X=4.13 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A2_M1007_g N_A_607_297#_c_428_n 0.0166903f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A2_c_323_n N_A_607_297#_c_428_n 5.21484e-19 $X=4.13 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A2_c_324_n N_A_607_297#_c_428_n 0.0413838f $X=4.13 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A2_c_323_n N_VGND_c_453_n 9.87152e-19 $X=4.13 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A2_c_324_n N_VGND_c_453_n 0.028757f $X=4.13 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A2_c_325_n N_VGND_c_453_n 0.0155601f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_325_n N_VGND_c_459_n 0.00541287f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A2_c_325_n N_VGND_c_461_n 0.0109563f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_242 N_VPWR_c_351_n N_X_M1005_s 0.00321211f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_243 N_VPWR_c_358_n N_X_c_407_n 0.0115784f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_351_n N_X_c_407_n 0.0105011f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_245 N_VPWR_c_351_n A_427_297# 0.0049004f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_246 N_VPWR_c_351_n A_499_297# 0.00848418f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_247 N_VPWR_c_351_n N_A_607_297#_M1010_d 0.00445292f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_248 N_VPWR_c_351_n N_A_607_297#_M1007_d 0.00213418f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_356_n N_A_607_297#_c_442_n 0.0208881f $X=3.59 $Y=2.72 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_351_n N_A_607_297#_c_442_n 0.0125525f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_251 N_VPWR_M1000_d N_A_607_297#_c_428_n 0.00962523f $X=3.575 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_355_n N_A_607_297#_c_428_n 0.021058f $X=3.755 $Y=2.34 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_356_n N_A_607_297#_c_428_n 0.00282957f $X=3.59 $Y=2.72 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_359_n N_A_607_297#_c_428_n 0.0299351f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_351_n N_A_607_297#_c_428_n 0.0261948f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_256 N_X_c_407_n N_VGND_c_450_n 0.048663f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_257 N_X_c_407_n N_VGND_c_458_n 0.017735f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_258 N_X_M1004_d N_VGND_c_461_n 0.00379452f $X=0.66 $Y=0.235 $X2=0 $Y2=0
cc_259 N_X_c_407_n N_VGND_c_461_n 0.010772f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_260 N_VGND_c_461_n A_715_47# 0.00315916f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__sdfrtp_1.spice
* Created: Thu Aug 27 14:46:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfrtp_1.spice.pex"
.subckt sky130_fd_sc_hd__sdfrtp_1  VNB VPB CLK D SCE SCD RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* SCD	SCD
* SCE	SCE
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1032 N_VGND_M1032_d N_CLK_M1032_g N_A_27_47#_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1020 N_A_193_47#_M1020_d N_A_27_47#_M1020_g N_VGND_M1032_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_SCE_M1022_g N_A_299_66#_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_569_119# N_A_299_66#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1016 N_A_620_389#_M1016_d N_D_M1016_g A_569_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.110275 AS=0.0441 PD=1.065 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 A_817_66# N_SCE_M1015_g N_A_620_389#_M1016_d VNB NSHORT L=0.5 W=0.42
+ AD=0.0441 AS=0.110275 PD=0.63 PS=1.065 NRD=14.28 NRS=59.292 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1027 N_VGND_M1027_d N_SCD_M1027_g A_817_66# VNB NSHORT L=0.18 W=0.42 AD=0.1176
+ AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.33333 SA=90001.2 SB=90000.2
+ A=0.0756 P=1.2 MULT=1
MM1021 N_A_1079_413#_M1021_d N_A_27_47#_M1021_g N_A_620_389#_M1021_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.063 AS=0.0936 PD=0.71 PS=1.24 NRD=24.996 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75004.9 A=0.054 P=1.02 MULT=1
MM1018 A_1187_47# N_A_193_47#_M1018_g N_A_1079_413#_M1021_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0700615 AS=0.063 PD=0.738462 PS=0.71 NRD=46.536 NRS=0 M=1 R=2.4
+ SA=75000.7 SB=75004.4 A=0.054 P=1.02 MULT=1
MM1009 A_1293_47# N_A_1245_303#_M1009_g A_1187_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0817385 PD=0.63 PS=0.861538 NRD=14.28 NRS=39.888 M=1 R=2.8
+ SA=75001.1 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_RESET_B_M1012_g A_1293_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.106664 AS=0.0441 PD=0.911321 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1034 N_A_1245_303#_M1034_d N_A_1079_413#_M1034_g N_VGND_M1012_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.11968 AS=0.162536 PD=1.2352 PS=1.38868 NRD=0 NRS=21.552 M=1
+ R=4.26667 SA=75001.4 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_1592_47#_M1013_d N_A_193_47#_M1013_g N_A_1245_303#_M1034_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0711 AS=0.06732 PD=0.755 PS=0.6948 NRD=23.328 NRS=16.656
+ M=1 R=2.4 SA=75002.7 SB=75002.4 A=0.054 P=1.02 MULT=1
MM1010 A_1701_47# N_A_27_47#_M1010_g N_A_1592_47#_M1013_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0618923 AS=0.0711 PD=0.692308 PS=0.755 NRD=38.964 NRS=14.988 M=1
+ R=2.4 SA=75003.3 SB=75001.8 A=0.054 P=1.02 MULT=1
MM1024 N_VGND_M1024_d N_A_1767_21#_M1024_g A_1701_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.12495 AS=0.0722077 PD=1.015 PS=0.807692 NRD=12.852 NRS=33.396 M=1 R=2.8
+ SA=75003.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 A_1946_47# N_RESET_B_M1000_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.05145 AS=0.12495 PD=0.665 PS=1.015 NRD=19.284 NRS=77.136 M=1 R=2.8
+ SA=75004 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_1767_21#_M1014_d N_A_1592_47#_M1014_g A_1946_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.05145 PD=1.4 PS=0.665 NRD=0 NRS=19.284 M=1 R=2.8
+ SA=75004.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_Q_M1017_d N_A_1767_21#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1026 N_VPWR_M1026_d N_CLK_M1026_g N_A_27_47#_M1026_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1425 AS=0.26 PD=1.285 PS=2.52 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1035 N_A_193_47#_M1035_d N_A_27_47#_M1035_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.1425 PD=2.53 PS=1.285 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_SCE_M1005_g N_A_299_66#_M1005_s VPB PHIGHVT L=0.15
+ W=0.54 AD=0.0729 AS=0.189 PD=0.81 PS=1.78 NRD=0 NRS=0 M=1 R=3.6 SA=75000.3
+ SB=75002.3 A=0.081 P=1.38 MULT=1
MM1002 A_538_389# N_SCE_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.54
+ AD=0.0702 AS=0.0729 PD=0.8 PS=0.81 NRD=27.3436 NRS=0 M=1 R=3.6 SA=75000.7
+ SB=75001.8 A=0.081 P=1.38 MULT=1
MM1023 N_A_620_389#_M1023_d N_D_M1023_g A_538_389# VPB PHIGHVT L=0.15 W=0.54
+ AD=0.1755 AS=0.0702 PD=1.19 PS=0.8 NRD=111.266 NRS=27.3436 M=1 R=3.6
+ SA=75001.1 SB=75001.4 A=0.081 P=1.38 MULT=1
MM1003 A_780_389# N_A_299_66#_M1003_g N_A_620_389#_M1023_d VPB PHIGHVT L=0.15
+ W=0.54 AD=0.0756 AS=0.1755 PD=0.82 PS=1.19 NRD=31.0078 NRS=23.6991 M=1 R=3.6
+ SA=75001.9 SB=75000.6 A=0.081 P=1.38 MULT=1
MM1031 N_VPWR_M1031_d N_SCD_M1031_g A_780_389# VPB PHIGHVT L=0.15 W=0.54
+ AD=0.1512 AS=0.0756 PD=1.64 PS=0.82 NRD=0 NRS=31.0078 M=1 R=3.6 SA=75002.3
+ SB=75000.2 A=0.081 P=1.38 MULT=1
MM1006 N_A_1079_413#_M1006_d N_A_193_47#_M1006_g N_A_620_389#_M1006_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0861 AS=0.1533 PD=0.83 PS=1.57 NRD=63.3158 NRS=0
+ M=1 R=2.8 SA=75000.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_1191_413#_M1004_d N_A_27_47#_M1004_g N_A_1079_413#_M1006_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0567 AS=0.0861 PD=0.69 PS=0.83 NRD=0 NRS=0 M=1
+ R=2.8 SA=75000.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1033 N_VPWR_M1033_d N_A_1245_303#_M1033_g N_A_1191_413#_M1004_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1007 AS=0.0567 PD=0.94 PS=0.69 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75001.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1030 N_A_1191_413#_M1030_d N_RESET_B_M1030_g N_VPWR_M1033_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1007 PD=1.36 PS=0.94 NRD=0 NRS=39.8531 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_1245_303#_M1019_d N_A_1079_413#_M1019_g N_VPWR_M1019_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.161 AS=0.2184 PD=1.55333 PS=2.2 NRD=7.0329 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_1592_47#_M1001_d N_A_27_47#_M1001_g N_A_1245_303#_M1019_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0805 PD=0.7 PS=0.776667 NRD=2.3443 NRS=7.0329 M=1
+ R=2.8 SA=75000.7 SB=75002 A=0.063 P=1.14 MULT=1
MM1028 A_1758_413# N_A_193_47#_M1028_g N_A_1592_47#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0546 AS=0.0588 PD=0.68 PS=0.7 NRD=35.1645 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_1767_21#_M1025_g A_1758_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0546 PD=0.8 PS=0.68 NRD=49.25 NRS=35.1645 M=1 R=2.8 SA=75001.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_A_1767_21#_M1011_d N_RESET_B_M1011_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0798 PD=0.69 PS=0.8 NRD=0 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_VPWR_M1029_d N_A_1592_47#_M1029_g N_A_1767_21#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_Q_M1007_d N_A_1767_21#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX36_noxref VNB VPB NWDIODE A=18.7752 P=27.21
c_127 VNB 0 1.58318e-19 $X=0.215 $Y=-0.01
c_256 VPB 0 3.75206e-19 $X=0.17 $Y=2.64
*
.include "sky130_fd_sc_hd__sdfrtp_1.spice.SKY130_FD_SC_HD__SDFRTP_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__mux2i_4.pex.spice
* Created: Thu Aug 27 14:28:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A0 1 3 6 8 10 13 15 17 20 22 24 27 29 30 40
+ 42
c64 30 0 1.39126e-19 $X=1.155 $Y=1.19
r65 39 40 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r66 38 42 3.34494 $w=3.3e-07 $l=8e-08 $layer=LI1_cond $X=0.985 $Y=1.16 $X2=0.905
+ $Y2=1.16
r67 37 39 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.985 $Y=1.16
+ $X2=1.31 $Y2=1.16
r68 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.985
+ $Y=1.16 $X2=0.985 $Y2=1.16
r69 35 37 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.985 $Y2=1.16
r70 33 35 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r71 30 38 7.56934 $w=2.74e-07 $l=1.7e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=0.985 $Y2=1.16
r72 29 42 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.905 $Y2=1.16
r73 25 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r74 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r75 22 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r76 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r77 18 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r78 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r79 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r80 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r81 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r82 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r83 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r84 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r85 4 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r86 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r87 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r88 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47
r71 45 47 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.26 $Y=1.16
+ $X2=3.41 $Y2=1.16
r72 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.26
+ $Y=1.16 $X2=3.26 $Y2=1.16
r73 43 45 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.26 $Y2=1.16
r74 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r75 40 42 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.24 $Y=1.16
+ $X2=2.57 $Y2=1.16
r76 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r77 37 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.15 $Y=1.16 $X2=2.24
+ $Y2=1.16
r78 32 46 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.26 $Y2=1.16
r79 31 46 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=3.26 $Y2=1.16
r80 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.995 $Y2=1.16
r81 30 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.24 $Y2=1.16
r82 29 41 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=1.16
+ $X2=2.24 $Y2=1.16
r83 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r85 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r87 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r89 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r91 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r93 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r95 4 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r97 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%S 1 3 6 8 10 13 15 17 20 22 24 27 31 34 36
+ 40 41 43 44 45 46 47 64 67 69
r134 62 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.52 $Y=1.16 $X2=5.61
+ $Y2=1.16
r135 62 63 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.52
+ $Y=1.16 $X2=5.52 $Y2=1.16
r136 60 62 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=5.19 $Y=1.16
+ $X2=5.52 $Y2=1.16
r137 59 60 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16
+ $X2=5.19 $Y2=1.16
r138 58 59 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.35 $Y=1.16
+ $X2=4.77 $Y2=1.16
r139 55 58 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.16 $Y=1.16
+ $X2=4.35 $Y2=1.16
r140 55 56 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.16
+ $Y=1.16 $X2=4.16 $Y2=1.16
r141 47 86 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.845 $Y=1.19
+ $X2=5.845 $Y2=1.51
r142 47 69 0.521925 $w=1.68e-07 $l=8e-09 $layer=LI1_cond $X=5.845 $Y=1.19
+ $X2=5.845 $Y2=1.182
r143 47 69 1.87607 $w=2.13e-07 $l=3.5e-08 $layer=LI1_cond $X=5.725 $Y=1.182
+ $X2=5.76 $Y2=1.182
r144 47 63 10.9884 $w=2.13e-07 $l=2.05e-07 $layer=LI1_cond $X=5.725 $Y=1.182
+ $X2=5.52 $Y2=1.182
r145 46 63 10.9884 $w=2.13e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=1.182
+ $X2=5.52 $Y2=1.182
r146 45 46 24.6569 $w=2.13e-07 $l=4.6e-07 $layer=LI1_cond $X=4.855 $Y=1.182
+ $X2=5.315 $Y2=1.182
r147 44 45 24.6569 $w=2.13e-07 $l=4.6e-07 $layer=LI1_cond $X=4.395 $Y=1.182
+ $X2=4.855 $Y2=1.182
r148 44 56 12.5965 $w=2.13e-07 $l=2.35e-07 $layer=LI1_cond $X=4.395 $Y=1.182
+ $X2=4.16 $Y2=1.182
r149 43 56 12.0604 $w=2.13e-07 $l=2.25e-07 $layer=LI1_cond $X=3.935 $Y=1.182
+ $X2=4.16 $Y2=1.182
r150 41 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=1.16
+ $X2=7.765 $Y2=1.325
r151 41 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=1.16
+ $X2=7.765 $Y2=0.995
r152 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.765
+ $Y=1.16 $X2=7.765 $Y2=1.16
r153 38 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.765 $Y=1.425
+ $X2=7.765 $Y2=1.16
r154 37 86 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=1.51
+ $X2=5.845 $Y2=1.51
r155 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.68 $Y=1.51
+ $X2=7.765 $Y2=1.425
r156 36 37 114.171 $w=1.68e-07 $l=1.75e-06 $layer=LI1_cond $X=7.68 $Y=1.51
+ $X2=5.93 $Y2=1.51
r157 34 68 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.81 $Y=1.985
+ $X2=7.81 $Y2=1.325
r158 31 67 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.81 $Y=0.56
+ $X2=7.81 $Y2=0.995
r159 25 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.16
r160 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.985
r161 22 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r162 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r163 18 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.16
r164 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.985
r165 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r166 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r167 11 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.16
r168 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.985
r169 8 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.16
r170 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r171 4 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.16
r172 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.985
r173 1 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.16
r174 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A_1191_21# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 35 41 42 43 46 48 50 54 55 61
c111 21 0 3.76464e-19 $X=6.87 $Y=0.995
r112 58 59 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.87 $Y2=1.16
r113 56 58 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.03 $Y=1.16
+ $X2=6.45 $Y2=1.16
r114 52 54 4.18896 $w=2.17e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.107 $Y=0.825
+ $X2=8.065 $Y2=0.74
r115 52 55 61.4753 $w=1.73e-07 $l=9.7e-07 $layer=LI1_cond $X=8.107 $Y=0.825
+ $X2=8.107 $Y2=1.795
r116 48 55 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=8.065 $Y=1.925
+ $X2=8.065 $Y2=1.795
r117 48 50 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=8.065 $Y=1.925
+ $X2=8.065 $Y2=1.96
r118 44 54 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=0.655
+ $X2=8.065 $Y2=0.74
r119 44 46 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=8.065 $Y=0.655
+ $X2=8.065 $Y2=0.42
r120 42 54 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.935 $Y=0.74
+ $X2=8.065 $Y2=0.74
r121 42 43 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.935 $Y=0.74
+ $X2=7.51 $Y2=0.74
r122 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.425 $Y=0.825
+ $X2=7.51 $Y2=0.74
r123 40 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.425 $Y=0.825
+ $X2=7.425 $Y2=1.075
r124 38 61 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.255 $Y=1.16
+ $X2=7.345 $Y2=1.16
r125 38 59 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=7.255 $Y=1.16
+ $X2=6.87 $Y2=1.16
r126 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.255
+ $Y=1.16 $X2=7.255 $Y2=1.16
r127 35 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.34 $Y=1.16
+ $X2=7.425 $Y2=1.075
r128 35 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=1.16
+ $X2=7.255 $Y2=1.16
r129 31 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.325
+ $X2=7.345 $Y2=1.16
r130 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.345 $Y=1.325
+ $X2=7.345 $Y2=1.985
r131 28 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=0.995
+ $X2=7.345 $Y2=1.16
r132 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.345 $Y=0.995
+ $X2=7.345 $Y2=0.56
r133 24 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.16
r134 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.985
r135 21 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=1.16
r136 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=0.56
r137 17 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r138 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r139 14 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r140 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r141 10 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r142 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r143 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r144 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
r145 2 50 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=1.96
r146 1 46 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%Y 1 2 3 4 5 6 7 8 9 10 39 41 44 45 46 47 48
+ 56 67 77
r71 75 77 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=2.34
+ $X2=3.62 $Y2=2.34
r72 73 75 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.94 $Y=2.34
+ $X2=2.78 $Y2=2.34
r73 70 73 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=2.34 $X2=1.94
+ $Y2=2.34
r74 56 67 2.30489 $w=2.23e-07 $l=4.5e-08 $layer=LI1_cond $X=0.207 $Y=2.255
+ $X2=0.207 $Y2=2.21
r75 48 56 3.00067 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.207 $Y=2.34
+ $X2=0.207 $Y2=2.255
r76 48 70 41.6297 $w=2.08e-07 $l=7.8e-07 $layer=LI1_cond $X=0.32 $Y=2.34 $X2=1.1
+ $Y2=2.34
r77 48 67 1.02439 $w=2.23e-07 $l=2e-08 $layer=LI1_cond $X=0.207 $Y=2.19
+ $X2=0.207 $Y2=2.21
r78 47 48 16.3903 $w=2.23e-07 $l=3.2e-07 $layer=LI1_cond $X=0.207 $Y=1.87
+ $X2=0.207 $Y2=2.19
r79 46 47 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.53
+ $X2=0.207 $Y2=1.87
r80 45 46 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r81 44 45 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=0.85
+ $X2=0.207 $Y2=1.19
r82 41 44 18.6952 $w=2.23e-07 $l=3.65e-07 $layer=LI1_cond $X=0.207 $Y=0.485
+ $X2=0.207 $Y2=0.85
r83 41 43 3.00067 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.207 $Y=0.485
+ $X2=0.207 $Y2=0.4
r84 37 39 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.4 $X2=3.62
+ $Y2=0.4
r85 35 37 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.94 $Y=0.4 $X2=2.78
+ $Y2=0.4
r86 33 35 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=0.4 $X2=1.94
+ $Y2=0.4
r87 31 43 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.32 $Y=0.4
+ $X2=0.207 $Y2=0.4
r88 31 33 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.32 $Y=0.4 $X2=1.1
+ $Y2=0.4
r89 10 77 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2.34
r90 9 75 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.34
r91 8 73 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.34
r92 7 70 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r93 6 48 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r94 5 39 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.4
r95 4 37 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.4
r96 3 35 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.4
r97 2 33 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r98 1 43 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A_109_297# 1 2 3 4 21
r42 19 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=1.66 $X2=5.4
+ $Y2=1.66
r43 17 19 198.332 $w=1.68e-07 $l=3.04e-06 $layer=LI1_cond $X=1.52 $Y=1.66
+ $X2=4.56 $Y2=1.66
r44 14 17 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.68 $Y=1.66
+ $X2=1.52 $Y2=1.66
r45 4 21 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.66
r46 3 19 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.66
r47 2 17 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r48 1 14 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A_445_297# 1 2 3 4 13 21 23 25 27 30
r54 25 32 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.08 $Y=2.085
+ $X2=7.08 $Y2=1.94
r55 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.08 $Y=2.085
+ $X2=7.08 $Y2=2.3
r56 24 30 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=6.325 $Y=2
+ $X2=6.24 $Y2=1.94
r57 23 32 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=6.995 $Y=2
+ $X2=7.08 $Y2=1.94
r58 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.995 $Y=2 $X2=6.325
+ $Y2=2
r59 19 30 1.34256 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.24 $Y=2.085
+ $X2=6.24 $Y2=1.94
r60 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.24 $Y=2.085
+ $X2=6.24 $Y2=2.3
r61 15 18 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=2 $X2=3.2
+ $Y2=2
r62 13 30 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=6.155 $Y=2
+ $X2=6.24 $Y2=1.94
r63 13 18 192.786 $w=1.68e-07 $l=2.955e-06 $layer=LI1_cond $X=6.155 $Y=2 $X2=3.2
+ $Y2=2
r64 4 32 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=1.96
r65 4 27 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=2.3
r66 3 30 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.96
r67 3 21 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=2.3
r68 2 18 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2
r69 1 15 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 38 39 40 49
+ 54 59 66 67 70 73 76 79
r116 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r117 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r118 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r119 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r120 67 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r122 64 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=2.72
+ $X2=7.6 $Y2=2.72
r123 64 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.765 $Y=2.72
+ $X2=8.05 $Y2=2.72
r124 63 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r125 63 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r126 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r127 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=2.72
+ $X2=6.66 $Y2=2.72
r128 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.825 $Y=2.72
+ $X2=7.13 $Y2=2.72
r129 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=2.72
+ $X2=7.6 $Y2=2.72
r130 59 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.435 $Y=2.72
+ $X2=7.13 $Y2=2.72
r131 58 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r132 58 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r133 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r134 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=2.72
+ $X2=5.82 $Y2=2.72
r135 55 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.985 $Y=2.72
+ $X2=6.21 $Y2=2.72
r136 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=2.72
+ $X2=6.66 $Y2=2.72
r137 54 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.495 $Y=2.72
+ $X2=6.21 $Y2=2.72
r138 53 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r139 53 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r140 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r141 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=2.72
+ $X2=4.98 $Y2=2.72
r142 50 52 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.145 $Y=2.72
+ $X2=5.29 $Y2=2.72
r143 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=2.72
+ $X2=5.82 $Y2=2.72
r144 49 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.655 $Y=2.72
+ $X2=5.29 $Y2=2.72
r145 48 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 47 48 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r147 43 47 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r148 40 48 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r149 40 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r150 38 47 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=3.91 $Y2=2.72
r151 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=4.14 $Y2=2.72
r152 34 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=2.635 $X2=7.6
+ $Y2=2.72
r153 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.6 $Y=2.635
+ $X2=7.6 $Y2=2.34
r154 30 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2.72
r155 30 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2.34
r156 26 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r157 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.34
r158 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r159 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.34
r160 21 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.14 $Y2=2.72
r161 20 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=2.72
+ $X2=4.98 $Y2=2.72
r162 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.815 $Y=2.72
+ $X2=4.305 $Y2=2.72
r163 16 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.72
r164 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.34
r165 5 36 600 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=7.42
+ $Y=1.485 $X2=7.6 $Y2=2.34
r166 4 32 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=2.34
r167 3 28 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2.34
r168 2 24 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2.34
r169 1 18 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.485 $X2=4.14 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A_109_47# 1 2 3 4 19 21 24 28 29 35 39 40 45
c95 45 0 1.56989e-19 $X=6.45 $Y=0.825
c96 35 0 1.39226e-19 $X=6.235 $Y=0.85
c97 24 0 8.02492e-20 $X=7.08 $Y=0.675
r98 44 45 11.4037 $w=2.18e-07 $l=2.13e-07 $layer=LI1_cond $X=6.237 $Y=0.825
+ $X2=6.45 $Y2=0.825
r99 39 40 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0.795
+ $X2=1.355 $Y2=0.795
r100 36 44 0.104768 $w=2.18e-07 $l=2e-09 $layer=LI1_cond $X=6.235 $Y=0.825
+ $X2=6.237 $Y2=0.825
r101 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.235 $Y=0.85
+ $X2=6.235 $Y2=0.85
r102 31 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=0.85
+ $X2=1.615 $Y2=0.85
r103 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=0.85
+ $X2=1.615 $Y2=0.85
r104 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.09 $Y=0.85
+ $X2=6.235 $Y2=0.85
r105 28 29 5.3589 $w=1.4e-07 $l=4.33e-06 $layer=MET1_cond $X=6.09 $Y=0.85
+ $X2=1.76 $Y2=0.85
r106 24 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.08 $Y=0.675
+ $X2=7.08 $Y2=0.81
r107 21 26 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=0.81
+ $X2=7.08 $Y2=0.81
r108 21 45 31.8134 $w=1.88e-07 $l=5.45e-07 $layer=LI1_cond $X=6.995 $Y=0.81
+ $X2=6.45 $Y2=0.81
r109 17 44 2.10765 $w=1.75e-07 $l=1.1e-07 $layer=LI1_cond $X=6.237 $Y=0.715
+ $X2=6.237 $Y2=0.825
r110 17 19 18.6961 $w=1.73e-07 $l=2.95e-07 $layer=LI1_cond $X=6.237 $Y=0.715
+ $X2=6.237 $Y2=0.42
r111 15 40 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=1.355 $Y2=0.74
r112 4 24 182 $w=1.7e-07 $l=5.02991e-07 $layer=licon1_NDIFF $count=1 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.675
r113 3 19 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.42
r114 2 39 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.74
r115 1 15 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%A_445_47# 1 2 3 4 13 21 23 27 29
r49 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.4 $Y=0.655
+ $X2=5.4 $Y2=0.42
r50 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=0.74
+ $X2=4.56 $Y2=0.74
r51 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.315 $Y=0.74
+ $X2=5.4 $Y2=0.655
r52 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.315 $Y=0.74
+ $X2=4.645 $Y2=0.74
r53 19 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.655
+ $X2=4.56 $Y2=0.74
r54 19 21 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.56 $Y=0.655
+ $X2=4.56 $Y2=0.42
r55 15 18 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.74 $X2=3.2
+ $Y2=0.74
r56 13 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.74
+ $X2=4.56 $Y2=0.74
r57 13 18 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=4.475 $Y=0.74
+ $X2=3.2 $Y2=0.74
r58 4 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.42
r59 3 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.42
r60 2 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.74
r61 1 15 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_4%VGND 1 2 3 4 5 18 20 24 28 32 36 38 39 40 49
+ 54 59 66 67 70 73 76 79
r128 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r129 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r130 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r131 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r132 67 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=7.59
+ $Y2=0
r133 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r134 64 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0 $X2=7.6
+ $Y2=0
r135 64 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=8.05 $Y2=0
r136 63 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r137 63 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=6.67
+ $Y2=0
r138 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r139 60 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.795 $Y=0 $X2=6.67
+ $Y2=0
r140 60 62 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.795 $Y=0
+ $X2=7.13 $Y2=0
r141 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=0 $X2=7.6
+ $Y2=0
r142 59 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.435 $Y=0
+ $X2=7.13 $Y2=0
r143 58 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r144 58 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r145 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r146 55 73 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=5.98 $Y=0 $X2=5.817
+ $Y2=0
r147 55 57 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.98 $Y=0 $X2=6.21
+ $Y2=0
r148 54 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=0 $X2=6.67
+ $Y2=0
r149 54 57 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.21 $Y2=0
r150 53 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r151 53 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r152 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r153 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=4.98
+ $Y2=0
r154 50 52 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.145 $Y=0
+ $X2=5.29 $Y2=0
r155 49 73 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.817
+ $Y2=0
r156 49 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.655 $Y=0
+ $X2=5.29 $Y2=0
r157 48 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r158 47 48 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r159 43 47 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=3.91
+ $Y2=0
r160 40 48 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=3.91
+ $Y2=0
r161 40 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r162 38 47 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.91
+ $Y2=0
r163 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r164 34 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=0.085 $X2=7.6
+ $Y2=0
r165 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0.38
r166 30 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.67 $Y=0.085
+ $X2=6.67 $Y2=0
r167 30 32 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.67 $Y=0.085
+ $X2=6.67 $Y2=0.38
r168 26 73 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.817 $Y=0.085
+ $X2=5.817 $Y2=0
r169 26 28 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=5.817 $Y=0.085
+ $X2=5.817 $Y2=0.425
r170 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r171 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.38
r172 21 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r173 20 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.98
+ $Y2=0
r174 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.815 $Y=0
+ $X2=4.305 $Y2=0
r175 16 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r176 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.38
r177 5 36 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=7.42
+ $Y=0.235 $X2=7.6 $Y2=0.38
r178 4 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.38
r179 3 28 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.425
r180 2 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.38
r181 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o2111ai_4.pex.spice
* Created: Tue Sep  1 19:20:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2111AI_4%D1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 45
r62 43 45 26.4478 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=1.205
+ $X2=1.73 $Y2=1.205
r63 41 43 40.8738 $w=3.6e-07 $l=2.55e-07 $layer=POLY_cond $X=1.31 $Y=1.205
+ $X2=1.565 $Y2=1.205
r64 40 41 67.3216 $w=3.6e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.205
+ $X2=1.31 $Y2=1.205
r65 38 40 28.8521 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.71 $Y=1.205
+ $X2=0.89 $Y2=1.205
r66 35 38 38.4695 $w=3.6e-07 $l=2.4e-07 $layer=POLY_cond $X=0.47 $Y=1.205
+ $X2=0.71 $Y2=1.205
r67 31 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.16 $X2=1.565 $Y2=1.16
r68 30 31 17.5001 $w=2.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.155 $Y=1.21
+ $X2=1.565 $Y2=1.21
r69 29 30 19.6342 $w=2.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.21
+ $X2=1.155 $Y2=1.21
r70 29 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.16 $X2=0.71 $Y2=1.16
r71 26 45 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.73 $Y=1.385
+ $X2=1.73 $Y2=1.205
r72 26 28 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.73 $Y=1.385 $X2=1.73
+ $Y2=1.985
r73 22 45 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.205
r74 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r75 19 41 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.31 $Y=1.385
+ $X2=1.31 $Y2=1.205
r76 19 21 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.31 $Y=1.385 $X2=1.31
+ $Y2=1.985
r77 15 41 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.205
r78 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r79 12 40 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.89 $Y=1.385
+ $X2=0.89 $Y2=1.205
r80 12 14 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.89 $Y=1.385 $X2=0.89
+ $Y2=1.985
r81 8 40 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.205
r82 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r83 5 35 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.47 $Y=1.385
+ $X2=0.47 $Y2=1.205
r84 5 7 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.47 $Y=1.385 $X2=0.47
+ $Y2=1.985
r85 1 35 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.205
r86 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%C1 3 7 11 15 19 23 27 31 33 34 35 36 54
c74 36 0 1.77425e-19 $X=3.455 $Y=1.19
c75 3 0 7.52102e-20 $X=2.15 $Y=0.56
r76 52 54 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.26 $Y=1.16
+ $X2=3.41 $Y2=1.16
r77 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.16 $X2=3.26 $Y2=1.16
r78 50 52 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.26 $Y2=1.16
r79 48 50 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=2.92 $Y=1.16 $X2=2.99
+ $Y2=1.16
r80 46 48 77.7608 $w=2.7e-07 $l=3.5e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.92 $Y2=1.16
r81 44 46 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.24 $Y=1.16
+ $X2=2.57 $Y2=1.16
r82 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r83 41 44 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.15 $Y=1.16 $X2=2.24
+ $Y2=1.16
r84 36 53 8.3232 $w=2.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.455 $Y=1.21
+ $X2=3.26 $Y2=1.21
r85 35 53 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.92 $Y=1.21
+ $X2=3.26 $Y2=1.21
r86 35 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.92
+ $Y=1.16 $X2=2.92 $Y2=1.16
r87 34 35 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.535 $Y=1.21
+ $X2=2.92 $Y2=1.21
r88 34 45 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.535 $Y=1.21
+ $X2=2.24 $Y2=1.21
r89 33 45 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=1.21
+ $X2=2.24 $Y2=1.21
r90 29 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r91 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r92 25 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r93 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r94 21 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r95 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r96 17 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r97 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r98 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r99 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r100 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r101 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r102 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r103 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r104 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r105 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%B1 3 7 11 15 19 21 23 26 28 29 30 32 33 34
+ 35 36
c80 28 0 1.23236e-19 $X=5.535 $Y=1.035
c81 3 0 1.77425e-19 $X=4.035 $Y=1.985
r82 55 56 17.7579 $w=2.85e-07 $l=1.05e-07 $layer=POLY_cond $X=5.19 $Y=1.127
+ $X2=5.295 $Y2=1.127
r83 53 55 43.1263 $w=2.85e-07 $l=2.55e-07 $layer=POLY_cond $X=4.935 $Y=1.127
+ $X2=5.19 $Y2=1.127
r84 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.16 $X2=4.935 $Y2=1.16
r85 51 53 10.1474 $w=2.85e-07 $l=6e-08 $layer=POLY_cond $X=4.875 $Y=1.127
+ $X2=4.935 $Y2=1.127
r86 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.595
+ $Y=1.16 $X2=4.595 $Y2=1.16
r87 46 48 23.6772 $w=2.85e-07 $l=1.4e-07 $layer=POLY_cond $X=4.455 $Y=1.127
+ $X2=4.595 $Y2=1.127
r88 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.255
+ $Y=1.16 $X2=4.255 $Y2=1.16
r89 41 43 37.207 $w=2.85e-07 $l=2.2e-07 $layer=POLY_cond $X=4.035 $Y=1.127
+ $X2=4.255 $Y2=1.127
r90 36 54 15.1525 $w=2.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.29 $Y=1.21
+ $X2=4.935 $Y2=1.21
r91 35 54 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.83 $Y=1.21
+ $X2=4.935 $Y2=1.21
r92 35 49 10.0305 $w=2.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.83 $Y=1.21
+ $X2=4.595 $Y2=1.21
r93 34 49 9.60369 $w=2.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.37 $Y=1.21
+ $X2=4.595 $Y2=1.21
r94 34 44 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.37 $Y=1.21
+ $X2=4.255 $Y2=1.21
r95 33 44 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.91 $Y=1.21
+ $X2=4.255 $Y2=1.21
r96 30 32 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.61 $Y=0.96 $X2=5.61
+ $Y2=0.56
r97 29 56 23.4449 $w=2.85e-07 $l=1.23952e-07 $layer=POLY_cond $X=5.37 $Y=1.035
+ $X2=5.295 $Y2=1.127
r98 28 30 31.2341 $w=1.29e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.535 $Y=1.035
+ $X2=5.61 $Y2=0.96
r99 28 29 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.035
+ $X2=5.37 $Y2=1.035
r100 24 56 17.7656 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=5.295 $Y=1.295
+ $X2=5.295 $Y2=1.127
r101 24 26 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.295 $Y=1.295
+ $X2=5.295 $Y2=1.985
r102 21 55 17.7656 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=5.19 $Y=0.96
+ $X2=5.19 $Y2=1.127
r103 21 23 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.19 $Y=0.96 $X2=5.19
+ $Y2=0.56
r104 17 51 17.7656 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=4.875 $Y=1.295
+ $X2=4.875 $Y2=1.127
r105 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.875 $Y=1.295
+ $X2=4.875 $Y2=1.985
r106 13 51 17.7579 $w=2.85e-07 $l=1.05e-07 $layer=POLY_cond $X=4.77 $Y=1.127
+ $X2=4.875 $Y2=1.127
r107 13 48 29.5965 $w=2.85e-07 $l=1.75e-07 $layer=POLY_cond $X=4.77 $Y=1.127
+ $X2=4.595 $Y2=1.127
r108 13 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.77 $Y=1.02
+ $X2=4.77 $Y2=0.56
r109 9 46 17.7656 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=4.455 $Y=1.295
+ $X2=4.455 $Y2=1.127
r110 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.455 $Y=1.295
+ $X2=4.455 $Y2=1.985
r111 5 46 17.7579 $w=2.85e-07 $l=1.05e-07 $layer=POLY_cond $X=4.35 $Y=1.127
+ $X2=4.455 $Y2=1.127
r112 5 43 16.0667 $w=2.85e-07 $l=9.5e-08 $layer=POLY_cond $X=4.35 $Y=1.127
+ $X2=4.255 $Y2=1.127
r113 5 7 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.35 $Y=1.02 $X2=4.35
+ $Y2=0.56
r114 1 41 17.7656 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=4.035 $Y=1.295
+ $X2=4.035 $Y2=1.127
r115 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.035 $Y=1.295
+ $X2=4.035 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%A2 1 3 4 5 8 10 12 15 19 23 25 27 31 33 34
+ 35
c89 35 0 2.34689e-19 $X=7.13 $Y=1.19
c90 19 0 1.02312e-19 $X=6.58 $Y=1.985
r91 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.995
+ $Y=1.16 $X2=6.995 $Y2=1.16
r92 46 48 13.2966 $w=2.9e-07 $l=8e-08 $layer=POLY_cond $X=6.915 $Y=1.217
+ $X2=6.995 $Y2=1.217
r93 42 44 26.5931 $w=2.9e-07 $l=1.6e-07 $layer=POLY_cond $X=6.315 $Y=1.217
+ $X2=6.475 $Y2=1.217
r94 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.315
+ $Y=1.16 $X2=6.315 $Y2=1.16
r95 40 42 25.7621 $w=2.9e-07 $l=1.55e-07 $layer=POLY_cond $X=6.16 $Y=1.217
+ $X2=6.315 $Y2=1.217
r96 39 40 17.4517 $w=2.9e-07 $l=1.05e-07 $layer=POLY_cond $X=6.055 $Y=1.217
+ $X2=6.16 $Y2=1.217
r97 35 49 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.13 $Y=1.21
+ $X2=6.995 $Y2=1.21
r98 34 49 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.67 $Y=1.21
+ $X2=6.995 $Y2=1.21
r99 34 43 15.1525 $w=2.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.67 $Y=1.21
+ $X2=6.315 $Y2=1.21
r100 33 43 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.21 $Y=1.21
+ $X2=6.315 $Y2=1.21
r101 29 51 18.1727 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.335 $Y=1.025
+ $X2=7.335 $Y2=1.217
r102 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.335 $Y=1.025
+ $X2=7.335 $Y2=0.56
r103 25 51 55.6793 $w=2.9e-07 $l=3.35e-07 $layer=POLY_cond $X=7 $Y=1.217
+ $X2=7.335 $Y2=1.217
r104 25 48 0.831034 $w=2.9e-07 $l=5e-09 $layer=POLY_cond $X=7 $Y=1.217 $X2=6.995
+ $Y2=1.217
r105 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7 $Y=1.295 $X2=7
+ $Y2=1.985
r106 21 46 18.1727 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.915 $Y=1.025
+ $X2=6.915 $Y2=1.217
r107 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.915 $Y=1.025
+ $X2=6.915 $Y2=0.56
r108 17 46 55.6793 $w=2.9e-07 $l=3.35e-07 $layer=POLY_cond $X=6.58 $Y=1.217
+ $X2=6.915 $Y2=1.217
r109 17 44 17.4517 $w=2.9e-07 $l=1.05e-07 $layer=POLY_cond $X=6.58 $Y=1.217
+ $X2=6.475 $Y2=1.217
r110 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.58 $Y=1.295
+ $X2=6.58 $Y2=1.985
r111 13 44 18.1727 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.475 $Y=1.025
+ $X2=6.475 $Y2=1.217
r112 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.475 $Y=1.025
+ $X2=6.475 $Y2=0.56
r113 10 40 18.1727 $w=1.5e-07 $l=1.93e-07 $layer=POLY_cond $X=6.16 $Y=1.41
+ $X2=6.16 $Y2=1.217
r114 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.16 $Y=1.41
+ $X2=6.16 $Y2=1.985
r115 6 39 18.1727 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.055 $Y=1.025
+ $X2=6.055 $Y2=1.217
r116 6 8 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.055 $Y=1.025
+ $X2=6.055 $Y2=0.56
r117 4 39 23.6571 $w=2.9e-07 $l=1.50911e-07 $layer=POLY_cond $X=5.98 $Y=1.335
+ $X2=6.055 $Y2=1.217
r118 4 5 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.98 $Y=1.335
+ $X2=5.815 $Y2=1.335
r119 1 5 31.7663 $w=1.27e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.74 $Y=1.41
+ $X2=5.815 $Y2=1.335
r120 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.74 $Y=1.41
+ $X2=5.74 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 58
r68 57 58 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=9.04 $Y=1.16
+ $X2=9.19 $Y2=1.16
r69 55 57 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=9.01 $Y=1.16 $X2=9.04
+ $Y2=1.16
r70 53 55 53.3217 $w=2.7e-07 $l=2.4e-07 $layer=POLY_cond $X=8.77 $Y=1.16
+ $X2=9.01 $Y2=1.16
r71 51 53 22.2174 $w=2.7e-07 $l=1e-07 $layer=POLY_cond $X=8.67 $Y=1.16 $X2=8.77
+ $Y2=1.16
r72 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.67
+ $Y=1.16 $X2=8.67 $Y2=1.16
r73 49 51 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=8.62 $Y=1.16 $X2=8.67
+ $Y2=1.16
r74 48 49 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=8.35 $Y=1.16
+ $X2=8.62 $Y2=1.16
r75 46 48 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=8.33 $Y=1.16 $X2=8.35
+ $Y2=1.16
r76 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.33
+ $Y=1.16 $X2=8.33 $Y2=1.16
r77 44 46 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=8.2 $Y=1.16 $X2=8.33
+ $Y2=1.16
r78 43 44 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=7.93 $Y=1.16 $X2=8.2
+ $Y2=1.16
r79 41 43 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=7.78 $Y=1.16
+ $X2=7.93 $Y2=1.16
r80 35 36 20.0047 $w=2.63e-07 $l=4.6e-07 $layer=LI1_cond $X=8.97 $Y=1.207
+ $X2=9.43 $Y2=1.207
r81 35 52 13.0465 $w=2.63e-07 $l=3e-07 $layer=LI1_cond $X=8.97 $Y=1.207 $X2=8.67
+ $Y2=1.207
r82 35 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.01
+ $Y=1.16 $X2=9.01 $Y2=1.16
r83 34 52 6.95815 $w=2.63e-07 $l=1.6e-07 $layer=LI1_cond $X=8.51 $Y=1.207
+ $X2=8.67 $Y2=1.207
r84 34 47 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=8.51 $Y=1.207
+ $X2=8.33 $Y2=1.207
r85 33 47 12.1768 $w=2.63e-07 $l=2.8e-07 $layer=LI1_cond $X=8.05 $Y=1.207
+ $X2=8.33 $Y2=1.207
r86 29 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.19 $Y=1.295
+ $X2=9.19 $Y2=1.16
r87 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.19 $Y=1.295
+ $X2=9.19 $Y2=1.985
r88 25 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.04 $Y=1.025
+ $X2=9.04 $Y2=1.16
r89 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.04 $Y=1.025
+ $X2=9.04 $Y2=0.56
r90 21 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.77 $Y=1.295
+ $X2=8.77 $Y2=1.16
r91 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.77 $Y=1.295
+ $X2=8.77 $Y2=1.985
r92 17 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.62 $Y=1.025
+ $X2=8.62 $Y2=1.16
r93 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.62 $Y=1.025
+ $X2=8.62 $Y2=0.56
r94 13 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.35 $Y=1.295
+ $X2=8.35 $Y2=1.16
r95 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.35 $Y=1.295
+ $X2=8.35 $Y2=1.985
r96 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.2 $Y=1.025 $X2=8.2
+ $Y2=1.16
r97 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.2 $Y=1.025 $X2=8.2
+ $Y2=0.56
r98 5 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.93 $Y=1.295
+ $X2=7.93 $Y2=1.16
r99 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.93 $Y=1.295 $X2=7.93
+ $Y2=1.985
r100 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.78 $Y=1.025
+ $X2=7.78 $Y2=1.16
r101 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.78 $Y=1.025
+ $X2=7.78 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%Y 1 2 3 4 5 6 7 8 9 10 11 38 40 44 46 50
+ 52 56 58 62 64 68 70 74 76 80 84 85 86 87 88 89 90 92 93 95 96 97 98 99 107
+ 110
c126 107 0 1.98909e-19 $X=0.23 $Y=0.815
c127 92 0 1.02312e-19 $X=7.21 $Y=1.63
c128 38 0 7.52102e-20 $X=1.52 $Y=0.73
r129 107 110 1.39088 $w=2.88e-07 $l=3.5e-08 $layer=LI1_cond $X=0.23 $Y=0.815
+ $X2=0.23 $Y2=0.85
r130 99 119 10.4768 $w=2.73e-07 $l=2.5e-07 $layer=LI1_cond $X=0.222 $Y=2.21
+ $X2=0.222 $Y2=1.96
r131 98 119 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=1.96
r132 98 115 7.7528 $w=2.73e-07 $l=1.85e-07 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=1.685
r133 97 108 3.32435 $w=2.82e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=1.6
+ $X2=0.23 $Y2=1.515
r134 97 115 3.32435 $w=2.82e-07 $l=8.89101e-08 $layer=LI1_cond $X=0.23 $Y=1.6
+ $X2=0.222 $Y2=1.685
r135 97 108 1.39088 $w=2.88e-07 $l=3.5e-08 $layer=LI1_cond $X=0.23 $Y=1.48
+ $X2=0.23 $Y2=1.515
r136 96 97 11.5244 $w=2.88e-07 $l=2.9e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.23 $Y2=1.48
r137 95 107 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=0.73
+ $X2=0.23 $Y2=0.815
r138 95 96 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=0.23 $Y=0.875
+ $X2=0.23 $Y2=1.19
r139 95 110 0.993485 $w=2.88e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=0.875
+ $X2=0.23 $Y2=0.85
r140 92 93 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.21 $Y=1.617
+ $X2=7.045 $Y2=1.617
r141 83 90 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=6.48 $Y=1.6
+ $X2=6.382 $Y2=1.6
r142 83 93 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.48 $Y=1.6
+ $X2=7.045 $Y2=1.6
r143 78 90 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.382 $Y=1.685
+ $X2=6.382 $Y2=1.6
r144 78 80 14.2191 $w=1.93e-07 $l=2.5e-07 $layer=LI1_cond $X=6.382 $Y=1.685
+ $X2=6.382 $Y2=1.935
r145 77 89 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.6 $Y=1.6 $X2=5.505
+ $Y2=1.6
r146 76 90 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=6.285 $Y=1.6
+ $X2=6.382 $Y2=1.6
r147 76 77 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.285 $Y=1.6
+ $X2=5.6 $Y2=1.6
r148 72 89 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=1.685
+ $X2=5.505 $Y2=1.6
r149 72 74 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=5.505 $Y=1.685
+ $X2=5.505 $Y2=1.96
r150 71 88 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.76 $Y=1.6
+ $X2=4.665 $Y2=1.6
r151 70 89 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.41 $Y=1.6
+ $X2=5.505 $Y2=1.6
r152 70 71 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.41 $Y=1.6
+ $X2=4.76 $Y2=1.6
r153 66 88 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=1.685
+ $X2=4.665 $Y2=1.6
r154 66 68 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=4.665 $Y=1.685
+ $X2=4.665 $Y2=1.96
r155 65 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.715 $Y=1.6
+ $X2=3.62 $Y2=1.6
r156 64 88 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.57 $Y=1.6
+ $X2=4.665 $Y2=1.6
r157 64 65 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.57 $Y=1.6
+ $X2=3.715 $Y2=1.6
r158 60 87 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.685
+ $X2=3.62 $Y2=1.6
r159 60 62 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=3.62 $Y=1.685
+ $X2=3.62 $Y2=1.96
r160 59 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.875 $Y=1.6
+ $X2=2.78 $Y2=1.6
r161 58 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.525 $Y=1.6
+ $X2=3.62 $Y2=1.6
r162 58 59 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.525 $Y=1.6
+ $X2=2.875 $Y2=1.6
r163 54 86 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=1.685
+ $X2=2.78 $Y2=1.6
r164 54 56 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=2.78 $Y=1.685
+ $X2=2.78 $Y2=1.96
r165 53 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.035 $Y=1.6
+ $X2=1.94 $Y2=1.6
r166 52 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.685 $Y=1.6
+ $X2=2.78 $Y2=1.6
r167 52 53 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.685 $Y=1.6
+ $X2=2.035 $Y2=1.6
r168 48 85 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=1.685
+ $X2=1.94 $Y2=1.6
r169 48 50 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.94 $Y=1.685
+ $X2=1.94 $Y2=1.96
r170 47 84 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.195 $Y=1.6 $X2=1.105
+ $Y2=1.6
r171 46 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.845 $Y=1.6
+ $X2=1.94 $Y2=1.6
r172 46 47 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.845 $Y=1.6
+ $X2=1.195 $Y2=1.6
r173 42 84 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=1.685
+ $X2=1.105 $Y2=1.6
r174 42 44 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.105 $Y=1.685
+ $X2=1.105 $Y2=1.96
r175 41 97 3.22099 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.375 $Y=1.6
+ $X2=0.23 $Y2=1.6
r176 40 84 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.015 $Y=1.6 $X2=1.105
+ $Y2=1.6
r177 40 41 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.015 $Y=1.6
+ $X2=0.375 $Y2=1.6
r178 36 38 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.68 $Y=0.73
+ $X2=1.52 $Y2=0.73
r179 34 95 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.375 $Y=0.73
+ $X2=0.23 $Y2=0.73
r180 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.375 $Y=0.73
+ $X2=0.68 $Y2=0.73
r181 11 92 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.075
+ $Y=1.485 $X2=7.21 $Y2=1.63
r182 10 80 600 $w=1.7e-07 $l=5.13079e-07 $layer=licon1_PDIFF $count=1 $X=6.235
+ $Y=1.485 $X2=6.37 $Y2=1.935
r183 9 74 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.37
+ $Y=1.485 $X2=5.505 $Y2=1.96
r184 8 68 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.53
+ $Y=1.485 $X2=4.665 $Y2=1.96
r185 7 62 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.96
r186 6 56 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.96
r187 5 50 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r188 4 44 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r189 3 119 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r190 2 38 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.73
r191 1 36 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 58 60 62 65 66 68 69 71 72 74 75 77 78 79 81 102 106 111 117 120 123 127
r157 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r158 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r159 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r160 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r161 115 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r162 115 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r163 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r164 112 123 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.72 $Y=2.72
+ $X2=8.565 $Y2=2.72
r165 112 114 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.72 $Y=2.72
+ $X2=8.97 $Y2=2.72
r166 111 126 4.6205 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.265 $Y=2.72
+ $X2=9.462 $Y2=2.72
r167 111 114 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.265 $Y=2.72
+ $X2=8.97 $Y2=2.72
r168 110 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r169 110 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r170 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r171 107 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.885 $Y=2.72
+ $X2=7.72 $Y2=2.72
r172 107 109 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.885 $Y=2.72
+ $X2=8.05 $Y2=2.72
r173 106 123 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.41 $Y=2.72
+ $X2=8.565 $Y2=2.72
r174 106 109 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.41 $Y=2.72
+ $X2=8.05 $Y2=2.72
r175 105 121 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.59 $Y2=2.72
r176 104 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r177 102 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.555 $Y=2.72
+ $X2=7.72 $Y2=2.72
r178 102 104 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=7.555 $Y=2.72
+ $X2=5.29 $Y2=2.72
r179 101 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r180 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r181 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r182 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r183 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r184 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r185 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r186 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r187 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r188 89 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r189 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r190 86 117 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.687 $Y2=2.72
r191 86 88 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r192 81 117 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.53 $Y=2.72
+ $X2=0.687 $Y2=2.72
r193 81 83 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.53 $Y=2.72 $X2=0.23
+ $Y2=2.72
r194 79 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r195 79 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r196 77 100 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.93 $Y=2.72
+ $X2=4.83 $Y2=2.72
r197 77 78 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.93 $Y=2.72
+ $X2=5.075 $Y2=2.72
r198 76 104 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.22 $Y=2.72
+ $X2=5.29 $Y2=2.72
r199 76 78 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.22 $Y=2.72
+ $X2=5.075 $Y2=2.72
r200 74 97 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.72
+ $X2=3.91 $Y2=2.72
r201 74 75 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=4.075 $Y=2.72
+ $X2=4.237 $Y2=2.72
r202 73 100 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.4 $Y=2.72
+ $X2=4.83 $Y2=2.72
r203 73 75 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.4 $Y=2.72
+ $X2=4.237 $Y2=2.72
r204 71 94 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.99 $Y2=2.72
r205 71 72 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.2 $Y2=2.72
r206 70 97 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.355 $Y=2.72
+ $X2=3.91 $Y2=2.72
r207 70 72 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.355 $Y=2.72
+ $X2=3.2 $Y2=2.72
r208 68 91 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.07 $Y2=2.72
r209 68 69 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.36 $Y2=2.72
r210 67 94 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.515 $Y=2.72
+ $X2=2.99 $Y2=2.72
r211 67 69 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.515 $Y=2.72
+ $X2=2.36 $Y2=2.72
r212 65 88 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.39 $Y=2.72
+ $X2=1.15 $Y2=2.72
r213 65 66 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.39 $Y=2.72
+ $X2=1.532 $Y2=2.72
r214 64 91 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.675 $Y=2.72
+ $X2=2.07 $Y2=2.72
r215 64 66 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.675 $Y=2.72
+ $X2=1.532 $Y2=2.72
r216 60 126 2.9787 $w=3.1e-07 $l=1.03899e-07 $layer=LI1_cond $X=9.42 $Y=2.635
+ $X2=9.462 $Y2=2.72
r217 60 62 23.6065 $w=3.08e-07 $l=6.35e-07 $layer=LI1_cond $X=9.42 $Y=2.635
+ $X2=9.42 $Y2=2
r218 56 123 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.565 $Y=2.635
+ $X2=8.565 $Y2=2.72
r219 56 58 22.863 $w=3.08e-07 $l=6.15e-07 $layer=LI1_cond $X=8.565 $Y=2.635
+ $X2=8.565 $Y2=2.02
r220 52 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.72 $Y=2.635
+ $X2=7.72 $Y2=2.72
r221 52 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.72 $Y=2.635
+ $X2=7.72 $Y2=2.34
r222 48 78 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=2.635
+ $X2=5.075 $Y2=2.72
r223 48 50 24.4397 $w=2.88e-07 $l=6.15e-07 $layer=LI1_cond $X=5.075 $Y=2.635
+ $X2=5.075 $Y2=2.02
r224 44 75 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.237 $Y=2.635
+ $X2=4.237 $Y2=2.72
r225 44 46 21.8078 $w=3.23e-07 $l=6.15e-07 $layer=LI1_cond $X=4.237 $Y=2.635
+ $X2=4.237 $Y2=2.02
r226 40 72 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.72
r227 40 42 22.863 $w=3.08e-07 $l=6.15e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.02
r228 36 69 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r229 36 38 22.863 $w=3.08e-07 $l=6.15e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.02
r230 32 66 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.532 $Y=2.635
+ $X2=1.532 $Y2=2.72
r231 32 34 24.8685 $w=2.83e-07 $l=6.15e-07 $layer=LI1_cond $X=1.532 $Y=2.635
+ $X2=1.532 $Y2=2.02
r232 28 117 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.687 $Y=2.635
+ $X2=0.687 $Y2=2.72
r233 28 30 22.5001 $w=3.13e-07 $l=6.15e-07 $layer=LI1_cond $X=0.687 $Y=2.635
+ $X2=0.687 $Y2=2.02
r234 9 62 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.265
+ $Y=1.485 $X2=9.4 $Y2=2
r235 8 58 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=8.425
+ $Y=1.485 $X2=8.56 $Y2=2.02
r236 7 54 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.595
+ $Y=2.2 $X2=7.72 $Y2=2.34
r237 6 50 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.485 $X2=5.085 $Y2=2.02
r238 5 46 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=4.11
+ $Y=1.485 $X2=4.245 $Y2=2.02
r239 4 42 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.02
r240 3 38 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.02
r241 2 34 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.02
r242 1 30 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%A_1163_297# 1 2 3 4 15 17 18 22 23 24 29
+ 31 32 35 38
r57 33 35 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=8.985 $Y=1.685
+ $X2=8.985 $Y2=1.96
r58 31 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.89 $Y=1.6
+ $X2=8.985 $Y2=1.685
r59 31 32 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.89 $Y=1.6
+ $X2=8.235 $Y2=1.6
r60 27 38 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=8.145 $Y=2.06
+ $X2=8.14 $Y2=1.975
r61 27 29 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=8.145 $Y=2.06
+ $X2=8.145 $Y2=2.3
r62 26 38 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.14 $Y=1.89
+ $X2=8.14 $Y2=1.975
r63 25 32 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.14 $Y=1.685
+ $X2=8.235 $Y2=1.6
r64 25 26 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=8.14 $Y=1.685
+ $X2=8.14 $Y2=1.89
r65 23 38 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.045 $Y=1.975
+ $X2=8.14 $Y2=1.975
r66 23 24 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=8.045 $Y=1.975
+ $X2=7.005 $Y2=1.975
r67 20 22 5.37807 $w=2.98e-07 $l=1.4e-07 $layer=LI1_cond $X=6.855 $Y=2.27
+ $X2=6.855 $Y2=2.13
r68 19 24 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.855 $Y=2.06
+ $X2=7.005 $Y2=1.975
r69 19 22 2.68903 $w=2.98e-07 $l=7e-08 $layer=LI1_cond $X=6.855 $Y=2.06
+ $X2=6.855 $Y2=2.13
r70 17 20 7.22316 $w=1.95e-07 $l=1.92484e-07 $layer=LI1_cond $X=6.705 $Y=2.367
+ $X2=6.855 $Y2=2.27
r71 17 18 33.5571 $w=1.93e-07 $l=5.9e-07 $layer=LI1_cond $X=6.705 $Y=2.367
+ $X2=6.115 $Y2=2.367
r72 13 18 7.4197 $w=1.95e-07 $l=2.07918e-07 $layer=LI1_cond $X=5.95 $Y=2.27
+ $X2=6.115 $Y2=2.367
r73 13 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.95 $Y=2.27
+ $X2=5.95 $Y2=2.02
r74 4 35 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.845
+ $Y=1.485 $X2=8.98 $Y2=1.96
r75 3 38 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=8.005
+ $Y=1.485 $X2=8.14 $Y2=1.96
r76 3 29 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.005
+ $Y=1.485 $X2=8.14 $Y2=2.3
r77 2 22 600 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=1 $X=6.655
+ $Y=1.485 $X2=6.79 $Y2=2.13
r78 1 15 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.815
+ $Y=1.485 $X2=5.95 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%A_27_47# 1 2 3 4 5 16 26 30
r36 28 30 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.72
+ $X2=3.62 $Y2=0.72
r37 26 28 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.72
+ $X2=2.78 $Y2=0.72
r38 23 26 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.94 $Y=0.615
+ $X2=2.025 $Y2=0.72
r39 23 25 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.94 $Y=0.615
+ $X2=1.94 $Y2=0.56
r40 22 25 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.475
+ $X2=1.94 $Y2=0.56
r41 18 21 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=0.26 $Y=0.38 $X2=1.1
+ $Y2=0.38
r42 16 22 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.855 $Y=0.38
+ $X2=1.94 $Y2=0.475
r43 16 21 44.0718 $w=1.88e-07 $l=7.55e-07 $layer=LI1_cond $X=1.855 $Y=0.38
+ $X2=1.1 $Y2=0.38
r44 5 30 182 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.7
r45 4 28 182 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.7
r46 3 25 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.56
r47 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r48 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%A_445_47# 1 2 3 4 21
r30 19 21 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.35 $X2=5.4
+ $Y2=0.35
r31 17 19 79.3876 $w=1.88e-07 $l=1.36e-06 $layer=LI1_cond $X=3.2 $Y=0.35
+ $X2=4.56 $Y2=0.35
r32 14 17 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.35 $X2=3.2
+ $Y2=0.35
r33 4 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.36
r34 3 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.36
r35 2 17 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.36
r36 1 14 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%A_803_47# 1 2 3 4 5 6 7 36
r51 34 36 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=8.41 $Y=0.78
+ $X2=9.25 $Y2=0.78
r52 32 34 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=7.57 $Y=0.78
+ $X2=8.41 $Y2=0.78
r53 30 32 40.7965 $w=2.48e-07 $l=8.85e-07 $layer=LI1_cond $X=6.685 $Y=0.78
+ $X2=7.57 $Y2=0.78
r54 28 30 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=5.845 $Y=0.78
+ $X2=6.685 $Y2=0.78
r55 26 28 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=4.98 $Y=0.78
+ $X2=5.845 $Y2=0.78
r56 23 26 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.78
+ $X2=4.98 $Y2=0.78
r57 7 36 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=9.115
+ $Y=0.235 $X2=9.25 $Y2=0.74
r58 6 34 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=8.275
+ $Y=0.235 $X2=8.41 $Y2=0.74
r59 5 32 182 $w=1.7e-07 $l=5.79504e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.235 $X2=7.57 $Y2=0.74
r60 4 30 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=6.55
+ $Y=0.235 $X2=6.685 $Y2=0.74
r61 3 28 182 $w=1.7e-07 $l=5.79504e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.845 $Y2=0.74
r62 2 26 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.74
r63 1 23 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_4%VGND 1 2 3 4 15 19 23 27 30 31 32 34 42 47
+ 57 58 61 64 67
c109 34 0 1.98909e-19 $X=6.1 $Y=0
r110 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r111 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r112 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r113 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r114 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r115 55 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.05
+ $Y2=0
r116 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r117 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.155 $Y=0 $X2=7.99
+ $Y2=0
r118 52 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.155 $Y=0
+ $X2=8.51 $Y2=0
r119 51 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r120 51 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r121 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r122 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=7.125
+ $Y2=0
r123 48 50 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=7.59
+ $Y2=0
r124 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=0 $X2=7.99
+ $Y2=0
r125 47 50 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.825 $Y=0
+ $X2=7.59 $Y2=0
r126 46 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r127 46 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r128 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r129 43 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.43 $Y=0 $X2=6.265
+ $Y2=0
r130 43 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.43 $Y=0 $X2=6.67
+ $Y2=0
r131 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.125
+ $Y2=0
r132 42 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=6.67
+ $Y2=0
r133 41 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r134 40 41 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r135 36 40 360.128 $w=1.68e-07 $l=5.52e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=5.75
+ $Y2=0
r136 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.1 $Y=0 $X2=6.265
+ $Y2=0
r137 34 40 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.1 $Y=0 $X2=5.75
+ $Y2=0
r138 32 41 1.57067 $w=4.8e-07 $l=5.52e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=5.75
+ $Y2=0
r139 32 36 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r140 30 54 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.665 $Y=0
+ $X2=8.51 $Y2=0
r141 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=0 $X2=8.83
+ $Y2=0
r142 29 57 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.995 $Y=0
+ $X2=9.43 $Y2=0
r143 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.995 $Y=0 $X2=8.83
+ $Y2=0
r144 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.83 $Y=0.085
+ $X2=8.83 $Y2=0
r145 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.83 $Y=0.085
+ $X2=8.83 $Y2=0.36
r146 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=0.085
+ $X2=7.99 $Y2=0
r147 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.99 $Y=0.085
+ $X2=7.99 $Y2=0.36
r148 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=0.085
+ $X2=7.125 $Y2=0
r149 17 19 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.125 $Y=0.085
+ $X2=7.125 $Y2=0.365
r150 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.265 $Y=0.085
+ $X2=6.265 $Y2=0
r151 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.265 $Y=0.085
+ $X2=6.265 $Y2=0.38
r152 4 27 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=8.695
+ $Y=0.235 $X2=8.83 $Y2=0.36
r153 3 23 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.855
+ $Y=0.235 $X2=7.99 $Y2=0.36
r154 2 19 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=6.99
+ $Y=0.235 $X2=7.125 $Y2=0.365
r155 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.13
+ $Y=0.235 $X2=6.265 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a32oi_4.pxi.spice
* Created: Tue Sep  1 18:56:05 2020
* 
x_PM_SKY130_FD_SC_HD__A32OI_4%B2 N_B2_c_105_n N_B2_M1014_g N_B2_M1002_g
+ N_B2_c_106_n N_B2_M1021_g N_B2_M1005_g N_B2_c_107_n N_B2_M1025_g N_B2_M1027_g
+ N_B2_c_108_n N_B2_M1038_g N_B2_M1034_g B2 B2 B2 B2 B2 B2 N_B2_c_109_n
+ N_B2_c_110_n PM_SKY130_FD_SC_HD__A32OI_4%B2
x_PM_SKY130_FD_SC_HD__A32OI_4%B1 N_B1_c_184_n N_B1_M1022_g N_B1_M1000_g
+ N_B1_c_185_n N_B1_M1028_g N_B1_M1006_g N_B1_c_186_n N_B1_M1032_g N_B1_M1031_g
+ N_B1_c_187_n N_B1_M1033_g N_B1_M1035_g B1 B1 N_B1_c_189_n
+ PM_SKY130_FD_SC_HD__A32OI_4%B1
x_PM_SKY130_FD_SC_HD__A32OI_4%A1 N_A1_M1004_g N_A1_M1008_g N_A1_c_262_n
+ N_A1_M1013_g N_A1_M1012_g N_A1_c_263_n N_A1_M1015_g N_A1_c_264_n N_A1_M1023_g
+ N_A1_M1039_g N_A1_c_265_n N_A1_M1029_g A1 A1 A1 A1 N_A1_c_267_n
+ PM_SKY130_FD_SC_HD__A32OI_4%A1
x_PM_SKY130_FD_SC_HD__A32OI_4%A2 N_A2_c_328_n N_A2_M1016_g N_A2_M1003_g
+ N_A2_c_329_n N_A2_M1018_g N_A2_M1024_g N_A2_c_330_n N_A2_M1026_g N_A2_M1036_g
+ N_A2_c_331_n N_A2_M1030_g N_A2_M1037_g A2 A2 A2 A2
+ PM_SKY130_FD_SC_HD__A32OI_4%A2
x_PM_SKY130_FD_SC_HD__A32OI_4%A3 N_A3_c_391_n N_A3_M1009_g N_A3_M1001_g
+ N_A3_c_392_n N_A3_M1011_g N_A3_M1007_g N_A3_c_393_n N_A3_M1017_g N_A3_M1010_g
+ N_A3_c_394_n N_A3_M1019_g N_A3_M1020_g A3 A3 A3 A3 A3 N_A3_c_396_n
+ N_A3_c_397_n N_A3_c_398_n PM_SKY130_FD_SC_HD__A32OI_4%A3
x_PM_SKY130_FD_SC_HD__A32OI_4%A_27_297# N_A_27_297#_M1002_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1034_s N_A_27_297#_M1006_s N_A_27_297#_M1035_s
+ N_A_27_297#_M1008_d N_A_27_297#_M1039_d N_A_27_297#_M1024_s
+ N_A_27_297#_M1037_s N_A_27_297#_M1007_d N_A_27_297#_M1020_d
+ N_A_27_297#_c_461_n N_A_27_297#_c_473_n N_A_27_297#_c_474_n
+ N_A_27_297#_c_472_n N_A_27_297#_c_533_p N_A_27_297#_c_478_n
+ N_A_27_297#_c_485_n N_A_27_297#_c_486_n N_A_27_297#_c_537_p
+ N_A_27_297#_c_490_n N_A_27_297#_c_497_n N_A_27_297#_c_498_n
+ N_A_27_297#_c_545_p N_A_27_297#_c_502_n N_A_27_297#_c_546_p
+ N_A_27_297#_c_482_n N_A_27_297#_c_484_n N_A_27_297#_c_494_n
+ N_A_27_297#_c_496_n N_A_27_297#_c_507_n PM_SKY130_FD_SC_HD__A32OI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A32OI_4%Y N_Y_M1022_d N_Y_M1032_d N_Y_M1013_d N_Y_M1023_d
+ N_Y_M1002_d N_Y_M1027_d N_Y_M1000_d N_Y_M1031_d N_Y_c_571_n N_Y_c_575_n
+ N_Y_c_594_n N_Y_c_566_n N_Y_c_600_n N_Y_c_577_n N_Y_c_583_n N_Y_c_605_n Y Y Y
+ Y Y N_Y_c_569_n PM_SKY130_FD_SC_HD__A32OI_4%Y
x_PM_SKY130_FD_SC_HD__A32OI_4%VPWR N_VPWR_M1004_s N_VPWR_M1012_s N_VPWR_M1003_d
+ N_VPWR_M1036_d N_VPWR_M1001_s N_VPWR_M1010_s N_VPWR_c_670_n N_VPWR_c_671_n
+ N_VPWR_c_672_n N_VPWR_c_673_n N_VPWR_c_674_n N_VPWR_c_675_n N_VPWR_c_676_n
+ N_VPWR_c_677_n N_VPWR_c_678_n N_VPWR_c_679_n VPWR N_VPWR_c_680_n
+ N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_669_n N_VPWR_c_685_n
+ N_VPWR_c_686_n N_VPWR_c_687_n N_VPWR_c_688_n N_VPWR_c_689_n
+ PM_SKY130_FD_SC_HD__A32OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A32OI_4%A_27_47# N_A_27_47#_M1014_d N_A_27_47#_M1021_d
+ N_A_27_47#_M1038_d N_A_27_47#_M1028_s N_A_27_47#_M1033_s N_A_27_47#_c_828_p
+ N_A_27_47#_c_795_n N_A_27_47#_c_799_n N_A_27_47#_c_831_p N_A_27_47#_c_802_n
+ N_A_27_47#_c_826_p N_A_27_47#_c_794_n N_A_27_47#_c_806_n
+ PM_SKY130_FD_SC_HD__A32OI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__A32OI_4%VGND N_VGND_M1014_s N_VGND_M1025_s N_VGND_M1009_d
+ N_VGND_M1011_d N_VGND_M1019_d N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n
+ N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n VGND
+ N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n
+ PM_SKY130_FD_SC_HD__A32OI_4%VGND
x_PM_SKY130_FD_SC_HD__A32OI_4%A_803_47# N_A_803_47#_M1013_s N_A_803_47#_M1015_s
+ N_A_803_47#_M1029_s N_A_803_47#_M1018_d N_A_803_47#_M1030_d
+ N_A_803_47#_c_977_n PM_SKY130_FD_SC_HD__A32OI_4%A_803_47#
x_PM_SKY130_FD_SC_HD__A32OI_4%A_1249_47# N_A_1249_47#_M1016_s
+ N_A_1249_47#_M1026_s N_A_1249_47#_M1009_s N_A_1249_47#_M1017_s
+ N_A_1249_47#_c_1006_n N_A_1249_47#_c_1031_n N_A_1249_47#_c_1015_n
+ N_A_1249_47#_c_1038_n N_A_1249_47#_c_1019_n
+ PM_SKY130_FD_SC_HD__A32OI_4%A_1249_47#
cc_1 VNB N_B2_c_105_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_106_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_B2_c_107_n 0.0157099f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_B2_c_108_n 0.0159385f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_B2_c_109_n 0.0874061f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_6 VNB N_B2_c_110_n 0.00936732f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.305
cc_7 VNB N_B1_c_184_n 0.0156371f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B1_c_185_n 0.0159777f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_9 VNB N_B1_c_186_n 0.0160026f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_10 VNB N_B1_c_187_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_11 VNB B1 0.00328581f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_12 VNB N_B1_c_189_n 0.061374f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_13 VNB N_A1_c_262_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_14 VNB N_A1_c_263_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_15 VNB N_A1_c_264_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_16 VNB N_A1_c_265_n 0.0182888f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_17 VNB A1 0.00147415f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_18 VNB N_A1_c_267_n 0.0946662f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_19 VNB N_A2_c_328_n 0.0174381f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A2_c_329_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_21 VNB N_A2_c_330_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_22 VNB N_A2_c_331_n 0.0922932f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_23 VNB A2 0.00975135f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_24 VNB N_A3_c_391_n 0.0210871f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_25 VNB N_A3_c_392_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_26 VNB N_A3_c_393_n 0.0157748f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_27 VNB N_A3_c_394_n 0.0183607f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_28 VNB A3 0.00570534f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_29 VNB N_A3_c_396_n 0.0922167f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_30 VNB N_A3_c_397_n 0.00332226f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_31 VNB N_A3_c_398_n 0.00834913f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.19
cc_32 VNB N_Y_c_566_n 0.00751058f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_33 VNB Y 0.00292839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB Y 7.84964e-19 $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.19
cc_35 VNB N_Y_c_569_n 9.73907e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_669_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_794_n 0.00216815f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_38 VNB N_VGND_c_845_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_39 VNB N_VGND_c_846_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_40 VNB N_VGND_c_847_n 0.147234f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_41 VNB N_VGND_c_848_n 0.00551074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_849_n 3.03604e-19 $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_43 VNB N_VGND_c_850_n 0.0105543f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_44 VNB N_VGND_c_851_n 0.0131974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_852_n 0.0151407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_853_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_47 VNB N_VGND_c_854_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_48 VNB N_VGND_c_855_n 0.0120461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_856_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_857_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_858_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_859_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_860_n 0.473164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_803_47#_c_977_n 0.00430013f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_55 VNB N_A_1249_47#_c_1006_n 0.0140526f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_56 VPB N_B2_M1002_g 0.0218881f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_57 VPB N_B2_M1005_g 0.0185002f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_58 VPB N_B2_M1027_g 0.0185036f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_59 VPB N_B2_M1034_g 0.018798f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_60 VPB B2 0.0257322f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_61 VPB N_B2_c_109_n 0.0202562f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_62 VPB N_B1_M1000_g 0.0172006f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_63 VPB N_B1_M1006_g 0.0184662f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_64 VPB N_B1_M1031_g 0.0185026f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_65 VPB N_B1_M1035_g 0.0190626f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_66 VPB B1 0.00230149f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_67 VPB N_B1_c_189_n 0.0105074f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_68 VPB N_A1_M1004_g 0.017785f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_69 VPB N_A1_M1008_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A1_M1012_g 0.0208556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A1_M1039_g 0.0232143f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_72 VPB N_A1_c_267_n 0.0303494f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_73 VPB N_A2_M1003_g 0.0196624f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_74 VPB N_A2_M1024_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_75 VPB N_A2_M1036_g 0.0172788f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_76 VPB N_A2_c_331_n 0.0160578f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_77 VPB N_A2_M1037_g 0.0241559f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_78 VPB N_A3_M1001_g 0.025757f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_79 VPB N_A3_M1007_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_80 VPB N_A3_M1010_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_81 VPB N_A3_M1020_g 0.025757f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_82 VPB N_A3_c_396_n 0.020695f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_83 VPB N_A_27_297#_c_461_n 0.00821562f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_84 VPB Y 0.00357195f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.19
cc_85 VPB N_VPWR_c_670_n 4.01796e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_671_n 0.0146009f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_87 VPB N_VPWR_c_672_n 0.00681796f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_88 VPB N_VPWR_c_673_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.785
cc_89 VPB N_VPWR_c_674_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_90 VPB N_VPWR_c_675_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_676_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_92 VPB N_VPWR_c_677_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_93 VPB N_VPWR_c_678_n 0.0219711f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.16
cc_94 VPB N_VPWR_c_679_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.16
cc_95 VPB N_VPWR_c_680_n 0.0936941f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.305
cc_96 VPB N_VPWR_c_681_n 0.0290389f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.19
cc_97 VPB N_VPWR_c_682_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_683_n 0.0165408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_669_n 0.0480211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_685_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_686_n 0.0128614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_687_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_688_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_689_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 N_B2_c_108_n N_B1_c_184_n 0.0274585f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_106 N_B2_M1034_g N_B1_M1000_g 0.0274585f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_107 B2 N_B1_c_189_n 2.26828e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B2_c_109_n N_B1_c_189_n 0.0274585f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_109 B2 N_A_27_297#_M1002_s 0.0121542f $X=0.15 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_110 N_B2_M1002_g N_A_27_297#_c_461_n 0.0115553f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_111 N_B2_M1005_g N_A_27_297#_c_461_n 0.00922647f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B2_M1027_g N_A_27_297#_c_461_n 0.00922647f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B2_M1034_g N_A_27_297#_c_461_n 0.00922647f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_114 B2 N_A_27_297#_c_461_n 0.0106869f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_115 N_B2_M1005_g N_Y_c_571_n 0.00889401f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B2_M1027_g N_Y_c_571_n 0.00889401f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_117 B2 N_Y_c_571_n 0.0221146f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B2_c_109_n N_Y_c_571_n 0.00192838f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B2_M1034_g N_Y_c_575_n 0.00970434f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_120 B2 N_Y_c_575_n 0.00309329f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_121 N_B2_M1002_g N_Y_c_577_n 0.0105959f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B2_M1005_g N_Y_c_577_n 0.00727492f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B2_M1027_g N_Y_c_577_n 9.97172e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_124 B2 N_Y_c_577_n 0.0282162f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_125 B2 N_Y_c_577_n 0.0144995f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B2_c_109_n N_Y_c_577_n 0.00200399f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B2_M1005_g N_Y_c_583_n 9.97172e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B2_M1027_g N_Y_c_583_n 0.00727492f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B2_M1034_g N_Y_c_583_n 0.00582938f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_130 B2 N_Y_c_583_n 0.0144995f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B2_c_109_n N_Y_c_583_n 0.00200399f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B2_c_108_n Y 0.00353901f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_133 B2 Y 0.0156534f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B2_M1034_g Y 0.00641082f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B2_c_109_n Y 0.00353901f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B2_c_108_n N_Y_c_569_n 9.17572e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B2_M1002_g N_VPWR_c_680_n 0.00366111f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B2_M1005_g N_VPWR_c_680_n 0.00366111f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B2_M1027_g N_VPWR_c_680_n 0.00366111f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B2_M1034_g N_VPWR_c_680_n 0.00366111f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B2_M1002_g N_VPWR_c_669_n 0.00619429f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B2_M1005_g N_VPWR_c_669_n 0.00524008f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B2_M1027_g N_VPWR_c_669_n 0.00524008f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B2_M1034_g N_VPWR_c_669_n 0.00526729f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B2_c_105_n N_A_27_47#_c_795_n 0.0132392f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B2_c_106_n N_A_27_47#_c_795_n 0.0119869f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_147 B2 N_A_27_47#_c_795_n 0.0274913f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_148 N_B2_c_109_n N_A_27_47#_c_795_n 0.00207061f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_149 B2 N_A_27_47#_c_799_n 5.91515e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_150 N_B2_c_109_n N_A_27_47#_c_799_n 0.00385879f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_151 N_B2_c_110_n N_A_27_47#_c_799_n 0.00931777f $X=0.22 $Y=1.305 $X2=0 $Y2=0
cc_152 N_B2_c_107_n N_A_27_47#_c_802_n 0.0119869f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B2_c_108_n N_A_27_47#_c_802_n 0.0128313f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_154 B2 N_A_27_47#_c_802_n 0.0236275f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_155 N_B2_c_109_n N_A_27_47#_c_802_n 0.00207061f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_156 B2 N_A_27_47#_c_806_n 0.0090006f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_157 N_B2_c_109_n N_A_27_47#_c_806_n 0.00216182f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B2_c_105_n N_VGND_c_845_n 0.00834749f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B2_c_106_n N_VGND_c_845_n 0.00664421f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_107_n N_VGND_c_845_n 5.08801e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_106_n N_VGND_c_846_n 5.08801e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B2_c_107_n N_VGND_c_846_n 0.00664421f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B2_c_108_n N_VGND_c_846_n 0.00815339f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_108_n N_VGND_c_847_n 0.00339367f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_165 N_B2_c_105_n N_VGND_c_852_n 0.00339367f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_166 N_B2_c_106_n N_VGND_c_853_n 0.00339367f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B2_c_107_n N_VGND_c_853_n 0.00339367f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B2_c_105_n N_VGND_c_860_n 0.00489827f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B2_c_106_n N_VGND_c_860_n 0.00394406f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B2_c_107_n N_VGND_c_860_n 0.00394406f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B2_c_108_n N_VGND_c_860_n 0.00401529f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_M1035_g N_A1_M1004_g 0.0258389f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_173 B1 A1 0.015263f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_174 N_B1_c_189_n A1 2.33231e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_175 B1 N_A1_c_267_n 0.0041816f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_176 N_B1_c_189_n N_A1_c_267_n 0.0258389f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B1_M1000_g N_A_27_297#_c_461_n 0.00788535f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_178 N_B1_M1006_g N_A_27_297#_c_461_n 0.00922647f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_179 N_B1_M1031_g N_A_27_297#_c_461_n 0.00918232f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1035_g N_A_27_297#_c_461_n 0.0115553f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_181 B1 N_A_27_297#_c_472_n 0.00107674f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_182 N_B1_M1000_g N_Y_c_575_n 2.32576e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_c_184_n N_Y_c_594_n 0.00217694f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_c_185_n N_Y_c_566_n 0.0111239f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B1_c_186_n N_Y_c_566_n 0.00847802f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_187_n N_Y_c_566_n 0.010581f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_187 B1 N_Y_c_566_n 0.0555522f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_188 N_B1_c_189_n N_Y_c_566_n 0.0054372f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B1_M1006_g N_Y_c_600_n 0.0110066f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B1_M1031_g N_Y_c_600_n 0.00880672f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_191 B1 N_Y_c_600_n 0.0211289f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_192 N_B1_c_189_n N_Y_c_600_n 0.00191112f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B1_M1000_g N_Y_c_583_n 3.18843e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B1_M1006_g N_Y_c_605_n 9.97172e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_M1031_g N_Y_c_605_n 0.00725326f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_M1035_g N_Y_c_605_n 0.00620391f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_197 B1 N_Y_c_605_n 0.0158881f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_198 N_B1_c_189_n N_Y_c_605_n 0.0019817f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_c_184_n Y 0.00330483f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_200 B1 Y 0.0215106f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_201 N_B1_c_189_n Y 0.0103741f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_M1000_g Y 0.0122558f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_M1006_g Y 0.00867382f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_204 N_B1_M1031_g Y 0.00107659f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B1_c_189_n Y 0.0015642f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B1_M1000_g Y 0.00603409f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1006_g Y 0.00601384f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_c_189_n Y 0.00803287f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_209 N_B1_c_184_n N_Y_c_569_n 0.00389039f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B1_c_185_n N_Y_c_569_n 0.00380472f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B1_M1035_g N_VPWR_c_670_n 0.00124093f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1000_g N_VPWR_c_680_n 0.00366111f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1006_g N_VPWR_c_680_n 0.00366111f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1031_g N_VPWR_c_680_n 0.00366111f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1035_g N_VPWR_c_680_n 0.00366111f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_M1000_g N_VPWR_c_669_n 0.00526729f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B1_M1006_g N_VPWR_c_669_n 0.00524008f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_M1031_g N_VPWR_c_669_n 0.00524008f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B1_M1035_g N_VPWR_c_669_n 0.00535777f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B1_c_184_n N_A_27_47#_c_794_n 0.00928405f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_185_n N_A_27_47#_c_794_n 0.00784733f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_186_n N_A_27_47#_c_794_n 0.00789149f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B1_c_187_n N_A_27_47#_c_794_n 0.00789149f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B1_c_189_n N_A_27_47#_c_794_n 2.21602e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_225 N_B1_c_184_n N_VGND_c_846_n 0.00127293f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B1_c_184_n N_VGND_c_847_n 0.00366111f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B1_c_185_n N_VGND_c_847_n 0.00366111f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_186_n N_VGND_c_847_n 0.00366111f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_187_n N_VGND_c_847_n 0.00366111f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_184_n N_VGND_c_860_n 0.00530732f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_185_n N_VGND_c_860_n 0.00524008f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B1_c_186_n N_VGND_c_860_n 0.00524008f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_187_n N_VGND_c_860_n 0.00656615f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A1_c_265_n N_A2_c_328_n 0.0170425f $X=5.61 $Y=1.01 $X2=-0.19 $Y2=-0.24
cc_235 N_A1_M1039_g N_A2_M1003_g 0.0100453f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A1_c_267_n N_A2_c_331_n 0.0270878f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_237 A1 A2 0.00588806f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_238 N_A1_c_267_n A2 0.00118416f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_239 N_A1_M1004_g N_A_27_297#_c_473_n 0.00562448f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A1_M1004_g N_A_27_297#_c_474_n 0.0144167f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A1_M1008_g N_A_27_297#_c_474_n 0.0147045f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_242 A1 N_A_27_297#_c_474_n 0.024622f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_243 N_A1_c_267_n N_A_27_297#_c_474_n 0.00201508f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_244 N_A1_M1012_g N_A_27_297#_c_478_n 0.0171984f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A1_M1039_g N_A_27_297#_c_478_n 0.0214679f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_246 A1 N_A_27_297#_c_478_n 0.0381823f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_247 N_A1_c_267_n N_A_27_297#_c_478_n 0.0124751f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_248 A1 N_A_27_297#_c_482_n 0.00861209f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_249 N_A1_c_267_n N_A_27_297#_c_482_n 0.0024041f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_250 N_A1_c_267_n N_A_27_297#_c_484_n 0.00184277f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_251 N_A1_c_262_n N_Y_c_566_n 0.0110355f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_263_n N_Y_c_566_n 0.00893253f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_264_n N_Y_c_566_n 0.00893253f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_265_n N_Y_c_566_n 0.00510026f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_255 A1 N_Y_c_566_n 0.074891f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_256 N_A1_c_267_n N_Y_c_566_n 0.0197771f $X=5.515 $Y=1.17 $X2=0 $Y2=0
cc_257 N_A1_M1004_g N_VPWR_c_670_n 0.0119706f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A1_M1008_g N_VPWR_c_670_n 0.0102769f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A1_M1012_g N_VPWR_c_670_n 6.23635e-19 $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A1_M1008_g N_VPWR_c_671_n 0.0046653f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A1_M1012_g N_VPWR_c_671_n 0.00585385f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A1_M1012_g N_VPWR_c_672_n 0.00224235f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_M1039_g N_VPWR_c_672_n 0.00394726f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A1_M1039_g N_VPWR_c_673_n 9.92594e-19 $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A1_M1039_g N_VPWR_c_678_n 0.00583607f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A1_M1004_g N_VPWR_c_680_n 0.0046653f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A1_M1004_g N_VPWR_c_669_n 0.00804636f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A1_M1008_g N_VPWR_c_669_n 0.00789179f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A1_M1012_g N_VPWR_c_669_n 0.0111738f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A1_M1039_g N_VPWR_c_669_n 0.0116498f $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A1_c_262_n N_VGND_c_847_n 0.00366111f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_c_263_n N_VGND_c_847_n 0.00366111f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_c_264_n N_VGND_c_847_n 0.00366111f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_c_265_n N_VGND_c_847_n 0.00366111f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_275 N_A1_c_262_n N_VGND_c_860_n 0.00656615f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A1_c_263_n N_VGND_c_860_n 0.00524008f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A1_c_264_n N_VGND_c_860_n 0.00524008f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A1_c_265_n N_VGND_c_860_n 0.00557302f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_279 N_A1_c_262_n N_A_803_47#_c_977_n 0.00789149f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A1_c_263_n N_A_803_47#_c_977_n 0.00789149f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A1_c_264_n N_A_803_47#_c_977_n 0.00789149f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A1_c_265_n N_A_803_47#_c_977_n 0.0115259f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_283 N_A1_c_265_n N_A_1249_47#_c_1006_n 5.26688e-19 $X=5.61 $Y=1.01 $X2=0
+ $Y2=0
cc_284 A2 N_A3_c_396_n 0.00189259f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_285 A2 N_A3_c_397_n 0.00693886f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_286 N_A2_M1003_g N_A_27_297#_c_485_n 0.00792986f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A2_M1003_g N_A_27_297#_c_486_n 0.0156926f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A2_M1024_g N_A_27_297#_c_486_n 0.0146685f $X=6.59 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A2_c_331_n N_A_27_297#_c_486_n 0.00200188f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_290 A2 N_A_27_297#_c_486_n 0.0258363f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_291 N_A2_M1036_g N_A_27_297#_c_490_n 0.0146685f $X=7.01 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A2_c_331_n N_A_27_297#_c_490_n 0.00198468f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_293 N_A2_M1037_g N_A_27_297#_c_490_n 0.0167715f $X=7.43 $Y=1.985 $X2=0 $Y2=0
cc_294 A2 N_A_27_297#_c_490_n 0.0272427f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_295 N_A2_c_331_n N_A_27_297#_c_494_n 0.00211036f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_296 A2 N_A_27_297#_c_494_n 0.00901315f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_297 A2 N_A_27_297#_c_496_n 0.00813047f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_298 N_A2_c_328_n N_Y_c_566_n 5.26688e-19 $X=6.17 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A2_M1003_g N_VPWR_c_673_n 0.0146506f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A2_M1024_g N_VPWR_c_673_n 0.0101939f $X=6.59 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A2_M1036_g N_VPWR_c_673_n 6.0901e-19 $X=7.01 $Y=1.985 $X2=0 $Y2=0
cc_302 N_A2_M1024_g N_VPWR_c_674_n 0.0046653f $X=6.59 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A2_M1036_g N_VPWR_c_674_n 0.0046653f $X=7.01 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A2_M1024_g N_VPWR_c_675_n 6.0901e-19 $X=6.59 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A2_M1036_g N_VPWR_c_675_n 0.0128916f $X=7.01 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A2_M1037_g N_VPWR_c_675_n 0.0147873f $X=7.43 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A2_M1003_g N_VPWR_c_678_n 0.0046653f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A2_M1037_g N_VPWR_c_681_n 0.0046653f $X=7.43 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A2_M1003_g N_VPWR_c_669_n 0.00848713f $X=6.17 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A2_M1024_g N_VPWR_c_669_n 0.00789179f $X=6.59 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A2_M1036_g N_VPWR_c_669_n 0.00789179f $X=7.01 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A2_M1037_g N_VPWR_c_669_n 0.00921786f $X=7.43 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A2_c_328_n N_VGND_c_847_n 0.00366111f $X=6.17 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A2_c_329_n N_VGND_c_847_n 0.00366111f $X=6.59 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_c_330_n N_VGND_c_847_n 0.00366111f $X=7.01 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A2_c_331_n N_VGND_c_847_n 0.00366111f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_317 N_A2_c_331_n N_VGND_c_848_n 0.00294182f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_318 N_A2_c_328_n N_VGND_c_860_n 0.00562481f $X=6.17 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A2_c_329_n N_VGND_c_860_n 0.00524008f $X=6.59 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A2_c_330_n N_VGND_c_860_n 0.00524008f $X=7.01 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A2_c_331_n N_VGND_c_860_n 0.00656615f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_322 N_A2_c_328_n N_A_803_47#_c_977_n 0.0122055f $X=6.17 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A2_c_329_n N_A_803_47#_c_977_n 0.00789149f $X=6.59 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A2_c_330_n N_A_803_47#_c_977_n 0.00789149f $X=7.01 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A2_c_331_n N_A_803_47#_c_977_n 0.00789149f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_326 A2 N_A_803_47#_c_977_n 0.00288497f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_327 N_A2_c_328_n N_A_1249_47#_c_1006_n 0.00432658f $X=6.17 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_A2_c_329_n N_A_1249_47#_c_1006_n 0.00893253f $X=6.59 $Y=0.995 $X2=0
+ $Y2=0
cc_329 N_A2_c_330_n N_A_1249_47#_c_1006_n 0.00893253f $X=7.01 $Y=0.995 $X2=0
+ $Y2=0
cc_330 N_A2_c_331_n N_A_1249_47#_c_1006_n 0.0172648f $X=7.43 $Y=1.01 $X2=0 $Y2=0
cc_331 A2 N_A_1249_47#_c_1006_n 0.0636236f $X=7.49 $Y=1.105 $X2=0 $Y2=0
cc_332 N_A3_M1001_g N_A_27_297#_c_497_n 0.016242f $X=8.37 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A3_M1001_g N_A_27_297#_c_498_n 0.0168781f $X=8.37 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A3_M1007_g N_A_27_297#_c_498_n 0.0147751f $X=8.79 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A3_c_396_n N_A_27_297#_c_498_n 0.0019496f $X=9.63 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A3_c_397_n N_A_27_297#_c_498_n 0.024239f $X=9.805 $Y=1.177 $X2=0 $Y2=0
cc_337 N_A3_M1010_g N_A_27_297#_c_502_n 0.0147309f $X=9.21 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A3_M1020_g N_A_27_297#_c_502_n 0.0159832f $X=9.63 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A3_c_396_n N_A_27_297#_c_502_n 0.00562831f $X=9.63 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A3_c_397_n N_A_27_297#_c_502_n 0.0277486f $X=9.805 $Y=1.177 $X2=0 $Y2=0
cc_341 N_A3_c_398_n N_A_27_297#_c_502_n 0.00669658f $X=9.895 $Y=1.075 $X2=0
+ $Y2=0
cc_342 N_A3_c_396_n N_A_27_297#_c_507_n 0.00206078f $X=9.63 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A3_c_397_n N_A_27_297#_c_507_n 0.00848579f $X=9.805 $Y=1.177 $X2=0
+ $Y2=0
cc_344 N_A3_M1001_g N_VPWR_c_676_n 0.0301025f $X=8.37 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A3_M1007_g N_VPWR_c_676_n 0.0101939f $X=8.79 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A3_M1010_g N_VPWR_c_676_n 6.0901e-19 $X=9.21 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A3_M1007_g N_VPWR_c_677_n 6.0901e-19 $X=8.79 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A3_M1010_g N_VPWR_c_677_n 0.0101939f $X=9.21 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A3_M1020_g N_VPWR_c_677_n 0.0120895f $X=9.63 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A3_M1001_g N_VPWR_c_681_n 0.0046653f $X=8.37 $Y=1.985 $X2=0 $Y2=0
cc_351 N_A3_M1007_g N_VPWR_c_682_n 0.0046653f $X=8.79 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A3_M1010_g N_VPWR_c_682_n 0.0046653f $X=9.21 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A3_M1020_g N_VPWR_c_683_n 0.0046653f $X=9.63 $Y=1.985 $X2=0 $Y2=0
cc_354 N_A3_M1001_g N_VPWR_c_669_n 0.00934473f $X=8.37 $Y=1.985 $X2=0 $Y2=0
cc_355 N_A3_M1007_g N_VPWR_c_669_n 0.00789179f $X=8.79 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A3_M1010_g N_VPWR_c_669_n 0.00789179f $X=9.21 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A3_M1020_g N_VPWR_c_669_n 0.00886468f $X=9.63 $Y=1.985 $X2=0 $Y2=0
cc_358 A3 N_VGND_M1019_d 0.00961608f $X=9.81 $Y=0.765 $X2=0 $Y2=0
cc_359 N_A3_c_391_n N_VGND_c_848_n 0.00774571f $X=8.37 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A3_c_392_n N_VGND_c_848_n 5.08801e-19 $X=8.79 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A3_c_391_n N_VGND_c_849_n 5.08801e-19 $X=8.37 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A3_c_392_n N_VGND_c_849_n 0.00664421f $X=8.79 $Y=0.995 $X2=0 $Y2=0
cc_363 N_A3_c_393_n N_VGND_c_849_n 0.00666824f $X=9.21 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A3_c_394_n N_VGND_c_849_n 5.13014e-19 $X=9.63 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A3_c_393_n N_VGND_c_851_n 5.04142e-19 $X=9.21 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A3_c_394_n N_VGND_c_851_n 0.00754737f $X=9.63 $Y=0.995 $X2=0 $Y2=0
cc_367 A3 N_VGND_c_851_n 0.00937686f $X=9.81 $Y=0.765 $X2=0 $Y2=0
cc_368 N_A3_c_396_n N_VGND_c_851_n 0.00233751f $X=9.63 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A3_c_397_n N_VGND_c_851_n 0.00240088f $X=9.805 $Y=1.177 $X2=0 $Y2=0
cc_370 N_A3_c_391_n N_VGND_c_854_n 0.00339367f $X=8.37 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A3_c_392_n N_VGND_c_854_n 0.00339367f $X=8.79 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A3_c_393_n N_VGND_c_855_n 0.00339367f $X=9.21 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A3_c_394_n N_VGND_c_855_n 0.00505556f $X=9.63 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A3_c_391_n N_VGND_c_860_n 0.00394406f $X=8.37 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A3_c_392_n N_VGND_c_860_n 0.00394406f $X=8.79 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A3_c_393_n N_VGND_c_860_n 0.00394406f $X=9.21 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A3_c_394_n N_VGND_c_860_n 0.00850607f $X=9.63 $Y=0.995 $X2=0 $Y2=0
cc_378 A3 N_VGND_c_860_n 9.42702e-19 $X=9.81 $Y=0.765 $X2=0 $Y2=0
cc_379 N_A3_c_391_n N_A_1249_47#_c_1006_n 0.0141341f $X=8.37 $Y=0.995 $X2=0
+ $Y2=0
cc_380 N_A3_c_397_n N_A_1249_47#_c_1006_n 0.00833304f $X=9.805 $Y=1.177 $X2=0
+ $Y2=0
cc_381 N_A3_c_392_n N_A_1249_47#_c_1015_n 0.0119869f $X=8.79 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A3_c_393_n N_A_1249_47#_c_1015_n 0.0115547f $X=9.21 $Y=0.995 $X2=0
+ $Y2=0
cc_383 N_A3_c_396_n N_A_1249_47#_c_1015_n 0.00423243f $X=9.63 $Y=1.16 $X2=0
+ $Y2=0
cc_384 N_A3_c_397_n N_A_1249_47#_c_1015_n 0.0361307f $X=9.805 $Y=1.177 $X2=0
+ $Y2=0
cc_385 N_A3_c_396_n N_A_1249_47#_c_1019_n 0.00216182f $X=9.63 $Y=1.16 $X2=0
+ $Y2=0
cc_386 N_A3_c_397_n N_A_1249_47#_c_1019_n 0.00892733f $X=9.805 $Y=1.177 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_461_n N_Y_M1002_d 0.00325424f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_388 N_A_27_297#_c_461_n N_Y_M1027_d 0.00325424f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_389 N_A_27_297#_c_461_n N_Y_M1000_d 0.00325424f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_390 N_A_27_297#_c_461_n N_Y_M1031_d 0.00325424f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_391 N_A_27_297#_M1005_s N_Y_c_571_n 0.00465037f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_392 N_A_27_297#_c_461_n N_Y_c_571_n 0.0115975f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_393 N_A_27_297#_M1034_s N_Y_c_575_n 0.00677304f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_394 N_A_27_297#_c_461_n N_Y_c_575_n 0.00692481f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_395 N_A_27_297#_M1006_s N_Y_c_600_n 0.00458867f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_396 N_A_27_297#_c_461_n N_Y_c_600_n 0.0116113f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_397 N_A_27_297#_c_461_n N_Y_c_577_n 0.0157268f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_398 N_A_27_297#_c_461_n N_Y_c_583_n 0.0157268f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_399 N_A_27_297#_c_461_n N_Y_c_605_n 0.0157268f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_400 N_A_27_297#_M1034_s Y 0.00388422f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_461_n Y 0.0278073f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_402 N_A_27_297#_M1034_s Y 0.0011411f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_403 N_A_27_297#_c_474_n N_VPWR_M1004_s 0.00351323f $X=4.395 $Y=1.66 $X2=-0.19
+ $Y2=1.305
cc_404 N_A_27_297#_c_478_n N_VPWR_M1012_s 0.0150542f $X=5.64 $Y=1.66 $X2=0 $Y2=0
cc_405 N_A_27_297#_c_486_n N_VPWR_M1003_d 0.0034684f $X=6.715 $Y=1.66 $X2=0
+ $Y2=0
cc_406 N_A_27_297#_c_490_n N_VPWR_M1036_d 0.0034684f $X=7.555 $Y=1.66 $X2=0
+ $Y2=0
cc_407 N_A_27_297#_c_498_n N_VPWR_M1001_s 0.0035361f $X=8.915 $Y=1.66 $X2=0
+ $Y2=0
cc_408 N_A_27_297#_c_502_n N_VPWR_M1010_s 0.0035361f $X=9.755 $Y=1.66 $X2=0
+ $Y2=0
cc_409 N_A_27_297#_c_473_n N_VPWR_c_670_n 0.0358854f $X=3.62 $Y=2.255 $X2=0
+ $Y2=0
cc_410 N_A_27_297#_c_474_n N_VPWR_c_670_n 0.0170259f $X=4.395 $Y=1.66 $X2=0
+ $Y2=0
cc_411 N_A_27_297#_c_533_p N_VPWR_c_671_n 0.0113958f $X=4.48 $Y=1.96 $X2=0 $Y2=0
cc_412 N_A_27_297#_c_478_n N_VPWR_c_672_n 0.0456421f $X=5.64 $Y=1.66 $X2=0 $Y2=0
cc_413 N_A_27_297#_c_485_n N_VPWR_c_673_n 0.0207852f $X=5.725 $Y=1.96 $X2=0
+ $Y2=0
cc_414 N_A_27_297#_c_486_n N_VPWR_c_673_n 0.0170259f $X=6.715 $Y=1.66 $X2=0
+ $Y2=0
cc_415 N_A_27_297#_c_537_p N_VPWR_c_674_n 0.0113958f $X=6.8 $Y=1.96 $X2=0 $Y2=0
cc_416 N_A_27_297#_c_490_n N_VPWR_c_675_n 0.0171101f $X=7.555 $Y=1.66 $X2=0
+ $Y2=0
cc_417 N_A_27_297#_c_498_n N_VPWR_c_676_n 0.0170259f $X=8.915 $Y=1.66 $X2=0
+ $Y2=0
cc_418 N_A_27_297#_c_502_n N_VPWR_c_677_n 0.0170259f $X=9.755 $Y=1.66 $X2=0
+ $Y2=0
cc_419 N_A_27_297#_c_485_n N_VPWR_c_678_n 0.0116048f $X=5.725 $Y=1.96 $X2=0
+ $Y2=0
cc_420 N_A_27_297#_c_461_n N_VPWR_c_680_n 0.15191f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_421 N_A_27_297#_c_473_n N_VPWR_c_680_n 0.00931283f $X=3.62 $Y=2.255 $X2=0
+ $Y2=0
cc_422 N_A_27_297#_c_497_n N_VPWR_c_681_n 0.0116048f $X=7.64 $Y=1.96 $X2=0 $Y2=0
cc_423 N_A_27_297#_c_545_p N_VPWR_c_682_n 0.0113958f $X=9 $Y=1.96 $X2=0 $Y2=0
cc_424 N_A_27_297#_c_546_p N_VPWR_c_683_n 0.0116048f $X=9.84 $Y=1.96 $X2=0 $Y2=0
cc_425 N_A_27_297#_M1002_s N_VPWR_c_669_n 0.00211652f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_426 N_A_27_297#_M1005_s N_VPWR_c_669_n 0.00217615f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_427 N_A_27_297#_M1034_s N_VPWR_c_669_n 0.00217615f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_428 N_A_27_297#_M1006_s N_VPWR_c_669_n 0.00217615f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_429 N_A_27_297#_M1035_s N_VPWR_c_669_n 0.00477801f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_430 N_A_27_297#_M1008_d N_VPWR_c_669_n 0.00562358f $X=4.345 $Y=1.485 $X2=0
+ $Y2=0
cc_431 N_A_27_297#_M1039_d N_VPWR_c_669_n 0.0157359f $X=5.59 $Y=1.485 $X2=0
+ $Y2=0
cc_432 N_A_27_297#_M1024_s N_VPWR_c_669_n 0.00562358f $X=6.665 $Y=1.485 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_M1037_s N_VPWR_c_669_n 0.0279663f $X=7.505 $Y=1.485 $X2=0
+ $Y2=0
cc_434 N_A_27_297#_M1007_d N_VPWR_c_669_n 0.00562358f $X=8.865 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_A_27_297#_M1020_d N_VPWR_c_669_n 0.00525232f $X=9.705 $Y=1.485 $X2=0
+ $Y2=0
cc_436 N_A_27_297#_c_461_n N_VPWR_c_669_n 0.11894f $X=3.535 $Y=2.34 $X2=0 $Y2=0
cc_437 N_A_27_297#_c_473_n N_VPWR_c_669_n 0.00641762f $X=3.62 $Y=2.255 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_c_533_p N_VPWR_c_669_n 0.00646998f $X=4.48 $Y=1.96 $X2=0
+ $Y2=0
cc_439 N_A_27_297#_c_485_n N_VPWR_c_669_n 0.00646998f $X=5.725 $Y=1.96 $X2=0
+ $Y2=0
cc_440 N_A_27_297#_c_537_p N_VPWR_c_669_n 0.00646998f $X=6.8 $Y=1.96 $X2=0 $Y2=0
cc_441 N_A_27_297#_c_497_n N_VPWR_c_669_n 0.00646998f $X=7.64 $Y=1.96 $X2=0
+ $Y2=0
cc_442 N_A_27_297#_c_545_p N_VPWR_c_669_n 0.00646998f $X=9 $Y=1.96 $X2=0 $Y2=0
cc_443 N_A_27_297#_c_546_p N_VPWR_c_669_n 0.00646998f $X=9.84 $Y=1.96 $X2=0
+ $Y2=0
cc_444 N_Y_M1002_d N_VPWR_c_669_n 0.00219239f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_445 N_Y_M1027_d N_VPWR_c_669_n 0.00219239f $X=1.385 $Y=1.485 $X2=0 $Y2=0
cc_446 N_Y_M1000_d N_VPWR_c_669_n 0.00219239f $X=2.225 $Y=1.485 $X2=0 $Y2=0
cc_447 N_Y_M1031_d N_VPWR_c_669_n 0.00219239f $X=3.065 $Y=1.485 $X2=0 $Y2=0
cc_448 N_Y_c_566_n N_A_27_47#_M1028_s 0.00312766f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_449 N_Y_c_566_n N_A_27_47#_M1033_s 0.0102196f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_450 Y N_A_27_47#_c_802_n 0.00386389f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_451 N_Y_M1022_d N_A_27_47#_c_794_n 0.00314796f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_452 N_Y_M1032_d N_A_27_47#_c_794_n 0.00315945f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_453 N_Y_c_594_n N_A_27_47#_c_794_n 0.00849635f $X=2.28 $Y=0.805 $X2=0 $Y2=0
cc_454 N_Y_c_566_n N_A_27_47#_c_794_n 0.0721087f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_455 Y N_A_27_47#_c_794_n 0.00467444f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_456 N_Y_c_566_n N_VGND_c_847_n 0.00347243f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_457 N_Y_M1022_d N_VGND_c_860_n 0.00219239f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_458 N_Y_M1032_d N_VGND_c_860_n 0.00219239f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_459 N_Y_M1013_d N_VGND_c_860_n 0.00219239f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_460 N_Y_M1023_d N_VGND_c_860_n 0.00219239f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_461 N_Y_c_566_n N_VGND_c_860_n 0.0108733f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_462 N_Y_c_566_n N_A_803_47#_M1013_s 0.00488547f $X=5.4 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_463 N_Y_c_566_n N_A_803_47#_M1015_s 0.00337959f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_464 N_Y_M1013_d N_A_803_47#_c_977_n 0.00315945f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_465 N_Y_M1023_d N_A_803_47#_c_977_n 0.00316323f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_466 N_Y_c_566_n N_A_803_47#_c_977_n 0.0797617f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_467 N_Y_c_566_n N_A_1249_47#_c_1006_n 0.00461841f $X=5.4 $Y=0.72 $X2=0 $Y2=0
cc_468 N_A_27_47#_c_795_n N_VGND_M1014_s 0.00337587f $X=1.015 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_469 N_A_27_47#_c_802_n N_VGND_M1025_s 0.00337587f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_795_n N_VGND_c_845_n 0.0159625f $X=1.015 $Y=0.72 $X2=0 $Y2=0
cc_471 N_A_27_47#_c_802_n N_VGND_c_846_n 0.0159625f $X=1.855 $Y=0.72 $X2=0 $Y2=0
cc_472 N_A_27_47#_c_802_n N_VGND_c_847_n 0.00243651f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_826_p N_VGND_c_847_n 0.00894629f $X=1.94 $Y=0.465 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_794_n N_VGND_c_847_n 0.0780741f $X=3.62 $Y=0.38 $X2=0 $Y2=0
cc_475 N_A_27_47#_c_828_p N_VGND_c_852_n 0.01143f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_795_n N_VGND_c_852_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_795_n N_VGND_c_853_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_831_p N_VGND_c_853_n 0.0112274f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_479 N_A_27_47#_c_802_n N_VGND_c_853_n 0.00244309f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_M1014_d N_VGND_c_860_n 0.00368727f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_M1021_d N_VGND_c_860_n 0.00249348f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_M1038_d N_VGND_c_860_n 0.00236972f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_M1028_s N_VGND_c_860_n 0.00217615f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_M1033_s N_VGND_c_860_n 0.00211652f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_828_p N_VGND_c_860_n 0.00643448f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_486 N_A_27_47#_c_795_n N_VGND_c_860_n 0.00984256f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_831_p N_VGND_c_860_n 0.00643448f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_488 N_A_27_47#_c_802_n N_VGND_c_860_n 0.00987412f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_826_p N_VGND_c_860_n 0.00636368f $X=1.94 $Y=0.465 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_794_n N_VGND_c_860_n 0.0609512f $X=3.62 $Y=0.38 $X2=0 $Y2=0
cc_491 N_A_27_47#_c_794_n N_A_803_47#_c_977_n 0.0145425f $X=3.62 $Y=0.38 $X2=0
+ $Y2=0
cc_492 N_VGND_c_860_n N_A_803_47#_M1013_s 0.00211652f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_493 N_VGND_c_860_n N_A_803_47#_M1015_s 0.00217615f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_494 N_VGND_c_860_n N_A_803_47#_M1029_s 0.00332948f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_495 N_VGND_c_860_n N_A_803_47#_M1018_d 0.00217615f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_860_n N_A_803_47#_M1030_d 0.00211652f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_847_n N_A_803_47#_c_977_n 0.171536f $X=7.995 $Y=0 $X2=0 $Y2=0
cc_498 N_VGND_c_848_n N_A_803_47#_c_977_n 0.0137364f $X=8.16 $Y=0.38 $X2=0 $Y2=0
cc_499 N_VGND_c_860_n N_A_803_47#_c_977_n 0.133125f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_500 N_VGND_c_860_n N_A_1249_47#_M1016_s 0.00219239f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_501 N_VGND_c_860_n N_A_1249_47#_M1026_s 0.00219239f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_c_860_n N_A_1249_47#_M1009_s 0.00249348f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_503 N_VGND_c_860_n N_A_1249_47#_M1017_s 0.00405853f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_504 N_VGND_M1009_d N_A_1249_47#_c_1006_n 0.0105655f $X=8.035 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_VGND_c_847_n N_A_1249_47#_c_1006_n 0.00346265f $X=7.995 $Y=0 $X2=0
+ $Y2=0
cc_506 N_VGND_c_848_n N_A_1249_47#_c_1006_n 0.0206068f $X=8.16 $Y=0.38 $X2=0
+ $Y2=0
cc_507 N_VGND_c_854_n N_A_1249_47#_c_1006_n 0.00244309f $X=8.835 $Y=0 $X2=0
+ $Y2=0
cc_508 N_VGND_c_860_n N_A_1249_47#_c_1006_n 0.013978f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_854_n N_A_1249_47#_c_1031_n 0.0112274f $X=8.835 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_860_n N_A_1249_47#_c_1031_n 0.00643448f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_M1011_d N_A_1249_47#_c_1015_n 0.00337587f $X=8.865 $Y=0.235 $X2=0
+ $Y2=0
cc_512 N_VGND_c_849_n N_A_1249_47#_c_1015_n 0.0159625f $X=9 $Y=0.38 $X2=0 $Y2=0
cc_513 N_VGND_c_854_n N_A_1249_47#_c_1015_n 0.00244309f $X=8.835 $Y=0 $X2=0
+ $Y2=0
cc_514 N_VGND_c_855_n N_A_1249_47#_c_1015_n 0.00244309f $X=9.685 $Y=0 $X2=0
+ $Y2=0
cc_515 N_VGND_c_860_n N_A_1249_47#_c_1015_n 0.00984256f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_855_n N_A_1249_47#_c_1038_n 0.0112274f $X=9.685 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_860_n N_A_1249_47#_c_1038_n 0.00643448f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_518 N_A_803_47#_c_977_n N_A_1249_47#_M1016_s 0.00315945f $X=7.64 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_519 N_A_803_47#_c_977_n N_A_1249_47#_M1026_s 0.00316323f $X=7.64 $Y=0.38
+ $X2=0 $Y2=0
cc_520 N_A_803_47#_M1018_d N_A_1249_47#_c_1006_n 0.00337959f $X=6.665 $Y=0.235
+ $X2=0 $Y2=0
cc_521 N_A_803_47#_M1030_d N_A_1249_47#_c_1006_n 0.00724259f $X=7.505 $Y=0.235
+ $X2=0 $Y2=0
cc_522 N_A_803_47#_c_977_n N_A_1249_47#_c_1006_n 0.0797617f $X=7.64 $Y=0.38
+ $X2=0 $Y2=0

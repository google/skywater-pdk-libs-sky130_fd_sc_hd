* File: sky130_fd_sc_hd__dfbbp_1.pxi.spice
* Created: Tue Sep  1 19:02:43 2020
* 
x_PM_SKY130_FD_SC_HD__DFBBP_1%CLK N_CLK_c_257_n N_CLK_c_252_n N_CLK_M1037_g
+ N_CLK_c_258_n N_CLK_M1013_g N_CLK_c_253_n N_CLK_c_259_n CLK CLK N_CLK_c_255_n
+ N_CLK_c_256_n PM_SKY130_FD_SC_HD__DFBBP_1%CLK
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_27_47# N_A_27_47#_M1037_s N_A_27_47#_M1013_s
+ N_A_27_47#_M1014_g N_A_27_47#_M1000_g N_A_27_47#_c_297_n N_A_27_47#_M1032_g
+ N_A_27_47#_M1012_g N_A_27_47#_M1031_g N_A_27_47#_c_298_n N_A_27_47#_c_299_n
+ N_A_27_47#_M1024_g N_A_27_47#_c_301_n N_A_27_47#_c_302_n N_A_27_47#_c_303_n
+ N_A_27_47#_c_313_n N_A_27_47#_c_421_p N_A_27_47#_c_304_n N_A_27_47#_c_305_n
+ N_A_27_47#_c_306_n N_A_27_47#_c_316_n N_A_27_47#_c_317_n N_A_27_47#_c_318_n
+ N_A_27_47#_c_319_n N_A_27_47#_c_320_n N_A_27_47#_c_321_n N_A_27_47#_c_307_n
+ N_A_27_47#_c_323_n N_A_27_47#_c_324_n N_A_27_47#_c_325_n N_A_27_47#_c_326_n
+ N_A_27_47#_c_327_n PM_SKY130_FD_SC_HD__DFBBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DFBBP_1%D N_D_M1006_g N_D_M1020_g D D N_D_c_546_n
+ N_D_c_547_n PM_SKY130_FD_SC_HD__DFBBP_1%D
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_193_47# N_A_193_47#_M1014_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1016_g N_A_193_47#_c_585_n N_A_193_47#_c_586_n
+ N_A_193_47#_M1026_g N_A_193_47#_c_588_n N_A_193_47#_c_589_n
+ N_A_193_47#_M1027_g N_A_193_47#_M1018_g N_A_193_47#_c_590_n
+ N_A_193_47#_c_591_n N_A_193_47#_c_592_n N_A_193_47#_c_607_n
+ N_A_193_47#_c_608_n N_A_193_47#_c_593_n N_A_193_47#_c_594_n
+ N_A_193_47#_c_595_n N_A_193_47#_c_596_n N_A_193_47#_c_597_n
+ N_A_193_47#_c_598_n N_A_193_47#_c_599_n N_A_193_47#_c_600_n
+ N_A_193_47#_c_601_n N_A_193_47#_c_602_n PM_SKY130_FD_SC_HD__DFBBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_648_21# N_A_648_21#_M1023_d N_A_648_21#_M1005_d
+ N_A_648_21#_M1002_g N_A_648_21#_M1021_g N_A_648_21#_M1030_g
+ N_A_648_21#_c_802_n N_A_648_21#_M1003_g N_A_648_21#_c_811_n
+ N_A_648_21#_c_858_p N_A_648_21#_c_824_n N_A_648_21#_c_803_n
+ N_A_648_21#_c_804_n N_A_648_21#_c_805_n N_A_648_21#_c_813_n
+ N_A_648_21#_c_814_n N_A_648_21#_c_829_n N_A_648_21#_c_806_n
+ N_A_648_21#_c_807_n PM_SKY130_FD_SC_HD__DFBBP_1%A_648_21#
x_PM_SKY130_FD_SC_HD__DFBBP_1%SET_B N_SET_B_c_947_n N_SET_B_M1005_g
+ N_SET_B_M1029_g N_SET_B_M1025_g N_SET_B_M1010_g SET_B N_SET_B_c_953_n
+ N_SET_B_c_954_n N_SET_B_c_955_n N_SET_B_c_956_n N_SET_B_c_957_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%SET_B
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_474_413# N_A_474_413#_M1032_d
+ N_A_474_413#_M1016_d N_A_474_413#_M1023_g N_A_474_413#_M1022_g
+ N_A_474_413#_c_1088_n N_A_474_413#_c_1094_n N_A_474_413#_c_1084_n
+ N_A_474_413#_c_1079_n N_A_474_413#_c_1080_n N_A_474_413#_c_1081_n
+ N_A_474_413#_c_1082_n PM_SKY130_FD_SC_HD__DFBBP_1%A_474_413#
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_942_21# N_A_942_21#_M1017_s N_A_942_21#_M1034_s
+ N_A_942_21#_M1019_g N_A_942_21#_M1015_g N_A_942_21#_M1007_g
+ N_A_942_21#_M1036_g N_A_942_21#_c_1185_n N_A_942_21#_c_1186_n
+ N_A_942_21#_c_1194_n N_A_942_21#_c_1195_n N_A_942_21#_c_1187_n
+ N_A_942_21#_c_1188_n N_A_942_21#_c_1189_n N_A_942_21#_c_1198_n
+ N_A_942_21#_c_1199_n N_A_942_21#_c_1200_n N_A_942_21#_c_1201_n
+ N_A_942_21#_c_1190_n N_A_942_21#_c_1191_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%A_942_21#
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_1429_21# N_A_1429_21#_M1028_d
+ N_A_1429_21#_M1010_d N_A_1429_21#_M1009_g N_A_1429_21#_M1001_g
+ N_A_1429_21#_c_1344_n N_A_1429_21#_M1035_g N_A_1429_21#_M1039_g
+ N_A_1429_21#_c_1345_n N_A_1429_21#_c_1346_n N_A_1429_21#_c_1347_n
+ N_A_1429_21#_c_1348_n N_A_1429_21#_c_1349_n N_A_1429_21#_M1011_g
+ N_A_1429_21#_c_1359_n N_A_1429_21#_M1008_g N_A_1429_21#_c_1350_n
+ N_A_1429_21#_c_1351_n N_A_1429_21#_c_1360_n N_A_1429_21#_c_1361_n
+ N_A_1429_21#_c_1362_n N_A_1429_21#_c_1363_n N_A_1429_21#_c_1418_p
+ N_A_1429_21#_c_1465_p N_A_1429_21#_c_1389_n N_A_1429_21#_c_1352_n
+ N_A_1429_21#_c_1365_n N_A_1429_21#_c_1366_n N_A_1429_21#_c_1406_n
+ N_A_1429_21#_c_1382_n N_A_1429_21#_c_1409_n N_A_1429_21#_c_1353_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%A_1429_21#
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_1255_47# N_A_1255_47#_M1027_d
+ N_A_1255_47#_M1031_d N_A_1255_47#_M1028_g N_A_1255_47#_M1004_g
+ N_A_1255_47#_c_1533_n N_A_1255_47#_c_1536_n N_A_1255_47#_c_1522_n
+ N_A_1255_47#_c_1528_n N_A_1255_47#_c_1523_n N_A_1255_47#_c_1524_n
+ N_A_1255_47#_c_1525_n N_A_1255_47#_c_1526_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%A_1255_47#
x_PM_SKY130_FD_SC_HD__DFBBP_1%RESET_B N_RESET_B_M1034_g N_RESET_B_M1017_g
+ RESET_B N_RESET_B_c_1622_n RESET_B PM_SKY130_FD_SC_HD__DFBBP_1%RESET_B
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_2136_47# N_A_2136_47#_M1011_s
+ N_A_2136_47#_M1008_s N_A_2136_47#_M1033_g N_A_2136_47#_M1038_g
+ N_A_2136_47#_c_1658_n N_A_2136_47#_c_1664_n N_A_2136_47#_c_1659_n
+ N_A_2136_47#_c_1660_n N_A_2136_47#_c_1661_n N_A_2136_47#_c_1662_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%A_2136_47#
x_PM_SKY130_FD_SC_HD__DFBBP_1%VPWR N_VPWR_M1013_d N_VPWR_M1020_s N_VPWR_M1021_d
+ N_VPWR_M1015_d N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_M1034_d N_VPWR_M1008_d
+ N_VPWR_c_1709_n N_VPWR_c_1710_n N_VPWR_c_1711_n N_VPWR_c_1712_n
+ N_VPWR_c_1713_n N_VPWR_c_1714_n N_VPWR_c_1715_n N_VPWR_c_1716_n
+ N_VPWR_c_1717_n VPWR VPWR N_VPWR_c_1718_n N_VPWR_c_1719_n N_VPWR_c_1720_n
+ N_VPWR_c_1721_n N_VPWR_c_1722_n N_VPWR_c_1723_n N_VPWR_c_1724_n
+ N_VPWR_c_1708_n N_VPWR_c_1726_n N_VPWR_c_1727_n N_VPWR_c_1728_n
+ N_VPWR_c_1729_n N_VPWR_c_1730_n N_VPWR_c_1731_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%VPWR
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_381_47# N_A_381_47#_M1006_d N_A_381_47#_M1020_d
+ N_A_381_47#_c_1892_n N_A_381_47#_c_1893_n N_A_381_47#_c_1894_n
+ N_A_381_47#_c_1896_n N_A_381_47#_c_1897_n N_A_381_47#_c_1905_n
+ N_A_381_47#_c_1898_n PM_SKY130_FD_SC_HD__DFBBP_1%A_381_47#
x_PM_SKY130_FD_SC_HD__DFBBP_1%Q_N N_Q_N_M1035_d N_Q_N_M1039_d N_Q_N_c_1970_n
+ N_Q_N_c_1967_n Q_N Q_N Q_N N_Q_N_c_1969_n Q_N PM_SKY130_FD_SC_HD__DFBBP_1%Q_N
x_PM_SKY130_FD_SC_HD__DFBBP_1%Q N_Q_M1033_d N_Q_M1038_d N_Q_c_1997_n
+ N_Q_c_2000_n N_Q_c_1998_n Q Q Q PM_SKY130_FD_SC_HD__DFBBP_1%Q
x_PM_SKY130_FD_SC_HD__DFBBP_1%VGND N_VGND_M1037_d N_VGND_M1006_s N_VGND_M1002_d
+ N_VGND_M1003_s N_VGND_M1009_d N_VGND_M1017_d N_VGND_M1011_d N_VGND_c_2013_n
+ N_VGND_c_2014_n N_VGND_c_2015_n N_VGND_c_2016_n N_VGND_c_2017_n
+ N_VGND_c_2018_n N_VGND_c_2019_n N_VGND_c_2020_n N_VGND_c_2021_n
+ N_VGND_c_2022_n N_VGND_c_2023_n N_VGND_c_2024_n N_VGND_c_2025_n VGND VGND
+ N_VGND_c_2026_n N_VGND_c_2027_n N_VGND_c_2028_n N_VGND_c_2029_n
+ N_VGND_c_2030_n N_VGND_c_2031_n N_VGND_c_2032_n N_VGND_c_2033_n
+ N_VGND_c_2034_n N_VGND_c_2035_n PM_SKY130_FD_SC_HD__DFBBP_1%VGND
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_788_47# N_A_788_47#_M1029_d N_A_788_47#_M1019_d
+ N_A_788_47#_c_2201_n N_A_788_47#_c_2204_n N_A_788_47#_c_2211_n
+ PM_SKY130_FD_SC_HD__DFBBP_1%A_788_47#
x_PM_SKY130_FD_SC_HD__DFBBP_1%A_1545_47# N_A_1545_47#_M1025_d
+ N_A_1545_47#_M1036_d N_A_1545_47#_c_2236_n N_A_1545_47#_c_2232_n
+ N_A_1545_47#_c_2237_n PM_SKY130_FD_SC_HD__DFBBP_1%A_1545_47#
cc_1 VNB N_CLK_c_252_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_253_n 0.0229857f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK 0.0161955f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_CLK_c_255_n 0.0197972f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_CLK_c_256_n 0.0141141f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1014_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_297_n 0.01789f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_8 VNB N_A_27_47#_c_298_n 0.0124337f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.19
cc_9 VNB N_A_27_47#_c_299_n 0.00338665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1024_g 0.0470935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_301_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_302_n 0.00174761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_303_n 0.00789919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_304_n 0.00246672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_305_n 0.00418425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_306_n 0.0307531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_307_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_D_M1006_g 0.033904f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_19 VNB N_D_c_546_n 0.025724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_c_547_n 0.00418405f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_21 VNB N_A_193_47#_c_585_n 0.0133502f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_22 VNB N_A_193_47#_c_586_n 0.0045891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_193_47#_M1026_g 0.0197935f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_24 VNB N_A_193_47#_c_588_n 0.00878653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_c_589_n 0.018063f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB N_A_193_47#_c_590_n 0.00302353f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.19
cc_27 VNB N_A_193_47#_c_591_n 0.0315468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_592_n 0.00458399f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_29 VNB N_A_193_47#_c_593_n 0.0192255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_594_n 0.00568423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_595_n 0.00124359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_596_n 0.0216332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_597_n 0.00235584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_598_n 0.00201153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_599_n 0.00492219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_600_n 0.00147534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_601_n 0.0249207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_602_n 0.0159168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_648_21#_M1002_g 0.0393082f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_40 VNB N_A_648_21#_c_802_n 0.0192786f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_41 VNB N_A_648_21#_c_803_n 0.00190301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_648_21#_c_804_n 0.00419895f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_43 VNB N_A_648_21#_c_805_n 0.0116425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_648_21#_c_806_n 0.00589338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_648_21#_c_807_n 0.0321818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_SET_B_c_947_n 0.031114f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_47 VNB N_SET_B_M1005_g 0.00696335f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_48 VNB N_SET_B_M1029_g 0.0204338f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_49 VNB N_SET_B_M1025_g 0.0200444f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_50 VNB N_SET_B_M1010_g 0.00793898f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_51 VNB SET_B 0.00769431f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_52 VNB N_SET_B_c_953_n 0.0153139f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_53 VNB N_SET_B_c_954_n 0.00178135f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_54 VNB N_SET_B_c_955_n 0.00209085f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_55 VNB N_SET_B_c_956_n 0.00538514f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_56 VNB N_SET_B_c_957_n 0.0316983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_474_413#_M1023_g 0.0259951f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_58 VNB N_A_474_413#_c_1079_n 0.00755759f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_59 VNB N_A_474_413#_c_1080_n 0.00778508f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_60 VNB N_A_474_413#_c_1081_n 0.0040045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_474_413#_c_1082_n 0.0141708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_942_21#_M1019_g 0.0293266f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_63 VNB N_A_942_21#_M1036_g 0.0282197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_942_21#_c_1185_n 0.011477f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_65 VNB N_A_942_21#_c_1186_n 0.0020589f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_66 VNB N_A_942_21#_c_1187_n 0.00678122f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_67 VNB N_A_942_21#_c_1188_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_942_21#_c_1189_n 0.0214041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_942_21#_c_1190_n 0.0199031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_942_21#_c_1191_n 0.00545043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1429_21#_M1009_g 0.0441996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_72 VNB N_A_1429_21#_c_1344_n 0.0203843f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_73 VNB N_A_1429_21#_c_1345_n 0.0533873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1429_21#_c_1346_n 0.0159756f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_75 VNB N_A_1429_21#_c_1347_n 0.0081567f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_76 VNB N_A_1429_21#_c_1348_n 4.83176e-19 $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_77 VNB N_A_1429_21#_c_1349_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.19
cc_78 VNB N_A_1429_21#_c_1350_n 0.0183891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1429_21#_c_1351_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1429_21#_c_1352_n 0.00321658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1429_21#_c_1353_n 0.00364581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1255_47#_M1028_g 0.0224258f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_83 VNB N_A_1255_47#_c_1522_n 0.0117849f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_84 VNB N_A_1255_47#_c_1523_n 0.0114143f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_85 VNB N_A_1255_47#_c_1524_n 4.91252e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1255_47#_c_1525_n 0.00186712f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.53
cc_87 VNB N_A_1255_47#_c_1526_n 0.017672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_RESET_B_M1017_g 0.0348106f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_89 VNB RESET_B 0.00369111f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_90 VNB N_RESET_B_c_1622_n 0.0249908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_2136_47#_c_1658_n 0.00730219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2136_47#_c_1659_n 0.0051319f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_93 VNB N_A_2136_47#_c_1660_n 0.0256194f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_94 VNB N_A_2136_47#_c_1661_n 2.9362e-19 $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_95 VNB N_A_2136_47#_c_1662_n 0.0201161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VPWR_c_1708_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_381_47#_c_1892_n 0.0095618f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_98 VNB N_A_381_47#_c_1893_n 0.00434373f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_99 VNB N_A_381_47#_c_1894_n 0.00304926f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_100 VNB N_Q_N_c_1967_n 0.00373782f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_101 VNB Q_N 0.00139223f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_102 VNB N_Q_N_c_1969_n 0.00364683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_Q_c_1997_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_104 VNB N_Q_c_1998_n 0.0230748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB Q 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_106 VNB N_VGND_c_2013_n 4.09336e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_107 VNB N_VGND_c_2014_n 0.00527676f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.19
cc_108 VNB N_VGND_c_2015_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2016_n 0.00562135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2017_n 0.0024154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2018_n 0.00601958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2019_n 0.00262354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2020_n 0.0440436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2021_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2022_n 0.0391628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2023_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2024_n 0.0404697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2025_n 0.00372951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2026_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2027_n 0.0157985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2028_n 0.0537804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2029_n 0.0287938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2030_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2031_n 0.560087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2032_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2033_n 0.00545594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2034_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2035_n 0.00440331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VPB N_CLK_c_257_n 0.0118724f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_130 VPB N_CLK_c_258_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_131 VPB N_CLK_c_259_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_132 VPB CLK 0.0152683f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_133 VPB N_CLK_c_255_n 0.0102819f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_134 VPB N_A_27_47#_M1000_g 0.0364682f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_135 VPB N_A_27_47#_M1012_g 0.0215877f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_136 VPB N_A_27_47#_M1031_g 0.020906f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_137 VPB N_A_27_47#_c_298_n 0.0178865f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.19
cc_138 VPB N_A_27_47#_c_299_n 0.00403646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_313_n 0.00121034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_304_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_305_n 0.00245106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_316_n 0.0299356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_317_n 0.0135949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_318_n 0.00241912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_319_n 0.00875464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_320_n 0.00166365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_321_n 0.00361706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_27_47#_c_307_n 0.0115872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_323_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_27_47#_c_324_n 0.00575214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_27_47#_c_325_n 0.0282388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_27_47#_c_326_n 0.00514398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_27_47#_c_327_n 0.0125285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_D_M1020_g 0.05617f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_155 VPB N_D_c_546_n 0.00528891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_D_c_547_n 0.0069609f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_157 VPB N_A_193_47#_M1016_g 0.0461312f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_158 VPB N_A_193_47#_c_585_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_159 VPB N_A_193_47#_c_586_n 0.00324503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_193_47#_M1018_g 0.0222026f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_161 VPB N_A_193_47#_c_607_n 0.00384216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_193_47#_c_608_n 0.0287783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_193_47#_c_600_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_193_47#_c_602_n 0.0180923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_648_21#_M1002_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_166 VPB N_A_648_21#_M1021_g 0.0210587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_167 VPB N_A_648_21#_M1030_g 0.0317411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_168 VPB N_A_648_21#_c_811_n 0.0055347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_648_21#_c_804_n 0.00619168f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.53
cc_170 VPB N_A_648_21#_c_813_n 0.00575673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_648_21#_c_814_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_648_21#_c_807_n 0.00659461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_SET_B_M1005_g 0.0508831f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_174 VPB N_SET_B_M1010_g 0.0496547f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_175 VPB N_A_474_413#_M1022_g 0.0203673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_176 VPB N_A_474_413#_c_1084_n 0.0121994f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_177 VPB N_A_474_413#_c_1080_n 0.00799914f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_178 VPB N_A_474_413#_c_1081_n 0.00260739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_474_413#_c_1082_n 0.0165426f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_942_21#_M1015_g 0.0205161f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_181 VPB N_A_942_21#_M1007_g 0.0210664f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_182 VPB N_A_942_21#_c_1194_n 0.00188964f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_183 VPB N_A_942_21#_c_1195_n 0.0051323f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_184 VPB N_A_942_21#_c_1188_n 0.00162652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_942_21#_c_1189_n 0.0228551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_942_21#_c_1198_n 0.0329117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_942_21#_c_1199_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_942_21#_c_1200_n 0.00737873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_942_21#_c_1201_n 0.0033154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_942_21#_c_1190_n 0.026124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_942_21#_c_1191_n 0.00364078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1429_21#_M1009_g 0.0159543f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_193 VPB N_A_1429_21#_M1001_g 0.021027f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_194 VPB N_A_1429_21#_M1039_g 0.0245199f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_195 VPB N_A_1429_21#_c_1346_n 0.00445201f $X=-0.19 $Y=1.305 $X2=0.242
+ $Y2=1.235
cc_196 VPB N_A_1429_21#_c_1348_n 0.0132086f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_197 VPB N_A_1429_21#_c_1359_n 0.0188726f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.53
cc_198 VPB N_A_1429_21#_c_1360_n 0.0184285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1429_21#_c_1361_n 0.00421617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1429_21#_c_1362_n 0.0324865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1429_21#_c_1363_n 0.00304218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1429_21#_c_1352_n 0.00331499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1429_21#_c_1365_n 0.00717262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1429_21#_c_1366_n 0.0015513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1255_47#_M1004_g 0.021833f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_206 VPB N_A_1255_47#_c_1528_n 0.0118251f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_207 VPB N_A_1255_47#_c_1523_n 0.00584496f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_208 VPB N_A_1255_47#_c_1524_n 7.62954e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_1255_47#_c_1525_n 0.00126723f $X=-0.19 $Y=1.305 $X2=0.262
+ $Y2=1.53
cc_210 VPB N_A_1255_47#_c_1526_n 0.00899175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_RESET_B_M1034_g 0.0248365f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_212 VPB RESET_B 8.96726e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_213 VPB N_RESET_B_c_1622_n 0.00713638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_2136_47#_M1038_g 0.0243069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_A_2136_47#_c_1664_n 0.0133005f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_216 VPB N_A_2136_47#_c_1659_n 0.00518989f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_217 VPB N_A_2136_47#_c_1660_n 0.00561003f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_218 VPB N_VPWR_c_1709_n 0.00105566f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_219 VPB N_VPWR_c_1710_n 0.00617748f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.53
cc_220 VPB N_VPWR_c_1711_n 0.00313724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1712_n 0.00562862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1713_n 0.00361128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1714_n 0.0292737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1715_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1716_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1717_n 0.022998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1718_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1719_n 0.0156708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1720_n 0.0410023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1721_n 0.0591311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1722_n 0.0304826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1723_n 0.0291788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1724_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1708_n 0.0642133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1726_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1727_n 0.00546299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1728_n 0.00609488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1729_n 0.00928062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1730_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1731_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_381_47#_c_1892_n 0.00987822f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_242 VPB N_A_381_47#_c_1896_n 0.00977754f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=0.805
cc_243 VPB N_A_381_47#_c_1897_n 0.0033348f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_A_381_47#_c_1898_n 0.00183028f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_245 VPB N_Q_N_c_1970_n 0.00136543f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_246 VPB N_Q_N_c_1967_n 0.0037728f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_247 VPB Q_N 0.00756399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_Q_c_2000_n 0.00617439f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_249 VPB N_Q_c_1998_n 0.00721226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB Q 0.0341455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 N_CLK_c_252_n N_A_27_47#_M1014_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_252 CLK N_A_27_47#_M1014_g 3.10561e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_253 N_CLK_c_256_n N_A_27_47#_M1014_g 0.00508036f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_254 N_CLK_c_259_n N_A_27_47#_M1000_g 0.0276478f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_255 CLK N_A_27_47#_M1000_g 5.74563e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_256 N_CLK_c_255_n N_A_27_47#_M1000_g 0.00530931f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_257 N_CLK_c_252_n N_A_27_47#_c_302_n 0.00695828f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_258 N_CLK_c_253_n N_A_27_47#_c_302_n 0.00787672f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_259 CLK N_A_27_47#_c_302_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_260 N_CLK_c_253_n N_A_27_47#_c_303_n 0.00615556f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_261 CLK N_A_27_47#_c_303_n 0.0224836f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_262 N_CLK_c_255_n N_A_27_47#_c_303_n 7.46966e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_263 N_CLK_c_258_n N_A_27_47#_c_313_n 0.0128417f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_264 N_CLK_c_259_n N_A_27_47#_c_313_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_265 CLK N_A_27_47#_c_313_n 0.00728212f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_266 N_CLK_c_253_n N_A_27_47#_c_304_n 0.00189711f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_267 N_CLK_c_259_n N_A_27_47#_c_304_n 0.00440146f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_268 CLK N_A_27_47#_c_304_n 0.0517716f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_269 N_CLK_c_255_n N_A_27_47#_c_304_n 9.99163e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_270 N_CLK_c_256_n N_A_27_47#_c_304_n 0.00246927f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_271 N_CLK_c_258_n N_A_27_47#_c_316_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_272 N_CLK_c_259_n N_A_27_47#_c_316_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_273 CLK N_A_27_47#_c_316_n 0.0236377f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_274 N_CLK_c_255_n N_A_27_47#_c_316_n 5.90345e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_275 N_CLK_c_258_n N_A_27_47#_c_318_n 0.00103212f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_276 CLK N_A_27_47#_c_307_n 0.00162113f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_277 N_CLK_c_255_n N_A_27_47#_c_307_n 0.0169711f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_278 N_CLK_c_258_n N_VPWR_c_1709_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_279 N_CLK_c_258_n N_VPWR_c_1718_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_280 N_CLK_c_258_n N_VPWR_c_1708_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_281 N_CLK_c_252_n N_VGND_c_2013_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_282 N_CLK_c_252_n N_VGND_c_2026_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_283 N_CLK_c_253_n N_VGND_c_2026_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_284 N_CLK_c_252_n N_VGND_c_2031_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_297_n N_D_M1006_g 0.0212406f $X=2.305 $Y=0.705 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_305_n N_D_M1006_g 0.00124452f $X=2.415 $Y=0.87 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_324_n N_D_M1020_g 0.00106311f $X=2.745 $Y=1.74 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_305_n N_D_c_546_n 0.0010622f $X=2.415 $Y=0.87 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_306_n N_D_c_546_n 0.00140034f $X=2.415 $Y=0.87 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_305_n N_D_c_547_n 0.0453933f $X=2.415 $Y=0.87 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_306_n N_D_c_547_n 2.35131e-19 $X=2.415 $Y=0.87 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_317_n N_D_c_547_n 0.00488305f $X=2.39 $Y=1.87 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_324_n N_D_c_547_n 0.00408526f $X=2.745 $Y=1.74 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_317_n N_A_193_47#_M1000_d 6.81311e-19 $X=2.39 $Y=1.87 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1012_g N_A_193_47#_M1016_g 0.0190634f $X=2.715 $Y=2.275 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_305_n N_A_193_47#_M1016_g 0.00533835f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_317_n N_A_193_47#_M1016_g 0.00694689f $X=2.39 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_320_n N_A_193_47#_M1016_g 5.24592e-19 $X=2.68 $Y=1.87 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_323_n N_A_193_47#_M1016_g 0.0174486f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_324_n N_A_193_47#_M1016_g 0.01034f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_305_n N_A_193_47#_c_585_n 0.010154f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_319_n N_A_193_47#_c_585_n 3.83457e-19 $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_323_n N_A_193_47#_c_585_n 0.0212215f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_324_n N_A_193_47#_c_585_n 0.00655916f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_305_n N_A_193_47#_c_586_n 0.00203988f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_306_n N_A_193_47#_c_586_n 0.0224511f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_297_n N_A_193_47#_M1026_g 0.00868479f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_305_n N_A_193_47#_M1026_g 4.48322e-19 $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_306_n N_A_193_47#_M1026_g 0.021346f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1024_g N_A_193_47#_c_589_n 0.0129153f $X=6.745 $Y=0.415 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_321_n N_A_193_47#_M1018_g 0.00133927f $X=6.215 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_325_n N_A_193_47#_M1018_g 0.0192968f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_326_n N_A_193_47#_M1018_g 6.52047e-19 $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_299_n N_A_193_47#_c_590_n 2.62384e-19 $X=6.285 $Y=1.32 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_M1024_g N_A_193_47#_c_590_n 0.00307377f $X=6.745 $Y=0.415
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_299_n N_A_193_47#_c_591_n 0.0209335f $X=6.285 $Y=1.32 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_M1024_g N_A_193_47#_c_591_n 0.021369f $X=6.745 $Y=0.415 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_298_n N_A_193_47#_c_592_n 0.0110561f $X=6.67 $Y=1.32 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_299_n N_A_193_47#_c_592_n 0.00356667f $X=6.285 $Y=1.32 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_M1024_g N_A_193_47#_c_592_n 0.00622479f $X=6.745 $Y=0.415
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_326_n N_A_193_47#_c_592_n 0.00682571f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_298_n N_A_193_47#_c_607_n 0.00853911f $X=6.67 $Y=1.32 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_321_n N_A_193_47#_c_607_n 0.00483121f $X=6.215 $Y=1.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_325_n N_A_193_47#_c_607_n 5.88448e-19 $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_326_n N_A_193_47#_c_607_n 0.0168759f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_327_n N_A_193_47#_c_607_n 0.00347329f $X=6.15 $Y=1.575 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_298_n N_A_193_47#_c_608_n 0.0216716f $X=6.67 $Y=1.32 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_321_n N_A_193_47#_c_608_n 0.00219663f $X=6.215 $Y=1.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_325_n N_A_193_47#_c_608_n 0.0169266f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_326_n N_A_193_47#_c_608_n 0.00153059f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_305_n N_A_193_47#_c_593_n 0.0172997f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_306_n N_A_193_47#_c_593_n 0.00499487f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_M1014_g N_A_193_47#_c_594_n 0.00654297f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_302_n N_A_193_47#_c_594_n 0.00215463f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_304_n N_A_193_47#_c_594_n 0.00507209f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_305_n N_A_193_47#_c_595_n 0.00927819f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_325_n N_A_193_47#_c_596_n 2.37019e-19 $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_319_n N_A_193_47#_c_597_n 0.111198f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_305_n N_A_193_47#_c_598_n 4.97018e-19 $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_297_n N_A_193_47#_c_599_n 5.18238e-19 $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_305_n N_A_193_47#_c_599_n 0.020859f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_306_n N_A_193_47#_c_599_n 0.00153447f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_323_n N_A_193_47#_c_599_n 3.19045e-19 $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_324_n N_A_193_47#_c_599_n 0.00336529f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_298_n N_A_193_47#_c_600_n 3.23054e-19 $X=6.67 $Y=1.32 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_299_n N_A_193_47#_c_600_n 9.01357e-19 $X=6.285 $Y=1.32 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_326_n N_A_193_47#_c_600_n 0.00149027f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_305_n N_A_193_47#_c_601_n 0.00673428f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_M1014_g N_A_193_47#_c_602_n 0.0272829f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_302_n N_A_193_47#_c_602_n 0.0119128f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_421_p N_A_193_47#_c_602_n 0.00826951f $X=0.725 $Y=1.795
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_304_n N_A_193_47#_c_602_n 0.0701354f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_317_n N_A_193_47#_c_602_n 0.0245972f $X=2.39 $Y=1.87 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_318_n N_A_193_47#_c_602_n 0.00185693f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_305_n N_A_648_21#_M1002_g 5.35023e-19 $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_319_n N_A_648_21#_M1021_g 0.00197541f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_M1031_g N_A_648_21#_M1030_g 0.0164618f $X=6.21 $Y=2.275 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_299_n N_A_648_21#_M1030_g 0.00557961f $X=6.285 $Y=1.32 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_319_n N_A_648_21#_M1030_g 0.00750594f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_325_n N_A_648_21#_M1030_g 0.00910409f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_326_n N_A_648_21#_M1030_g 0.00264318f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_319_n N_A_648_21#_c_811_n 0.0240118f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_319_n N_A_648_21#_c_824_n 0.0279846f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_319_n N_A_648_21#_c_813_n 0.0141612f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_M1012_g N_A_648_21#_c_814_n 0.0161827f $X=2.715 $Y=2.275 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_319_n N_A_648_21#_c_814_n 0.00193898f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_323_n N_A_648_21#_c_814_n 0.00927772f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_319_n N_A_648_21#_c_829_n 0.00959465f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_299_n N_A_648_21#_c_807_n 0.00272432f $X=6.285 $Y=1.32 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1024_g N_SET_B_c_953_n 0.00574501f $X=6.745 $Y=0.415 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_M1012_g N_A_474_413#_c_1088_n 0.0091014f $X=2.715 $Y=2.275
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_317_n N_A_474_413#_c_1088_n 2.09728e-19 $X=2.39 $Y=1.87
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_319_n N_A_474_413#_c_1088_n 0.00506942f $X=6.07 $Y=1.87
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_320_n N_A_474_413#_c_1088_n 0.00303545f $X=2.68 $Y=1.87
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_323_n N_A_474_413#_c_1088_n 0.00186639f $X=2.745 $Y=1.74
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_324_n N_A_474_413#_c_1088_n 0.0152514f $X=2.745 $Y=1.74
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_305_n N_A_474_413#_c_1094_n 0.00631717f $X=2.415 $Y=0.87
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_306_n N_A_474_413#_c_1094_n 8.71498e-19 $X=2.415 $Y=0.87
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_M1012_g N_A_474_413#_c_1084_n 0.00650943f $X=2.715 $Y=2.275
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_305_n N_A_474_413#_c_1084_n 0.00666284f $X=2.415 $Y=0.87
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_319_n N_A_474_413#_c_1084_n 0.013911f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_320_n N_A_474_413#_c_1084_n 0.00149623f $X=2.68 $Y=1.87
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_323_n N_A_474_413#_c_1084_n 0.00203066f $X=2.745 $Y=1.74
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_324_n N_A_474_413#_c_1084_n 0.0282877f $X=2.745 $Y=1.74
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_c_319_n N_A_474_413#_c_1080_n 0.00350894f $X=6.07 $Y=1.87
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_305_n N_A_474_413#_c_1081_n 0.00728836f $X=2.415 $Y=0.87
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_319_n N_A_474_413#_c_1081_n 0.00456412f $X=6.07 $Y=1.87
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_319_n N_A_942_21#_M1015_g 0.00576309f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_319_n N_A_942_21#_c_1188_n 0.00477237f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_319_n N_A_942_21#_c_1189_n 3.78923e-19 $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_298_n N_A_942_21#_c_1198_n 0.00389341f $X=6.67 $Y=1.32 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_319_n N_A_942_21#_c_1198_n 0.0139809f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_321_n N_A_942_21#_c_1198_n 0.0255925f $X=6.215 $Y=1.87 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_325_n N_A_942_21#_c_1198_n 0.00176885f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_326_n N_A_942_21#_c_1198_n 0.00661378f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_327_n N_A_942_21#_c_1198_n 0.00371524f $X=6.15 $Y=1.575
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_319_n N_A_942_21#_c_1199_n 0.0264578f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_325_n N_A_942_21#_c_1199_n 7.96394e-19 $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_326_n N_A_942_21#_c_1199_n 0.00130051f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_327_n N_A_942_21#_c_1199_n 7.27878e-19 $X=6.15 $Y=1.575
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_319_n N_A_942_21#_c_1200_n 0.020032f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_325_n N_A_942_21#_c_1200_n 6.45403e-19 $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_326_n N_A_942_21#_c_1200_n 0.00461622f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_327_n N_A_942_21#_c_1200_n 0.00148716f $X=6.15 $Y=1.575
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_M1024_g N_A_1429_21#_M1009_g 0.0428045f $X=6.745 $Y=0.415
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_M1031_g N_A_1255_47#_c_1533_n 0.00496872f $X=6.21 $Y=2.275
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_321_n N_A_1255_47#_c_1533_n 0.00187313f $X=6.215 $Y=1.87
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_326_n N_A_1255_47#_c_1533_n 0.00141396f $X=6.15 $Y=1.74
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_M1024_g N_A_1255_47#_c_1536_n 0.0096406f $X=6.745 $Y=0.415
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_M1024_g N_A_1255_47#_c_1522_n 0.010696f $X=6.745 $Y=0.415
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_321_n N_A_1255_47#_c_1528_n 0.00214622f $X=6.215 $Y=1.87
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_326_n N_A_1255_47#_c_1528_n 0.0013353f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_M1024_g N_A_1255_47#_c_1524_n 0.00156831f $X=6.745 $Y=0.415
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_421_p N_VPWR_M1013_d 6.91013e-19 $X=0.725 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_415 N_A_27_47#_c_318_n N_VPWR_M1013_d 0.00195102f $X=0.84 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_416 N_A_27_47#_c_319_n N_VPWR_M1015_d 0.00670518f $X=6.07 $Y=1.87 $X2=0 $Y2=0
cc_417 N_A_27_47#_M1000_g N_VPWR_c_1709_n 0.00824303f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_313_n N_VPWR_c_1709_n 0.00355272f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_421_p N_VPWR_c_1709_n 0.0133497f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_316_n N_VPWR_c_1709_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_421 N_A_27_47#_c_318_n N_VPWR_c_1709_n 0.00347913f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1000_g N_VPWR_c_1710_n 0.00192109f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_317_n N_VPWR_c_1710_n 0.00177243f $X=2.39 $Y=1.87 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_319_n N_VPWR_c_1711_n 0.00160449f $X=6.07 $Y=1.87 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_319_n N_VPWR_c_1712_n 0.0137399f $X=6.07 $Y=1.87 $X2=0 $Y2=0
cc_426 N_A_27_47#_c_313_n N_VPWR_c_1718_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_427 N_A_27_47#_c_316_n N_VPWR_c_1718_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_428 N_A_27_47#_M1000_g N_VPWR_c_1719_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_M1012_g N_VPWR_c_1720_n 0.00367119f $X=2.715 $Y=2.275 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_M1031_g N_VPWR_c_1721_n 0.00424681f $X=6.21 $Y=2.275 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_326_n N_VPWR_c_1721_n 0.00254851f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1000_g N_VPWR_c_1708_n 0.00536257f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_M1012_g N_VPWR_c_1708_n 0.00562272f $X=2.715 $Y=2.275 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_M1031_g N_VPWR_c_1708_n 0.0061745f $X=6.21 $Y=2.275 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_313_n N_VPWR_c_1708_n 0.00396423f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_316_n N_VPWR_c_1708_n 0.00993215f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_317_n N_VPWR_c_1708_n 0.072214f $X=2.39 $Y=1.87 $X2=0 $Y2=0
cc_438 N_A_27_47#_c_318_n N_VPWR_c_1708_n 0.0144757f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_439 N_A_27_47#_c_319_n N_VPWR_c_1708_n 0.159156f $X=6.07 $Y=1.87 $X2=0 $Y2=0
cc_440 N_A_27_47#_c_320_n N_VPWR_c_1708_n 0.0160117f $X=2.68 $Y=1.87 $X2=0 $Y2=0
cc_441 N_A_27_47#_c_321_n N_VPWR_c_1708_n 0.0148451f $X=6.215 $Y=1.87 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_324_n N_VPWR_c_1708_n 3.19863e-19 $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_325_n N_VPWR_c_1708_n 3.05853e-19 $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_326_n N_VPWR_c_1708_n 0.00131252f $X=6.15 $Y=1.74 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_297_n N_A_381_47#_c_1893_n 0.00218515f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_305_n N_A_381_47#_c_1893_n 0.00795457f $X=2.415 $Y=0.87
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_c_317_n N_A_381_47#_c_1896_n 0.0306489f $X=2.39 $Y=1.87 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_320_n N_A_381_47#_c_1896_n 7.03109e-19 $X=2.68 $Y=1.87 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_324_n N_A_381_47#_c_1896_n 0.0093841f $X=2.745 $Y=1.74 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_317_n N_A_381_47#_c_1897_n 0.0155962f $X=2.39 $Y=1.87 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_297_n N_A_381_47#_c_1905_n 0.00395861f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_320_n N_A_381_47#_c_1898_n 8.67219e-19 $X=2.68 $Y=1.87 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_319_n A_892_329# 0.00105375f $X=6.07 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_454 N_A_27_47#_c_319_n A_1113_329# 0.00532504f $X=6.07 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_455 N_A_27_47#_c_302_n N_VGND_M1037_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_456 N_A_27_47#_M1014_g N_VGND_c_2013_n 0.00780198f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_302_n N_VGND_c_2013_n 0.0170164f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_458 N_A_27_47#_c_307_n N_VGND_c_2013_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_M1014_g N_VGND_c_2014_n 0.00303061f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_297_n N_VGND_c_2014_n 0.0012123f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_M1024_g N_VGND_c_2017_n 0.00126137f $X=6.745 $Y=0.415 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_297_n N_VGND_c_2020_n 0.00536249f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_305_n N_VGND_c_2020_n 0.00113905f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_M1024_g N_VGND_c_2024_n 0.00359964f $X=6.745 $Y=0.415 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_301_n N_VGND_c_2026_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_466 N_A_27_47#_c_302_n N_VGND_c_2026_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_M1014_g N_VGND_c_2027_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_M1037_s N_VGND_c_2031_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1014_g N_VGND_c_2031_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_297_n N_VGND_c_2031_n 0.00659009f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_M1024_g N_VGND_c_2031_n 0.00564067f $X=6.745 $Y=0.415 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_301_n N_VGND_c_2031_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_302_n N_VGND_c_2031_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_305_n N_VGND_c_2031_n 0.00119206f $X=2.415 $Y=0.87 $X2=0
+ $Y2=0
cc_475 N_D_M1020_g N_A_193_47#_c_586_n 0.0330166f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_476 N_D_c_546_n N_A_193_47#_c_586_n 0.00467503f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_477 N_D_c_547_n N_A_193_47#_c_586_n 0.00322877f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_478 N_D_M1006_g N_A_193_47#_c_593_n 0.00346149f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_479 N_D_c_546_n N_A_193_47#_c_593_n 0.00129446f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_480 N_D_c_547_n N_A_193_47#_c_593_n 0.0120982f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_481 N_D_M1006_g N_A_193_47#_c_602_n 0.00368527f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_482 N_D_M1020_g N_A_193_47#_c_602_n 0.00470206f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_483 N_D_M1020_g N_VPWR_c_1710_n 0.0117242f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_484 N_D_M1020_g N_VPWR_c_1720_n 0.0035268f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_485 N_D_M1020_g N_VPWR_c_1708_n 0.00398394f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_486 N_D_M1006_g N_A_381_47#_c_1892_n 0.00541608f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_487 N_D_M1020_g N_A_381_47#_c_1892_n 0.00781219f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_488 N_D_c_546_n N_A_381_47#_c_1892_n 0.00753248f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_489 N_D_c_547_n N_A_381_47#_c_1892_n 0.0486092f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_490 N_D_M1006_g N_A_381_47#_c_1893_n 0.0125506f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_491 N_D_c_546_n N_A_381_47#_c_1893_n 0.00213787f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_492 N_D_c_547_n N_A_381_47#_c_1893_n 0.0242664f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_493 N_D_M1020_g N_A_381_47#_c_1896_n 0.0130388f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_494 N_D_c_546_n N_A_381_47#_c_1896_n 0.00165939f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_495 N_D_c_547_n N_A_381_47#_c_1896_n 0.0285608f $X=1.835 $Y=1.17 $X2=0 $Y2=0
cc_496 N_D_M1020_g N_A_381_47#_c_1898_n 0.00259685f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_497 N_D_M1006_g N_VGND_c_2014_n 0.00945348f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_498 N_D_M1006_g N_VGND_c_2020_n 0.00339367f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_499 N_D_M1006_g N_VGND_c_2031_n 0.00393034f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_500 N_A_193_47#_M1026_g N_A_648_21#_M1002_g 0.0243315f $X=2.835 $Y=0.415
+ $X2=0 $Y2=0
cc_501 N_A_193_47#_c_588_n N_A_648_21#_M1002_g 0.0102862f $X=2.835 $Y=1.245
+ $X2=0 $Y2=0
cc_502 N_A_193_47#_c_599_n N_A_648_21#_M1002_g 0.0010488f $X=2.975 $Y=0.85 $X2=0
+ $Y2=0
cc_503 N_A_193_47#_c_601_n N_A_648_21#_M1002_g 0.021533f $X=2.895 $Y=0.93 $X2=0
+ $Y2=0
cc_504 N_A_193_47#_c_589_n N_A_648_21#_c_802_n 0.0187265f $X=6.2 $Y=0.705 $X2=0
+ $Y2=0
cc_505 N_A_193_47#_c_590_n N_A_648_21#_c_802_n 0.001702f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_506 N_A_193_47#_c_596_n N_A_648_21#_c_811_n 0.00196084f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_507 N_A_193_47#_c_596_n N_A_648_21#_c_824_n 0.00348372f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_508 N_A_193_47#_c_596_n N_A_648_21#_c_803_n 0.00165548f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_509 N_A_193_47#_c_596_n N_A_648_21#_c_804_n 0.016449f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_510 N_A_193_47#_c_596_n N_A_648_21#_c_805_n 0.00907541f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_511 N_A_193_47#_c_596_n N_A_648_21#_c_813_n 8.24776e-19 $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_512 N_A_193_47#_c_596_n N_A_648_21#_c_829_n 6.83984e-19 $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_513 N_A_193_47#_c_590_n N_A_648_21#_c_806_n 0.0111636f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_514 N_A_193_47#_c_591_n N_A_648_21#_c_806_n 9.14426e-19 $X=6.325 $Y=0.87
+ $X2=0 $Y2=0
cc_515 N_A_193_47#_c_592_n N_A_648_21#_c_806_n 0.00462764f $X=6.642 $Y=1.305
+ $X2=0 $Y2=0
cc_516 N_A_193_47#_c_596_n N_A_648_21#_c_806_n 0.0153364f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_517 N_A_193_47#_c_600_n N_A_648_21#_c_806_n 0.00129536f $X=6.215 $Y=1.19
+ $X2=0 $Y2=0
cc_518 N_A_193_47#_c_590_n N_A_648_21#_c_807_n 5.13187e-19 $X=6.325 $Y=0.87
+ $X2=0 $Y2=0
cc_519 N_A_193_47#_c_591_n N_A_648_21#_c_807_n 0.0187265f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_520 N_A_193_47#_c_592_n N_A_648_21#_c_807_n 0.00174717f $X=6.642 $Y=1.305
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_c_596_n N_A_648_21#_c_807_n 0.00365485f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_522 N_A_193_47#_c_600_n N_A_648_21#_c_807_n 6.8647e-19 $X=6.215 $Y=1.19 $X2=0
+ $Y2=0
cc_523 N_A_193_47#_c_596_n N_SET_B_c_947_n 0.00392015f $X=6.07 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_524 N_A_193_47#_c_596_n N_SET_B_M1005_g 0.0011704f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_525 N_A_193_47#_c_596_n SET_B 0.00590244f $X=6.07 $Y=1.19 $X2=0 $Y2=0
cc_526 N_A_193_47#_c_590_n N_SET_B_c_953_n 0.0194369f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_c_591_n N_SET_B_c_953_n 0.0023282f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_528 N_A_193_47#_c_592_n N_SET_B_c_953_n 0.0053562f $X=6.642 $Y=1.305 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_c_596_n N_SET_B_c_953_n 0.158115f $X=6.07 $Y=1.19 $X2=0 $Y2=0
cc_530 N_A_193_47#_c_600_n N_SET_B_c_953_n 0.0254944f $X=6.215 $Y=1.19 $X2=0
+ $Y2=0
cc_531 N_A_193_47#_c_596_n N_SET_B_c_954_n 0.0265121f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_532 N_A_193_47#_c_596_n N_A_474_413#_M1023_g 0.00188875f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_533 N_A_193_47#_M1016_g N_A_474_413#_c_1088_n 0.00277448f $X=2.295 $Y=2.275
+ $X2=0 $Y2=0
cc_534 N_A_193_47#_M1026_g N_A_474_413#_c_1094_n 0.00882839f $X=2.835 $Y=0.415
+ $X2=0 $Y2=0
cc_535 N_A_193_47#_c_593_n N_A_474_413#_c_1094_n 0.00575474f $X=2.83 $Y=0.85
+ $X2=0 $Y2=0
cc_536 N_A_193_47#_c_598_n N_A_474_413#_c_1094_n 0.00258895f $X=2.975 $Y=0.85
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_c_599_n N_A_474_413#_c_1094_n 0.0182033f $X=2.975 $Y=0.85
+ $X2=0 $Y2=0
cc_538 N_A_193_47#_c_601_n N_A_474_413#_c_1094_n 5.24271e-19 $X=2.895 $Y=0.93
+ $X2=0 $Y2=0
cc_539 N_A_193_47#_M1016_g N_A_474_413#_c_1084_n 8.73767e-19 $X=2.295 $Y=2.275
+ $X2=0 $Y2=0
cc_540 N_A_193_47#_c_597_n N_A_474_413#_c_1084_n 3.06883e-19 $X=3.12 $Y=1.19
+ $X2=0 $Y2=0
cc_541 N_A_193_47#_M1026_g N_A_474_413#_c_1079_n 2.58936e-19 $X=2.835 $Y=0.415
+ $X2=0 $Y2=0
cc_542 N_A_193_47#_c_588_n N_A_474_413#_c_1079_n 0.00144384f $X=2.835 $Y=1.245
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_c_596_n N_A_474_413#_c_1079_n 0.0152458f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_544 N_A_193_47#_c_598_n N_A_474_413#_c_1079_n 0.0143395f $X=2.975 $Y=0.85
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_599_n N_A_474_413#_c_1079_n 0.0251282f $X=2.975 $Y=0.85
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_601_n N_A_474_413#_c_1079_n 0.00218717f $X=2.895 $Y=0.93
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_c_596_n N_A_474_413#_c_1080_n 0.0384689f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_c_588_n N_A_474_413#_c_1081_n 0.00268821f $X=2.835 $Y=1.245
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_596_n N_A_474_413#_c_1081_n 0.0110554f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_550 N_A_193_47#_c_597_n N_A_474_413#_c_1081_n 0.0060147f $X=3.12 $Y=1.19
+ $X2=0 $Y2=0
cc_551 N_A_193_47#_c_599_n N_A_474_413#_c_1081_n 0.00391072f $X=2.975 $Y=0.85
+ $X2=0 $Y2=0
cc_552 N_A_193_47#_c_601_n N_A_474_413#_c_1081_n 5.70501e-19 $X=2.895 $Y=0.93
+ $X2=0 $Y2=0
cc_553 N_A_193_47#_c_596_n N_A_474_413#_c_1082_n 0.00386813f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_554 N_A_193_47#_c_596_n N_A_942_21#_M1019_g 0.00150073f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_555 N_A_193_47#_c_596_n N_A_942_21#_c_1188_n 0.0122882f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_556 N_A_193_47#_c_596_n N_A_942_21#_c_1189_n 0.00603655f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_557 N_A_193_47#_c_592_n N_A_942_21#_c_1198_n 0.00715591f $X=6.642 $Y=1.305
+ $X2=0 $Y2=0
cc_558 N_A_193_47#_c_607_n N_A_942_21#_c_1198_n 0.0157692f $X=6.66 $Y=1.74 $X2=0
+ $Y2=0
cc_559 N_A_193_47#_c_608_n N_A_942_21#_c_1198_n 0.00184742f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_560 N_A_193_47#_c_596_n N_A_942_21#_c_1198_n 0.014133f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_561 N_A_193_47#_c_600_n N_A_942_21#_c_1198_n 0.027417f $X=6.215 $Y=1.19 $X2=0
+ $Y2=0
cc_562 N_A_193_47#_c_596_n N_A_942_21#_c_1199_n 0.0276968f $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_563 N_A_193_47#_c_607_n N_A_942_21#_c_1200_n 0.00264766f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_564 N_A_193_47#_c_596_n N_A_942_21#_c_1200_n 0.00618009f $X=6.07 $Y=1.19
+ $X2=0 $Y2=0
cc_565 N_A_193_47#_c_607_n N_A_1429_21#_M1009_g 3.51933e-19 $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_566 N_A_193_47#_M1018_g N_A_1429_21#_c_1362_n 0.0162278f $X=6.63 $Y=2.275
+ $X2=0 $Y2=0
cc_567 N_A_193_47#_c_608_n N_A_1429_21#_c_1362_n 0.00879184f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_568 N_A_193_47#_M1018_g N_A_1255_47#_c_1533_n 0.00935459f $X=6.63 $Y=2.275
+ $X2=0 $Y2=0
cc_569 N_A_193_47#_c_607_n N_A_1255_47#_c_1533_n 0.00669245f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_570 N_A_193_47#_c_608_n N_A_1255_47#_c_1533_n 0.0028948f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_571 N_A_193_47#_c_590_n N_A_1255_47#_c_1536_n 0.00390894f $X=6.325 $Y=0.87
+ $X2=0 $Y2=0
cc_572 N_A_193_47#_c_591_n N_A_1255_47#_c_1536_n 0.00184507f $X=6.325 $Y=0.87
+ $X2=0 $Y2=0
cc_573 N_A_193_47#_c_592_n N_A_1255_47#_c_1536_n 0.00315233f $X=6.642 $Y=1.305
+ $X2=0 $Y2=0
cc_574 N_A_193_47#_c_590_n N_A_1255_47#_c_1522_n 0.0117718f $X=6.325 $Y=0.87
+ $X2=0 $Y2=0
cc_575 N_A_193_47#_c_592_n N_A_1255_47#_c_1522_n 0.00837612f $X=6.642 $Y=1.305
+ $X2=0 $Y2=0
cc_576 N_A_193_47#_c_600_n N_A_1255_47#_c_1522_n 6.65017e-19 $X=6.215 $Y=1.19
+ $X2=0 $Y2=0
cc_577 N_A_193_47#_M1018_g N_A_1255_47#_c_1528_n 0.00655877f $X=6.63 $Y=2.275
+ $X2=0 $Y2=0
cc_578 N_A_193_47#_c_607_n N_A_1255_47#_c_1528_n 0.0359925f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_579 N_A_193_47#_c_608_n N_A_1255_47#_c_1528_n 0.00212049f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_580 N_A_193_47#_c_592_n N_A_1255_47#_c_1524_n 0.00588724f $X=6.642 $Y=1.305
+ $X2=0 $Y2=0
cc_581 N_A_193_47#_c_607_n N_A_1255_47#_c_1524_n 0.00820578f $X=6.66 $Y=1.74
+ $X2=0 $Y2=0
cc_582 N_A_193_47#_c_600_n N_A_1255_47#_c_1524_n 2.68785e-19 $X=6.215 $Y=1.19
+ $X2=0 $Y2=0
cc_583 N_A_193_47#_c_602_n N_VPWR_c_1709_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_584 N_A_193_47#_M1016_g N_VPWR_c_1710_n 0.00112467f $X=2.295 $Y=2.275 $X2=0
+ $Y2=0
cc_585 N_A_193_47#_c_602_n N_VPWR_c_1710_n 0.0243614f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_586 N_A_193_47#_c_602_n N_VPWR_c_1719_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_587 N_A_193_47#_M1016_g N_VPWR_c_1720_n 0.00541732f $X=2.295 $Y=2.275 $X2=0
+ $Y2=0
cc_588 N_A_193_47#_M1018_g N_VPWR_c_1721_n 0.00367119f $X=6.63 $Y=2.275 $X2=0
+ $Y2=0
cc_589 N_A_193_47#_M1016_g N_VPWR_c_1708_n 0.00622656f $X=2.295 $Y=2.275 $X2=0
+ $Y2=0
cc_590 N_A_193_47#_M1018_g N_VPWR_c_1708_n 0.00567418f $X=6.63 $Y=2.275 $X2=0
+ $Y2=0
cc_591 N_A_193_47#_c_602_n N_VPWR_c_1708_n 0.00409094f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_592 N_A_193_47#_c_593_n N_A_381_47#_c_1892_n 0.0148981f $X=2.83 $Y=0.85 $X2=0
+ $Y2=0
cc_593 N_A_193_47#_c_594_n N_A_381_47#_c_1892_n 0.00137704f $X=1.3 $Y=0.85 $X2=0
+ $Y2=0
cc_594 N_A_193_47#_c_602_n N_A_381_47#_c_1892_n 0.0733768f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_595 N_A_193_47#_c_593_n N_A_381_47#_c_1893_n 0.0206043f $X=2.83 $Y=0.85 $X2=0
+ $Y2=0
cc_596 N_A_193_47#_c_599_n N_A_381_47#_c_1893_n 0.00215645f $X=2.975 $Y=0.85
+ $X2=0 $Y2=0
cc_597 N_A_193_47#_c_593_n N_A_381_47#_c_1894_n 0.00431451f $X=2.83 $Y=0.85
+ $X2=0 $Y2=0
cc_598 N_A_193_47#_c_594_n N_A_381_47#_c_1894_n 0.00142577f $X=1.3 $Y=0.85 $X2=0
+ $Y2=0
cc_599 N_A_193_47#_c_602_n N_A_381_47#_c_1894_n 0.0152139f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_600 N_A_193_47#_M1016_g N_A_381_47#_c_1896_n 0.00141994f $X=2.295 $Y=2.275
+ $X2=0 $Y2=0
cc_601 N_A_193_47#_c_602_n N_A_381_47#_c_1897_n 0.0127262f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_602 N_A_193_47#_M1016_g N_A_381_47#_c_1898_n 0.00735844f $X=2.295 $Y=2.275
+ $X2=0 $Y2=0
cc_603 N_A_193_47#_c_593_n N_VGND_c_2014_n 0.00130587f $X=2.83 $Y=0.85 $X2=0
+ $Y2=0
cc_604 N_A_193_47#_c_602_n N_VGND_c_2014_n 0.00885868f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_605 N_A_193_47#_c_596_n N_VGND_c_2015_n 9.89759e-19 $X=6.07 $Y=1.19 $X2=0
+ $Y2=0
cc_606 N_A_193_47#_c_589_n N_VGND_c_2016_n 0.00174046f $X=6.2 $Y=0.705 $X2=0
+ $Y2=0
cc_607 N_A_193_47#_M1026_g N_VGND_c_2020_n 0.00359964f $X=2.835 $Y=0.415 $X2=0
+ $Y2=0
cc_608 N_A_193_47#_c_589_n N_VGND_c_2024_n 0.00435972f $X=6.2 $Y=0.705 $X2=0
+ $Y2=0
cc_609 N_A_193_47#_c_590_n N_VGND_c_2024_n 0.00288727f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_610 N_A_193_47#_c_591_n N_VGND_c_2024_n 2.15978e-19 $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_611 N_A_193_47#_c_602_n N_VGND_c_2027_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_612 N_A_193_47#_M1014_d N_VGND_c_2031_n 0.0033946f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_613 N_A_193_47#_M1026_g N_VGND_c_2031_n 0.00559644f $X=2.835 $Y=0.415 $X2=0
+ $Y2=0
cc_614 N_A_193_47#_c_589_n N_VGND_c_2031_n 0.00616197f $X=6.2 $Y=0.705 $X2=0
+ $Y2=0
cc_615 N_A_193_47#_c_590_n N_VGND_c_2031_n 0.00224883f $X=6.325 $Y=0.87 $X2=0
+ $Y2=0
cc_616 N_A_193_47#_c_593_n N_VGND_c_2031_n 0.0709836f $X=2.83 $Y=0.85 $X2=0
+ $Y2=0
cc_617 N_A_193_47#_c_594_n N_VGND_c_2031_n 0.0151433f $X=1.3 $Y=0.85 $X2=0 $Y2=0
cc_618 N_A_193_47#_c_598_n N_VGND_c_2031_n 0.015297f $X=2.975 $Y=0.85 $X2=0
+ $Y2=0
cc_619 N_A_193_47#_c_602_n N_VGND_c_2031_n 0.00372614f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_620 N_A_193_47#_c_599_n A_582_47# 8.80342e-19 $X=2.975 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_621 N_A_648_21#_M1002_g N_SET_B_c_947_n 0.0190011f $X=3.315 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_622 N_A_648_21#_M1002_g N_SET_B_M1005_g 0.0137896f $X=3.315 $Y=0.445 $X2=0
+ $Y2=0
cc_623 N_A_648_21#_M1021_g N_SET_B_M1005_g 0.0101628f $X=3.315 $Y=2.275 $X2=0
+ $Y2=0
cc_624 N_A_648_21#_c_811_n N_SET_B_M1005_g 0.0159332f $X=4.09 $Y=1.91 $X2=0
+ $Y2=0
cc_625 N_A_648_21#_c_858_p N_SET_B_M1005_g 0.00507112f $X=4.175 $Y=2.21 $X2=0
+ $Y2=0
cc_626 N_A_648_21#_c_813_n N_SET_B_M1005_g 0.00473578f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_627 N_A_648_21#_c_814_n N_SET_B_M1005_g 0.020182f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_628 N_A_648_21#_M1002_g N_SET_B_M1029_g 0.0156014f $X=3.315 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_A_648_21#_c_803_n N_SET_B_M1029_g 5.56585e-19 $X=4.605 $Y=1.065 $X2=0
+ $Y2=0
cc_630 N_A_648_21#_M1002_g SET_B 0.00118793f $X=3.315 $Y=0.445 $X2=0 $Y2=0
cc_631 N_A_648_21#_c_803_n SET_B 0.00825406f $X=4.605 $Y=1.065 $X2=0 $Y2=0
cc_632 N_A_648_21#_M1023_d N_SET_B_c_953_n 5.1491e-19 $X=4.44 $Y=0.235 $X2=0
+ $Y2=0
cc_633 N_A_648_21#_c_802_n N_SET_B_c_953_n 0.00507207f $X=5.725 $Y=0.985 $X2=0
+ $Y2=0
cc_634 N_A_648_21#_c_803_n N_SET_B_c_953_n 0.0208059f $X=4.605 $Y=1.065 $X2=0
+ $Y2=0
cc_635 N_A_648_21#_c_805_n N_SET_B_c_953_n 0.0214137f $X=5.5 $Y=0.98 $X2=0 $Y2=0
cc_636 N_A_648_21#_c_806_n N_SET_B_c_953_n 0.0108883f $X=5.665 $Y=0.98 $X2=0
+ $Y2=0
cc_637 N_A_648_21#_c_803_n N_SET_B_c_954_n 0.00230334f $X=4.605 $Y=1.065 $X2=0
+ $Y2=0
cc_638 N_A_648_21#_c_803_n N_A_474_413#_M1023_g 0.00722888f $X=4.605 $Y=1.065
+ $X2=0 $Y2=0
cc_639 N_A_648_21#_c_804_n N_A_474_413#_M1023_g 0.00191659f $X=4.605 $Y=1.785
+ $X2=0 $Y2=0
cc_640 N_A_648_21#_c_824_n N_A_474_413#_M1022_g 0.0126303f $X=4.52 $Y=1.91 $X2=0
+ $Y2=0
cc_641 N_A_648_21#_M1021_g N_A_474_413#_c_1088_n 0.00191115f $X=3.315 $Y=2.275
+ $X2=0 $Y2=0
cc_642 N_A_648_21#_M1002_g N_A_474_413#_c_1094_n 0.00797698f $X=3.315 $Y=0.445
+ $X2=0 $Y2=0
cc_643 N_A_648_21#_M1002_g N_A_474_413#_c_1084_n 0.0154362f $X=3.315 $Y=0.445
+ $X2=0 $Y2=0
cc_644 N_A_648_21#_c_813_n N_A_474_413#_c_1084_n 0.0330453f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_645 N_A_648_21#_M1002_g N_A_474_413#_c_1079_n 0.0153158f $X=3.315 $Y=0.445
+ $X2=0 $Y2=0
cc_646 N_A_648_21#_c_811_n N_A_474_413#_c_1080_n 0.0141289f $X=4.09 $Y=1.91
+ $X2=0 $Y2=0
cc_647 N_A_648_21#_c_824_n N_A_474_413#_c_1080_n 0.00218253f $X=4.52 $Y=1.91
+ $X2=0 $Y2=0
cc_648 N_A_648_21#_c_804_n N_A_474_413#_c_1080_n 0.0246731f $X=4.605 $Y=1.785
+ $X2=0 $Y2=0
cc_649 N_A_648_21#_c_829_n N_A_474_413#_c_1080_n 0.00650509f $X=4.175 $Y=1.87
+ $X2=0 $Y2=0
cc_650 N_A_648_21#_M1002_g N_A_474_413#_c_1081_n 0.0106244f $X=3.315 $Y=0.445
+ $X2=0 $Y2=0
cc_651 N_A_648_21#_c_813_n N_A_474_413#_c_1081_n 0.0169621f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_652 N_A_648_21#_c_814_n N_A_474_413#_c_1081_n 0.00119732f $X=3.425 $Y=1.74
+ $X2=0 $Y2=0
cc_653 N_A_648_21#_c_804_n N_A_474_413#_c_1082_n 0.0092978f $X=4.605 $Y=1.785
+ $X2=0 $Y2=0
cc_654 N_A_648_21#_c_829_n N_A_474_413#_c_1082_n 9.09922e-19 $X=4.175 $Y=1.87
+ $X2=0 $Y2=0
cc_655 N_A_648_21#_c_803_n N_A_942_21#_M1019_g 0.00955091f $X=4.605 $Y=1.065
+ $X2=0 $Y2=0
cc_656 N_A_648_21#_c_804_n N_A_942_21#_M1019_g 0.00587629f $X=4.605 $Y=1.785
+ $X2=0 $Y2=0
cc_657 N_A_648_21#_c_805_n N_A_942_21#_M1019_g 0.00930678f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_658 N_A_648_21#_c_806_n N_A_942_21#_M1019_g 0.00136887f $X=5.665 $Y=0.98
+ $X2=0 $Y2=0
cc_659 N_A_648_21#_c_807_n N_A_942_21#_M1019_g 0.00197459f $X=5.665 $Y=1.15
+ $X2=0 $Y2=0
cc_660 N_A_648_21#_M1030_g N_A_942_21#_M1015_g 0.0153539f $X=5.49 $Y=2.065 $X2=0
+ $Y2=0
cc_661 N_A_648_21#_c_824_n N_A_942_21#_M1015_g 0.00219889f $X=4.52 $Y=1.91 $X2=0
+ $Y2=0
cc_662 N_A_648_21#_c_804_n N_A_942_21#_M1015_g 0.00171343f $X=4.605 $Y=1.785
+ $X2=0 $Y2=0
cc_663 N_A_648_21#_M1030_g N_A_942_21#_c_1188_n 2.86505e-19 $X=5.49 $Y=2.065
+ $X2=0 $Y2=0
cc_664 N_A_648_21#_c_804_n N_A_942_21#_c_1188_n 0.0309285f $X=4.605 $Y=1.785
+ $X2=0 $Y2=0
cc_665 N_A_648_21#_c_805_n N_A_942_21#_c_1188_n 0.0205705f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_666 N_A_648_21#_c_807_n N_A_942_21#_c_1188_n 0.00382982f $X=5.665 $Y=1.15
+ $X2=0 $Y2=0
cc_667 N_A_648_21#_c_805_n N_A_942_21#_c_1189_n 0.00594187f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_668 N_A_648_21#_c_806_n N_A_942_21#_c_1189_n 7.54142e-19 $X=5.665 $Y=0.98
+ $X2=0 $Y2=0
cc_669 N_A_648_21#_c_807_n N_A_942_21#_c_1189_n 0.0166765f $X=5.665 $Y=1.15
+ $X2=0 $Y2=0
cc_670 N_A_648_21#_c_806_n N_A_942_21#_c_1199_n 9.59092e-19 $X=5.665 $Y=0.98
+ $X2=0 $Y2=0
cc_671 N_A_648_21#_c_807_n N_A_942_21#_c_1199_n 0.00358318f $X=5.665 $Y=1.15
+ $X2=0 $Y2=0
cc_672 N_A_648_21#_M1030_g N_A_942_21#_c_1200_n 0.0143059f $X=5.49 $Y=2.065
+ $X2=0 $Y2=0
cc_673 N_A_648_21#_c_805_n N_A_942_21#_c_1200_n 0.00760725f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_674 N_A_648_21#_c_806_n N_A_942_21#_c_1200_n 0.0207118f $X=5.665 $Y=0.98
+ $X2=0 $Y2=0
cc_675 N_A_648_21#_c_807_n N_A_942_21#_c_1200_n 0.00632961f $X=5.665 $Y=1.15
+ $X2=0 $Y2=0
cc_676 N_A_648_21#_M1030_g N_A_1255_47#_c_1533_n 7.04843e-19 $X=5.49 $Y=2.065
+ $X2=0 $Y2=0
cc_677 N_A_648_21#_M1021_g N_VPWR_c_1711_n 0.00326498f $X=3.315 $Y=2.275 $X2=0
+ $Y2=0
cc_678 N_A_648_21#_c_811_n N_VPWR_c_1711_n 0.0124698f $X=4.09 $Y=1.91 $X2=0
+ $Y2=0
cc_679 N_A_648_21#_c_858_p N_VPWR_c_1711_n 0.00820313f $X=4.175 $Y=2.21 $X2=0
+ $Y2=0
cc_680 N_A_648_21#_c_813_n N_VPWR_c_1711_n 0.0125544f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_681 N_A_648_21#_c_814_n N_VPWR_c_1711_n 7.62241e-19 $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_682 N_A_648_21#_M1030_g N_VPWR_c_1712_n 0.0163458f $X=5.49 $Y=2.065 $X2=0
+ $Y2=0
cc_683 N_A_648_21#_c_824_n N_VPWR_c_1712_n 0.0048929f $X=4.52 $Y=1.91 $X2=0
+ $Y2=0
cc_684 N_A_648_21#_c_811_n N_VPWR_c_1714_n 0.00474052f $X=4.09 $Y=1.91 $X2=0
+ $Y2=0
cc_685 N_A_648_21#_c_858_p N_VPWR_c_1714_n 0.00725778f $X=4.175 $Y=2.21 $X2=0
+ $Y2=0
cc_686 N_A_648_21#_c_824_n N_VPWR_c_1714_n 0.00598455f $X=4.52 $Y=1.91 $X2=0
+ $Y2=0
cc_687 N_A_648_21#_M1021_g N_VPWR_c_1720_n 0.00535335f $X=3.315 $Y=2.275 $X2=0
+ $Y2=0
cc_688 N_A_648_21#_c_813_n N_VPWR_c_1720_n 0.00111392f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_689 N_A_648_21#_M1030_g N_VPWR_c_1721_n 0.00585385f $X=5.49 $Y=2.065 $X2=0
+ $Y2=0
cc_690 N_A_648_21#_M1005_d N_VPWR_c_1708_n 0.0031612f $X=3.92 $Y=2.065 $X2=0
+ $Y2=0
cc_691 N_A_648_21#_M1021_g N_VPWR_c_1708_n 0.00664368f $X=3.315 $Y=2.275 $X2=0
+ $Y2=0
cc_692 N_A_648_21#_M1030_g N_VPWR_c_1708_n 0.00762825f $X=5.49 $Y=2.065 $X2=0
+ $Y2=0
cc_693 N_A_648_21#_c_811_n N_VPWR_c_1708_n 0.00386836f $X=4.09 $Y=1.91 $X2=0
+ $Y2=0
cc_694 N_A_648_21#_c_858_p N_VPWR_c_1708_n 0.0029026f $X=4.175 $Y=2.21 $X2=0
+ $Y2=0
cc_695 N_A_648_21#_c_824_n N_VPWR_c_1708_n 0.00505387f $X=4.52 $Y=1.91 $X2=0
+ $Y2=0
cc_696 N_A_648_21#_c_813_n N_VPWR_c_1708_n 0.00128163f $X=3.425 $Y=1.74 $X2=0
+ $Y2=0
cc_697 N_A_648_21#_c_824_n A_892_329# 0.00339576f $X=4.52 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_698 N_A_648_21#_c_804_n A_892_329# 0.00178287f $X=4.605 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_699 N_A_648_21#_M1002_g N_VGND_c_2015_n 0.00372247f $X=3.315 $Y=0.445 $X2=0
+ $Y2=0
cc_700 N_A_648_21#_c_802_n N_VGND_c_2016_n 0.0111314f $X=5.725 $Y=0.985 $X2=0
+ $Y2=0
cc_701 N_A_648_21#_c_805_n N_VGND_c_2016_n 0.00387395f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_702 N_A_648_21#_c_806_n N_VGND_c_2016_n 0.00379129f $X=5.665 $Y=0.98 $X2=0
+ $Y2=0
cc_703 N_A_648_21#_c_807_n N_VGND_c_2016_n 8.52393e-19 $X=5.665 $Y=1.15 $X2=0
+ $Y2=0
cc_704 N_A_648_21#_M1002_g N_VGND_c_2020_n 0.00359757f $X=3.315 $Y=0.445 $X2=0
+ $Y2=0
cc_705 N_A_648_21#_c_802_n N_VGND_c_2024_n 0.0046653f $X=5.725 $Y=0.985 $X2=0
+ $Y2=0
cc_706 N_A_648_21#_M1023_d N_VGND_c_2031_n 0.00178362f $X=4.44 $Y=0.235 $X2=0
+ $Y2=0
cc_707 N_A_648_21#_M1002_g N_VGND_c_2031_n 0.00576589f $X=3.315 $Y=0.445 $X2=0
+ $Y2=0
cc_708 N_A_648_21#_c_802_n N_VGND_c_2031_n 0.00460207f $X=5.725 $Y=0.985 $X2=0
+ $Y2=0
cc_709 N_A_648_21#_M1023_d N_A_788_47#_c_2201_n 0.0030477f $X=4.44 $Y=0.235
+ $X2=0 $Y2=0
cc_710 N_A_648_21#_c_803_n N_A_788_47#_c_2201_n 0.0147704f $X=4.605 $Y=1.065
+ $X2=0 $Y2=0
cc_711 N_A_648_21#_c_805_n N_A_788_47#_c_2201_n 0.00259503f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_712 N_A_648_21#_c_802_n N_A_788_47#_c_2204_n 0.00441801f $X=5.725 $Y=0.985
+ $X2=0 $Y2=0
cc_713 N_A_648_21#_c_805_n N_A_788_47#_c_2204_n 0.0106429f $X=5.5 $Y=0.98 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_947_n N_A_474_413#_M1023_g 0.00619508f $X=3.845 $Y=1.145 $X2=0
+ $Y2=0
cc_715 N_SET_B_M1029_g N_A_474_413#_M1023_g 0.0234092f $X=3.865 $Y=0.445 $X2=0
+ $Y2=0
cc_716 SET_B N_A_474_413#_M1023_g 0.0018678f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_717 N_SET_B_c_953_n N_A_474_413#_M1023_g 0.00496613f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_954_n N_A_474_413#_M1023_g 0.00135305f $X=4.06 $Y=0.85 $X2=0
+ $Y2=0
cc_719 N_SET_B_M1005_g N_A_474_413#_M1022_g 0.0228864f $X=3.845 $Y=2.275 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_947_n N_A_474_413#_c_1079_n 0.00214594f $X=3.845 $Y=1.145 $X2=0
+ $Y2=0
cc_721 N_SET_B_M1005_g N_A_474_413#_c_1079_n 5.82142e-19 $X=3.845 $Y=2.275 $X2=0
+ $Y2=0
cc_722 N_SET_B_M1029_g N_A_474_413#_c_1079_n 0.0018137f $X=3.865 $Y=0.445 $X2=0
+ $Y2=0
cc_723 SET_B N_A_474_413#_c_1079_n 0.0221461f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_724 N_SET_B_c_954_n N_A_474_413#_c_1079_n 0.00112047f $X=4.06 $Y=0.85 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_947_n N_A_474_413#_c_1080_n 0.00299221f $X=3.845 $Y=1.145 $X2=0
+ $Y2=0
cc_726 N_SET_B_M1005_g N_A_474_413#_c_1080_n 0.0131452f $X=3.845 $Y=2.275 $X2=0
+ $Y2=0
cc_727 SET_B N_A_474_413#_c_1080_n 0.024648f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_728 N_SET_B_c_953_n N_A_474_413#_c_1080_n 0.00284271f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_954_n N_A_474_413#_c_1080_n 6.67689e-19 $X=4.06 $Y=0.85 $X2=0
+ $Y2=0
cc_730 N_SET_B_M1005_g N_A_474_413#_c_1081_n 4.98733e-19 $X=3.845 $Y=2.275 $X2=0
+ $Y2=0
cc_731 N_SET_B_M1005_g N_A_474_413#_c_1082_n 0.021088f $X=3.845 $Y=2.275 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_953_n N_A_942_21#_M1019_g 0.00317213f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_953_n N_A_942_21#_c_1188_n 5.29205e-19 $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_734 N_SET_B_M1010_g N_A_942_21#_c_1198_n 0.00583258f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_953_n N_A_942_21#_c_1198_n 0.0486538f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_SET_B_c_955_n N_A_942_21#_c_1198_n 0.0135087f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_737 N_SET_B_M1025_g N_A_1429_21#_M1009_g 0.0180201f $X=7.65 $Y=0.445 $X2=0
+ $Y2=0
cc_738 N_SET_B_M1010_g N_A_1429_21#_M1009_g 0.0136409f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_739 N_SET_B_c_953_n N_A_1429_21#_M1009_g 0.00627116f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_740 N_SET_B_c_955_n N_A_1429_21#_M1009_g 0.00136404f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_741 N_SET_B_c_956_n N_A_1429_21#_M1009_g 0.00227945f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_742 N_SET_B_c_957_n N_A_1429_21#_M1009_g 0.020875f $X=7.64 $Y=0.98 $X2=0
+ $Y2=0
cc_743 N_SET_B_M1010_g N_A_1429_21#_M1001_g 0.0109753f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_744 N_SET_B_M1010_g N_A_1429_21#_c_1361_n 0.00710111f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_745 N_SET_B_M1010_g N_A_1429_21#_c_1362_n 0.019738f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_746 N_SET_B_M1010_g N_A_1429_21#_c_1363_n 0.0136222f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_956_n N_A_1429_21#_c_1352_n 0.00828511f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_748 N_SET_B_M1025_g N_A_1429_21#_c_1382_n 6.74813e-19 $X=7.65 $Y=0.445 $X2=0
+ $Y2=0
cc_749 N_SET_B_c_955_n N_A_1429_21#_c_1382_n 2.37563e-19 $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_750 N_SET_B_c_956_n N_A_1429_21#_c_1382_n 0.00144717f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_751 N_SET_B_M1025_g N_A_1255_47#_M1028_g 0.0175593f $X=7.65 $Y=0.445 $X2=0
+ $Y2=0
cc_752 N_SET_B_c_956_n N_A_1255_47#_M1028_g 0.00170408f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_753 N_SET_B_c_957_n N_A_1255_47#_M1028_g 0.009306f $X=7.64 $Y=0.98 $X2=0
+ $Y2=0
cc_754 N_SET_B_M1010_g N_A_1255_47#_M1004_g 0.0325064f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_755 N_SET_B_c_953_n N_A_1255_47#_c_1536_n 0.00883541f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_756 N_SET_B_c_953_n N_A_1255_47#_c_1522_n 0.017797f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_757 N_SET_B_c_955_n N_A_1255_47#_c_1522_n 0.0022902f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_758 N_SET_B_c_956_n N_A_1255_47#_c_1522_n 0.0118231f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_759 N_SET_B_M1010_g N_A_1255_47#_c_1523_n 0.0117331f $X=7.76 $Y=2.275 $X2=0
+ $Y2=0
cc_760 N_SET_B_c_953_n N_A_1255_47#_c_1523_n 0.00876649f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_SET_B_c_955_n N_A_1255_47#_c_1523_n 0.00124273f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_762 N_SET_B_c_956_n N_A_1255_47#_c_1523_n 0.0248283f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_763 N_SET_B_c_957_n N_A_1255_47#_c_1523_n 0.00490678f $X=7.64 $Y=0.98 $X2=0
+ $Y2=0
cc_764 N_SET_B_c_957_n N_A_1255_47#_c_1525_n 0.00111089f $X=7.64 $Y=0.98 $X2=0
+ $Y2=0
cc_765 N_SET_B_c_957_n N_A_1255_47#_c_1526_n 0.0212822f $X=7.64 $Y=0.98 $X2=0
+ $Y2=0
cc_766 N_SET_B_M1005_g N_VPWR_c_1711_n 0.0094739f $X=3.845 $Y=2.275 $X2=0 $Y2=0
cc_767 N_SET_B_M1005_g N_VPWR_c_1714_n 0.00373914f $X=3.845 $Y=2.275 $X2=0 $Y2=0
cc_768 N_SET_B_M1010_g N_VPWR_c_1717_n 0.00368415f $X=7.76 $Y=2.275 $X2=0 $Y2=0
cc_769 N_SET_B_M1005_g N_VPWR_c_1708_n 0.00439789f $X=3.845 $Y=2.275 $X2=0 $Y2=0
cc_770 N_SET_B_M1010_g N_VPWR_c_1708_n 0.00444663f $X=7.76 $Y=2.275 $X2=0 $Y2=0
cc_771 N_SET_B_M1010_g N_VPWR_c_1729_n 0.00857728f $X=7.76 $Y=2.275 $X2=0 $Y2=0
cc_772 N_SET_B_c_953_n N_VGND_M1003_s 0.00213341f $X=7.45 $Y=0.85 $X2=0 $Y2=0
cc_773 N_SET_B_c_947_n N_VGND_c_2015_n 7.32772e-19 $X=3.845 $Y=1.145 $X2=0 $Y2=0
cc_774 N_SET_B_M1029_g N_VGND_c_2015_n 0.00287306f $X=3.865 $Y=0.445 $X2=0 $Y2=0
cc_775 SET_B N_VGND_c_2015_n 0.00971383f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_776 N_SET_B_c_953_n N_VGND_c_2016_n 0.00404506f $X=7.45 $Y=0.85 $X2=0 $Y2=0
cc_777 N_SET_B_M1025_g N_VGND_c_2017_n 0.00282278f $X=7.65 $Y=0.445 $X2=0 $Y2=0
cc_778 N_SET_B_c_953_n N_VGND_c_2017_n 0.00604269f $X=7.45 $Y=0.85 $X2=0 $Y2=0
cc_779 N_SET_B_c_955_n N_VGND_c_2017_n 7.41662e-19 $X=7.595 $Y=0.85 $X2=0 $Y2=0
cc_780 N_SET_B_c_956_n N_VGND_c_2017_n 0.00350326f $X=7.595 $Y=0.85 $X2=0 $Y2=0
cc_781 N_SET_B_M1029_g N_VGND_c_2022_n 0.00423333f $X=3.865 $Y=0.445 $X2=0 $Y2=0
cc_782 SET_B N_VGND_c_2022_n 0.00223437f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_783 N_SET_B_M1025_g N_VGND_c_2028_n 0.00439071f $X=7.65 $Y=0.445 $X2=0 $Y2=0
cc_784 N_SET_B_c_956_n N_VGND_c_2028_n 0.00352663f $X=7.595 $Y=0.85 $X2=0 $Y2=0
cc_785 N_SET_B_M1029_g N_VGND_c_2031_n 0.00593301f $X=3.865 $Y=0.445 $X2=0 $Y2=0
cc_786 N_SET_B_M1025_g N_VGND_c_2031_n 0.00595177f $X=7.65 $Y=0.445 $X2=0 $Y2=0
cc_787 SET_B N_VGND_c_2031_n 0.00248323f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_788 N_SET_B_c_953_n N_VGND_c_2031_n 0.165461f $X=7.45 $Y=0.85 $X2=0 $Y2=0
cc_789 N_SET_B_c_954_n N_VGND_c_2031_n 0.014763f $X=4.06 $Y=0.85 $X2=0 $Y2=0
cc_790 N_SET_B_c_955_n N_VGND_c_2031_n 0.0141642f $X=7.595 $Y=0.85 $X2=0 $Y2=0
cc_791 N_SET_B_c_956_n N_VGND_c_2031_n 0.00284893f $X=7.595 $Y=0.85 $X2=0 $Y2=0
cc_792 N_SET_B_c_953_n N_A_788_47#_M1029_d 0.00177886f $X=7.45 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_793 N_SET_B_c_954_n N_A_788_47#_M1029_d 6.34838e-19 $X=4.06 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_794 N_SET_B_c_953_n N_A_788_47#_M1019_d 0.00215149f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_795 N_SET_B_c_953_n N_A_788_47#_c_2201_n 0.00611167f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_796 N_SET_B_c_953_n N_A_788_47#_c_2204_n 0.00234876f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_797 N_SET_B_M1029_g N_A_788_47#_c_2211_n 0.0039841f $X=3.865 $Y=0.445 $X2=0
+ $Y2=0
cc_798 SET_B N_A_788_47#_c_2211_n 0.00361223f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_799 N_SET_B_c_953_n N_A_788_47#_c_2211_n 0.00386944f $X=7.45 $Y=0.85 $X2=0
+ $Y2=0
cc_800 N_SET_B_c_954_n N_A_788_47#_c_2211_n 0.00238177f $X=4.06 $Y=0.85 $X2=0
+ $Y2=0
cc_801 N_SET_B_c_953_n A_1160_47# 0.00369541f $X=7.45 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_802 N_SET_B_M1025_g N_A_1545_47#_c_2232_n 0.00349862f $X=7.65 $Y=0.445 $X2=0
+ $Y2=0
cc_803 N_SET_B_c_956_n N_A_1545_47#_c_2232_n 0.00344477f $X=7.595 $Y=0.85 $X2=0
+ $Y2=0
cc_804 N_SET_B_c_957_n N_A_1545_47#_c_2232_n 2.8008e-19 $X=7.64 $Y=0.98 $X2=0
+ $Y2=0
cc_805 N_A_474_413#_M1023_g N_A_942_21#_M1019_g 0.0306362f $X=4.365 $Y=0.555
+ $X2=0 $Y2=0
cc_806 N_A_474_413#_M1022_g N_A_942_21#_M1015_g 0.0493171f $X=4.385 $Y=2.065
+ $X2=0 $Y2=0
cc_807 N_A_474_413#_c_1082_n N_A_942_21#_c_1189_n 0.0167931f $X=4.265 $Y=1.32
+ $X2=0 $Y2=0
cc_808 N_A_474_413#_M1022_g N_VPWR_c_1711_n 0.00136797f $X=4.385 $Y=2.065 $X2=0
+ $Y2=0
cc_809 N_A_474_413#_M1022_g N_VPWR_c_1714_n 0.00432313f $X=4.385 $Y=2.065 $X2=0
+ $Y2=0
cc_810 N_A_474_413#_c_1088_n N_VPWR_c_1720_n 0.0377433f $X=3 $Y=2.335 $X2=0
+ $Y2=0
cc_811 N_A_474_413#_M1016_d N_VPWR_c_1708_n 0.00173085f $X=2.37 $Y=2.065 $X2=0
+ $Y2=0
cc_812 N_A_474_413#_M1022_g N_VPWR_c_1708_n 0.00600471f $X=4.385 $Y=2.065 $X2=0
+ $Y2=0
cc_813 N_A_474_413#_c_1088_n N_VPWR_c_1708_n 0.0132511f $X=3 $Y=2.335 $X2=0
+ $Y2=0
cc_814 N_A_474_413#_c_1088_n N_A_381_47#_c_1898_n 0.0110044f $X=3 $Y=2.335 $X2=0
+ $Y2=0
cc_815 N_A_474_413#_c_1088_n A_558_413# 0.00858887f $X=3 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_816 N_A_474_413#_c_1084_n A_558_413# 0.00579571f $X=3.085 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_817 N_A_474_413#_c_1094_n N_VGND_c_2020_n 0.0544815f $X=3.23 $Y=0.365 $X2=0
+ $Y2=0
cc_818 N_A_474_413#_M1023_g N_VGND_c_2022_n 0.00357877f $X=4.365 $Y=0.555 $X2=0
+ $Y2=0
cc_819 N_A_474_413#_M1032_d N_VGND_c_2031_n 0.00255824f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_820 N_A_474_413#_M1023_g N_VGND_c_2031_n 0.00545888f $X=4.365 $Y=0.555 $X2=0
+ $Y2=0
cc_821 N_A_474_413#_c_1094_n N_VGND_c_2031_n 0.021542f $X=3.23 $Y=0.365 $X2=0
+ $Y2=0
cc_822 N_A_474_413#_c_1094_n A_582_47# 0.00625863f $X=3.23 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_823 N_A_474_413#_M1023_g N_A_788_47#_c_2201_n 0.00927812f $X=4.365 $Y=0.555
+ $X2=0 $Y2=0
cc_824 N_A_474_413#_c_1080_n N_A_788_47#_c_2211_n 0.00119392f $X=4.1 $Y=1.32
+ $X2=0 $Y2=0
cc_825 N_A_474_413#_c_1082_n N_A_788_47#_c_2211_n 5.73033e-19 $X=4.265 $Y=1.32
+ $X2=0 $Y2=0
cc_826 N_A_942_21#_c_1198_n N_A_1429_21#_M1009_g 0.00413345f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_827 N_A_942_21#_c_1198_n N_A_1429_21#_c_1361_n 0.015309f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_828 N_A_942_21#_c_1198_n N_A_1429_21#_c_1362_n 0.00677286f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_829 N_A_942_21#_c_1198_n N_A_1429_21#_c_1363_n 0.010417f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_830 N_A_942_21#_c_1198_n N_A_1429_21#_c_1389_n 0.00964432f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_831 N_A_942_21#_M1007_g N_A_1429_21#_c_1352_n 0.0128951f $X=8.6 $Y=2.065
+ $X2=0 $Y2=0
cc_832 N_A_942_21#_M1036_g N_A_1429_21#_c_1352_n 0.0062981f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_833 N_A_942_21#_c_1186_n N_A_1429_21#_c_1352_n 0.00727045f $X=9.06 $Y=0.84
+ $X2=0 $Y2=0
cc_834 N_A_942_21#_c_1194_n N_A_1429_21#_c_1352_n 0.0130479f $X=9.06 $Y=1.66
+ $X2=0 $Y2=0
cc_835 N_A_942_21#_c_1198_n N_A_1429_21#_c_1352_n 0.0270698f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_836 N_A_942_21#_c_1201_n N_A_1429_21#_c_1352_n 5.62937e-19 $X=8.975 $Y=1.53
+ $X2=0 $Y2=0
cc_837 N_A_942_21#_c_1190_n N_A_1429_21#_c_1352_n 0.00937037f $X=8.66 $Y=1.32
+ $X2=0 $Y2=0
cc_838 N_A_942_21#_c_1191_n N_A_1429_21#_c_1352_n 0.046128f $X=8.87 $Y=1.32
+ $X2=0 $Y2=0
cc_839 N_A_942_21#_M1034_s N_A_1429_21#_c_1365_n 0.00489108f $X=9.255 $Y=1.505
+ $X2=0 $Y2=0
cc_840 N_A_942_21#_M1007_g N_A_1429_21#_c_1365_n 0.00712539f $X=8.6 $Y=2.065
+ $X2=0 $Y2=0
cc_841 N_A_942_21#_c_1194_n N_A_1429_21#_c_1365_n 0.0212381f $X=9.06 $Y=1.66
+ $X2=0 $Y2=0
cc_842 N_A_942_21#_c_1195_n N_A_1429_21#_c_1365_n 0.0310528f $X=9.38 $Y=1.66
+ $X2=0 $Y2=0
cc_843 N_A_942_21#_c_1198_n N_A_1429_21#_c_1365_n 0.00648571f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_844 N_A_942_21#_c_1201_n N_A_1429_21#_c_1365_n 0.00170504f $X=8.975 $Y=1.53
+ $X2=0 $Y2=0
cc_845 N_A_942_21#_c_1190_n N_A_1429_21#_c_1365_n 0.0026574f $X=8.66 $Y=1.32
+ $X2=0 $Y2=0
cc_846 N_A_942_21#_c_1195_n N_A_1429_21#_c_1366_n 0.00819527f $X=9.38 $Y=1.66
+ $X2=0 $Y2=0
cc_847 N_A_942_21#_c_1198_n N_A_1429_21#_c_1406_n 0.00453864f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_848 N_A_942_21#_M1036_g N_A_1429_21#_c_1382_n 0.00422152f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_849 N_A_942_21#_c_1187_n N_A_1429_21#_c_1382_n 0.00455062f $X=9.39 $Y=0.43
+ $X2=0 $Y2=0
cc_850 N_A_942_21#_M1007_g N_A_1429_21#_c_1409_n 0.00499743f $X=8.6 $Y=2.065
+ $X2=0 $Y2=0
cc_851 N_A_942_21#_M1036_g N_A_1255_47#_M1028_g 0.0191895f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_852 N_A_942_21#_M1007_g N_A_1255_47#_M1004_g 0.039703f $X=8.6 $Y=2.065 $X2=0
+ $Y2=0
cc_853 N_A_942_21#_c_1198_n N_A_1255_47#_M1004_g 0.00713863f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_854 N_A_942_21#_c_1198_n N_A_1255_47#_c_1528_n 0.0219541f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_855 N_A_942_21#_c_1198_n N_A_1255_47#_c_1523_n 0.0228947f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_856 N_A_942_21#_M1036_g N_A_1255_47#_c_1525_n 2.36981e-19 $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_857 N_A_942_21#_c_1198_n N_A_1255_47#_c_1525_n 0.00714757f $X=8.83 $Y=1.53
+ $X2=0 $Y2=0
cc_858 N_A_942_21#_c_1190_n N_A_1255_47#_c_1526_n 0.0588925f $X=8.66 $Y=1.32
+ $X2=0 $Y2=0
cc_859 N_A_942_21#_c_1195_n N_RESET_B_M1034_g 0.00322142f $X=9.38 $Y=1.66 $X2=0
+ $Y2=0
cc_860 N_A_942_21#_c_1201_n N_RESET_B_M1034_g 0.00265509f $X=8.975 $Y=1.53 $X2=0
+ $Y2=0
cc_861 N_A_942_21#_c_1190_n N_RESET_B_M1034_g 0.00254673f $X=8.66 $Y=1.32 $X2=0
+ $Y2=0
cc_862 N_A_942_21#_c_1191_n N_RESET_B_M1034_g 0.0031169f $X=8.87 $Y=1.32 $X2=0
+ $Y2=0
cc_863 N_A_942_21#_c_1185_n N_RESET_B_M1017_g 0.00680458f $X=9.24 $Y=0.84 $X2=0
+ $Y2=0
cc_864 N_A_942_21#_c_1187_n N_RESET_B_M1017_g 0.00288605f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_865 N_A_942_21#_c_1191_n N_RESET_B_M1017_g 0.00236652f $X=8.87 $Y=1.32 $X2=0
+ $Y2=0
cc_866 N_A_942_21#_c_1185_n RESET_B 0.0133113f $X=9.24 $Y=0.84 $X2=0 $Y2=0
cc_867 N_A_942_21#_c_1195_n RESET_B 0.0108125f $X=9.38 $Y=1.66 $X2=0 $Y2=0
cc_868 N_A_942_21#_c_1190_n RESET_B 6.14512e-19 $X=8.66 $Y=1.32 $X2=0 $Y2=0
cc_869 N_A_942_21#_c_1191_n RESET_B 0.0142997f $X=8.87 $Y=1.32 $X2=0 $Y2=0
cc_870 N_A_942_21#_M1036_g N_RESET_B_c_1622_n 0.00156948f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_871 N_A_942_21#_c_1185_n N_RESET_B_c_1622_n 0.00294469f $X=9.24 $Y=0.84 $X2=0
+ $Y2=0
cc_872 N_A_942_21#_c_1195_n N_RESET_B_c_1622_n 0.0032113f $X=9.38 $Y=1.66 $X2=0
+ $Y2=0
cc_873 N_A_942_21#_c_1190_n N_RESET_B_c_1622_n 0.0062814f $X=8.66 $Y=1.32 $X2=0
+ $Y2=0
cc_874 N_A_942_21#_c_1191_n N_RESET_B_c_1622_n 0.00312615f $X=8.87 $Y=1.32 $X2=0
+ $Y2=0
cc_875 N_A_942_21#_c_1188_n N_VPWR_M1015_d 0.00297048f $X=5.025 $Y=1.32 $X2=0
+ $Y2=0
cc_876 N_A_942_21#_c_1200_n N_VPWR_M1015_d 0.00221014f $X=5.755 $Y=1.53 $X2=0
+ $Y2=0
cc_877 N_A_942_21#_c_1194_n N_VPWR_M1007_d 0.00311394f $X=9.06 $Y=1.66 $X2=0
+ $Y2=0
cc_878 N_A_942_21#_M1015_g N_VPWR_c_1712_n 0.00353361f $X=4.805 $Y=2.065 $X2=0
+ $Y2=0
cc_879 N_A_942_21#_c_1188_n N_VPWR_c_1712_n 0.011531f $X=5.025 $Y=1.32 $X2=0
+ $Y2=0
cc_880 N_A_942_21#_c_1189_n N_VPWR_c_1712_n 0.00111411f $X=5.025 $Y=1.32 $X2=0
+ $Y2=0
cc_881 N_A_942_21#_c_1200_n N_VPWR_c_1712_n 7.83548e-19 $X=5.755 $Y=1.53 $X2=0
+ $Y2=0
cc_882 N_A_942_21#_M1015_g N_VPWR_c_1714_n 0.00583607f $X=4.805 $Y=2.065 $X2=0
+ $Y2=0
cc_883 N_A_942_21#_M1007_g N_VPWR_c_1716_n 0.0111257f $X=8.6 $Y=2.065 $X2=0
+ $Y2=0
cc_884 N_A_942_21#_M1007_g N_VPWR_c_1717_n 0.00339278f $X=8.6 $Y=2.065 $X2=0
+ $Y2=0
cc_885 N_A_942_21#_M1015_g N_VPWR_c_1708_n 0.00670824f $X=4.805 $Y=2.065 $X2=0
+ $Y2=0
cc_886 N_A_942_21#_M1007_g N_VPWR_c_1708_n 0.0038354f $X=8.6 $Y=2.065 $X2=0
+ $Y2=0
cc_887 N_A_942_21#_c_1200_n A_1113_329# 0.00272182f $X=5.755 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_888 N_A_942_21#_M1019_g N_VGND_c_2016_n 0.00318127f $X=4.785 $Y=0.555 $X2=0
+ $Y2=0
cc_889 N_A_942_21#_c_1185_n N_VGND_c_2018_n 0.00363139f $X=9.24 $Y=0.84 $X2=0
+ $Y2=0
cc_890 N_A_942_21#_c_1187_n N_VGND_c_2018_n 0.00656552f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_891 N_A_942_21#_M1019_g N_VGND_c_2022_n 0.00357877f $X=4.785 $Y=0.555 $X2=0
+ $Y2=0
cc_892 N_A_942_21#_M1036_g N_VGND_c_2028_n 0.00357877f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_893 N_A_942_21#_c_1185_n N_VGND_c_2028_n 0.00257748f $X=9.24 $Y=0.84 $X2=0
+ $Y2=0
cc_894 N_A_942_21#_c_1186_n N_VGND_c_2028_n 0.00167617f $X=9.06 $Y=0.84 $X2=0
+ $Y2=0
cc_895 N_A_942_21#_c_1187_n N_VGND_c_2028_n 0.0152007f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_896 N_A_942_21#_M1017_s N_VGND_c_2031_n 0.00383158f $X=9.265 $Y=0.235 $X2=0
+ $Y2=0
cc_897 N_A_942_21#_M1019_g N_VGND_c_2031_n 0.00661646f $X=4.785 $Y=0.555 $X2=0
+ $Y2=0
cc_898 N_A_942_21#_M1036_g N_VGND_c_2031_n 0.00657041f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_899 N_A_942_21#_c_1185_n N_VGND_c_2031_n 0.00463666f $X=9.24 $Y=0.84 $X2=0
+ $Y2=0
cc_900 N_A_942_21#_c_1186_n N_VGND_c_2031_n 0.00329575f $X=9.06 $Y=0.84 $X2=0
+ $Y2=0
cc_901 N_A_942_21#_c_1187_n N_VGND_c_2031_n 0.00892354f $X=9.39 $Y=0.43 $X2=0
+ $Y2=0
cc_902 N_A_942_21#_M1019_g N_A_788_47#_c_2201_n 0.0105472f $X=4.785 $Y=0.555
+ $X2=0 $Y2=0
cc_903 N_A_942_21#_c_1186_n N_A_1545_47#_M1036_d 0.00393453f $X=9.06 $Y=0.84
+ $X2=0 $Y2=0
cc_904 N_A_942_21#_M1036_g N_A_1545_47#_c_2236_n 0.0112006f $X=8.66 $Y=0.555
+ $X2=0 $Y2=0
cc_905 N_A_942_21#_c_1186_n N_A_1545_47#_c_2237_n 0.0133877f $X=9.06 $Y=0.84
+ $X2=0 $Y2=0
cc_906 N_A_942_21#_c_1187_n N_A_1545_47#_c_2237_n 0.0167873f $X=9.39 $Y=0.43
+ $X2=0 $Y2=0
cc_907 N_A_942_21#_c_1190_n N_A_1545_47#_c_2237_n 5.38954e-19 $X=8.66 $Y=1.32
+ $X2=0 $Y2=0
cc_908 N_A_1429_21#_c_1352_n N_A_1255_47#_M1028_g 0.0153921f $X=8.525 $Y=1.915
+ $X2=0 $Y2=0
cc_909 N_A_1429_21#_c_1382_n N_A_1255_47#_M1028_g 0.00536261f $X=8.525 $Y=0.687
+ $X2=0 $Y2=0
cc_910 N_A_1429_21#_c_1389_n N_A_1255_47#_M1004_g 0.0118664f $X=8.435 $Y=2 $X2=0
+ $Y2=0
cc_911 N_A_1429_21#_M1001_g N_A_1255_47#_c_1533_n 0.00204127f $X=7.22 $Y=2.275
+ $X2=0 $Y2=0
cc_912 N_A_1429_21#_M1009_g N_A_1255_47#_c_1536_n 0.0017558f $X=7.22 $Y=0.445
+ $X2=0 $Y2=0
cc_913 N_A_1429_21#_M1009_g N_A_1255_47#_c_1522_n 0.0128435f $X=7.22 $Y=0.445
+ $X2=0 $Y2=0
cc_914 N_A_1429_21#_M1009_g N_A_1255_47#_c_1528_n 0.0148682f $X=7.22 $Y=0.445
+ $X2=0 $Y2=0
cc_915 N_A_1429_21#_c_1361_n N_A_1255_47#_c_1528_n 0.0248026f $X=7.34 $Y=1.74
+ $X2=0 $Y2=0
cc_916 N_A_1429_21#_c_1418_p N_A_1255_47#_c_1528_n 0.0135579f $X=7.505 $Y=2
+ $X2=0 $Y2=0
cc_917 N_A_1429_21#_M1009_g N_A_1255_47#_c_1523_n 0.0115171f $X=7.22 $Y=0.445
+ $X2=0 $Y2=0
cc_918 N_A_1429_21#_c_1361_n N_A_1255_47#_c_1523_n 0.0154844f $X=7.34 $Y=1.74
+ $X2=0 $Y2=0
cc_919 N_A_1429_21#_c_1362_n N_A_1255_47#_c_1523_n 0.00126891f $X=7.34 $Y=1.74
+ $X2=0 $Y2=0
cc_920 N_A_1429_21#_c_1363_n N_A_1255_47#_c_1523_n 0.00635717f $X=7.945 $Y=2
+ $X2=0 $Y2=0
cc_921 N_A_1429_21#_c_1406_n N_A_1255_47#_c_1523_n 0.00162703f $X=8.03 $Y=2
+ $X2=0 $Y2=0
cc_922 N_A_1429_21#_c_1389_n N_A_1255_47#_c_1525_n 0.00158774f $X=8.435 $Y=2
+ $X2=0 $Y2=0
cc_923 N_A_1429_21#_c_1352_n N_A_1255_47#_c_1525_n 0.0241621f $X=8.525 $Y=1.915
+ $X2=0 $Y2=0
cc_924 N_A_1429_21#_c_1406_n N_A_1255_47#_c_1525_n 9.97507e-19 $X=8.03 $Y=2
+ $X2=0 $Y2=0
cc_925 N_A_1429_21#_c_1406_n N_A_1255_47#_c_1526_n 4.0151e-19 $X=8.03 $Y=2 $X2=0
+ $Y2=0
cc_926 N_A_1429_21#_M1039_g N_RESET_B_M1034_g 0.0287825f $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_927 N_A_1429_21#_c_1365_n N_RESET_B_M1034_g 0.0143706f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_928 N_A_1429_21#_c_1366_n N_RESET_B_M1034_g 0.00950142f $X=9.945 $Y=1.915
+ $X2=0 $Y2=0
cc_929 N_A_1429_21#_c_1344_n N_RESET_B_M1017_g 0.0197762f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_930 N_A_1429_21#_c_1346_n N_RESET_B_M1017_g 0.00112281f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_931 N_A_1429_21#_c_1353_n N_RESET_B_M1017_g 4.21417e-19 $X=10.025 $Y=1.16
+ $X2=0 $Y2=0
cc_932 N_A_1429_21#_c_1346_n RESET_B 7.11667e-19 $X=10.15 $Y=1.16 $X2=0 $Y2=0
cc_933 N_A_1429_21#_c_1365_n RESET_B 0.00333663f $X=9.86 $Y=2 $X2=0 $Y2=0
cc_934 N_A_1429_21#_c_1353_n RESET_B 0.0188593f $X=10.025 $Y=1.16 $X2=0 $Y2=0
cc_935 N_A_1429_21#_M1039_g N_RESET_B_c_1622_n 6.96081e-19 $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_936 N_A_1429_21#_c_1346_n N_RESET_B_c_1622_n 0.0199816f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_937 N_A_1429_21#_c_1353_n N_RESET_B_c_1622_n 0.00289174f $X=10.025 $Y=1.16
+ $X2=0 $Y2=0
cc_938 N_A_1429_21#_c_1348_n N_A_2136_47#_M1038_g 0.00455389f $X=10.885 $Y=1.535
+ $X2=0 $Y2=0
cc_939 N_A_1429_21#_c_1360_n N_A_2136_47#_M1038_g 0.0111821f $X=11.015 $Y=1.61
+ $X2=0 $Y2=0
cc_940 N_A_1429_21#_c_1347_n N_A_2136_47#_c_1658_n 0.00389093f $X=10.885
+ $Y=1.025 $X2=0 $Y2=0
cc_941 N_A_1429_21#_c_1349_n N_A_2136_47#_c_1658_n 0.00966775f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_942 N_A_1429_21#_c_1350_n N_A_2136_47#_c_1658_n 0.00992783f $X=11.015
+ $Y=0.805 $X2=0 $Y2=0
cc_943 N_A_1429_21#_c_1348_n N_A_2136_47#_c_1664_n 0.00716207f $X=10.885
+ $Y=1.535 $X2=0 $Y2=0
cc_944 N_A_1429_21#_c_1359_n N_A_2136_47#_c_1664_n 0.0105544f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_945 N_A_1429_21#_c_1360_n N_A_2136_47#_c_1664_n 0.0103307f $X=11.015 $Y=1.61
+ $X2=0 $Y2=0
cc_946 N_A_1429_21#_c_1350_n N_A_2136_47#_c_1659_n 0.00384385f $X=11.015
+ $Y=0.805 $X2=0 $Y2=0
cc_947 N_A_1429_21#_c_1360_n N_A_2136_47#_c_1659_n 0.0033881f $X=11.015 $Y=1.61
+ $X2=0 $Y2=0
cc_948 N_A_1429_21#_c_1347_n N_A_2136_47#_c_1660_n 0.0131369f $X=10.885 $Y=1.025
+ $X2=0 $Y2=0
cc_949 N_A_1429_21#_c_1345_n N_A_2136_47#_c_1661_n 0.0110113f $X=10.81 $Y=1.16
+ $X2=0 $Y2=0
cc_950 N_A_1429_21#_c_1347_n N_A_2136_47#_c_1661_n 0.00117559f $X=10.885
+ $Y=1.025 $X2=0 $Y2=0
cc_951 N_A_1429_21#_c_1348_n N_A_2136_47#_c_1661_n 0.00117559f $X=10.885
+ $Y=1.535 $X2=0 $Y2=0
cc_952 N_A_1429_21#_c_1351_n N_A_2136_47#_c_1661_n 0.00732445f $X=10.885 $Y=1.16
+ $X2=0 $Y2=0
cc_953 N_A_1429_21#_c_1347_n N_A_2136_47#_c_1662_n 0.00248624f $X=10.885
+ $Y=1.025 $X2=0 $Y2=0
cc_954 N_A_1429_21#_c_1349_n N_A_2136_47#_c_1662_n 0.0159717f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_955 N_A_1429_21#_c_1363_n N_VPWR_M1001_d 0.00124767f $X=7.945 $Y=2 $X2=0
+ $Y2=0
cc_956 N_A_1429_21#_c_1418_p N_VPWR_M1001_d 0.00160397f $X=7.505 $Y=2 $X2=0
+ $Y2=0
cc_957 N_A_1429_21#_c_1365_n N_VPWR_M1007_d 0.0044189f $X=9.86 $Y=2 $X2=0 $Y2=0
cc_958 N_A_1429_21#_c_1365_n N_VPWR_M1034_d 0.00750664f $X=9.86 $Y=2 $X2=0 $Y2=0
cc_959 N_A_1429_21#_c_1366_n N_VPWR_M1034_d 0.00490342f $X=9.945 $Y=1.915 $X2=0
+ $Y2=0
cc_960 N_A_1429_21#_c_1359_n N_VPWR_c_1713_n 0.00451861f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_961 N_A_1429_21#_c_1365_n N_VPWR_c_1716_n 0.0840165f $X=9.86 $Y=2 $X2=0 $Y2=0
cc_962 N_A_1429_21#_c_1363_n N_VPWR_c_1717_n 0.00359839f $X=7.945 $Y=2 $X2=0
+ $Y2=0
cc_963 N_A_1429_21#_c_1465_p N_VPWR_c_1717_n 0.00713694f $X=8.03 $Y=2.21 $X2=0
+ $Y2=0
cc_964 N_A_1429_21#_c_1389_n N_VPWR_c_1717_n 0.00458994f $X=8.435 $Y=2 $X2=0
+ $Y2=0
cc_965 N_A_1429_21#_c_1365_n N_VPWR_c_1717_n 4.74543e-19 $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_966 N_A_1429_21#_c_1409_n N_VPWR_c_1717_n 0.00279601f $X=8.525 $Y=2 $X2=0
+ $Y2=0
cc_967 N_A_1429_21#_M1001_g N_VPWR_c_1721_n 0.00542601f $X=7.22 $Y=2.275 $X2=0
+ $Y2=0
cc_968 N_A_1429_21#_c_1418_p N_VPWR_c_1721_n 9.91118e-19 $X=7.505 $Y=2 $X2=0
+ $Y2=0
cc_969 N_A_1429_21#_M1039_g N_VPWR_c_1723_n 0.0046653f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_970 N_A_1429_21#_c_1359_n N_VPWR_c_1723_n 0.00471278f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_971 N_A_1429_21#_M1010_d N_VPWR_c_1708_n 0.00327257f $X=7.835 $Y=2.065 $X2=0
+ $Y2=0
cc_972 N_A_1429_21#_M1001_g N_VPWR_c_1708_n 0.00997697f $X=7.22 $Y=2.275 $X2=0
+ $Y2=0
cc_973 N_A_1429_21#_M1039_g N_VPWR_c_1708_n 0.00929621f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_974 N_A_1429_21#_c_1359_n N_VPWR_c_1708_n 0.00941266f $X=11.015 $Y=1.685
+ $X2=0 $Y2=0
cc_975 N_A_1429_21#_c_1363_n N_VPWR_c_1708_n 0.00704318f $X=7.945 $Y=2 $X2=0
+ $Y2=0
cc_976 N_A_1429_21#_c_1418_p N_VPWR_c_1708_n 0.00270501f $X=7.505 $Y=2 $X2=0
+ $Y2=0
cc_977 N_A_1429_21#_c_1465_p N_VPWR_c_1708_n 0.00608739f $X=8.03 $Y=2.21 $X2=0
+ $Y2=0
cc_978 N_A_1429_21#_c_1389_n N_VPWR_c_1708_n 0.00829558f $X=8.435 $Y=2 $X2=0
+ $Y2=0
cc_979 N_A_1429_21#_c_1365_n N_VPWR_c_1708_n 0.00687203f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_980 N_A_1429_21#_c_1409_n N_VPWR_c_1708_n 0.0049407f $X=8.525 $Y=2 $X2=0
+ $Y2=0
cc_981 N_A_1429_21#_M1001_g N_VPWR_c_1729_n 0.00321606f $X=7.22 $Y=2.275 $X2=0
+ $Y2=0
cc_982 N_A_1429_21#_c_1362_n N_VPWR_c_1729_n 7.01948e-19 $X=7.34 $Y=1.74 $X2=0
+ $Y2=0
cc_983 N_A_1429_21#_c_1363_n N_VPWR_c_1729_n 0.0106677f $X=7.945 $Y=2 $X2=0
+ $Y2=0
cc_984 N_A_1429_21#_c_1418_p N_VPWR_c_1729_n 0.0126362f $X=7.505 $Y=2 $X2=0
+ $Y2=0
cc_985 N_A_1429_21#_c_1465_p N_VPWR_c_1729_n 0.00687131f $X=8.03 $Y=2.21 $X2=0
+ $Y2=0
cc_986 N_A_1429_21#_M1039_g N_VPWR_c_1730_n 0.0100464f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_987 N_A_1429_21#_c_1365_n N_VPWR_c_1730_n 0.00915613f $X=9.86 $Y=2 $X2=0
+ $Y2=0
cc_988 N_A_1429_21#_c_1389_n A_1663_329# 0.00202121f $X=8.435 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_989 N_A_1429_21#_c_1352_n A_1663_329# 0.00305059f $X=8.525 $Y=1.915 $X2=-0.19
+ $Y2=-0.24
cc_990 N_A_1429_21#_c_1409_n A_1663_329# 5.84995e-19 $X=8.525 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_991 N_A_1429_21#_c_1345_n N_Q_N_c_1970_n 0.00146072f $X=10.81 $Y=1.16 $X2=0
+ $Y2=0
cc_992 N_A_1429_21#_c_1359_n N_Q_N_c_1970_n 0.00128303f $X=11.015 $Y=1.685 $X2=0
+ $Y2=0
cc_993 N_A_1429_21#_c_1360_n N_Q_N_c_1970_n 5.65205e-19 $X=11.015 $Y=1.61 $X2=0
+ $Y2=0
cc_994 N_A_1429_21#_c_1344_n N_Q_N_c_1967_n 0.00606471f $X=10.075 $Y=0.995 $X2=0
+ $Y2=0
cc_995 N_A_1429_21#_c_1345_n N_Q_N_c_1967_n 0.0224186f $X=10.81 $Y=1.16 $X2=0
+ $Y2=0
cc_996 N_A_1429_21#_c_1346_n N_Q_N_c_1967_n 0.00356142f $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_997 N_A_1429_21#_c_1348_n N_Q_N_c_1967_n 5.65205e-19 $X=10.885 $Y=1.535 $X2=0
+ $Y2=0
cc_998 N_A_1429_21#_c_1350_n N_Q_N_c_1967_n 8.50428e-19 $X=11.015 $Y=0.805 $X2=0
+ $Y2=0
cc_999 N_A_1429_21#_c_1366_n N_Q_N_c_1967_n 0.0163486f $X=9.945 $Y=1.915 $X2=0
+ $Y2=0
cc_1000 N_A_1429_21#_c_1353_n N_Q_N_c_1967_n 0.0236073f $X=10.025 $Y=1.16 $X2=0
+ $Y2=0
cc_1001 N_A_1429_21#_c_1345_n Q_N 0.00141867f $X=10.81 $Y=1.16 $X2=0 $Y2=0
cc_1002 N_A_1429_21#_c_1359_n Q_N 8.69219e-19 $X=11.015 $Y=1.685 $X2=0 $Y2=0
cc_1003 N_A_1429_21#_c_1349_n N_Q_N_c_1969_n 0.00102311f $X=11.015 $Y=0.73 $X2=0
+ $Y2=0
cc_1004 N_A_1429_21#_M1009_g N_VGND_c_2017_n 0.00846638f $X=7.22 $Y=0.445 $X2=0
+ $Y2=0
cc_1005 N_A_1429_21#_c_1344_n N_VGND_c_2018_n 0.0149376f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1006 N_A_1429_21#_c_1346_n N_VGND_c_2018_n 6.74137e-19 $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_1007 N_A_1429_21#_c_1353_n N_VGND_c_2018_n 0.0111532f $X=10.025 $Y=1.16 $X2=0
+ $Y2=0
cc_1008 N_A_1429_21#_c_1349_n N_VGND_c_2019_n 0.00420958f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_1009 N_A_1429_21#_M1009_g N_VGND_c_2024_n 0.0046653f $X=7.22 $Y=0.445 $X2=0
+ $Y2=0
cc_1010 N_A_1429_21#_c_1344_n N_VGND_c_2029_n 0.0046653f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1011 N_A_1429_21#_c_1349_n N_VGND_c_2029_n 0.00541359f $X=11.015 $Y=0.73
+ $X2=0 $Y2=0
cc_1012 N_A_1429_21#_c_1350_n N_VGND_c_2029_n 2.96334e-19 $X=11.015 $Y=0.805
+ $X2=0 $Y2=0
cc_1013 N_A_1429_21#_M1028_d N_VGND_c_2031_n 0.00216833f $X=8.315 $Y=0.235 $X2=0
+ $Y2=0
cc_1014 N_A_1429_21#_M1009_g N_VGND_c_2031_n 0.00460207f $X=7.22 $Y=0.445 $X2=0
+ $Y2=0
cc_1015 N_A_1429_21#_c_1344_n N_VGND_c_2031_n 0.00934473f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1016 N_A_1429_21#_c_1349_n N_VGND_c_2031_n 0.0110992f $X=11.015 $Y=0.73 $X2=0
+ $Y2=0
cc_1017 N_A_1429_21#_M1028_d N_A_1545_47#_c_2236_n 0.00312752f $X=8.315 $Y=0.235
+ $X2=0 $Y2=0
cc_1018 N_A_1429_21#_c_1382_n N_A_1545_47#_c_2236_n 0.0145304f $X=8.525 $Y=0.687
+ $X2=0 $Y2=0
cc_1019 N_A_1255_47#_M1004_g N_VPWR_c_1716_n 0.00209073f $X=8.24 $Y=2.065 $X2=0
+ $Y2=0
cc_1020 N_A_1255_47#_M1004_g N_VPWR_c_1717_n 0.00425094f $X=8.24 $Y=2.065 $X2=0
+ $Y2=0
cc_1021 N_A_1255_47#_c_1533_n N_VPWR_c_1721_n 0.0377433f $X=6.915 $Y=2.335 $X2=0
+ $Y2=0
cc_1022 N_A_1255_47#_M1031_d N_VPWR_c_1708_n 0.00205544f $X=6.285 $Y=2.065 $X2=0
+ $Y2=0
cc_1023 N_A_1255_47#_M1004_g N_VPWR_c_1708_n 0.00591666f $X=8.24 $Y=2.065 $X2=0
+ $Y2=0
cc_1024 N_A_1255_47#_c_1533_n N_VPWR_c_1708_n 0.0272797f $X=6.915 $Y=2.335 $X2=0
+ $Y2=0
cc_1025 N_A_1255_47#_M1004_g N_VPWR_c_1729_n 0.00144209f $X=8.24 $Y=2.065 $X2=0
+ $Y2=0
cc_1026 N_A_1255_47#_c_1533_n A_1341_413# 0.0111731f $X=6.915 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1027 N_A_1255_47#_c_1528_n A_1341_413# 0.00577347f $X=7 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1028 N_A_1255_47#_c_1536_n N_VGND_c_2017_n 0.0155419f $X=6.915 $Y=0.365 $X2=0
+ $Y2=0
cc_1029 N_A_1255_47#_c_1522_n N_VGND_c_2017_n 0.00412668f $X=7 $Y=1.235 $X2=0
+ $Y2=0
cc_1030 N_A_1255_47#_c_1536_n N_VGND_c_2024_n 0.0433655f $X=6.915 $Y=0.365 $X2=0
+ $Y2=0
cc_1031 N_A_1255_47#_M1028_g N_VGND_c_2028_n 0.00357877f $X=8.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1032 N_A_1255_47#_M1027_d N_VGND_c_2031_n 0.00272713f $X=6.275 $Y=0.235 $X2=0
+ $Y2=0
cc_1033 N_A_1255_47#_M1028_g N_VGND_c_2031_n 0.00569618f $X=8.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1034 N_A_1255_47#_c_1536_n N_VGND_c_2031_n 0.0129183f $X=6.915 $Y=0.365 $X2=0
+ $Y2=0
cc_1035 N_A_1255_47#_c_1536_n A_1364_47# 0.0053026f $X=6.915 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1036 N_A_1255_47#_c_1522_n A_1364_47# 0.00495481f $X=7 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_1037 N_A_1255_47#_M1028_g N_A_1545_47#_c_2236_n 0.0110234f $X=8.24 $Y=0.555
+ $X2=0 $Y2=0
cc_1038 N_A_1255_47#_c_1525_n N_A_1545_47#_c_2236_n 0.00293167f $X=8.18 $Y=1.24
+ $X2=0 $Y2=0
cc_1039 N_A_1255_47#_c_1525_n N_A_1545_47#_c_2232_n 0.00206243f $X=8.18 $Y=1.24
+ $X2=0 $Y2=0
cc_1040 N_A_1255_47#_c_1526_n N_A_1545_47#_c_2232_n 3.6952e-19 $X=8.18 $Y=1.24
+ $X2=0 $Y2=0
cc_1041 N_RESET_B_M1034_g N_VPWR_c_1722_n 0.00655753f $X=9.59 $Y=1.825 $X2=0
+ $Y2=0
cc_1042 N_RESET_B_M1017_g N_VGND_c_2018_n 0.00494061f $X=9.6 $Y=0.445 $X2=0
+ $Y2=0
cc_1043 N_RESET_B_M1017_g N_VGND_c_2028_n 0.00585385f $X=9.6 $Y=0.445 $X2=0
+ $Y2=0
cc_1044 N_RESET_B_M1017_g N_VGND_c_2031_n 0.0119571f $X=9.6 $Y=0.445 $X2=0 $Y2=0
cc_1045 N_A_2136_47#_M1038_g N_VPWR_c_1713_n 0.0147323f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1046 N_A_2136_47#_c_1664_n N_VPWR_c_1713_n 0.0477132f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1047 N_A_2136_47#_c_1659_n N_VPWR_c_1713_n 0.010742f $X=11.405 $Y=1.16 $X2=0
+ $Y2=0
cc_1048 N_A_2136_47#_c_1660_n N_VPWR_c_1713_n 0.00259291f $X=11.405 $Y=1.16
+ $X2=0 $Y2=0
cc_1049 N_A_2136_47#_c_1664_n N_VPWR_c_1723_n 0.0169454f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1050 N_A_2136_47#_M1038_g N_VPWR_c_1724_n 0.0046653f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1051 N_A_2136_47#_M1038_g N_VPWR_c_1708_n 0.00895857f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1052 N_A_2136_47#_c_1664_n N_VPWR_c_1708_n 0.0116159f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1053 N_A_2136_47#_c_1664_n N_Q_N_c_1967_n 0.088721f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1054 N_A_2136_47#_c_1661_n N_Q_N_c_1967_n 0.0259687f $X=10.812 $Y=1.16 $X2=0
+ $Y2=0
cc_1055 N_A_2136_47#_c_1658_n N_Q_N_c_1969_n 0.060049f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1056 N_A_2136_47#_M1038_g N_Q_c_2000_n 0.00595806f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_1057 N_A_2136_47#_c_1664_n N_Q_c_2000_n 0.00487713f $X=10.805 $Y=1.91 $X2=0
+ $Y2=0
cc_1058 N_A_2136_47#_c_1659_n N_Q_c_1998_n 0.0266603f $X=11.405 $Y=1.16 $X2=0
+ $Y2=0
cc_1059 N_A_2136_47#_c_1662_n N_Q_c_1998_n 0.0189779f $X=11.417 $Y=0.995 $X2=0
+ $Y2=0
cc_1060 N_A_2136_47#_c_1658_n N_VGND_c_2019_n 0.0212808f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1061 N_A_2136_47#_c_1659_n N_VGND_c_2019_n 0.0104995f $X=11.405 $Y=1.16 $X2=0
+ $Y2=0
cc_1062 N_A_2136_47#_c_1660_n N_VGND_c_2019_n 0.00255976f $X=11.405 $Y=1.16
+ $X2=0 $Y2=0
cc_1063 N_A_2136_47#_c_1662_n N_VGND_c_2019_n 0.00941229f $X=11.417 $Y=0.995
+ $X2=0 $Y2=0
cc_1064 N_A_2136_47#_c_1658_n N_VGND_c_2029_n 0.0199954f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1065 N_A_2136_47#_c_1662_n N_VGND_c_2030_n 0.0046653f $X=11.417 $Y=0.995
+ $X2=0 $Y2=0
cc_1066 N_A_2136_47#_M1011_s N_VGND_c_2031_n 0.00210122f $X=10.68 $Y=0.235 $X2=0
+ $Y2=0
cc_1067 N_A_2136_47#_c_1658_n N_VGND_c_2031_n 0.0119216f $X=10.805 $Y=0.51 $X2=0
+ $Y2=0
cc_1068 N_A_2136_47#_c_1662_n N_VGND_c_2031_n 0.00895857f $X=11.417 $Y=0.995
+ $X2=0 $Y2=0
cc_1069 N_VPWR_c_1708_n N_A_381_47#_M1020_d 0.00295021f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1070 N_VPWR_c_1710_n N_A_381_47#_c_1896_n 0.0123761f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_1071 N_VPWR_c_1720_n N_A_381_47#_c_1896_n 0.00221328f $X=3.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1072 N_VPWR_c_1708_n N_A_381_47#_c_1896_n 0.00203369f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1073 N_VPWR_c_1710_n N_A_381_47#_c_1897_n 0.0116826f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_1074 N_VPWR_c_1719_n N_A_381_47#_c_1897_n 3.86777e-19 $X=1.435 $Y=2.72 $X2=0
+ $Y2=0
cc_1075 N_VPWR_c_1708_n N_A_381_47#_c_1897_n 7.1462e-19 $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1076 N_VPWR_c_1720_n N_A_381_47#_c_1898_n 0.0115924f $X=3.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1077 N_VPWR_c_1708_n N_A_381_47#_c_1898_n 0.00307944f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_1078 N_VPWR_c_1708_n A_558_413# 0.00355877f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1079 N_VPWR_c_1708_n A_892_329# 0.0026811f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1080 N_VPWR_c_1708_n A_1113_329# 0.00777501f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1081 N_VPWR_c_1708_n A_1341_413# 0.00566996f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1082 N_VPWR_c_1708_n A_1663_329# 0.00245111f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1083 N_VPWR_c_1708_n N_Q_N_M1039_d 0.00387172f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1084 N_VPWR_c_1713_n Q_N 0.00155557f $X=11.28 $Y=1.94 $X2=0 $Y2=0
cc_1085 N_VPWR_c_1723_n Q_N 0.0197934f $X=11.15 $Y=2.72 $X2=0 $Y2=0
cc_1086 N_VPWR_c_1708_n Q_N 0.0108988f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1087 N_VPWR_c_1708_n N_Q_M1038_d 0.00387172f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1088 N_VPWR_c_1724_n Q 0.018001f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1089 N_VPWR_c_1708_n Q 0.00993603f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_1090 N_A_381_47#_c_1893_n N_VGND_M1006_s 0.00120065f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1091 N_A_381_47#_c_1894_n N_VGND_M1006_s 9.93425e-19 $X=1.58 $Y=0.73 $X2=0
+ $Y2=0
cc_1092 N_A_381_47#_c_1893_n N_VGND_c_2014_n 0.0102636f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1093 N_A_381_47#_c_1894_n N_VGND_c_2014_n 0.0115074f $X=1.58 $Y=0.73 $X2=0
+ $Y2=0
cc_1094 N_A_381_47#_c_1893_n N_VGND_c_2020_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1095 N_A_381_47#_c_1905_n N_VGND_c_2020_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1096 N_A_381_47#_c_1894_n N_VGND_c_2027_n 4.97798e-19 $X=1.58 $Y=0.73 $X2=0
+ $Y2=0
cc_1097 N_A_381_47#_M1006_d N_VGND_c_2031_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1098 N_A_381_47#_c_1893_n N_VGND_c_2031_n 0.00238237f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1099 N_A_381_47#_c_1894_n N_VGND_c_2031_n 8.52239e-19 $X=1.58 $Y=0.73 $X2=0
+ $Y2=0
cc_1100 N_A_381_47#_c_1905_n N_VGND_c_2031_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1101 N_Q_N_c_1967_n N_VGND_c_2018_n 0.00498262f $X=10.342 $Y=1.63 $X2=0 $Y2=0
cc_1102 N_Q_N_c_1969_n N_VGND_c_2029_n 0.0196502f $X=10.342 $Y=0.573 $X2=0 $Y2=0
cc_1103 N_Q_N_M1035_d N_VGND_c_2031_n 0.00387172f $X=10.15 $Y=0.235 $X2=0 $Y2=0
cc_1104 N_Q_N_c_1969_n N_VGND_c_2031_n 0.0108686f $X=10.342 $Y=0.573 $X2=0 $Y2=0
cc_1105 Q N_VGND_c_2030_n 0.0179668f $X=11.64 $Y=0.425 $X2=0 $Y2=0
cc_1106 N_Q_M1033_d N_VGND_c_2031_n 0.00387172f $X=11.565 $Y=0.235 $X2=0 $Y2=0
cc_1107 Q N_VGND_c_2031_n 0.00992828f $X=11.64 $Y=0.425 $X2=0 $Y2=0
cc_1108 N_VGND_c_2031_n A_582_47# 0.00230551f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1109 N_VGND_c_2031_n N_A_788_47#_M1029_d 0.00227745f $X=11.73 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1110 N_VGND_c_2031_n N_A_788_47#_M1019_d 0.00204204f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1111 N_VGND_c_2016_n N_A_788_47#_c_2201_n 0.010563f $X=5.515 $Y=0.38 $X2=0
+ $Y2=0
cc_1112 N_VGND_c_2022_n N_A_788_47#_c_2201_n 0.0472843f $X=5.35 $Y=0 $X2=0 $Y2=0
cc_1113 N_VGND_c_2031_n N_A_788_47#_c_2201_n 0.01386f $X=11.73 $Y=0 $X2=0 $Y2=0
cc_1114 N_VGND_c_2016_n N_A_788_47#_c_2204_n 0.0022149f $X=5.515 $Y=0.38 $X2=0
+ $Y2=0
cc_1115 N_VGND_c_2022_n N_A_788_47#_c_2211_n 0.0197166f $X=5.35 $Y=0 $X2=0 $Y2=0
cc_1116 N_VGND_c_2031_n N_A_788_47#_c_2211_n 0.00556798f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1117 N_VGND_c_2031_n A_1160_47# 0.00467499f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1118 N_VGND_c_2031_n A_1364_47# 0.00261578f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1119 N_VGND_c_2031_n N_A_1545_47#_M1025_d 0.00378249f $X=11.73 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1120 N_VGND_c_2031_n N_A_1545_47#_M1036_d 0.00230679f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1121 N_VGND_c_2028_n N_A_1545_47#_c_2236_n 0.0358653f $X=9.7 $Y=0 $X2=0 $Y2=0
cc_1122 N_VGND_c_2031_n N_A_1545_47#_c_2236_n 0.0235203f $X=11.73 $Y=0 $X2=0
+ $Y2=0
cc_1123 N_VGND_c_2028_n N_A_1545_47#_c_2232_n 0.0215241f $X=9.7 $Y=0 $X2=0 $Y2=0
cc_1124 N_VGND_c_2031_n N_A_1545_47#_c_2232_n 0.01237f $X=11.73 $Y=0 $X2=0 $Y2=0
cc_1125 N_VGND_c_2028_n N_A_1545_47#_c_2237_n 0.0110309f $X=9.7 $Y=0 $X2=0 $Y2=0
cc_1126 N_VGND_c_2031_n N_A_1545_47#_c_2237_n 0.0063548f $X=11.73 $Y=0 $X2=0
+ $Y2=0

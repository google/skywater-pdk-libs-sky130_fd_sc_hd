* File: sky130_fd_sc_hd__probec_p_8.spice.SKY130_FD_SC_HD__PROBEC_P_8.pxi
* Created: Thu Aug 27 14:45:03 2020
* 
x_PM_SKY130_FD_SC_HD__PROBEC_P_8%A N_A_M1007_g N_A_M1002_g N_A_M1012_g
+ N_A_M1004_g N_A_c_148_n N_A_M1021_g N_A_M1013_g A A A
+ PM_SKY130_FD_SC_HD__PROBEC_P_8%A
x_PM_SKY130_FD_SC_HD__PROBEC_P_8%A_27_47# N_A_27_47#_M1007_d N_A_27_47#_M1012_d
+ N_A_27_47#_M1002_s N_A_27_47#_M1004_s N_A_27_47#_M1000_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1003_g N_A_27_47#_M1005_g N_A_27_47#_M1009_g N_A_27_47#_M1006_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1008_g N_A_27_47#_M1014_g N_A_27_47#_M1011_g
+ N_A_27_47#_M1016_g N_A_27_47#_M1015_g N_A_27_47#_M1017_g N_A_27_47#_M1019_g
+ N_A_27_47#_M1018_g N_A_27_47#_M1020_g N_A_27_47#_c_264_n N_A_27_47#_c_273_n
+ N_A_27_47#_c_247_n N_A_27_47#_c_248_n N_A_27_47#_c_265_n N_A_27_47#_c_266_n
+ N_A_27_47#_c_287_n N_A_27_47#_c_290_n N_A_27_47#_c_249_n N_A_27_47#_c_250_n
+ N_A_27_47#_c_251_n N_A_27_47#_c_252_n N_A_27_47#_c_268_n N_A_27_47#_c_253_n
+ N_A_27_47#_c_254_n N_A_27_47#_c_255_n PM_SKY130_FD_SC_HD__PROBEC_P_8%A_27_47#
x_PM_SKY130_FD_SC_HD__PROBEC_P_8%VPWR N_VPWR_M1002_d N_VPWR_M1013_d
+ N_VPWR_M1005_d N_VPWR_M1008_d N_VPWR_M1015_d N_VPWR_M1020_d N_VPWR_c_553_n
+ N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n
+ N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n VPWR VPWR
+ N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_R25_noxref_neg N_VPWR_c_571_n
+ N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_549_n N_VPWR_c_550_n
+ N_VPWR_c_551_n N_VPWR_c_552_n PM_SKY130_FD_SC_HD__PROBEC_P_8%VPWR
x_PM_SKY130_FD_SC_HD__PROBEC_P_8%noxref_6 N_noxref_6_M1000_d N_noxref_6_M1009_d
+ N_noxref_6_M1014_d N_noxref_6_M1017_d N_noxref_6_M1001_s N_noxref_6_M1006_s
+ N_noxref_6_M1011_s N_noxref_6_M1019_s N_noxref_6_c_717_n N_noxref_6_c_720_n
+ N_noxref_6_c_684_n N_noxref_6_c_685_n N_noxref_6_c_697_n N_noxref_6_c_698_n
+ N_noxref_6_c_739_n N_noxref_6_c_740_n N_noxref_6_c_686_n N_noxref_6_c_699_n
+ N_noxref_6_c_898_p N_noxref_6_c_859_n N_noxref_6_c_687_n N_noxref_6_c_700_n
+ N_noxref_6_c_688_n N_noxref_6_c_761_n N_noxref_6_c_763_n N_noxref_6_c_689_n
+ N_noxref_6_c_701_n N_noxref_6_c_690_n N_noxref_6_c_702_n N_noxref_6_c_691_n
+ N_noxref_6_c_703_n N_noxref_6_c_779_n N_noxref_6_c_704_n N_noxref_6_c_785_n
+ N_noxref_6_c_692_n N_noxref_6_c_693_n N_noxref_6_c_706_n N_noxref_6_c_710_n
+ N_noxref_6_c_694_n N_noxref_6_c_695_n N_noxref_6_R23_noxref_neg
+ N_noxref_6_c_696_n PM_SKY130_FD_SC_HD__PROBEC_P_8%noxref_6
x_PM_SKY130_FD_SC_HD__PROBEC_P_8%VGND N_VGND_M1007_s N_VGND_M1021_s
+ N_VGND_M1003_s N_VGND_M1010_s N_VGND_M1016_s N_VGND_M1018_s N_VGND_c_935_n
+ N_VGND_c_936_n N_VGND_c_937_n N_VGND_c_938_n N_VGND_c_939_n N_VGND_c_940_n
+ N_VGND_c_941_n N_VGND_c_942_n N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n
+ N_VGND_c_946_n N_VGND_c_947_n VGND VGND N_VGND_c_948_n N_VGND_c_949_n
+ N_VGND_R24_noxref_neg N_VGND_c_951_n VGND N_VGND_c_952_n N_VGND_c_953_n
+ N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n N_VGND_c_957_n N_VGND_c_958_n
+ N_VGND_c_959_n N_VGND_c_960_n PM_SKY130_FD_SC_HD__PROBEC_P_8%VGND
x_PM_SKY130_FD_SC_HD__PROBEC_P_8%X X N_X_c_1086_n N_X_c_1087_n
+ N_X_R23_noxref_pos PM_SKY130_FD_SC_HD__PROBEC_P_8%X
cc_1 VNB N_A_M1007_g 0.0222825f $X=-1.26 $Y=-1.17 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1012_g 0.0165644f $X=-1.26 $Y=-1.17 $X2=0.89 $Y2=0.56
cc_3 VNB N_A_M1004_g 4.12819e-19 $X=-1.26 $Y=-1.17 $X2=0.89 $Y2=1.985
cc_4 VNB N_A_c_148_n 0.0750715f $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=1.025
cc_5 VNB N_A_M1021_g 0.016794f $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=0.56
cc_6 VNB N_A_M1013_g 4.29284e-19 $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=1.985
cc_7 VNB A 0.00614839f $X=-1.26 $Y=-1.17 $X2=1.07 $Y2=1.105
cc_8 VNB N_A_27_47#_M1000_g 0.016824f $X=-1.26 $Y=-1.17 $X2=0.89 $Y2=1.985
cc_9 VNB N_A_27_47#_M1001_g 4.20085e-19 $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=0.56
cc_10 VNB N_A_27_47#_M1003_g 0.0164556f $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=1.985
cc_11 VNB N_A_27_47#_M1005_g 3.77304e-19 $X=-1.26 $Y=-1.17 $X2=1.07 $Y2=1.105
cc_12 VNB N_A_27_47#_M1009_g 0.0165247f $X=-1.26 $Y=-1.17 $X2=0.305 $Y2=1.16
cc_13 VNB N_A_27_47#_M1006_g 3.77304e-19 $X=-1.26 $Y=-1.17 $X2=0.89 $Y2=1.16
cc_14 VNB N_A_27_47#_M1010_g 0.0170779f $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=1.16
cc_15 VNB N_A_27_47#_M1008_g 4.5018e-19 $X=-1.26 $Y=-1.17 $X2=0.695 $Y2=1.175
cc_16 VNB N_A_27_47#_M1014_g 0.0170779f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_M1011_g 4.50211e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_M1016_g 0.0170518f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_M1015_g 4.49527e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_M1017_g 0.0165623f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_M1019_g 4.12504e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_M1018_g 0.0233974f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1020_g 5.16789e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_247_n 0.00250573f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_248_n 0.00172634f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_249_n 8.4101e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_250_n 0.00933312f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_251_n 0.00270733f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_252_n 0.00211055f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_253_n 0.00106925f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_254_n 0.00144525f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_255_n 0.137686f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_546_n 0.0363973f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_547_n 0.00928873f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_35 VNB N_VPWR_R25_noxref_neg 0.166954f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_549_n 0.00750641f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_550_n 0.00738469f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_551_n 0.00770441f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_552_n 0.190605f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_40 VNB N_noxref_6_c_684_n 0.00226675f $X=-1.26 $Y=-1.17 $X2=0.305 $Y2=1.16
cc_41 VNB N_noxref_6_c_685_n 0.00109487f $X=-1.26 $Y=-1.17 $X2=0.47 $Y2=1.16
cc_42 VNB N_noxref_6_c_686_n 0.00255676f $X=-1.26 $Y=-1.17 $X2=0.985 $Y2=1.175
cc_43 VNB N_noxref_6_c_687_n 0.00245814f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_44 VNB N_noxref_6_c_688_n 0.00113458f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_45 VNB N_noxref_6_c_689_n 0.00104218f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_46 VNB N_noxref_6_c_690_n 0.00105525f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_47 VNB N_noxref_6_c_691_n 2.04274e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_48 VNB N_noxref_6_c_692_n 0.0095583f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_49 VNB N_noxref_6_c_693_n 0.00482224f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_50 VNB N_noxref_6_c_694_n 0.218494f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_51 VNB N_noxref_6_c_695_n 0.0025284f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_52 VNB N_noxref_6_c_696_n 2.37651e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_935_n 3.95446e-19 $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=1.295
cc_54 VNB N_VGND_c_936_n 3.01744e-19 $X=-1.26 $Y=-1.17 $X2=0.15 $Y2=1.105
cc_55 VNB N_VGND_c_937_n 3.01744e-19 $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_938_n 3.01744e-19 $X=-1.26 $Y=-1.17 $X2=0.305 $Y2=1.16
cc_57 VNB N_VGND_c_939_n 0.0112357f $X=-1.26 $Y=-1.17 $X2=0.89 $Y2=1.16
cc_58 VNB N_VGND_c_940_n 3.01744e-19 $X=-1.26 $Y=-1.17 $X2=1.31 $Y2=1.16
cc_59 VNB N_VGND_c_941_n 0.0285416f $X=-1.26 $Y=-1.17 $X2=0.695 $Y2=1.175
cc_60 VNB N_VGND_c_942_n 0.0112511f $X=-1.26 $Y=-1.17 $X2=1.155 $Y2=1.175
cc_61 VNB N_VGND_c_943_n 0.00436716f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_944_n 0.0118508f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_945_n 0.00436716f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_946_n 0.0112357f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_947_n 0.00436716f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_948_n 0.0434956f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_949_n 0.0139421f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_68 VNB N_VGND_R24_noxref_neg 0.170589f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_951_n 0.0152765f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_952_n 0.011863f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_953_n 0.0172331f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_954_n 0.00436716f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_955_n 0.00436716f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_956_n 0.00510472f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_957_n 0.0175422f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_958_n 0.0126802f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_959_n 0.0119695f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_960_n 0.219484f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_79 VNB N_X_c_1086_n 0.0380493f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_80 VNB N_X_c_1087_n 0.028536f $X=-1.26 $Y=-1.17 $X2=0 $Y2=0
cc_81 VNB N_X_R23_noxref_pos 0.147985f $X=-1.26 $Y=-1.17 $X2=0.89 $Y2=0.56
cc_82 VNB noxref_9 8.97967e-19 $X=-1.26 $Y=-1.17 $X2=0.47 $Y2=1.015
cc_83 VNB noxref_10 8.97967e-19 $X=-1.26 $Y=-1.17 $X2=0.47 $Y2=1.015
cc_84 VPB N_A_M1002_g 0.025885f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_85 VPB N_A_M1004_g 0.0185877f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_86 VPB N_A_c_148_n 0.0115707f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_87 VPB N_A_M1013_g 0.0189023f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_88 VPB N_A_27_47#_M1001_g 0.0189935f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_89 VPB N_A_27_47#_M1005_g 0.0181316f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_90 VPB N_A_27_47#_M1006_g 0.0181875f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_91 VPB N_A_27_47#_M1008_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_92 VPB N_A_27_47#_M1011_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_27_47#_M1015_g 0.0189506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_47#_M1019_g 0.0183706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_M1020_g 0.0264665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_27_47#_c_264_n 0.0290878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_47#_c_265_n 0.00183845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_27_47#_c_266_n 0.00864366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_47#_c_251_n 0.00792443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_c_268_n 0.00258557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_553_n 0.00410835f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.295
cc_102 VPB N_VPWR_c_554_n 0.00354062f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_103 VPB N_VPWR_c_555_n 3.15634e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_556_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.16
cc_105 VPB N_VPWR_c_557_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_106 VPB N_VPWR_c_558_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_107 VPB N_VPWR_c_559_n 0.0420863f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_108 VPB N_VPWR_c_560_n 0.0178658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_561_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_562_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_563_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_564_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_565_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_566_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_567_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_546_n 0.00709828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_547_n 0.00465337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_R25_noxref_neg 0.00363507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_571_n 0.0124659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_572_n 0.0172331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_573_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_574_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_549_n 0.0100358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_550_n 0.00529549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_551_n 0.00426506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_552_n 0.0282636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_noxref_6_c_697_n 0.0024464f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_128 VPB N_noxref_6_c_698_n 0.0013946f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_129 VPB N_noxref_6_c_699_n 0.00265147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_noxref_6_c_700_n 0.00248955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_noxref_6_c_701_n 0.00111186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_noxref_6_c_702_n 0.00111344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_noxref_6_c_703_n 0.00163765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_noxref_6_c_704_n 3.76364e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_noxref_6_c_693_n 0.00329673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_noxref_6_c_706_n 0.00422453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_noxref_6_c_694_n 0.00318712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_noxref_6_c_695_n 0.00761317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_noxref_6_c_696_n 0.00586934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_X_c_1086_n 0.0088462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_X_c_1087_n 0.00425834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_X_R23_noxref_pos 0.00880667f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_143 N_A_M1021_g N_A_27_47#_M1000_g 0.0260985f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A_M1013_g N_A_27_47#_M1001_g 0.0260985f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1002_g N_A_27_47#_c_264_n 0.0102175f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1004_g N_A_27_47#_c_264_n 0.00137214f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1007_g N_A_27_47#_c_273_n 0.00288541f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A_M1007_g N_A_27_47#_c_247_n 0.0121062f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_M1012_g N_A_27_47#_c_247_n 0.0109514f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_150 N_A_c_148_n N_A_27_47#_c_247_n 0.00319624f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_151 A N_A_27_47#_c_247_n 0.0488982f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A_c_148_n N_A_27_47#_c_248_n 0.00407757f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_153 A N_A_27_47#_c_248_n 0.0138782f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_A_27_47#_c_265_n 0.0100894f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1004_g N_A_27_47#_c_265_n 0.0100894f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_c_148_n N_A_27_47#_c_265_n 0.00196335f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_157 A N_A_27_47#_c_265_n 0.0595979f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A_M1002_g N_A_27_47#_c_266_n 0.0016057f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_c_148_n N_A_27_47#_c_266_n 0.00590258f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_160 A N_A_27_47#_c_266_n 0.0231973f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A_M1002_g N_A_27_47#_c_287_n 0.00137472f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_M1004_g N_A_27_47#_c_287_n 0.0102727f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_M1013_g N_A_27_47#_c_287_n 0.0102952f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1012_g N_A_27_47#_c_290_n 0.00119913f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A_M1021_g N_A_27_47#_c_290_n 0.00163022f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A_M1021_g N_A_27_47#_c_249_n 0.0120698f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_167 A N_A_27_47#_c_249_n 0.00405505f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A_M1021_g N_A_27_47#_c_250_n 0.00423626f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A_c_148_n N_A_27_47#_c_251_n 0.00451329f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_170 A N_A_27_47#_c_251_n 0.00219565f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A_M1004_g N_A_27_47#_c_268_n 0.0012801f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_c_148_n N_A_27_47#_c_268_n 0.00198167f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_173 N_A_M1013_g N_A_27_47#_c_268_n 0.012524f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_c_148_n N_A_27_47#_c_253_n 0.00213249f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_175 A N_A_27_47#_c_253_n 0.013829f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A_c_148_n N_A_27_47#_c_254_n 0.00171222f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_177 A N_A_27_47#_c_254_n 0.0141446f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A_c_148_n N_A_27_47#_c_255_n 0.0260985f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_179 A N_A_27_47#_c_255_n 2.88051e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_180 N_A_M1002_g N_VPWR_c_553_n 0.00314797f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_M1004_g N_VPWR_c_553_n 0.00192522f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1013_g N_VPWR_c_554_n 0.00242503f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1002_g N_VPWR_c_560_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_M1004_g N_VPWR_c_562_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_M1013_g N_VPWR_c_562_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_M1002_g N_VPWR_c_552_n 0.0102459f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_M1004_g N_VPWR_c_552_n 0.00929169f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_M1013_g N_VPWR_c_552_n 0.00901183f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_M1021_g N_noxref_6_c_710_n 0.00128153f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_190 A N_noxref_6_c_710_n 0.00109767f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A_c_148_n N_noxref_6_c_694_n 4.40213e-19 $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_192 N_A_M1021_g N_noxref_6_c_694_n 3.94565e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_M1013_g N_noxref_6_c_694_n 5.16911e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_194 A N_noxref_6_c_694_n 4.60477e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_195 A N_noxref_6_c_695_n 0.0010351f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_196 N_A_M1007_g N_VGND_c_935_n 0.00936627f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A_M1012_g N_VGND_c_935_n 0.00764412f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_M1021_g N_VGND_c_935_n 5.94015e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_M1012_g N_VGND_c_936_n 8.30543e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_M1021_g N_VGND_c_936_n 0.00731257f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_M1012_g N_VGND_c_942_n 0.00350562f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_M1021_g N_VGND_c_942_n 0.00350562f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_M1007_g N_VGND_c_951_n 0.00350562f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_204 N_A_M1007_g N_VGND_c_960_n 0.00511162f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A_M1012_g N_VGND_c_960_n 0.00412071f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_M1021_g N_VGND_c_960_n 0.0066984f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_M1007_g N_X_c_1086_n 7.41006e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_M1002_g N_X_c_1086_n 6.3996e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_M1002_g N_X_c_1087_n 5.19434e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_c_148_n N_X_c_1087_n 0.00125134f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_211 A N_X_c_1087_n 0.00432327f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_212 N_A_M1007_g N_X_R23_noxref_pos 0.00248103f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_213 N_A_M1002_g N_X_R23_noxref_pos 0.00273386f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_M1012_g N_X_R23_noxref_pos 0.00201108f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A_M1004_g N_X_R23_noxref_pos 0.00213402f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_c_148_n N_X_R23_noxref_pos 0.00363346f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_217 A N_X_R23_noxref_pos 0.00321318f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_265_n N_VPWR_M1002_d 0.00150139f $X=0.935 $Y=1.53 $X2=-1.26
+ $Y2=-1.17
cc_219 N_A_27_47#_c_268_n N_VPWR_M1013_d 0.00282822f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_264_n N_VPWR_c_553_n 0.0301045f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_265_n N_VPWR_c_553_n 0.0108584f $X=0.935 $Y=1.53 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_287_n N_VPWR_c_553_n 0.0301045f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_223 N_A_27_47#_M1001_g N_VPWR_c_554_n 0.00269948f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_287_n N_VPWR_c_554_n 0.0361719f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_252_n N_VPWR_c_554_n 2.25712e-19 $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_268_n N_VPWR_c_554_n 0.0103956f $X=1.507 $Y=1.53 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1001_g N_VPWR_c_555_n 0.00115389f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1005_g N_VPWR_c_555_n 0.0104957f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_27_47#_M1006_g N_VPWR_c_555_n 0.0103055f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_27_47#_M1008_g N_VPWR_c_555_n 0.00111773f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1006_g N_VPWR_c_556_n 6.71865e-19 $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1008_g N_VPWR_c_556_n 0.0110857f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A_27_47#_M1011_g N_VPWR_c_556_n 0.0110857f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_27_47#_M1015_g N_VPWR_c_556_n 6.72101e-19 $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_M1011_g N_VPWR_c_557_n 0.0046653f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_27_47#_M1015_g N_VPWR_c_557_n 0.0046653f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_27_47#_M1011_g N_VPWR_c_558_n 6.72101e-19 $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1015_g N_VPWR_c_558_n 0.0110857f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A_27_47#_M1019_g N_VPWR_c_558_n 0.0110857f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_27_47#_M1020_g N_VPWR_c_558_n 6.71865e-19 $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1019_g N_VPWR_c_559_n 0.00104017f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1020_g N_VPWR_c_559_n 0.0154568f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_264_n N_VPWR_c_560_n 0.0210382f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_287_n N_VPWR_c_562_n 0.0206903f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_245 N_A_27_47#_M1001_g N_VPWR_c_564_n 0.00585385f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_M1005_g N_VPWR_c_564_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1006_g N_VPWR_c_566_n 0.0046653f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_27_47#_M1008_g N_VPWR_c_566_n 0.0046653f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_27_47#_M1019_g N_VPWR_R25_noxref_neg 0.00210746f $X=4.25 $Y=1.985
+ $X2=0 $Y2=0
cc_250 N_A_27_47#_M1020_g N_VPWR_R25_noxref_neg 0.00103574f $X=4.67 $Y=1.985
+ $X2=0 $Y2=0
cc_251 N_A_27_47#_M1019_g N_VPWR_c_571_n 0.0046653f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1020_g N_VPWR_c_571_n 0.0046653f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1002_s N_VPWR_c_552_n 0.00200771f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1004_s N_VPWR_c_552_n 0.00386179f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1001_g N_VPWR_c_552_n 0.00907721f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1005_g N_VPWR_c_552_n 0.0066984f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A_27_47#_M1006_g N_VPWR_c_552_n 0.0066984f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_27_47#_M1008_g N_VPWR_c_552_n 0.00796766f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1011_g N_VPWR_c_552_n 0.00796766f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1015_g N_VPWR_c_552_n 0.00796766f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1019_g N_VPWR_c_552_n 0.00796766f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1020_g N_VPWR_c_552_n 0.0066984f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_264_n N_VPWR_c_552_n 0.0124268f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_287_n N_VPWR_c_552_n 0.0121942f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_265 N_A_27_47#_M1000_g N_noxref_6_c_717_n 0.00165817f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1003_g N_noxref_6_c_717_n 0.00165817f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_290_n N_noxref_6_c_717_n 0.00240618f $X=1.1 $Y=0.56 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1001_g N_noxref_6_c_720_n 0.00268077f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1005_g N_noxref_6_c_720_n 0.00239846f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_287_n N_noxref_6_c_720_n 0.00454491f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1003_g N_noxref_6_c_684_n 0.0105025f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1009_g N_noxref_6_c_684_n 0.0108845f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_252_n N_noxref_6_c_684_n 0.0469989f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_255_n N_noxref_6_c_684_n 0.00196874f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1000_g N_noxref_6_c_685_n 0.00113835f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_249_n N_noxref_6_c_685_n 0.00848213f $X=1.42 $Y=0.82 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_252_n N_noxref_6_c_685_n 0.0137916f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_255_n N_noxref_6_c_685_n 0.00203093f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1005_g N_noxref_6_c_697_n 0.0122351f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1006_g N_noxref_6_c_697_n 0.0123598f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_252_n N_noxref_6_c_697_n 0.0402184f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_255_n N_noxref_6_c_697_n 0.00158708f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1001_g N_noxref_6_c_698_n 0.0010746f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_252_n N_noxref_6_c_698_n 0.0120326f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_268_n N_noxref_6_c_698_n 0.00870005f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_255_n N_noxref_6_c_698_n 0.00189899f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1009_g N_noxref_6_c_739_n 0.00165817f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1006_g N_noxref_6_c_740_n 0.00239917f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_M1010_g N_noxref_6_c_686_n 0.0114673f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1014_g N_noxref_6_c_686_n 0.0114673f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_252_n N_noxref_6_c_686_n 0.0426017f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_255_n N_noxref_6_c_686_n 0.00205431f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1008_g N_noxref_6_c_699_n 0.0135372f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1011_g N_noxref_6_c_699_n 0.0135372f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_252_n N_noxref_6_c_699_n 0.0344123f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_255_n N_noxref_6_c_699_n 0.00201555f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1016_g N_noxref_6_c_687_n 0.0114232f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1017_g N_noxref_6_c_687_n 0.00889009f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_252_n N_noxref_6_c_687_n 0.0216261f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_255_n N_noxref_6_c_687_n 0.00222173f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1015_g N_noxref_6_c_700_n 0.0135372f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1019_g N_noxref_6_c_700_n 0.0112272f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_252_n N_noxref_6_c_700_n 0.0174698f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_255_n N_noxref_6_c_700_n 0.00215943f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1016_g N_noxref_6_c_688_n 5.93233e-19 $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1017_g N_noxref_6_c_688_n 0.00320213f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1018_g N_noxref_6_c_688_n 0.00307239f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_255_n N_noxref_6_c_688_n 0.00541619f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1017_g N_noxref_6_c_761_n 8.85384e-19 $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1018_g N_noxref_6_c_761_n 8.91448e-19 $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_M1019_g N_noxref_6_c_763_n 9.47157e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_252_n N_noxref_6_c_689_n 0.0128734f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_255_n N_noxref_6_c_689_n 0.00212631f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_252_n N_noxref_6_c_701_n 0.0106074f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_255_n N_noxref_6_c_701_n 0.0021011f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_252_n N_noxref_6_c_690_n 0.0123225f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_255_n N_noxref_6_c_690_n 0.00213429f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_252_n N_noxref_6_c_702_n 0.0100399f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_255_n N_noxref_6_c_702_n 0.00211055f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_M1017_g N_noxref_6_c_691_n 0.00272967f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1018_g N_noxref_6_c_691_n 0.00114299f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_M1015_g N_noxref_6_c_703_n 8.70811e-19 $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1019_g N_noxref_6_c_703_n 0.00782978f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1020_g N_noxref_6_c_703_n 0.00568779f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_252_n N_noxref_6_c_703_n 0.00733409f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_255_n N_noxref_6_c_703_n 0.0119217f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_252_n N_noxref_6_c_779_n 0.042053f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_255_n N_noxref_6_c_779_n 0.0182561f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_M1006_g N_noxref_6_c_704_n 0.0020807f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_M1008_g N_noxref_6_c_704_n 3.01733e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_252_n N_noxref_6_c_704_n 0.00469235f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_255_n N_noxref_6_c_704_n 0.00328141f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_M1019_g N_noxref_6_c_785_n 5.67835e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_252_n N_noxref_6_c_785_n 0.00129742f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_255_n N_noxref_6_c_785_n 0.00248761f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_M1020_g N_noxref_6_c_693_n 0.00662372f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_255_n N_noxref_6_c_693_n 0.0168734f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_M1001_g N_noxref_6_c_706_n 3.14325e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_M1005_g N_noxref_6_c_706_n 0.00287285f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1006_g N_noxref_6_c_706_n 7.62036e-19 $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_250_n N_noxref_6_c_706_n 4.21355e-19 $X=1.507 $Y=1.075 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_251_n N_noxref_6_c_706_n 0.0022543f $X=1.507 $Y=1.445 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_252_n N_noxref_6_c_706_n 0.0182391f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_255_n N_noxref_6_c_706_n 0.0106133f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_M1000_g N_noxref_6_c_710_n 0.0021128f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_M1001_g N_noxref_6_c_710_n 0.00211985f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_M1003_g N_noxref_6_c_710_n 4.57766e-19 $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_M1005_g N_noxref_6_c_710_n 0.00200891f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_M1009_g N_noxref_6_c_710_n 0.0015196f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_M1006_g N_noxref_6_c_710_n 0.00640478f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_M1010_g N_noxref_6_c_710_n 5.23911e-19 $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_M1008_g N_noxref_6_c_710_n 3.97315e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_287_n N_noxref_6_c_710_n 0.0024401f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_249_n N_noxref_6_c_710_n 0.00363994f $X=1.42 $Y=0.82 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_250_n N_noxref_6_c_710_n 0.00338326f $X=1.507 $Y=1.075 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_251_n N_noxref_6_c_710_n 0.00406049f $X=1.507 $Y=1.445 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_252_n N_noxref_6_c_710_n 0.00230097f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_268_n N_noxref_6_c_710_n 0.00301616f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_254_n N_noxref_6_c_710_n 0.00187497f $X=1.507 $Y=1.16 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_255_n N_noxref_6_c_710_n 4.93702e-19 $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_M1012_d N_noxref_6_c_694_n 4.56111e-19 $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_M1004_s N_noxref_6_c_694_n 3.42391e-19 $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_M1000_g N_noxref_6_c_694_n 4.58397e-19 $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_M1003_g N_noxref_6_c_694_n 3.82902e-19 $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_M1010_g N_noxref_6_c_694_n 9.8258e-19 $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_M1008_g N_noxref_6_c_694_n 0.00120747f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_287_n N_noxref_6_c_694_n 0.00640715f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_290_n N_noxref_6_c_694_n 0.00582647f $X=1.1 $Y=0.56 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_249_n N_noxref_6_c_694_n 0.00138244f $X=1.42 $Y=0.82 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_250_n N_noxref_6_c_694_n 5.60679e-19 $X=1.507 $Y=1.075 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_251_n N_noxref_6_c_694_n 6.3334e-19 $X=1.507 $Y=1.445 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_252_n N_noxref_6_c_694_n 8.56901e-19 $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_268_n N_noxref_6_c_694_n 0.00146721f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_254_n N_noxref_6_c_694_n 2.91981e-19 $X=1.507 $Y=1.16 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_255_n N_noxref_6_c_694_n 0.00171247f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_M1001_g N_noxref_6_c_695_n 4.70964e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_M1005_g N_noxref_6_c_695_n 0.00224266f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_M1006_g N_noxref_6_c_695_n 0.00227359f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_M1008_g N_noxref_6_c_695_n 5.1822e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_250_n N_noxref_6_c_695_n 6.76651e-19 $X=1.507 $Y=1.075 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_251_n N_noxref_6_c_695_n 0.00161112f $X=1.507 $Y=1.445 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_252_n N_noxref_6_c_695_n 0.00384274f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_255_n N_noxref_6_c_695_n 0.0124694f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1001_g N_noxref_6_c_696_n 3.47972e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1005_g N_noxref_6_c_696_n 0.0022224f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_M1006_g N_noxref_6_c_696_n 0.00221683f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_250_n N_noxref_6_c_696_n 4.98958e-19 $X=1.507 $Y=1.075 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_251_n N_noxref_6_c_696_n 0.00179882f $X=1.507 $Y=1.445 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_252_n N_noxref_6_c_696_n 0.00383285f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_255_n N_noxref_6_c_696_n 0.013073f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_247_n N_VGND_M1007_s 0.00131614f $X=1.015 $Y=0.82 $X2=-1.26
+ $Y2=-1.17
cc_392 N_A_27_47#_c_249_n N_VGND_M1021_s 0.00295051f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_273_n N_VGND_c_935_n 0.0117314f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_247_n N_VGND_c_935_n 0.0220716f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_290_n N_VGND_c_935_n 0.0115438f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_396 N_A_27_47#_M1000_g N_VGND_c_936_n 0.00758618f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_397 N_A_27_47#_M1003_g N_VGND_c_936_n 8.11501e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_398 N_A_27_47#_c_290_n N_VGND_c_936_n 0.0175118f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_399 N_A_27_47#_c_249_n N_VGND_c_936_n 0.0182886f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_400 N_A_27_47#_c_252_n N_VGND_c_936_n 0.00255027f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_401 N_A_27_47#_M1000_g N_VGND_c_937_n 8.11501e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_402 N_A_27_47#_M1003_g N_VGND_c_937_n 0.00730885f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_403 N_A_27_47#_M1009_g N_VGND_c_937_n 0.00730885f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_404 N_A_27_47#_M1010_g N_VGND_c_937_n 8.11737e-19 $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_405 N_A_27_47#_M1009_g N_VGND_c_938_n 5.77551e-19 $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_406 N_A_27_47#_M1010_g N_VGND_c_938_n 0.00768852f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_407 N_A_27_47#_M1014_g N_VGND_c_938_n 0.00768852f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_408 N_A_27_47#_M1016_g N_VGND_c_938_n 5.77787e-19 $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_409 N_A_27_47#_M1014_g N_VGND_c_939_n 0.00350562f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_410 N_A_27_47#_M1016_g N_VGND_c_939_n 0.00350562f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_411 N_A_27_47#_M1014_g N_VGND_c_940_n 5.77787e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_412 N_A_27_47#_M1016_g N_VGND_c_940_n 0.00768852f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A_27_47#_M1017_g N_VGND_c_940_n 0.00768852f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_414 N_A_27_47#_M1018_g N_VGND_c_940_n 5.77551e-19 $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_415 N_A_27_47#_M1017_g N_VGND_c_941_n 9.61933e-19 $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_416 N_A_27_47#_M1018_g N_VGND_c_941_n 0.0118037f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_417 N_A_27_47#_c_247_n N_VGND_c_942_n 0.00295005f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_290_n N_VGND_c_942_n 0.0113055f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_419 N_A_27_47#_c_249_n N_VGND_c_942_n 0.00295005f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_420 N_A_27_47#_M1000_g N_VGND_c_944_n 0.0046653f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_421 N_A_27_47#_M1003_g N_VGND_c_944_n 0.00350562f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_422 N_A_27_47#_M1009_g N_VGND_c_946_n 0.00350562f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A_27_47#_M1010_g N_VGND_c_946_n 0.00350562f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_424 N_A_27_47#_M1017_g N_VGND_R24_noxref_neg 0.00214313f $X=4.25 $Y=0.56
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_M1018_g N_VGND_R24_noxref_neg 0.00102843f $X=4.67 $Y=0.56
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_273_n N_VGND_c_951_n 0.0115672f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_427 N_A_27_47#_c_247_n N_VGND_c_951_n 0.00295005f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_M1017_g N_VGND_c_952_n 0.0035053f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_429 N_A_27_47#_M1018_g N_VGND_c_952_n 0.0046653f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_430 N_A_27_47#_M1007_d N_VGND_c_960_n 0.00361805f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_M1012_d N_VGND_c_960_n 0.00410807f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1000_g N_VGND_c_960_n 0.0066984f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_433 N_A_27_47#_M1003_g N_VGND_c_960_n 0.0066984f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_434 N_A_27_47#_M1009_g N_VGND_c_960_n 0.0066984f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_435 N_A_27_47#_M1010_g N_VGND_c_960_n 0.00418574f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_436 N_A_27_47#_M1014_g N_VGND_c_960_n 0.00418574f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_437 N_A_27_47#_M1016_g N_VGND_c_960_n 0.00418574f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_438 N_A_27_47#_M1017_g N_VGND_c_960_n 0.00418516f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A_27_47#_M1018_g N_VGND_c_960_n 0.0066984f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A_27_47#_c_273_n N_VGND_c_960_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_441 N_A_27_47#_c_247_n N_VGND_c_960_n 0.00892758f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_290_n N_VGND_c_960_n 0.00642029f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_443 N_A_27_47#_c_249_n N_VGND_c_960_n 0.00669036f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_444 N_A_27_47#_c_264_n N_X_c_1086_n 0.00401157f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_445 N_A_27_47#_c_248_n N_X_c_1086_n 0.00176862f $X=0.345 $Y=0.82 $X2=0 $Y2=0
cc_446 N_A_27_47#_c_266_n N_X_c_1086_n 0.00228854f $X=0.425 $Y=1.53 $X2=0 $Y2=0
cc_447 N_A_27_47#_M1007_d N_X_R23_noxref_pos 0.00181957f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_M1012_d N_X_R23_noxref_pos 9.81339e-19 $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_264_n N_X_R23_noxref_pos 0.00954548f $X=0.26 $Y=1.63 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_273_n N_X_R23_noxref_pos 0.00389194f $X=0.26 $Y=0.56 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_247_n N_X_R23_noxref_pos 0.00150005f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_248_n N_X_R23_noxref_pos 0.00136491f $X=0.345 $Y=0.82 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_265_n N_X_R23_noxref_pos 0.00197585f $X=0.935 $Y=1.53 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_266_n N_X_R23_noxref_pos 0.00211114f $X=0.425 $Y=1.53 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_287_n N_X_R23_noxref_pos 0.00272412f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_290_n N_X_R23_noxref_pos 0.00114294f $X=1.1 $Y=0.56 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_268_n N_X_R23_noxref_pos 2.2498e-19 $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_552_n N_noxref_6_M1001_s 0.00851965f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_459 N_VPWR_c_552_n N_noxref_6_M1006_s 0.00664387f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_552_n N_noxref_6_M1011_s 0.00570907f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_461 N_VPWR_R25_noxref_neg N_noxref_6_M1019_s 0.00338561f $X=4.46 $Y=2.875
+ $X2=0 $Y2=0
cc_462 N_VPWR_c_552_n N_noxref_6_M1019_s 0.00891135f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_463 N_VPWR_c_554_n N_noxref_6_c_720_n 0.0184767f $X=1.52 $Y=2 $X2=0 $Y2=0
cc_464 N_VPWR_c_555_n N_noxref_6_c_720_n 0.0362016f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_465 N_VPWR_c_564_n N_noxref_6_c_720_n 0.0131197f $X=2.195 $Y=2.72 $X2=0 $Y2=0
cc_466 N_VPWR_c_552_n N_noxref_6_c_720_n 0.00629235f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_467 N_VPWR_M1005_d N_noxref_6_c_697_n 0.00138461f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_555_n N_noxref_6_c_697_n 0.0179526f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_469 N_VPWR_c_555_n N_noxref_6_c_740_n 0.0361787f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_470 N_VPWR_c_566_n N_noxref_6_c_740_n 0.012072f $X=3.035 $Y=2.72 $X2=0 $Y2=0
cc_471 N_VPWR_c_552_n N_noxref_6_c_740_n 0.00640231f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_472 N_VPWR_M1008_d N_noxref_6_c_699_n 0.00185611f $X=3.065 $Y=1.485 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_556_n N_noxref_6_c_699_n 0.0132093f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_474 N_VPWR_c_557_n N_noxref_6_c_859_n 0.0113958f $X=3.875 $Y=2.72 $X2=0 $Y2=0
cc_475 N_VPWR_c_552_n N_noxref_6_c_859_n 0.00646998f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_476 N_VPWR_M1015_d N_noxref_6_c_700_n 0.00185611f $X=3.905 $Y=1.485 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_558_n N_noxref_6_c_700_n 0.0132093f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_478 N_VPWR_c_558_n N_noxref_6_c_763_n 0.0295762f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_479 N_VPWR_c_559_n N_noxref_6_c_763_n 0.0428394f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_480 N_VPWR_R25_noxref_neg N_noxref_6_c_763_n 0.00230519f $X=4.46 $Y=2.875
+ $X2=0 $Y2=0
cc_481 N_VPWR_c_571_n N_noxref_6_c_763_n 0.0131197f $X=4.715 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_552_n N_noxref_6_c_763_n 0.00629235f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_c_559_n N_noxref_6_c_692_n 0.00215253f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_484 N_VPWR_R25_noxref_neg N_noxref_6_c_692_n 0.00486541f $X=4.46 $Y=2.875
+ $X2=0 $Y2=0
cc_485 N_VPWR_c_559_n N_noxref_6_c_693_n 0.00954751f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_486 N_VPWR_R25_noxref_neg N_noxref_6_c_693_n 0.00151646f $X=4.46 $Y=2.875
+ $X2=0 $Y2=0
cc_487 N_VPWR_M1013_d N_noxref_6_c_710_n 0.00303829f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_554_n N_noxref_6_c_710_n 0.00361827f $X=1.52 $Y=2 $X2=0 $Y2=0
cc_489 N_VPWR_c_555_n N_noxref_6_c_710_n 0.00485937f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_490 N_VPWR_c_552_n N_noxref_6_c_710_n 0.016322f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_491 N_VPWR_c_553_n N_noxref_6_c_694_n 0.00107119f $X=0.68 $Y=2 $X2=0 $Y2=0
cc_492 N_VPWR_c_554_n N_noxref_6_c_694_n 0.00215163f $X=1.52 $Y=2 $X2=0 $Y2=0
cc_493 N_VPWR_c_555_n N_noxref_6_c_694_n 0.00133918f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_494 N_VPWR_c_556_n N_noxref_6_c_694_n 0.00179516f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_495 N_VPWR_R25_noxref_neg N_noxref_6_c_694_n 0.102351f $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_552_n N_noxref_6_c_694_n 0.0544082f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_497 N_VPWR_c_559_n N_VGND_c_941_n 0.00566773f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_498 N_VPWR_R25_noxref_neg N_VGND_c_941_n 3.34522e-19 $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_499 N_VPWR_R25_noxref_neg N_VGND_c_948_n 0.0131744f $X=4.46 $Y=2.875 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_559_n N_VGND_R24_noxref_neg 4.04958e-19 $X=4.88 $Y=1.66 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_546_n N_VGND_R24_noxref_neg 0.0131744f $X=5.72 $Y=2.72 $X2=0
+ $Y2=0
cc_502 N_VPWR_R25_noxref_neg N_VGND_R24_noxref_neg 0.171841f $X=4.46 $Y=2.875
+ $X2=0 $Y2=0
cc_503 N_VPWR_c_552_n N_X_c_1086_n 8.18796e-19 $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_504 N_VPWR_M1002_d N_X_R23_noxref_pos 0.00196268f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_553_n N_X_R23_noxref_pos 0.00391339f $X=0.68 $Y=2 $X2=0 $Y2=0
cc_506 N_VPWR_c_552_n N_X_R23_noxref_pos 0.0196951f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_507 N_noxref_6_c_710_n N_VGND_M1021_s 6.80213e-19 $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_508 N_noxref_6_c_684_n N_VGND_M1003_s 0.00131614f $X=2.695 $Y=0.82 $X2=0
+ $Y2=0
cc_509 N_noxref_6_c_686_n N_VGND_M1010_s 0.00162006f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_510 N_noxref_6_c_687_n N_VGND_M1016_s 0.00162006f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_511 N_noxref_6_c_694_n N_VGND_c_935_n 0.00111839f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_512 N_noxref_6_c_717_n N_VGND_c_936_n 0.0177989f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_513 N_noxref_6_c_710_n N_VGND_c_936_n 0.00150511f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_514 N_noxref_6_c_694_n N_VGND_c_936_n 0.00139873f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_515 N_noxref_6_c_717_n N_VGND_c_937_n 0.0177989f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_516 N_noxref_6_c_684_n N_VGND_c_937_n 0.0220716f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_517 N_noxref_6_c_739_n N_VGND_c_937_n 0.0177989f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_518 N_noxref_6_c_710_n N_VGND_c_937_n 0.00185669f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_519 N_noxref_6_c_694_n N_VGND_c_937_n 0.00131357f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_520 N_noxref_6_c_686_n N_VGND_c_938_n 0.0158883f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_521 N_noxref_6_c_694_n N_VGND_c_938_n 8.07372e-19 $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_522 N_noxref_6_c_686_n N_VGND_c_939_n 0.00193763f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_523 N_noxref_6_c_898_p N_VGND_c_939_n 0.0113595f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_524 N_noxref_6_c_687_n N_VGND_c_939_n 0.00193763f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_525 N_noxref_6_c_687_n N_VGND_c_940_n 0.0158883f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_526 N_noxref_6_c_761_n N_VGND_c_940_n 0.0175691f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_527 N_noxref_6_c_761_n N_VGND_c_941_n 0.0240782f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_528 N_noxref_6_c_692_n N_VGND_c_941_n 0.00210597f $X=4.75 $Y=1.19 $X2=0 $Y2=0
cc_529 N_noxref_6_c_693_n N_VGND_c_941_n 0.00956372f $X=4.75 $Y=1.19 $X2=0 $Y2=0
cc_530 N_noxref_6_c_717_n N_VGND_c_944_n 0.013084f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_531 N_noxref_6_c_684_n N_VGND_c_944_n 0.00295005f $X=2.695 $Y=0.82 $X2=0
+ $Y2=0
cc_532 N_noxref_6_c_684_n N_VGND_c_946_n 0.00295005f $X=2.695 $Y=0.82 $X2=0
+ $Y2=0
cc_533 N_noxref_6_c_739_n N_VGND_c_946_n 0.0120358f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_534 N_noxref_6_c_686_n N_VGND_c_946_n 0.00193763f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_535 N_noxref_6_M1017_d N_VGND_R24_noxref_neg 0.00338189f $X=4.325 $Y=0.235
+ $X2=0 $Y2=0
cc_536 N_noxref_6_c_761_n N_VGND_R24_noxref_neg 0.00229539f $X=4.46 $Y=0.56
+ $X2=0 $Y2=0
cc_537 N_noxref_6_c_692_n N_VGND_R24_noxref_neg 0.00547878f $X=4.75 $Y=1.19
+ $X2=0 $Y2=0
cc_538 N_noxref_6_c_693_n N_VGND_R24_noxref_neg 0.00167545f $X=4.75 $Y=1.19
+ $X2=0 $Y2=0
cc_539 N_noxref_6_c_694_n N_VGND_R24_noxref_neg 0.102351f $X=2.05 $Y=1.36 $X2=0
+ $Y2=0
cc_540 N_noxref_6_c_687_n N_VGND_c_952_n 0.0011009f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_541 N_noxref_6_c_761_n N_VGND_c_952_n 0.0131197f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_542 N_noxref_6_c_691_n N_VGND_c_952_n 8.77886e-19 $X=4.417 $Y=0.82 $X2=0
+ $Y2=0
cc_543 N_noxref_6_M1000_d N_VGND_c_960_n 0.0084881f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_544 N_noxref_6_M1009_d N_VGND_c_960_n 0.00508982f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_545 N_noxref_6_M1014_d N_VGND_c_960_n 0.00266406f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_546 N_noxref_6_M1017_d N_VGND_c_960_n 0.00784344f $X=4.325 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_noxref_6_c_717_n N_VGND_c_960_n 0.00628629f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_548 N_noxref_6_c_684_n N_VGND_c_960_n 0.0113794f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_549 N_noxref_6_c_739_n N_VGND_c_960_n 0.00639525f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_550 N_noxref_6_c_686_n N_VGND_c_960_n 0.00895872f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_551 N_noxref_6_c_898_p N_VGND_c_960_n 0.0064623f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_552 N_noxref_6_c_687_n N_VGND_c_960_n 0.00691507f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_553 N_noxref_6_c_761_n N_VGND_c_960_n 0.00629235f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_554 N_noxref_6_c_691_n N_VGND_c_960_n 0.0021633f $X=4.417 $Y=0.82 $X2=0 $Y2=0
cc_555 N_noxref_6_c_710_n N_VGND_c_960_n 0.0157742f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_556 N_noxref_6_c_694_n N_VGND_c_960_n 0.0539201f $X=2.05 $Y=1.36 $X2=0 $Y2=0
cc_557 N_noxref_6_c_695_n N_VGND_c_960_n 0.0156542f $X=2.475 $Y=1.19 $X2=0 $Y2=0
cc_558 N_noxref_6_c_694_n noxref_9 0.00673347f $X=2.05 $Y=1.36 $X2=-1.26
+ $Y2=-1.17
cc_559 N_noxref_6_c_694_n noxref_10 0.00673347f $X=2.05 $Y=1.36 $X2=-1.26
+ $Y2=-1.17
cc_560 N_VGND_c_960_n N_X_c_1086_n 8.18796e-19 $X=5.28 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_960_n N_X_c_1087_n 0.00174134f $X=5.28 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_935_n N_X_R23_noxref_pos 0.00547012f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_563 N_VGND_c_960_n N_X_R23_noxref_pos 0.0196457f $X=5.28 $Y=0 $X2=0 $Y2=0

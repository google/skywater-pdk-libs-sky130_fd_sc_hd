* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_16.spice.pex
* Created: Thu Aug 27 14:23:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%A 3 7 11 15 19 23 27 31 35 39
+ 43 47 51 55 59 63 67 71 73 74 77 81 85 89 93 97 101 105 109 113 117 121 125
+ 129 133 137 141 145 149 153 157 161 163 165 170 171 172 174 212 213
r355 211 213 16.8304 $w=3.6e-07 $l=1.05e-07 $layer=POLY_cond $X=10.46 $Y=1.17
+ $X2=10.565 $Y2=1.17
r356 211 212 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.46
+ $Y=1.16 $X2=10.46 $Y2=1.16
r357 209 211 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=10.135 $Y=1.17
+ $X2=10.46 $Y2=1.17
r358 208 209 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=9.705 $Y=1.17
+ $X2=10.135 $Y2=1.17
r359 207 208 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=9.275 $Y=1.17
+ $X2=9.705 $Y2=1.17
r360 205 207 28.0507 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=9.1 $Y=1.17
+ $X2=9.275 $Y2=1.17
r361 205 206 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.1
+ $Y=1.16 $X2=9.1 $Y2=1.16
r362 203 205 40.8738 $w=3.6e-07 $l=2.55e-07 $layer=POLY_cond $X=8.845 $Y=1.17
+ $X2=9.1 $Y2=1.17
r363 202 203 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=8.415 $Y=1.17
+ $X2=8.845 $Y2=1.17
r364 201 202 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=7.985 $Y=1.17
+ $X2=8.415 $Y2=1.17
r365 200 201 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=7.555 $Y=1.17
+ $X2=7.985 $Y2=1.17
r366 199 200 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=7.125 $Y=1.17
+ $X2=7.555 $Y2=1.17
r367 198 199 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=6.695 $Y=1.17
+ $X2=7.125 $Y2=1.17
r368 197 198 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=6.265 $Y=1.17
+ $X2=6.695 $Y2=1.17
r369 196 197 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=5.835 $Y=1.17
+ $X2=6.265 $Y2=1.17
r370 195 196 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=5.405 $Y=1.17
+ $X2=5.835 $Y2=1.17
r371 193 194 74.5346 $w=3.6e-07 $l=4.65e-07 $layer=POLY_cond $X=4.355 $Y=1.17
+ $X2=4.82 $Y2=1.17
r372 192 193 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=3.925 $Y=1.17
+ $X2=4.355 $Y2=1.17
r373 191 192 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=3.495 $Y=1.17
+ $X2=3.925 $Y2=1.17
r374 190 191 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=3.065 $Y=1.17
+ $X2=3.495 $Y2=1.17
r375 189 190 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=2.635 $Y=1.17
+ $X2=3.065 $Y2=1.17
r376 188 189 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=2.205 $Y=1.17
+ $X2=2.635 $Y2=1.17
r377 186 188 40.8738 $w=3.6e-07 $l=2.55e-07 $layer=POLY_cond $X=1.95 $Y=1.17
+ $X2=2.205 $Y2=1.17
r378 184 186 28.0507 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=1.775 $Y=1.17
+ $X2=1.95 $Y2=1.17
r379 183 184 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=1.345 $Y=1.17
+ $X2=1.775 $Y2=1.17
r380 182 183 68.9245 $w=3.6e-07 $l=4.3e-07 $layer=POLY_cond $X=0.915 $Y=1.17
+ $X2=1.345 $Y2=1.17
r381 180 182 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=0.59 $Y=1.17
+ $X2=0.915 $Y2=1.17
r382 180 181 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r383 177 180 16.8304 $w=3.6e-07 $l=1.05e-07 $layer=POLY_cond $X=0.485 $Y=1.17
+ $X2=0.59 $Y2=1.17
r384 175 212 17.2866 $w=3.78e-07 $l=5.7e-07 $layer=LI1_cond $X=9.89 $Y=1.085
+ $X2=10.46 $Y2=1.085
r385 175 206 23.9587 $w=3.78e-07 $l=7.9e-07 $layer=LI1_cond $X=9.89 $Y=1.085
+ $X2=9.1 $Y2=1.085
r386 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=1.19
+ $X2=9.89 $Y2=1.19
r387 172 174 0.314386 $w=2.3e-07 $l=4.9e-07 $layer=MET1_cond $X=9.4 $Y=1.19
+ $X2=9.89 $Y2=1.19
r388 170 172 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.285 $Y=1.19
+ $X2=9.4 $Y2=1.19
r389 170 171 8.74998 $w=1.4e-07 $l=7.07e-06 $layer=MET1_cond $X=9.285 $Y=1.19
+ $X2=2.215 $Y2=1.19
r390 165 171 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=2.1 $Y=1.19
+ $X2=2.215 $Y2=1.19
r391 165 167 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=2.1 $Y=1.19
+ $X2=2.07 $Y2=1.19
r392 163 181 41.2453 $w=3.78e-07 $l=1.36e-06 $layer=LI1_cond $X=1.95 $Y=1.085
+ $X2=0.59 $Y2=1.085
r393 163 186 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r394 163 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.19
r395 159 213 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=10.565 $Y=1.35
+ $X2=10.565 $Y2=1.17
r396 159 161 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.565 $Y=1.35
+ $X2=10.565 $Y2=1.985
r397 155 209 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=10.135 $Y=1.35
+ $X2=10.135 $Y2=1.17
r398 155 157 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.135 $Y=1.35
+ $X2=10.135 $Y2=1.985
r399 151 208 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=9.705 $Y=1.35
+ $X2=9.705 $Y2=1.17
r400 151 153 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.705 $Y=1.35
+ $X2=9.705 $Y2=1.985
r401 147 207 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=9.275 $Y=1.35
+ $X2=9.275 $Y2=1.17
r402 147 149 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.275 $Y=1.35
+ $X2=9.275 $Y2=1.985
r403 143 203 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.845 $Y=1.35
+ $X2=8.845 $Y2=1.17
r404 143 145 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.845 $Y=1.35
+ $X2=8.845 $Y2=1.985
r405 139 203 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.845 $Y=0.99
+ $X2=8.845 $Y2=1.17
r406 139 141 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=8.845 $Y=0.99
+ $X2=8.845 $Y2=0.445
r407 135 202 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.415 $Y=1.35
+ $X2=8.415 $Y2=1.17
r408 135 137 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.415 $Y=1.35
+ $X2=8.415 $Y2=1.985
r409 131 202 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.415 $Y=0.99
+ $X2=8.415 $Y2=1.17
r410 131 133 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=8.415 $Y=0.99
+ $X2=8.415 $Y2=0.445
r411 127 201 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.985 $Y=1.35
+ $X2=7.985 $Y2=1.17
r412 127 129 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.985 $Y=1.35
+ $X2=7.985 $Y2=1.985
r413 123 201 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.985 $Y=0.99
+ $X2=7.985 $Y2=1.17
r414 123 125 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.985 $Y=0.99
+ $X2=7.985 $Y2=0.445
r415 119 200 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=1.17
r416 119 121 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=1.985
r417 115 200 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.555 $Y=0.99
+ $X2=7.555 $Y2=1.17
r418 115 117 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.555 $Y=0.99
+ $X2=7.555 $Y2=0.445
r419 111 199 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=1.17
r420 111 113 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=1.985
r421 107 199 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.125 $Y=0.99
+ $X2=7.125 $Y2=1.17
r422 107 109 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.125 $Y=0.99
+ $X2=7.125 $Y2=0.445
r423 103 198 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.17
r424 103 105 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.985
r425 99 198 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.695 $Y=0.99
+ $X2=6.695 $Y2=1.17
r426 99 101 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.695 $Y=0.99
+ $X2=6.695 $Y2=0.445
r427 95 197 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.17
r428 95 97 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.985
r429 91 197 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.265 $Y=0.99
+ $X2=6.265 $Y2=1.17
r430 91 93 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.265 $Y=0.99
+ $X2=6.265 $Y2=0.445
r431 87 196 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.17
r432 87 89 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.985
r433 83 196 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.835 $Y=0.99
+ $X2=5.835 $Y2=1.17
r434 83 85 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.835 $Y=0.99
+ $X2=5.835 $Y2=0.445
r435 79 195 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.17
r436 79 81 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.985
r437 75 195 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.405 $Y=0.99
+ $X2=5.405 $Y2=1.17
r438 75 77 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.405 $Y=0.99
+ $X2=5.405 $Y2=0.445
r439 74 194 12.0217 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=4.895 $Y=1.17
+ $X2=4.82 $Y2=1.17
r440 73 195 12.0217 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.17
+ $X2=5.405 $Y2=1.17
r441 73 74 69.7259 $w=3.6e-07 $l=4.35e-07 $layer=POLY_cond $X=5.33 $Y=1.17
+ $X2=4.895 $Y2=1.17
r442 69 194 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.82 $Y=1.35
+ $X2=4.82 $Y2=1.17
r443 69 71 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.82 $Y=1.35
+ $X2=4.82 $Y2=1.985
r444 65 194 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.82 $Y=0.99
+ $X2=4.82 $Y2=1.17
r445 65 67 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.82 $Y=0.99
+ $X2=4.82 $Y2=0.445
r446 61 193 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.355 $Y2=1.17
r447 61 63 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.355 $Y2=1.985
r448 57 193 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.355 $Y=0.99
+ $X2=4.355 $Y2=1.17
r449 57 59 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.355 $Y=0.99
+ $X2=4.355 $Y2=0.445
r450 53 192 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=1.17
r451 53 55 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=1.985
r452 49 192 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.925 $Y=0.99
+ $X2=3.925 $Y2=1.17
r453 49 51 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.925 $Y=0.99
+ $X2=3.925 $Y2=0.445
r454 45 191 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=1.17
r455 45 47 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=1.985
r456 41 191 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.495 $Y=0.99
+ $X2=3.495 $Y2=1.17
r457 41 43 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.495 $Y=0.99
+ $X2=3.495 $Y2=0.445
r458 37 190 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=1.17
r459 37 39 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=1.985
r460 33 190 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.065 $Y=0.99
+ $X2=3.065 $Y2=1.17
r461 33 35 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.065 $Y=0.99
+ $X2=3.065 $Y2=0.445
r462 29 189 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=1.17
r463 29 31 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=1.985
r464 25 189 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.635 $Y=0.99
+ $X2=2.635 $Y2=1.17
r465 25 27 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.635 $Y=0.99
+ $X2=2.635 $Y2=0.445
r466 21 188 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=1.17
r467 21 23 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=1.985
r468 17 188 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.205 $Y=0.99
+ $X2=2.205 $Y2=1.17
r469 17 19 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.205 $Y=0.99
+ $X2=2.205 $Y2=0.445
r470 13 184 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.775 $Y=1.35
+ $X2=1.775 $Y2=1.17
r471 13 15 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.775 $Y=1.35
+ $X2=1.775 $Y2=1.985
r472 9 183 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.345 $Y=1.35
+ $X2=1.345 $Y2=1.17
r473 9 11 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.345 $Y=1.35
+ $X2=1.345 $Y2=1.985
r474 5 182 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.915 $Y=1.35
+ $X2=0.915 $Y2=1.17
r475 5 7 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.915 $Y=1.35
+ $X2=0.915 $Y2=1.985
r476 1 177 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.485 $Y=1.35
+ $X2=0.485 $Y2=1.17
r477 1 3 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.485 $Y=1.35
+ $X2=0.485 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%KAPWR 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 62 67 68 72 73 77 78 81 82 83 86 87 88 92 93 97 98 102 103 107 108 112
+ 113 117 118 122 125 135 138 143 160 163 168 173 178 183 188 195
r245 125 128 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.275 $Y=1.66
+ $X2=0.275 $Y2=2.21
r246 122 195 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.215 $Y=2.21
+ $X2=0.36 $Y2=2.21
r247 122 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.215 $Y=2.21
+ $X2=0.215 $Y2=2.21
r248 121 188 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=10.775 $Y=2.21
+ $X2=10.775 $Y2=2
r249 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.805 $Y=2.21
+ $X2=10.805 $Y2=2.21
r250 116 183 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=9.92 $Y=2.21
+ $X2=9.92 $Y2=2
r251 115 118 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=9.905 $Y=2.21
+ $X2=10.05 $Y2=2.21
r252 115 117 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=9.905 $Y=2.21
+ $X2=9.76 $Y2=2.21
r253 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.905 $Y=2.21
+ $X2=9.905 $Y2=2.21
r254 113 117 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=9.19 $Y=2.24
+ $X2=9.76 $Y2=2.24
r255 111 178 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=9.06 $Y=2.21
+ $X2=9.06 $Y2=2
r256 110 113 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=9.045 $Y=2.21
+ $X2=9.19 $Y2=2.21
r257 110 112 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=9.045 $Y=2.21
+ $X2=8.9 $Y2=2.21
r258 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.045 $Y=2.21
+ $X2=9.045 $Y2=2.21
r259 108 112 0.414474 $w=2e-07 $l=5.4e-07 $layer=MET1_cond $X=8.36 $Y=2.24
+ $X2=8.9 $Y2=2.24
r260 106 173 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8.2 $Y=2.21
+ $X2=8.2 $Y2=2
r261 105 108 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=8.215 $Y=2.21
+ $X2=8.36 $Y2=2.21
r262 105 107 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=8.215 $Y=2.21
+ $X2=8.07 $Y2=2.21
r263 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.215 $Y=2.21
+ $X2=8.215 $Y2=2.21
r264 103 107 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=7.46 $Y=2.24
+ $X2=8.07 $Y2=2.24
r265 101 168 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.34 $Y=2.21
+ $X2=7.34 $Y2=2
r266 100 103 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.315 $Y=2.21
+ $X2=7.46 $Y2=2.21
r267 100 102 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=7.315 $Y=2.21
+ $X2=7.17 $Y2=2.21
r268 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.315 $Y=2.21
+ $X2=7.315 $Y2=2.21
r269 98 102 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=6.6 $Y=2.24
+ $X2=7.17 $Y2=2.24
r270 96 163 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.48 $Y=2.21
+ $X2=6.48 $Y2=2
r271 95 98 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=6.455 $Y=2.21
+ $X2=6.6 $Y2=2.21
r272 95 97 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=6.455 $Y=2.21
+ $X2=6.31 $Y2=2.21
r273 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.455 $Y=2.21
+ $X2=6.455 $Y2=2.21
r274 93 97 0.483553 $w=2e-07 $l=6.3e-07 $layer=MET1_cond $X=5.68 $Y=2.24
+ $X2=6.31 $Y2=2.24
r275 91 160 1.51883 $w=6.28e-07 $l=8e-08 $layer=LI1_cond $X=5.535 $Y=2.15
+ $X2=5.615 $Y2=2.15
r276 90 93 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.535 $Y=2.21
+ $X2=5.68 $Y2=2.21
r277 90 92 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.535 $Y=2.21
+ $X2=5.39 $Y2=2.21
r278 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.535 $Y=2.21
+ $X2=5.535 $Y2=2.21
r279 88 92 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=4.78 $Y=2.24
+ $X2=5.39 $Y2=2.24
r280 86 153 0.854342 $w=6.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.635 $Y=2.15
+ $X2=4.59 $Y2=2.15
r281 85 88 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.635 $Y=2.21
+ $X2=4.78 $Y2=2.21
r282 85 87 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.635 $Y=2.21
+ $X2=4.49 $Y2=2.21
r283 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=2.21
+ $X2=4.635 $Y2=2.21
r284 83 87 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=3.92 $Y=2.24
+ $X2=4.49 $Y2=2.24
r285 81 148 1.23405 $w=6.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.775 $Y=2.15
+ $X2=3.71 $Y2=2.15
r286 80 83 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.775 $Y=2.21
+ $X2=3.92 $Y2=2.21
r287 80 82 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.775 $Y=2.21
+ $X2=3.63 $Y2=2.21
r288 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.775 $Y=2.21
+ $X2=3.775 $Y2=2.21
r289 78 82 0.483553 $w=2e-07 $l=6.3e-07 $layer=MET1_cond $X=3 $Y=2.24 $X2=3.63
+ $Y2=2.24
r290 76 143 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=2.21
+ $X2=2.85 $Y2=2
r291 75 78 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.855 $Y=2.21
+ $X2=3 $Y2=2.21
r292 75 77 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.855 $Y=2.21
+ $X2=2.71 $Y2=2.21
r293 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.855 $Y=2.21
+ $X2=2.855 $Y2=2.21
r294 73 77 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=2.12 $Y=2.24
+ $X2=2.71 $Y2=2.24
r295 71 138 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.99 $Y=2.21
+ $X2=1.99 $Y2=2
r296 70 73 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=2.12 $Y2=2.21
r297 70 72 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=1.83 $Y2=2.21
r298 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.975 $Y=2.21
+ $X2=1.975 $Y2=2.21
r299 68 72 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=1.22 $Y=2.24
+ $X2=1.83 $Y2=2.24
r300 67 195 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=0.93 $Y=2.24
+ $X2=0.36 $Y2=2.24
r301 66 135 1.0442 $w=6.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.075 $Y=2.15
+ $X2=1.13 $Y2=2.15
r302 65 68 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.075 $Y=2.21
+ $X2=1.22 $Y2=2.21
r303 65 67 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.075 $Y=2.21
+ $X2=0.93 $Y2=2.21
r304 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.075 $Y=2.21
+ $X2=1.075 $Y2=2.21
r305 62 120 0.0771209 $w=2.56e-07 $l=1.59295e-07 $layer=MET1_cond $X=10.66
+ $Y=2.24 $X2=10.805 $Y2=2.21
r306 62 118 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=10.66 $Y=2.24
+ $X2=10.05 $Y2=2.24
r307 13 188 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=10.64
+ $Y=1.485 $X2=10.775 $Y2=2
r308 12 183 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=9.78
+ $Y=1.485 $X2=9.92 $Y2=2
r309 11 178 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=8.92
+ $Y=1.485 $X2=9.06 $Y2=2
r310 10 173 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=8.06
+ $Y=1.485 $X2=8.2 $Y2=2
r311 9 168 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=7.2
+ $Y=1.485 $X2=7.34 $Y2=2
r312 8 163 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=6.34
+ $Y=1.485 $X2=6.48 $Y2=2
r313 7 160 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.48
+ $Y=1.485 $X2=5.615 $Y2=2
r314 6 153 300 $w=1.7e-07 $l=5.89597e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.485 $X2=4.59 $Y2=2
r315 5 148 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=3.57
+ $Y=1.485 $X2=3.71 $Y2=2
r316 4 143 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=1.485 $X2=2.85 $Y2=2
r317 3 138 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1.85
+ $Y=1.485 $X2=1.99 $Y2=2
r318 2 135 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=0.99
+ $Y=1.485 $X2=1.13 $Y2=2
r319 1 128 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.34
r320 1 125 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%Y 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 18 19 20 61 63 65 69 73 77 81 85 89 93 97 103 107 111 115 119
+ 123 127 131 135 142 144 146 148 149 151 153 155 157 159 161 162 167
r354 165 167 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.255 $Y=1.54
+ $X2=5.29 $Y2=1.54
r355 162 165 3.17047 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=5.08 $Y=1.54
+ $X2=5.255 $Y2=1.54
r356 162 167 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=1.54
+ $X2=5.29 $Y2=1.54
r357 149 162 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=5.315 $Y2=1.54
r358 149 151 2.53577 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.925 $Y=1.54
+ $X2=6.05 $Y2=1.54
r359 136 159 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=1.56
+ $X2=9.49 $Y2=1.56
r360 135 161 3.16207 $w=2.1e-07 $l=1.07e-07 $layer=LI1_cond $X=10.265 $Y=1.56
+ $X2=10.372 $Y2=1.56
r361 135 136 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=10.265 $Y=1.56
+ $X2=9.575 $Y2=1.56
r362 132 157 2.77723 $w=2.1e-07 $l=1.34629e-07 $layer=LI1_cond $X=8.755 $Y=1.56
+ $X2=8.63 $Y2=1.54
r363 131 159 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.405 $Y=1.56
+ $X2=9.49 $Y2=1.56
r364 131 132 34.329 $w=2.08e-07 $l=6.5e-07 $layer=LI1_cond $X=9.405 $Y=1.56
+ $X2=8.755 $Y2=1.56
r365 125 157 3.33195 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.63 $Y=1.415
+ $X2=8.63 $Y2=1.54
r366 125 127 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=8.63 $Y=1.415
+ $X2=8.63 $Y2=0.445
r367 124 155 2.53577 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.895 $Y=1.54
+ $X2=7.77 $Y2=1.54
r368 123 157 2.77723 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.505 $Y=1.54
+ $X2=8.63 $Y2=1.54
r369 123 124 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=8.505 $Y=1.54
+ $X2=7.895 $Y2=1.54
r370 117 155 3.59786 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.77 $Y=1.415
+ $X2=7.77 $Y2=1.54
r371 117 119 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=7.77 $Y=1.415
+ $X2=7.77 $Y2=0.445
r372 116 153 2.53577 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.035 $Y=1.54
+ $X2=6.91 $Y2=1.54
r373 115 155 2.53577 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.645 $Y=1.54
+ $X2=7.77 $Y2=1.54
r374 115 116 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.645 $Y=1.54
+ $X2=7.035 $Y2=1.54
r375 109 153 3.59786 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.91 $Y=1.415
+ $X2=6.91 $Y2=1.54
r376 109 111 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=6.91 $Y=1.415
+ $X2=6.91 $Y2=0.445
r377 108 151 2.53577 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.175 $Y=1.54
+ $X2=6.05 $Y2=1.54
r378 107 153 2.53577 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=6.91 $Y2=1.54
r379 107 108 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=6.175 $Y2=1.54
r380 101 151 3.59786 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.05 $Y=1.415
+ $X2=6.05 $Y2=1.54
r381 101 103 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=6.05 $Y=1.415
+ $X2=6.05 $Y2=0.445
r382 95 162 2.93124 $w=3.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.08 $Y=1.415
+ $X2=5.08 $Y2=1.54
r383 95 97 31.9391 $w=3.48e-07 $l=9.7e-07 $layer=LI1_cond $X=5.08 $Y=1.415
+ $X2=5.08 $Y2=0.445
r384 94 148 2.46758 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.255 $Y=1.54
+ $X2=4.135 $Y2=1.54
r385 93 162 3.17047 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=5.08 $Y2=1.54
r386 93 94 29.9635 $w=2.48e-07 $l=6.5e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=4.255 $Y2=1.54
r387 87 148 3.67597 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=4.135 $Y=1.415
+ $X2=4.135 $Y2=1.54
r388 87 89 46.5779 $w=2.38e-07 $l=9.7e-07 $layer=LI1_cond $X=4.135 $Y=1.415
+ $X2=4.135 $Y2=0.445
r389 86 146 2.56953 $w=2.5e-07 $l=1.28e-07 $layer=LI1_cond $X=3.41 $Y=1.54
+ $X2=3.282 $Y2=1.54
r390 85 148 2.46758 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.015 $Y=1.54
+ $X2=4.135 $Y2=1.54
r391 85 86 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=4.015 $Y=1.54
+ $X2=3.41 $Y2=1.54
r392 79 146 3.55971 $w=2.55e-07 $l=1.25e-07 $layer=LI1_cond $X=3.282 $Y=1.415
+ $X2=3.282 $Y2=1.54
r393 79 81 43.838 $w=2.53e-07 $l=9.7e-07 $layer=LI1_cond $X=3.282 $Y=1.415
+ $X2=3.282 $Y2=0.445
r394 78 144 2.5987 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=2.55 $Y=1.54
+ $X2=2.437 $Y2=1.54
r395 77 146 2.56953 $w=2.5e-07 $l=1.27e-07 $layer=LI1_cond $X=3.155 $Y=1.54
+ $X2=3.282 $Y2=1.54
r396 77 78 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=3.155 $Y=1.54
+ $X2=2.55 $Y2=1.54
r397 71 144 3.527 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=2.437 $Y=1.415
+ $X2=2.437 $Y2=1.54
r398 71 73 49.6831 $w=2.23e-07 $l=9.7e-07 $layer=LI1_cond $X=2.437 $Y=1.415
+ $X2=2.437 $Y2=0.445
r399 70 142 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.56
+ $X2=1.56 $Y2=1.56
r400 69 144 2.5987 $w=2.1e-07 $l=1.21589e-07 $layer=LI1_cond $X=2.325 $Y=1.56
+ $X2=2.437 $Y2=1.54
r401 69 70 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=2.325 $Y=1.56
+ $X2=1.645 $Y2=1.56
r402 66 140 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=1.56
+ $X2=0.7 $Y2=1.56
r403 65 142 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.56
+ $X2=1.56 $Y2=1.56
r404 65 66 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.475 $Y=1.56
+ $X2=0.785 $Y2=1.56
r405 61 140 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.7 $Y=1.665
+ $X2=0.7 $Y2=1.56
r406 61 63 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=1.665
+ $X2=0.7 $Y2=2.3
r407 20 161 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=10.21
+ $Y=1.485 $X2=10.35 $Y2=1.62
r408 19 159 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=9.35
+ $Y=1.485 $X2=9.49 $Y2=1.62
r409 18 157 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=1.485 $X2=8.63 $Y2=1.62
r410 17 155 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=7.63
+ $Y=1.485 $X2=7.77 $Y2=1.62
r411 16 153 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=6.77
+ $Y=1.485 $X2=6.91 $Y2=1.62
r412 15 151 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.485 $X2=6.05 $Y2=1.62
r413 14 162 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.485 $X2=5.165 $Y2=1.62
r414 13 148 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=4
+ $Y=1.485 $X2=4.14 $Y2=1.62
r415 12 146 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=3.14
+ $Y=1.485 $X2=3.28 $Y2=1.62
r416 11 144 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=2.28
+ $Y=1.485 $X2=2.42 $Y2=1.62
r417 10 142 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=1.42
+ $Y=1.485 $X2=1.56 $Y2=1.62
r418 9 140 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.7 $Y2=1.62
r419 9 63 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.7 $Y2=2.3
r420 8 127 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.49
+ $Y=0.235 $X2=8.63 $Y2=0.445
r421 7 119 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.63
+ $Y=0.235 $X2=7.77 $Y2=0.445
r422 6 111 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.235 $X2=6.91 $Y2=0.445
r423 5 103 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.235 $X2=6.05 $Y2=0.445
r424 4 97 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=4.895
+ $Y=0.235 $X2=5.065 $Y2=0.445
r425 3 89 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.235 $X2=4.14 $Y2=0.445
r426 2 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.14
+ $Y=0.235 $X2=3.28 $Y2=0.445
r427 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.42 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%VGND 1 2 3 4 5 6 7 8 9 30 34
+ 38 42 46 50 54 58 60 64 67 68 70 71 73 74 76 77 79 80 82 83 85 86 87 88 89 124
+ 125 128
r121 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r122 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r123 122 125 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r124 122 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r125 121 124 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r126 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r127 119 128 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.062 $Y2=0
r128 119 121 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.43 $Y2=0
r129 118 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r130 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r131 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r132 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r133 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r134 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r135 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r136 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r137 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r138 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r139 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r140 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r141 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r142 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r143 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r144 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r145 92 96 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r146 89 97 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.61 $Y2=0
r147 89 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r148 87 117 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.05
+ $Y2=0
r149 87 88 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.202
+ $Y2=0
r150 85 114 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.21 $Y=0 $X2=7.13
+ $Y2=0
r151 85 86 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.21 $Y=0 $X2=7.342
+ $Y2=0
r152 84 117 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=8.05 $Y2=0
r153 84 86 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.342 $Y2=0
r154 82 111 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.35 $Y=0 $X2=6.21
+ $Y2=0
r155 82 83 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=6.35 $Y=0 $X2=6.462
+ $Y2=0
r156 81 114 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=7.13 $Y2=0
r157 81 83 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.462 $Y2=0
r158 79 108 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.49 $Y=0 $X2=5.29
+ $Y2=0
r159 79 80 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.49 $Y=0 $X2=5.622
+ $Y2=0
r160 78 111 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=6.21 $Y2=0
r161 78 80 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.622 $Y2=0
r162 76 105 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.37 $Y2=0
r163 76 77 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.597 $Y2=0
r164 75 108 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=5.29
+ $Y2=0
r165 75 77 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.597
+ $Y2=0
r166 73 102 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.45
+ $Y2=0
r167 73 74 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.712
+ $Y2=0
r168 72 105 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.845 $Y=0
+ $X2=4.37 $Y2=0
r169 72 74 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.845 $Y=0
+ $X2=3.712 $Y2=0
r170 70 99 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.53
+ $Y2=0
r171 70 71 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.852
+ $Y2=0
r172 69 102 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=3.45 $Y2=0
r173 69 71 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=2.852 $Y2=0
r174 67 96 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r175 67 68 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.99
+ $Y2=0
r176 66 99 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=0
+ $X2=2.53 $Y2=0
r177 66 68 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.99
+ $Y2=0
r178 62 128 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=9.062 $Y=0.085
+ $X2=9.062 $Y2=0
r179 62 64 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=9.062 $Y=0.085
+ $X2=9.062 $Y2=0.445
r180 61 88 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.335 $Y=0
+ $X2=8.202 $Y2=0
r181 60 128 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.93 $Y=0
+ $X2=9.062 $Y2=0
r182 60 61 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=8.93 $Y=0
+ $X2=8.335 $Y2=0
r183 56 88 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=8.202 $Y=0.085
+ $X2=8.202 $Y2=0
r184 56 58 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=8.202 $Y=0.085
+ $X2=8.202 $Y2=0.445
r185 52 86 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.342 $Y=0.085
+ $X2=7.342 $Y2=0
r186 52 54 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=7.342 $Y=0.085
+ $X2=7.342 $Y2=0.445
r187 48 83 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=6.462 $Y=0.085
+ $X2=6.462 $Y2=0
r188 48 50 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=6.462 $Y=0.085
+ $X2=6.462 $Y2=0.445
r189 44 80 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.622 $Y=0.085
+ $X2=5.622 $Y2=0
r190 44 46 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=5.622 $Y=0.085
+ $X2=5.622 $Y2=0.445
r191 40 77 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.597 $Y=0.085
+ $X2=4.597 $Y2=0
r192 40 42 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=4.597 $Y=0.085
+ $X2=4.597 $Y2=0.445
r193 36 74 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.712 $Y=0.085
+ $X2=3.712 $Y2=0
r194 36 38 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=3.712 $Y=0.085
+ $X2=3.712 $Y2=0.445
r195 32 71 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.852 $Y=0.085
+ $X2=2.852 $Y2=0
r196 32 34 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=2.852 $Y=0.085
+ $X2=2.852 $Y2=0.445
r197 28 68 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r198 28 30 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.445
r199 9 64 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.92
+ $Y=0.235 $X2=9.06 $Y2=0.445
r200 8 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.06
+ $Y=0.235 $X2=8.2 $Y2=0.445
r201 7 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.235 $X2=7.34 $Y2=0.445
r202 6 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.48 $Y2=0.445
r203 5 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.235 $X2=5.62 $Y2=0.445
r204 4 42 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.235 $X2=4.595 $Y2=0.445
r205 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.445
r206 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.85 $Y2=0.445
r207 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.235 $X2=1.99 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%VPWR 1 8 9
r146 8 9 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r147 4 8 690.246 $w=1.68e-07 $l=1.058e-05 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=10.81 $Y2=2.72
r148 1 9 3.01045 $w=4.8e-07 $l=1.058e-05 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=10.81 $Y2=2.72
r149 1 4 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


* File: sky130_fd_sc_hd__a22oi_2.pxi.spice
* Created: Thu Aug 27 14:02:57 2020
* 
x_PM_SKY130_FD_SC_HD__A22OI_2%B2 N_B2_c_66_n N_B2_M1005_g N_B2_M1001_g
+ N_B2_c_67_n N_B2_M1015_g N_B2_M1012_g B2 B2 N_B2_c_69_n
+ PM_SKY130_FD_SC_HD__A22OI_2%B2
x_PM_SKY130_FD_SC_HD__A22OI_2%B1 N_B1_c_106_n N_B1_M1010_g N_B1_M1000_g
+ N_B1_c_107_n N_B1_M1011_g N_B1_M1014_g B1 B1 N_B1_c_109_n
+ PM_SKY130_FD_SC_HD__A22OI_2%B1
x_PM_SKY130_FD_SC_HD__A22OI_2%A1 N_A1_c_152_n N_A1_M1006_g N_A1_M1004_g
+ N_A1_c_153_n N_A1_M1007_g N_A1_M1008_g A1 A1 N_A1_c_155_n
+ PM_SKY130_FD_SC_HD__A22OI_2%A1
x_PM_SKY130_FD_SC_HD__A22OI_2%A2 N_A2_c_201_n N_A2_M1002_g N_A2_M1009_g
+ N_A2_c_202_n N_A2_M1003_g N_A2_M1013_g A2 A2 N_A2_c_204_n
+ PM_SKY130_FD_SC_HD__A22OI_2%A2
x_PM_SKY130_FD_SC_HD__A22OI_2%Y N_Y_M1010_s N_Y_M1006_s N_Y_M1001_d N_Y_M1012_d
+ N_Y_M1014_s N_Y_c_243_n N_Y_c_249_n N_Y_c_244_n N_Y_c_255_n N_Y_c_260_n
+ N_Y_c_264_n N_Y_c_245_n Y Y Y Y Y N_Y_c_248_n N_Y_c_242_n
+ PM_SKY130_FD_SC_HD__A22OI_2%Y
x_PM_SKY130_FD_SC_HD__A22OI_2%A_109_297# N_A_109_297#_M1001_s
+ N_A_109_297#_M1000_d N_A_109_297#_M1004_d N_A_109_297#_M1008_d
+ N_A_109_297#_M1013_d N_A_109_297#_c_325_n N_A_109_297#_c_326_n
+ N_A_109_297#_c_327_n N_A_109_297#_c_361_n N_A_109_297#_c_320_n
+ N_A_109_297#_c_331_n N_A_109_297#_c_330_n N_A_109_297#_c_334_n
+ N_A_109_297#_c_321_n N_A_109_297#_c_341_n N_A_109_297#_c_322_n
+ N_A_109_297#_c_323_n N_A_109_297#_c_376_p N_A_109_297#_c_324_n
+ PM_SKY130_FD_SC_HD__A22OI_2%A_109_297#
x_PM_SKY130_FD_SC_HD__A22OI_2%VPWR N_VPWR_M1004_s N_VPWR_M1009_s N_VPWR_c_393_n
+ N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n
+ VPWR VPWR N_VPWR_c_399_n N_VPWR_c_392_n PM_SKY130_FD_SC_HD__A22OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A22OI_2%A_27_47# N_A_27_47#_M1005_d N_A_27_47#_M1015_d
+ N_A_27_47#_M1011_d N_A_27_47#_c_449_n N_A_27_47#_c_452_n N_A_27_47#_c_450_n
+ N_A_27_47#_c_473_p N_A_27_47#_c_451_n PM_SKY130_FD_SC_HD__A22OI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__A22OI_2%VGND N_VGND_M1005_s N_VGND_M1002_s N_VGND_c_486_n
+ N_VGND_c_487_n N_VGND_c_488_n VGND VGND N_VGND_c_490_n N_VGND_c_491_n
+ N_VGND_c_492_n N_VGND_c_493_n PM_SKY130_FD_SC_HD__A22OI_2%VGND
x_PM_SKY130_FD_SC_HD__A22OI_2%A_467_47# N_A_467_47#_M1006_d N_A_467_47#_M1007_d
+ N_A_467_47#_M1003_d N_A_467_47#_c_548_n N_A_467_47#_c_549_n
+ N_A_467_47#_c_561_n N_A_467_47#_c_550_n PM_SKY130_FD_SC_HD__A22OI_2%A_467_47#
cc_1 VNB N_B2_c_66_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_67_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB B2 0.0104987f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_B2_c_69_n 0.0455434f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B1_c_106_n 0.0162451f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B1_c_107_n 0.0191733f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_7 VNB B1 0.00499541f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_B1_c_109_n 0.0349812f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_9 VNB N_A1_c_152_n 0.0197855f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_A1_c_153_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_11 VNB A1 0.00245458f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_12 VNB N_A1_c_155_n 0.041881f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_13 VNB N_A2_c_201_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A2_c_202_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_15 VNB A2 0.0307193f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_16 VNB N_A2_c_204_n 0.0373358f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_17 VNB Y 0.00170628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.0120018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_242_n 0.0092054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_392_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_449_n 0.0161681f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_22 VNB N_A_27_47#_c_450_n 0.00783052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_451_n 0.00289148f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_24 VNB N_VGND_c_486_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_25 VNB N_VGND_c_487_n 0.0609027f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_26 VNB N_VGND_c_488_n 0.00436419f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_27 VNB VGND 0.00436419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_490_n 0.0144524f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_29 VNB N_VGND_c_491_n 0.0201583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_492_n 0.247386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_493_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_467_47#_c_548_n 0.00289221f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_33 VNB N_A_467_47#_c_549_n 0.00874558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_467_47#_c_550_n 0.0182437f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_35 VPB N_B2_M1001_g 0.0259042f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB N_B2_M1012_g 0.0187854f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_37 VPB N_B2_c_69_n 0.00800353f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_38 VPB N_B1_M1000_g 0.0187792f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB N_B1_M1014_g 0.0218338f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_40 VPB N_B1_c_109_n 0.00436553f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_41 VPB N_A1_M1004_g 0.0227213f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_42 VPB N_A1_M1008_g 0.0187854f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_43 VPB N_A1_c_155_n 0.00752771f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_44 VPB N_A2_M1009_g 0.0187854f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB N_A2_M1013_g 0.0259042f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_46 VPB N_A2_c_204_n 0.00484244f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_47 VPB N_Y_c_243_n 0.0305923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_Y_c_244_n 0.00977933f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_49 VPB N_Y_c_245_n 0.00190014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB Y 0.00201265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB Y 0.0051823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_Y_c_248_n 0.00596724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_109_297#_c_320_n 0.0105087f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_54 VPB N_A_109_297#_c_321_n 0.00190103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_109_297#_c_322_n 0.00963526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_109_297#_c_323_n 0.0316012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_109_297#_c_324_n 0.00262948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_393_n 0.00410284f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_59 VPB N_VPWR_c_394_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_60 VPB N_VPWR_c_395_n 0.0683005f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_61 VPB N_VPWR_c_396_n 0.00323699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_397_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_63 VPB N_VPWR_c_398_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_64 VPB N_VPWR_c_399_n 0.0242302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_392_n 0.0551673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_B2_c_67_n N_B1_c_106_n 0.0234841f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_67 N_B2_M1012_g N_B1_M1000_g 0.0234841f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_68 B2 B1 0.0116776f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_69 N_B2_c_69_n B1 0.00211269f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B2_c_69_n N_B1_c_109_n 0.0234841f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B2_M1001_g N_Y_c_249_n 0.0147047f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_72 N_B2_M1012_g N_Y_c_249_n 0.0105288f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 B2 N_Y_c_249_n 0.0219027f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_74 N_B2_c_69_n N_Y_c_249_n 0.00208466f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 B2 N_Y_c_244_n 0.0134456f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_76 N_B2_c_69_n N_Y_c_244_n 0.00167075f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B2_M1001_g N_Y_c_255_n 4.72397e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B2_M1012_g N_Y_c_255_n 0.00668438f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B2_M1012_g N_Y_c_245_n 0.00130065f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_80 N_B2_M1001_g N_A_109_297#_c_325_n 0.00556147f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_81 N_B2_M1012_g N_A_109_297#_c_326_n 0.00929389f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_82 N_B2_M1001_g N_A_109_297#_c_327_n 0.00211624f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_83 N_B2_M1001_g N_VPWR_c_395_n 0.00539841f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_84 N_B2_M1012_g N_VPWR_c_395_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_85 N_B2_M1001_g N_VPWR_c_392_n 0.0106541f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_86 N_B2_M1012_g N_VPWR_c_392_n 0.00525341f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_87 N_B2_c_66_n N_A_27_47#_c_452_n 0.0116039f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B2_c_67_n N_A_27_47#_c_452_n 0.0125251f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_89 B2 N_A_27_47#_c_452_n 0.0207498f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B2_c_69_n N_A_27_47#_c_452_n 0.00213849f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_91 B2 N_A_27_47#_c_450_n 0.0126462f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_92 N_B2_c_69_n N_A_27_47#_c_450_n 0.00170625f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B2_c_67_n N_VGND_c_487_n 0.00344532f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B2_c_66_n N_VGND_c_490_n 0.00344532f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B2_c_66_n N_VGND_c_492_n 0.00506656f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B2_c_67_n N_VGND_c_492_n 0.00410391f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B2_c_66_n N_VGND_c_493_n 0.00884363f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B2_c_67_n N_VGND_c_493_n 0.00829944f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_99 N_B1_c_109_n N_A1_c_155_n 0.00368839f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B1_M1000_g N_Y_c_255_n 0.00646869f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B1_M1014_g N_Y_c_255_n 5.43689e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_M1000_g N_Y_c_260_n 0.00900429f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_M1014_g N_Y_c_260_n 0.00992317f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_104 B1 N_Y_c_260_n 0.0223034f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_105 N_B1_c_109_n N_Y_c_260_n 0.00208466f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B1_c_106_n N_Y_c_264_n 0.00257667f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_c_107_n N_Y_c_264_n 0.0120416f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_108 B1 N_Y_c_264_n 0.01589f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B1_c_109_n N_Y_c_264_n 0.00213103f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B1_M1000_g N_Y_c_245_n 9.16882e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_111 B1 N_Y_c_245_n 0.0115197f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B1_M1014_g Y 0.00123943f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B1_c_107_n Y 0.0198608f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_114 B1 Y 0.0163566f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B1_M1000_g N_Y_c_248_n 5.4283e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_M1014_g N_Y_c_248_n 0.00646869f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B1_M1000_g N_A_109_297#_c_326_n 0.00929389f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_B1_M1014_g N_A_109_297#_c_320_n 0.011441f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B1_M1014_g N_A_109_297#_c_330_n 0.00322581f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_B1_M1000_g N_VPWR_c_395_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B1_M1014_g N_VPWR_c_395_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1000_g N_VPWR_c_392_n 0.00525341f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1014_g N_VPWR_c_392_n 0.00660224f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_124 B1 N_A_27_47#_c_452_n 0.00751874f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_125 N_B1_c_106_n N_A_27_47#_c_451_n 0.0123283f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_c_107_n N_A_27_47#_c_451_n 0.00964167f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_127 B1 N_A_27_47#_c_451_n 0.00395343f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_c_106_n N_VGND_c_487_n 0.00357877f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B1_c_107_n N_VGND_c_487_n 0.00357877f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_106_n N_VGND_c_492_n 0.0052923f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_107_n N_VGND_c_492_n 0.00655123f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_106_n N_VGND_c_493_n 0.00126885f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_c_153_n N_A2_c_201_n 0.0190775f $X=3.09 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 N_A1_M1008_g N_A2_M1009_g 0.0190775f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_135 A1 A2 0.0117884f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A1_c_155_n A2 0.00169621f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_137 A1 N_A2_c_204_n 2.11825e-19 $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A1_c_155_n N_A2_c_204_n 0.0190775f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A1_c_152_n Y 0.00411248f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_M1004_g Y 0.00437571f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_141 A1 Y 0.0120635f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_142 N_A1_c_155_n Y 0.0040481f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A1_c_152_n N_Y_c_242_n 0.0108195f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_153_n N_Y_c_242_n 0.00257667f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_145 A1 N_Y_c_242_n 0.0284641f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A1_c_155_n N_Y_c_242_n 0.00480091f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A1_M1004_g N_A_109_297#_c_331_n 0.00202914f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A1_M1004_g N_A_109_297#_c_330_n 0.00783241f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A1_M1008_g N_A_109_297#_c_330_n 5.95406e-19 $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A1_M1004_g N_A_109_297#_c_334_n 0.0109098f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A1_M1008_g N_A_109_297#_c_334_n 0.0118495f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_152 A1 N_A_109_297#_c_334_n 0.024622f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A1_c_155_n N_A_109_297#_c_334_n 0.00208466f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A1_M1004_g N_A_109_297#_c_321_n 9.34284e-19 $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_155 A1 N_A_109_297#_c_321_n 0.0100173f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_155_n N_A_109_297#_c_321_n 0.00269419f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_M1004_g N_A_109_297#_c_341_n 6.43898e-19 $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A1_M1008_g N_A_109_297#_c_341_n 0.00985568f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A1_M1008_g N_A_109_297#_c_324_n 0.00196977f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A1_M1004_g N_VPWR_c_393_n 0.00268723f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A1_M1008_g N_VPWR_c_393_n 0.00146448f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A1_M1004_g N_VPWR_c_395_n 0.00539841f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A1_M1008_g N_VPWR_c_397_n 0.00541359f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A1_M1004_g N_VPWR_c_392_n 0.0107906f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A1_M1008_g N_VPWR_c_392_n 0.00952874f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A1_c_153_n N_VGND_c_486_n 0.00126885f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_c_152_n N_VGND_c_487_n 0.00357877f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_153_n N_VGND_c_487_n 0.00357877f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_152_n N_VGND_c_492_n 0.00655123f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_153_n N_VGND_c_492_n 0.0052923f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_152_n N_A_467_47#_c_548_n 0.00964167f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A1_c_153_n N_A_467_47#_c_548_n 0.0135572f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_173 A1 N_A_467_47#_c_548_n 0.00143613f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A2_M1009_g N_A_109_297#_c_341_n 0.00985568f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A2_M1013_g N_A_109_297#_c_341_n 6.43898e-19 $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A2_M1009_g N_A_109_297#_c_322_n 0.0109098f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1013_g N_A_109_297#_c_322_n 0.0118441f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_178 A2 N_A_109_297#_c_322_n 0.0479471f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A2_c_204_n N_A_109_297#_c_322_n 0.00208466f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A2_M1009_g N_A_109_297#_c_323_n 6.43898e-19 $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A2_M1013_g N_A_109_297#_c_323_n 0.00985568f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A2_M1009_g N_A_109_297#_c_324_n 9.34284e-19 $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_183 A2 N_A_109_297#_c_324_n 0.00341698f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A2_M1009_g N_VPWR_c_394_n 0.00146448f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A2_M1013_g N_VPWR_c_394_n 0.00268723f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A2_M1009_g N_VPWR_c_397_n 0.00541359f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_M1013_g N_VPWR_c_399_n 0.00541359f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_M1009_g N_VPWR_c_392_n 0.00952874f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A2_M1013_g N_VPWR_c_392_n 0.0106001f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A2_c_201_n N_VGND_c_486_n 0.00829944f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_c_202_n N_VGND_c_486_n 0.00884363f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_201_n N_VGND_c_487_n 0.00344532f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_202_n N_VGND_c_491_n 0.00344532f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_201_n N_VGND_c_492_n 0.00410391f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_202_n N_VGND_c_492_n 0.00521643f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_201_n N_A_467_47#_c_549_n 0.0106913f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_202_n N_A_467_47#_c_549_n 0.0116873f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_198 A2 N_A_467_47#_c_549_n 0.0531444f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A2_c_204_n N_A_467_47#_c_549_n 0.00213849f $X=3.93 $Y=1.16 $X2=0 $Y2=0
cc_200 N_Y_c_249_n N_A_109_297#_M1001_s 0.00324353f $X=0.935 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_201 N_Y_c_260_n N_A_109_297#_M1000_d 0.00324353f $X=1.775 $Y=1.57 $X2=0 $Y2=0
cc_202 N_Y_c_249_n N_A_109_297#_c_325_n 0.0147854f $X=0.935 $Y=1.57 $X2=0 $Y2=0
cc_203 N_Y_M1012_d N_A_109_297#_c_326_n 0.00312348f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_Y_c_249_n N_A_109_297#_c_326_n 0.00267672f $X=0.935 $Y=1.57 $X2=0 $Y2=0
cc_205 N_Y_c_255_n N_A_109_297#_c_326_n 0.0158744f $X=1.1 $Y=1.66 $X2=0 $Y2=0
cc_206 N_Y_c_260_n N_A_109_297#_c_326_n 0.00267672f $X=1.775 $Y=1.57 $X2=0 $Y2=0
cc_207 N_Y_c_260_n N_A_109_297#_c_361_n 0.0126293f $X=1.775 $Y=1.57 $X2=0 $Y2=0
cc_208 N_Y_M1014_s N_A_109_297#_c_320_n 0.00480843f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_209 N_Y_c_260_n N_A_109_297#_c_320_n 0.00267672f $X=1.775 $Y=1.57 $X2=0 $Y2=0
cc_210 N_Y_c_248_n N_A_109_297#_c_320_n 0.0249213f $X=1.94 $Y=1.66 $X2=0 $Y2=0
cc_211 N_Y_c_248_n N_A_109_297#_c_330_n 0.0321241f $X=1.94 $Y=1.66 $X2=0 $Y2=0
cc_212 Y N_A_109_297#_c_321_n 0.0131731f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_213 N_Y_c_242_n N_A_109_297#_c_321_n 0.00209868f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_214 N_Y_c_243_n N_VPWR_c_395_n 0.0172841f $X=0.26 $Y=1.8 $X2=0 $Y2=0
cc_215 N_Y_M1001_d N_VPWR_c_392_n 0.00387172f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_216 N_Y_M1012_d N_VPWR_c_392_n 0.00216833f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_217 N_Y_M1014_s N_VPWR_c_392_n 0.00210147f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_218 N_Y_c_243_n N_VPWR_c_392_n 0.00955092f $X=0.26 $Y=1.8 $X2=0 $Y2=0
cc_219 N_Y_c_264_n N_A_27_47#_M1011_d 2.08474e-19 $X=1.87 $Y=0.76 $X2=0 $Y2=0
cc_220 Y N_A_27_47#_M1011_d 0.00284805f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_221 Y N_A_27_47#_M1011_d 6.30938e-19 $X=2.075 $Y=0.85 $X2=0 $Y2=0
cc_222 N_Y_c_249_n N_A_27_47#_c_452_n 0.00270783f $X=0.935 $Y=1.57 $X2=0 $Y2=0
cc_223 N_Y_c_245_n N_A_27_47#_c_452_n 0.00232109f $X=1.1 $Y=1.57 $X2=0 $Y2=0
cc_224 N_Y_c_244_n N_A_27_47#_c_450_n 0.00196792f $X=0.345 $Y=1.57 $X2=0 $Y2=0
cc_225 N_Y_M1010_s N_A_27_47#_c_451_n 0.00305418f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_226 N_Y_c_264_n N_A_27_47#_c_451_n 0.0236342f $X=1.87 $Y=0.76 $X2=0 $Y2=0
cc_227 Y N_A_27_47#_c_451_n 0.0188217f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_228 Y N_VGND_c_487_n 0.00103015f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_229 N_Y_c_242_n N_VGND_c_487_n 0.00226279f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_230 N_Y_M1010_s N_VGND_c_492_n 0.00216833f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_231 N_Y_M1006_s N_VGND_c_492_n 0.00216833f $X=2.745 $Y=0.235 $X2=0 $Y2=0
cc_232 Y N_VGND_c_492_n 0.00216666f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_233 N_Y_c_242_n N_VGND_c_492_n 0.00499764f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_234 N_Y_c_242_n N_A_467_47#_M1006_d 0.00676128f $X=2.88 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_235 N_Y_M1006_s N_A_467_47#_c_548_n 0.00305418f $X=2.745 $Y=0.235 $X2=0 $Y2=0
cc_236 N_Y_c_242_n N_A_467_47#_c_548_n 0.0405898f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_237 N_A_109_297#_c_334_n N_VPWR_M1004_s 0.00324353f $X=3.135 $Y=1.57
+ $X2=-0.19 $Y2=1.305
cc_238 N_A_109_297#_c_322_n N_VPWR_M1009_s 0.00324353f $X=3.975 $Y=1.57 $X2=0
+ $Y2=0
cc_239 N_A_109_297#_c_334_n N_VPWR_c_393_n 0.0126919f $X=3.135 $Y=1.57 $X2=0
+ $Y2=0
cc_240 N_A_109_297#_c_322_n N_VPWR_c_394_n 0.0126919f $X=3.975 $Y=1.57 $X2=0
+ $Y2=0
cc_241 N_A_109_297#_c_326_n N_VPWR_c_395_n 0.0358391f $X=1.435 $Y=2.38 $X2=0
+ $Y2=0
cc_242 N_A_109_297#_c_327_n N_VPWR_c_395_n 0.0151638f $X=0.765 $Y=2.38 $X2=0
+ $Y2=0
cc_243 N_A_109_297#_c_320_n N_VPWR_c_395_n 0.0457462f $X=2.375 $Y=2.38 $X2=0
+ $Y2=0
cc_244 N_A_109_297#_c_331_n N_VPWR_c_395_n 0.0154974f $X=2.5 $Y=2.295 $X2=0
+ $Y2=0
cc_245 N_A_109_297#_c_376_p N_VPWR_c_395_n 0.0114181f $X=1.52 $Y=2.38 $X2=0
+ $Y2=0
cc_246 N_A_109_297#_c_341_n N_VPWR_c_397_n 0.0189039f $X=3.3 $Y=1.66 $X2=0 $Y2=0
cc_247 N_A_109_297#_c_323_n N_VPWR_c_399_n 0.0210382f $X=4.14 $Y=1.66 $X2=0
+ $Y2=0
cc_248 N_A_109_297#_M1001_s N_VPWR_c_392_n 0.00215206f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_249 N_A_109_297#_M1000_d N_VPWR_c_392_n 0.0021521f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_250 N_A_109_297#_M1004_d N_VPWR_c_392_n 0.00209323f $X=2.335 $Y=1.485 $X2=0
+ $Y2=0
cc_251 N_A_109_297#_M1008_d N_VPWR_c_392_n 0.00215201f $X=3.165 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_109_297#_M1013_d N_VPWR_c_392_n 0.00209319f $X=4.005 $Y=1.485 $X2=0
+ $Y2=0
cc_253 N_A_109_297#_c_326_n N_VPWR_c_392_n 0.0234424f $X=1.435 $Y=2.38 $X2=0
+ $Y2=0
cc_254 N_A_109_297#_c_327_n N_VPWR_c_392_n 0.0093986f $X=0.765 $Y=2.38 $X2=0
+ $Y2=0
cc_255 N_A_109_297#_c_320_n N_VPWR_c_392_n 0.027919f $X=2.375 $Y=2.38 $X2=0
+ $Y2=0
cc_256 N_A_109_297#_c_331_n N_VPWR_c_392_n 0.00941829f $X=2.5 $Y=2.295 $X2=0
+ $Y2=0
cc_257 N_A_109_297#_c_341_n N_VPWR_c_392_n 0.0122217f $X=3.3 $Y=1.66 $X2=0 $Y2=0
cc_258 N_A_109_297#_c_323_n N_VPWR_c_392_n 0.0124268f $X=4.14 $Y=1.66 $X2=0
+ $Y2=0
cc_259 N_A_109_297#_c_376_p N_VPWR_c_392_n 0.00653671f $X=1.52 $Y=2.38 $X2=0
+ $Y2=0
cc_260 N_A_109_297#_c_324_n N_A_467_47#_c_561_n 0.00514931f $X=3.3 $Y=1.57 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_452_n N_VGND_M1005_s 0.00323654f $X=1.015 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_262 N_A_27_47#_c_452_n N_VGND_c_487_n 0.00219298f $X=1.015 $Y=0.765 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_473_p N_VGND_c_487_n 0.0113602f $X=1.185 $Y=0.38 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_451_n N_VGND_c_487_n 0.0527078f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_449_n N_VGND_c_490_n 0.0171173f $X=0.22 $Y=0.68 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_452_n N_VGND_c_490_n 0.00219298f $X=1.015 $Y=0.765 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_M1005_d N_VGND_c_492_n 0.00230841f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1015_d N_VGND_c_492_n 0.00238334f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1011_d N_VGND_c_492_n 0.00209344f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_449_n N_VGND_c_492_n 0.00951769f $X=0.22 $Y=0.68 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_452_n N_VGND_c_492_n 0.00946308f $X=1.015 $Y=0.765 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_473_p N_VGND_c_492_n 0.00652422f $X=1.185 $Y=0.38 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_451_n N_VGND_c_492_n 0.0331126f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_452_n N_VGND_c_493_n 0.0161795f $X=1.015 $Y=0.765 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_451_n N_A_467_47#_c_548_n 0.0214676f $X=1.94 $Y=0.42 $X2=0
+ $Y2=0
cc_276 N_VGND_c_492_n N_A_467_47#_M1006_d 0.00209344f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_277 N_VGND_c_492_n N_A_467_47#_M1007_d 0.00238334f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_492_n N_A_467_47#_M1003_d 0.00230841f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_487_n N_A_467_47#_c_548_n 0.0640679f $X=3.555 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_492_n N_A_467_47#_c_548_n 0.0396369f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_M1002_s N_A_467_47#_c_549_n 0.00323654f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_282 N_VGND_c_486_n N_A_467_47#_c_549_n 0.0161795f $X=3.72 $Y=0.4 $X2=0 $Y2=0
cc_283 N_VGND_c_487_n N_A_467_47#_c_549_n 0.00219298f $X=3.555 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_491_n N_A_467_47#_c_549_n 0.00219298f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_492_n N_A_467_47#_c_549_n 0.00946308f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_491_n N_A_467_47#_c_550_n 0.0220856f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_492_n N_A_467_47#_c_550_n 0.0122041f $X=4.37 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o2111a_1.spice.pex
* Created: Thu Aug 27 14:33:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2111A_1%A_79_21# 1 2 3 12 15 18 19 20 23 27 29 35
+ 36 38 40 42
c68 36 0 1.18508e-19 $X=0.78 $Y=1.115
r69 35 43 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.16
+ $X2=0.57 $Y2=1.325
r70 35 42 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.16
+ $X2=0.57 $Y2=0.995
r71 34 36 7.22648 $w=2.87e-07 $l=1.7e-07 $layer=LI1_cond $X=0.61 $Y=1.115
+ $X2=0.78 $Y2=1.115
r72 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.16 $X2=0.61 $Y2=1.16
r73 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r74 29 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.93 $Y=1.58
+ $X2=3.055 $Y2=1.58
r75 29 30 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=2.93 $Y=1.58
+ $X2=1.835 $Y2=1.58
r76 25 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r77 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.96
r78 21 36 17.6411 $w=2.87e-07 $l=5.74391e-07 $layer=LI1_cond $X=1.195 $Y=0.735
+ $X2=0.78 $Y2=1.115
r79 21 23 12.0329 $w=3.38e-07 $l=3.55e-07 $layer=LI1_cond $X=1.195 $Y=0.735
+ $X2=1.195 $Y2=0.38
r80 19 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r81 19 20 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.865 $Y2=1.58
r82 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.78 $Y=1.495
+ $X2=0.865 $Y2=1.58
r83 17 36 3.80104 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.78 $Y=1.325
+ $X2=0.78 $Y2=1.115
r84 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.78 $Y=1.325
+ $X2=0.78 $Y2=1.495
r85 15 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r86 12 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
r87 3 40 300 $w=1.7e-07 $l=3.67219e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=3.095 $Y2=1.66
r88 2 27 300 $w=1.7e-07 $l=5.70417e-07 $layer=licon1_PDIFF $count=2 $X=1.46
+ $Y=1.485 $X2=1.67 $Y2=1.96
r89 1 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%D1 3 7 9 10 11 16 28
c40 3 0 1.41804e-19 $X=1.385 $Y=1.985
r41 20 28 1.75975 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.64 $Y=1.075
+ $X2=1.64 $Y2=1.2
r42 16 19 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.43 $Y2=1.295
r43 16 18 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.43 $Y2=1.025
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.16 $X2=1.43 $Y2=1.16
r45 11 20 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=1.64 $Y=0.85
+ $X2=1.64 $Y2=1.075
r46 10 11 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.64 $Y=0.51
+ $X2=1.64 $Y2=0.85
r47 9 28 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=1.64
+ $Y2=1.2
r48 9 17 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=1.43
+ $Y2=1.2
r49 7 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.455 $Y=0.56
+ $X2=1.455 $Y2=1.025
r50 3 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.385 $Y=1.985
+ $X2=1.385 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%C1 3 7 9 10 11 16
c37 9 0 1.06898e-19 $X=2.07 $Y=0.51
c38 7 0 9.34721e-20 $X=1.97 $Y=1.985
r39 16 19 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.03 $Y=1.16
+ $X2=2.03 $Y2=1.295
r40 16 18 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.03 $Y=1.16
+ $X2=2.03 $Y2=1.025
r41 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.16 $X2=2.03 $Y2=1.16
r42 10 11 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.06 $Y=0.85
+ $X2=2.06 $Y2=1.16
r43 9 10 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.06 $Y=0.51 $X2=2.06
+ $Y2=0.85
r44 7 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.97 $Y=1.985
+ $X2=1.97 $Y2=1.295
r45 3 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.97 $Y=0.56
+ $X2=1.97 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%B1 3 7 9 10 11 19 20
c41 19 0 1.18418e-19 $X=2.62 $Y=1.16
c42 7 0 8.36011e-20 $X=2.73 $Y=1.985
r43 19 27 7.36562 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=1.16
+ $X2=2.575 $Y2=0.995
r44 18 20 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=2.62 $Y=1.16
+ $X2=2.73 $Y2=1.16
r45 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.16 $X2=2.62 $Y2=1.16
r46 15 18 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.485 $Y=1.16
+ $X2=2.62 $Y2=1.16
r47 11 19 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=2.575 $Y=1.19
+ $X2=2.575 $Y2=1.16
r48 10 27 6.82058 $w=2.43e-07 $l=1.45e-07 $layer=LI1_cond $X=2.567 $Y=0.85
+ $X2=2.567 $Y2=0.995
r49 9 10 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=2.567 $Y=0.51
+ $X2=2.567 $Y2=0.85
r50 5 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.73 $Y=1.295
+ $X2=2.73 $Y2=1.16
r51 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.73 $Y=1.295 $X2=2.73
+ $Y2=1.985
r52 1 15 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.485 $Y=1.025
+ $X2=2.485 $Y2=1.16
r53 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.485 $Y=1.025
+ $X2=2.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%A2 3 7 9 12 14 15 16 17 25
c44 25 0 1.11775e-19 $X=3.442 $Y=1.325
c45 7 0 2.4946e-20 $X=3.305 $Y=1.985
r46 16 17 20.3833 $w=1.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.442 $Y=1.87
+ $X2=3.442 $Y2=2.21
r47 15 16 20.3833 $w=1.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.442 $Y=1.53
+ $X2=3.442 $Y2=1.87
r48 15 25 12.2899 $w=1.83e-07 $l=2.05e-07 $layer=LI1_cond $X=3.442 $Y=1.53
+ $X2=3.442 $Y2=1.325
r49 14 25 4.04167 $w=1.85e-07 $l=1.25e-07 $layer=LI1_cond $X=3.442 $Y=1.2
+ $X2=3.442 $Y2=1.325
r50 12 24 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.215 $Y=1.16
+ $X2=3.215 $Y2=1.295
r51 12 23 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.215 $Y=1.16
+ $X2=3.215 $Y2=1.025
r52 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.16 $X2=3.215 $Y2=1.16
r53 9 14 2.97467 $w=2.5e-07 $l=9.2e-08 $layer=LI1_cond $X=3.35 $Y=1.2 $X2=3.442
+ $Y2=1.2
r54 9 11 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.35 $Y=1.2
+ $X2=3.215 $Y2=1.2
r55 7 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.305 $Y=1.985
+ $X2=3.305 $Y2=1.295
r56 3 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.245 $Y=0.56
+ $X2=3.245 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%A1 3 7 9 10 16
r25 13 16 42.4045 $w=2.9e-07 $l=2.05e-07 $layer=POLY_cond $X=3.665 $Y=1.16
+ $X2=3.87 $Y2=1.16
r26 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.87 $Y=1.16 $X2=3.87
+ $Y2=1.53
r27 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=1.16 $X2=3.87 $Y2=1.16
r28 5 13 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.665 $Y=1.305
+ $X2=3.665 $Y2=1.16
r29 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.665 $Y=1.305
+ $X2=3.665 $Y2=1.985
r30 1 13 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.665 $Y=1.015
+ $X2=3.665 $Y2=1.16
r31 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.665 $Y=1.015
+ $X2=3.665 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%X 1 2 7 8 9 10 11 12 20
r11 12 33 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.225 $Y=2.21
+ $X2=0.225 $Y2=1.96
r12 11 33 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.96
r13 10 11 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=1.53
+ $X2=0.225 $Y2=1.87
r14 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=1.19
+ $X2=0.225 $Y2=1.53
r15 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=0.85
+ $X2=0.225 $Y2=1.19
r16 7 8 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=0.51
+ $X2=0.225 $Y2=0.85
r17 7 20 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=0.225 $Y=0.51 $X2=0.225
+ $Y2=0.42
r18 2 33 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r19 1 20 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%VPWR 1 2 3 10 14 16 18 20 22 27 33 40 46
r57 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 41 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 40 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 37 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 33 36 10.6318 $w=8.08e-07 $l=7.2e-07 $layer=LI1_cond $X=0.93 $Y=2 $X2=0.93
+ $Y2=2.72
r64 31 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 31 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r66 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 28 40 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=2.76 $Y=2.72 $X2=2.39
+ $Y2=2.72
r68 28 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.76 $Y=2.72 $X2=3.45
+ $Y2=2.72
r69 27 45 4.75502 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.935 $Y2=2.72
r70 27 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r71 22 36 10.2922 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.93 $Y2=2.72
r72 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 20 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 20 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r75 16 45 2.96899 $w=3.25e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.935 $Y2=2.72
r76 16 18 22.517 $w=3.23e-07 $l=6.35e-07 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.892 $Y2=2
r77 12 40 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=2.635
+ $X2=2.39 $Y2=2.72
r78 12 14 10.2636 $w=7.38e-07 $l=6.35e-07 $layer=LI1_cond $X=2.39 $Y=2.635
+ $X2=2.39 $Y2=2
r79 11 36 10.2922 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=0.93 $Y2=2.72
r80 10 40 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=2.02 $Y=2.72 $X2=2.39
+ $Y2=2.72
r81 10 11 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.02 $Y=2.72
+ $X2=1.335 $Y2=2.72
r82 3 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.74
+ $Y=1.485 $X2=3.875 $Y2=2
r83 2 14 150 $w=1.7e-07 $l=7.14038e-07 $layer=licon1_PDIFF $count=4 $X=2.045
+ $Y=1.485 $X2=2.52 $Y2=2
r84 1 33 150 $w=1.7e-07 $l=8.44097e-07 $layer=licon1_PDIFF $count=4 $X=0.545
+ $Y=1.485 $X2=1.17 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r55 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r58 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r59 30 39 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.475
+ $Y2=0
r60 30 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.91
+ $Y2=0
r61 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r62 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r63 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r64 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r65 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r66 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 23 36 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.69
+ $Y2=0
r68 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r69 22 39 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.475
+ $Y2=0
r70 22 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=2.99
+ $Y2=0
r71 17 36 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.69
+ $Y2=0
r72 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.23
+ $Y2=0
r73 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r74 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 11 39 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.085
+ $X2=3.475 $Y2=0
r76 11 13 11.3257 $w=2.88e-07 $l=2.85e-07 $layer=LI1_cond $X=3.475 $Y=0.085
+ $X2=3.475 $Y2=0.37
r77 7 36 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r78 7 9 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r79 2 13 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.455 $Y2=0.37
r80 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_1%A_512_47# 1 2 9 11 12 15
r29 13 15 12.3942 $w=2.63e-07 $l=2.85e-07 $layer=LI1_cond $X=3.922 $Y=0.705
+ $X2=3.922 $Y2=0.42
r30 11 13 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.79 $Y=0.79
+ $X2=3.922 $Y2=0.705
r31 11 12 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.79 $Y=0.79
+ $X2=3.16 $Y2=0.79
r32 7 12 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.015 $Y=0.705
+ $X2=3.16 $Y2=0.79
r33 7 9 11.3257 $w=2.88e-07 $l=2.85e-07 $layer=LI1_cond $X=3.015 $Y=0.705
+ $X2=3.015 $Y2=0.42
r34 2 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.74
+ $Y=0.235 $X2=3.875 $Y2=0.42
r35 1 9 91 $w=1.7e-07 $l=5.59911e-07 $layer=licon1_NDIFF $count=2 $X=2.56
+ $Y=0.235 $X2=3.035 $Y2=0.42
.ends


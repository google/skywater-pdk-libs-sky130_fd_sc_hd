* File: sky130_fd_sc_hd__or2_2.pex.spice
* Created: Thu Aug 27 14:42:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR2_2%B 3 7 9 10 18
r27 17 18 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.53
+ $Y2=1.16
r28 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r29 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r30 9 10 17.6317 $w=1.93e-07 $l=3.1e-07 $layer=LI1_cond $X=0.247 $Y=0.85
+ $X2=0.247 $Y2=1.16
r31 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.325
+ $X2=0.53 $Y2=1.16
r32 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.53 $Y=1.325 $X2=0.53
+ $Y2=1.695
r33 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r34 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_2%A 3 7 9 10 14
r35 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=1.325
r36 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=0.995
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r38 10 15 0.843251 $w=4.08e-07 $l=3e-08 $layer=LI1_cond $X=1.07 $Y=1.19 $X2=1.07
+ $Y2=1.16
r39 9 15 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=1.07 $Y=0.85 $X2=1.07
+ $Y2=1.16
r40 7 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.89 $Y=1.695
+ $X2=0.89 $Y2=1.325
r41 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_2%A_39_297# 1 2 7 9 12 14 16 19 22 23 24 27 34
+ 40
c66 27 0 7.42925e-20 $X=1.53 $Y=1.16
c67 24 0 1.40438e-19 $X=0.695 $Y=1.58
c68 22 0 1.02064e-19 $X=0.605 $Y=1.495
r69 34 36 8.20519 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.66 $Y=0.43
+ $X2=0.66 $Y2=0.595
r70 28 40 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.53 $Y=1.16
+ $X2=1.815 $Y2=1.16
r71 28 37 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.53 $Y=1.16
+ $X2=1.395 $Y2=1.16
r72 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.53
+ $Y=1.16 $X2=1.53 $Y2=1.16
r73 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.53 $Y=1.495
+ $X2=1.53 $Y2=1.16
r74 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.445 $Y=1.58
+ $X2=1.53 $Y2=1.495
r75 23 24 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.445 $Y=1.58
+ $X2=0.695 $Y2=1.58
r76 22 24 5.83001 $w=2.86e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.695 $Y2=1.58
r77 22 31 12.1573 $w=2.86e-07 $l=3.60895e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.32 $Y2=1.667
r78 22 36 55.4545 $w=1.78e-07 $l=9e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.605 $Y2=0.595
r79 17 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.16
r80 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.985
r81 14 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r82 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=0.56
r83 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.16
r84 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.985
r85 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=1.16
r86 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=0.56
r87 2 31 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.485 $X2=0.32 $Y2=1.66
r88 1 34 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_2%VPWR 1 2 9 11 13 15 17 22 28 32
c29 9 0 1.40438e-19 $X=1.185 $Y=2.01
r30 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r31 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r32 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r33 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r35 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.72
+ $X2=1.185 $Y2=2.72
r36 23 25 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.27 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 22 31 3.40825 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.94 $Y=2.72 $X2=2.12
+ $Y2=2.72
r38 22 25 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=1.61 $Y2=2.72
r39 17 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.72 $X2=1.185
+ $Y2=2.72
r40 17 19 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.1 $Y=2.72 $X2=0.23
+ $Y2=2.72
r41 15 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 15 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r43 11 31 3.40825 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.025 $Y=2.635
+ $X2=2.12 $Y2=2.72
r44 11 13 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.025 $Y=2.635
+ $X2=2.025 $Y2=2.34
r45 7 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=2.72
r46 7 9 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=2.01
r47 2 13 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.025 $Y2=2.34
r48 1 9 300 $w=1.7e-07 $l=6.254e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.185 $Y2=2.01
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_2%X 1 2 10 13 19
c32 2 0 7.42925e-20 $X=1.47 $Y=1.485
r33 16 19 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2 $Y=1.92 $X2=1.605
+ $Y2=1.92
r34 13 16 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.075 $Y=1.92 $X2=2
+ $Y2=1.92
r35 13 16 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2 $Y=1.81 $X2=2
+ $Y2=1.835
r36 12 13 26.399 $w=4.28e-07 $l=9.85e-07 $layer=LI1_cond $X=2 $Y=0.825 $X2=2
+ $Y2=1.81
r37 10 12 20.4195 $w=2.36e-07 $l=3.95e-07 $layer=LI1_cond $X=1.605 $Y=0.655
+ $X2=2 $Y2=0.655
r38 2 19 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=1.485 $X2=1.605 $Y2=2
r39 1 10 182 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_NDIFF $count=1 $X=1.47
+ $Y=0.235 $X2=1.605 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_2%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r40 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r41 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r42 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r43 33 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r44 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r45 30 38 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.192
+ $Y2=0
r46 30 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.61
+ $Y2=0
r47 29 41 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.08
+ $Y2=0
r48 29 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.61
+ $Y2=0
r49 28 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r50 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 25 35 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r52 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r53 24 38 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.192
+ $Y2=0
r54 24 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r55 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r56 22 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r57 18 41 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.08 $Y2=0
r58 18 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.39
r59 14 38 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.192 $Y=0.085
+ $X2=1.192 $Y2=0
r60 14 16 12.622 $w=3.13e-07 $l=3.45e-07 $layer=LI1_cond $X=1.192 $Y=0.085
+ $X2=1.192 $Y2=0.43
r61 10 35 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r62 10 12 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.43
r63 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.235 $X2=2.025 $Y2=0.39
r64 2 16 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.18 $Y2=0.43
r65 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends


* File: sky130_fd_sc_hd__nor4bb_2.spice.pex
* Created: Thu Aug 27 14:33:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%D_N 3 5 7 8 9 13 14
c34 14 0 3.191e-20 $X=0.51 $Y=1.16
c35 13 0 5.30499e-20 $X=0.51 $Y=1.16
r36 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r38 8 9 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.602 $Y=1.19
+ $X2=0.602 $Y2=1.53
r39 8 14 0.973895 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=0.602 $Y=1.19
+ $X2=0.602 $Y2=1.16
r40 5 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=1.16
r41 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.51 $Y=0.995 $X2=0.51
+ $Y2=0.675
r42 3 15 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.47 $Y=2.26
+ $X2=0.47 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%C_N 3 6 8 11 13 19
r36 11 14 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.027 $Y=1.16
+ $X2=1.027 $Y2=1.325
r37 11 13 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.027 $Y=1.16
+ $X2=1.027 $Y2=0.995
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r39 8 19 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.155
+ $Y2=1.16
r40 8 12 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.035 $Y2=1.16
r41 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.955 $Y=1.695
+ $X2=0.955 $Y2=1.325
r42 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.93 $Y=0.675
+ $X2=0.93 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%A_201_93# 1 2 7 9 12 14 16 19 21 26 28 31
+ 35 37 41
c85 31 0 1.23788e-19 $X=2.225 $Y=1.16
c86 26 0 3.191e-20 $X=1.49 $Y=1.075
r87 35 36 17.3577 $w=2.46e-07 $l=3.5e-07 $layer=LI1_cond $X=1.14 $Y=0.655
+ $X2=1.49 $Y2=0.655
r88 32 41 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.435 $Y2=1.16
r89 32 38 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.015 $Y2=1.16
r90 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.225
+ $Y=1.16 $X2=2.225 $Y2=1.16
r91 29 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=1.16
+ $X2=1.49 $Y2=1.16
r92 29 31 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.575 $Y=1.16
+ $X2=2.225 $Y2=1.16
r93 27 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.245
+ $X2=1.49 $Y2=1.16
r94 27 28 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.49 $Y=1.245
+ $X2=1.49 $Y2=1.525
r95 26 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.075
+ $X2=1.49 $Y2=1.16
r96 25 36 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.49 $Y2=0.655
r97 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.49 $Y2=1.075
r98 21 28 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.405 $Y=1.62
+ $X2=1.49 $Y2=1.525
r99 21 23 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=1.405 $Y=1.62
+ $X2=1.165 $Y2=1.62
r100 17 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.325
+ $X2=2.435 $Y2=1.16
r101 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.435 $Y=1.325
+ $X2=2.435 $Y2=1.985
r102 14 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.435 $Y2=1.16
r103 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.435 $Y2=0.56
r104 10 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.325
+ $X2=2.015 $Y2=1.16
r105 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.015 $Y=1.325
+ $X2=2.015 $Y2=1.985
r106 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=1.16
r107 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
r108 2 23 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.63
r109 1 35 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.465 $X2=1.14 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%A_27_410# 1 2 7 9 12 14 16 19 22 25 27 30
+ 31 32 34 35 37 43 45 49
c106 49 0 1.23788e-19 $X=3.275 $Y=1.16
r107 40 43 3.99514 $w=3.73e-07 $l=1.3e-07 $layer=LI1_cond $X=0.17 $Y=0.637
+ $X2=0.3 $Y2=0.637
r108 38 49 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.24 $Y=1.16
+ $X2=3.275 $Y2=1.16
r109 38 46 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=3.24 $Y=1.16
+ $X2=2.855 $Y2=1.16
r110 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.24
+ $Y=1.16 $X2=3.24 $Y2=1.16
r111 35 37 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=2.73 $Y=1.175
+ $X2=3.24 $Y2=1.175
r112 33 35 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.645 $Y=1.275
+ $X2=2.73 $Y2=1.175
r113 33 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.645 $Y=1.275
+ $X2=2.645 $Y2=1.415
r114 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=1.5
+ $X2=2.645 $Y2=1.415
r115 31 32 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.56 $Y=1.5
+ $X2=1.915 $Y2=1.5
r116 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.83 $Y=1.585
+ $X2=1.915 $Y2=1.5
r117 29 30 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.83 $Y=1.585
+ $X2=1.83 $Y2=1.885
r118 28 45 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.97
+ $X2=0.215 $Y2=1.97
r119 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=1.97
+ $X2=1.83 $Y2=1.885
r120 27 28 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.745 $Y=1.97
+ $X2=0.345 $Y2=1.97
r121 23 45 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.055
+ $X2=0.215 $Y2=1.97
r122 23 25 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=0.215 $Y=2.055
+ $X2=0.215 $Y2=2.29
r123 22 45 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.17 $Y=1.885
+ $X2=0.215 $Y2=1.97
r124 21 40 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.637
r125 21 22 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.885
r126 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.325
+ $X2=3.275 $Y2=1.16
r127 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.275 $Y=1.325
+ $X2=3.275 $Y2=1.985
r128 14 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=0.995
+ $X2=3.275 $Y2=1.16
r129 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.275 $Y=0.995
+ $X2=3.275 $Y2=0.56
r130 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.325
+ $X2=2.855 $Y2=1.16
r131 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.855 $Y=1.325
+ $X2=2.855 $Y2=1.985
r132 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=0.995
+ $X2=2.855 $Y2=1.16
r133 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.855 $Y=0.995
+ $X2=2.855 $Y2=0.56
r134 2 25 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r135 1 43 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.465 $X2=0.3 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%B 1 3 6 8 10 13 15 21 22
c47 22 0 1.40616e-19 $X=4.655 $Y=1.16
r48 20 22 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.655 $Y2=1.16
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r50 17 20 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.235 $Y=1.16
+ $X2=4.46 $Y2=1.16
r51 15 21 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=4.37 $Y=1.175 $X2=4.46
+ $Y2=1.175
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.325
+ $X2=4.655 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.655 $Y=1.325
+ $X2=4.655 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=0.995
+ $X2=4.655 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.655 $Y=0.995
+ $X2=4.655 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.325
+ $X2=4.235 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.235 $Y=1.325
+ $X2=4.235 $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=0.995
+ $X2=4.235 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.235 $Y=0.995
+ $X2=4.235 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%A 1 3 6 8 10 13 15 22
c38 15 0 1.40616e-19 $X=5.29 $Y=1.19
c39 6 0 6.26685e-20 $X=5.075 $Y=1.985
r40 20 22 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=5.295 $Y=1.16
+ $X2=5.495 $Y2=1.16
r41 17 20 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.075 $Y=1.16
+ $X2=5.295 $Y2=1.16
r42 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.295
+ $Y=1.16 $X2=5.295 $Y2=1.16
r43 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.495 $Y=1.325
+ $X2=5.495 $Y2=1.16
r44 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.495 $Y=1.325
+ $X2=5.495 $Y2=1.985
r45 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.495 $Y=0.995
+ $X2=5.495 $Y2=1.16
r46 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.495 $Y=0.995
+ $X2=5.495 $Y2=0.56
r47 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.075 $Y=1.325
+ $X2=5.075 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.075 $Y=1.325
+ $X2=5.075 $Y2=1.985
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.075 $Y=0.995
+ $X2=5.075 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.075 $Y=0.995
+ $X2=5.075 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r60 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r62 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r63 30 31 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r64 28 31 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r65 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 27 30 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r67 27 28 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r69 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r71 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 16 30 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.16 $Y=2.72
+ $X2=4.83 $Y2=2.72
r75 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.16 $Y=2.72
+ $X2=5.265 $Y2=2.72
r76 15 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.37 $Y=2.72
+ $X2=5.75 $Y2=2.72
r77 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.37 $Y=2.72
+ $X2=5.265 $Y2=2.72
r78 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.265 $Y=2.635
+ $X2=5.265 $Y2=2.72
r79 11 13 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=5.265 $Y=2.635
+ $X2=5.265 $Y2=1.96
r80 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r81 7 9 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.325
r82 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.15
+ $Y=1.485 $X2=5.285 $Y2=1.96
r83 1 9 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.05 $X2=0.68 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%A_336_297# 1 2 3 12 16 21 22
r31 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.97 $Y=2.38
+ $X2=2.48 $Y2=2.38
r32 19 21 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=2.345
+ $X2=1.97 $Y2=2.345
r33 14 16 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=2.645 $Y=2.34
+ $X2=3.485 $Y2=2.34
r34 12 22 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.605 $Y=2.34
+ $X2=2.48 $Y2=2.34
r35 12 14 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=2.605 $Y=2.34
+ $X2=2.645 $Y2=2.34
r36 3 16 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=1.485 $X2=3.485 $Y2=2.3
r37 2 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=1.485 $X2=2.645 $Y2=2.3
r38 1 19 600 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.485 $X2=1.805 $Y2=2.31
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%A_418_297# 1 2 7 9 11 14
c35 11 0 6.26685e-20 $X=4.445 $Y=1.62
r36 9 18 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=1.875
+ $X2=4.465 $Y2=1.96
r37 9 11 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=4.465 $Y=1.875
+ $X2=4.465 $Y2=1.62
r38 8 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=1.96
+ $X2=2.225 $Y2=1.96
r39 7 18 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.32 $Y=1.96
+ $X2=4.465 $Y2=1.96
r40 7 8 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=4.32 $Y=1.96 $X2=2.31
+ $Y2=1.96
r41 2 18 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.485 $X2=4.445 $Y2=1.96
r42 2 11 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.485 $X2=4.445 $Y2=1.62
r43 1 14 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.485 $X2=2.225 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%Y 1 2 3 4 5 18 20 21 24 26 28 32 34 38 40
+ 42 43 44 45 49
r114 45 49 4.52065 $w=2.6e-07 $l=2.1e-07 $layer=LI1_cond $X=3.785 $Y=1.575
+ $X2=3.575 $Y2=1.575
r115 44 49 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=3.45 $Y=1.575
+ $X2=3.575 $Y2=1.575
r116 44 51 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.45 $Y=1.575
+ $X2=3.065 $Y2=1.575
r117 41 45 11.9572 $w=5.88e-07 $l=5.4e-07 $layer=LI1_cond $X=3.785 $Y=0.905
+ $X2=3.785 $Y2=1.445
r118 41 42 1.44414 $w=4.2e-07 $l=9e-08 $layer=LI1_cond $X=3.785 $Y=0.905
+ $X2=3.785 $Y2=0.815
r119 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.285 $Y=0.725
+ $X2=5.285 $Y2=0.39
r120 35 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.61 $Y=0.815
+ $X2=4.445 $Y2=0.815
r121 34 36 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.12 $Y=0.815
+ $X2=5.285 $Y2=0.725
r122 34 35 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.12 $Y=0.815
+ $X2=4.61 $Y2=0.815
r123 30 43 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.445 $Y=0.725
+ $X2=4.445 $Y2=0.815
r124 30 32 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.445 $Y=0.725
+ $X2=4.445 $Y2=0.39
r125 29 42 9.75736 $w=1.8e-07 $l=2.1e-07 $layer=LI1_cond $X=3.995 $Y=0.815
+ $X2=3.785 $Y2=0.815
r126 28 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.28 $Y=0.815
+ $X2=4.445 $Y2=0.815
r127 28 29 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=4.28 $Y=0.815
+ $X2=3.995 $Y2=0.815
r128 27 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=0.815
+ $X2=3.065 $Y2=0.815
r129 26 42 9.75736 $w=1.8e-07 $l=2.1e-07 $layer=LI1_cond $X=3.575 $Y=0.815
+ $X2=3.785 $Y2=0.815
r130 26 27 21.2576 $w=1.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.575 $Y=0.815
+ $X2=3.23 $Y2=0.815
r131 22 40 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.065 $Y=0.725
+ $X2=3.065 $Y2=0.815
r132 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.065 $Y=0.725
+ $X2=3.065 $Y2=0.39
r133 20 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=0.815
+ $X2=3.065 $Y2=0.815
r134 20 21 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.9 $Y=0.815
+ $X2=2.39 $Y2=0.815
r135 16 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.39 $Y2=0.815
r136 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.225 $Y=0.725
+ $X2=2.225 $Y2=0.39
r137 5 51 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.485 $X2=3.065 $Y2=1.62
r138 4 38 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.15
+ $Y=0.235 $X2=5.285 $Y2=0.39
r139 3 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.235 $X2=4.445 $Y2=0.39
r140 2 24 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.93
+ $Y=0.235 $X2=3.065 $Y2=0.39
r141 1 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.09
+ $Y=0.235 $X2=2.225 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%A_776_297# 1 2 3 10 14 15 16 20
r34 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.705 $Y=1.63
+ $X2=5.705 $Y2=2.31
r35 18 20 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=5.705 $Y=1.625
+ $X2=5.705 $Y2=1.63
r36 17 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.99 $Y=1.54
+ $X2=4.885 $Y2=1.54
r37 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.54 $Y=1.54
+ $X2=5.705 $Y2=1.625
r38 16 17 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.54 $Y=1.54
+ $X2=4.99 $Y2=1.54
r39 15 27 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=2.215
+ $X2=4.885 $Y2=2.34
r40 14 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=1.625
+ $X2=4.885 $Y2=1.54
r41 14 15 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.885 $Y=1.625
+ $X2=4.885 $Y2=2.215
r42 10 27 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.78 $Y=2.34
+ $X2=4.885 $Y2=2.34
r43 10 12 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=4.78 $Y=2.34
+ $X2=4.025 $Y2=2.34
r44 3 22 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.485 $X2=5.705 $Y2=2.31
r45 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.485 $X2=5.705 $Y2=1.63
r46 2 27 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.73
+ $Y=1.485 $X2=4.865 $Y2=2.3
r47 2 25 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.73
+ $Y=1.485 $X2=4.865 $Y2=1.62
r48 1 12 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.485 $X2=4.025 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_2%VGND 1 2 3 4 5 6 7 26 28 32 36 40 44 46 48
+ 50 51 52 58 64 67 72 80 82 86
c94 26 0 5.30499e-20 $X=0.72 $Y=0.66
r95 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r96 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r97 79 80 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=0.235
+ $X2=4.11 $Y2=0.235
r98 77 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r99 76 79 2.1492 $w=6.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.91 $Y=0.235
+ $X2=4.025 $Y2=0.235
r100 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r101 74 76 7.94271 $w=6.38e-07 $l=4.25e-07 $layer=LI1_cond $X=3.485 $Y=0.235
+ $X2=3.91 $Y2=0.235
r102 71 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r103 70 74 0.654105 $w=6.38e-07 $l=3.5e-08 $layer=LI1_cond $X=3.45 $Y=0.235
+ $X2=3.485 $Y2=0.235
r104 70 72 8.26766 $w=6.38e-07 $l=5e-08 $layer=LI1_cond $X=3.45 $Y=0.235 $X2=3.4
+ $Y2=0.235
r105 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r106 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r107 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r108 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r109 62 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r110 62 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r111 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r112 59 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=0 $X2=4.865
+ $Y2=0
r113 59 61 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=0 $X2=5.29
+ $Y2=0
r114 58 85 4.27912 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.62 $Y=0 $X2=5.8
+ $Y2=0
r115 58 61 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.62 $Y=0 $X2=5.29
+ $Y2=0
r116 57 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r117 57 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r118 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r119 54 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.725
+ $Y2=0
r120 54 56 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.53
+ $Y2=0
r121 52 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r122 50 56 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.53
+ $Y2=0
r123 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.645
+ $Y2=0
r124 46 85 3.04293 $w=2.75e-07 $l=1.04307e-07 $layer=LI1_cond $X=5.757 $Y=0.085
+ $X2=5.8 $Y2=0
r125 46 48 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=5.757 $Y=0.085
+ $X2=5.757 $Y2=0.39
r126 42 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=0.085
+ $X2=4.865 $Y2=0
r127 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.865 $Y=0.085
+ $X2=4.865 $Y2=0.39
r128 40 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=0 $X2=4.865
+ $Y2=0
r129 40 80 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.78 $Y=0 $X2=4.11
+ $Y2=0
r130 39 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.645
+ $Y2=0
r131 39 72 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=3.4
+ $Y2=0
r132 34 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0
r133 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0.39
r134 30 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0
r135 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0.39
r136 29 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.72
+ $Y2=0
r137 28 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.725
+ $Y2=0
r138 28 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.56 $Y=0
+ $X2=0.805 $Y2=0
r139 24 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r140 24 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.66
r141 7 48 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.57
+ $Y=0.235 $X2=5.705 $Y2=0.39
r142 6 44 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.73
+ $Y=0.235 $X2=4.865 $Y2=0.39
r143 5 79 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=3.88
+ $Y=0.235 $X2=4.025 $Y2=0.39
r144 4 74 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.235 $X2=3.485 $Y2=0.39
r145 3 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.235 $X2=2.645 $Y2=0.39
r146 2 32 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.6
+ $Y=0.235 $X2=1.725 $Y2=0.39
r147 1 26 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.465 $X2=0.72 $Y2=0.66
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__and4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.330000 1.635000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 0.765000 4.175000 1.305000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 0.420000 3.175000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.425000 3.655000 1.405000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.545000 1.320000 1.715000 ;
        RECT 1.015000 0.255000 1.240000 1.545000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.410000  0.085000 1.740000 0.465000 ;
        RECT 3.835000  0.085000 4.085000 0.585000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.515000 2.255000 0.845000 2.635000 ;
        RECT 1.490000 2.255000 2.160000 2.635000 ;
        RECT 2.735000 2.255000 3.075000 2.635000 ;
        RECT 3.755000 2.255000 4.085000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.255000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.670000 0.805000 ;
      RECT 0.175000 1.885000 1.925000 2.055000 ;
      RECT 0.175000 2.055000 0.345000 2.465000 ;
      RECT 0.500000 0.805000 0.670000 1.885000 ;
      RECT 1.415000 0.635000 2.405000 0.805000 ;
      RECT 1.415000 0.805000 1.585000 1.325000 ;
      RECT 1.755000 0.995000 2.065000 1.325000 ;
      RECT 1.755000 1.325000 1.925000 1.885000 ;
      RECT 2.010000 0.255000 2.180000 0.635000 ;
      RECT 2.235000 0.805000 2.405000 1.915000 ;
      RECT 2.235000 1.915000 3.415000 2.085000 ;
      RECT 2.395000 2.085000 2.565000 2.465000 ;
      RECT 2.575000 1.400000 2.745000 1.575000 ;
      RECT 2.575000 1.575000 3.755000 1.745000 ;
      RECT 3.245000 2.085000 3.415000 2.465000 ;
      RECT 3.585000 1.745000 3.755000 1.915000 ;
      RECT 3.585000 1.915000 4.515000 2.085000 ;
      RECT 4.255000 0.255000 4.515000 0.585000 ;
      RECT 4.255000 2.085000 4.515000 2.465000 ;
      RECT 4.345000 0.585000 4.515000 1.915000 ;
  END
END sky130_fd_sc_hd__and4bb_2

* File: sky130_fd_sc_hd__o211ai_4.spice
* Created: Thu Aug 27 14:35:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o211ai_4.pex.spice"
.subckt sky130_fd_sc_hd__o211ai_4  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM0_noxref N_VGND_M0_noxref_d N_A1_M0_noxref_g N_noxref_10_M0_noxref_s VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1_noxref N_noxref_10_M1_noxref_d N_A1_M1_noxref_g N_VGND_M0_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75000.6 SB=75006.4 A=0.0975 P=1.6 MULT=1
MM2_noxref N_VGND_M2_noxref_d N_A1_M2_noxref_g N_noxref_10_M1_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75001.1 SB=75005.9 A=0.0975 P=1.6 MULT=1
MM3_noxref N_noxref_10_M3_noxref_d N_A2_M3_noxref_g N_VGND_M2_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75001.5 SB=75005.5 A=0.0975 P=1.6 MULT=1
MM4_noxref N_VGND_M4_noxref_d N_A2_M4_noxref_g N_noxref_10_M3_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75001.9 SB=75005.1 A=0.0975 P=1.6 MULT=1
MM5_noxref N_noxref_10_M5_noxref_d N_A2_M5_noxref_g N_VGND_M4_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75002.3 SB=75004.7 A=0.0975 P=1.6 MULT=1
MM6_noxref N_VGND_M6_noxref_d N_A2_M6_noxref_g N_noxref_10_M5_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.09425 AS=0.091 PD=0.94 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75002.8 SB=75004.2 A=0.0975 P=1.6 MULT=1
MM7_noxref N_noxref_10_M7_noxref_d N_A1_M7_noxref_g N_VGND_M6_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.10075 AS=0.09425 PD=0.96 PS=0.94 NRD=1.836 NRS=1.836
+ M=1 R=4.33333 SA=75003.2 SB=75003.8 A=0.0975 P=1.6 MULT=1
MM8_noxref N_noxref_12_M8_noxref_d N_B1_M8_noxref_g N_noxref_10_M7_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.10075 PD=0.93 PS=0.96 NRD=0 NRS=3.684 M=1
+ R=4.33333 SA=75003.7 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM9_noxref N_noxref_10_M9_noxref_d N_B1_M9_noxref_g N_noxref_12_M8_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75004.1 SB=75002.9 A=0.0975 P=1.6 MULT=1
MM10_noxref noxref_13 N_B1_M10_noxref_g N_noxref_10_M9_noxref_d VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.091 PD=0.92 PS=0.93 NRD=14.76 NRS=0 M=1
+ R=4.33333 SA=75004.5 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM11_noxref N_Y_M11_noxref_d N_C1_M11_noxref_g noxref_13 VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333
+ SA=75004.9 SB=75002 A=0.0975 P=1.6 MULT=1
MM12_noxref N_noxref_12_M12_noxref_d N_C1_M12_noxref_g N_Y_M11_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75005.4 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM13_noxref N_Y_M13_noxref_d N_C1_M13_noxref_g N_noxref_12_M12_noxref_d VNB
+ NSHORT L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.33333 SA=75005.8 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM14_noxref noxref_14 N_C1_M14_noxref_g N_Y_M13_noxref_d VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=19.38 NRS=0 M=1 R=4.33333
+ SA=75006.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM15_noxref N_noxref_10_M15_noxref_d N_B1_M15_noxref_g noxref_14 VNB NSHORT
+ L=0.15 W=0.65 AD=0.25675 AS=0.104 PD=2.09 PS=0.97 NRD=0 NRS=19.38 M=1
+ R=4.33333 SA=75006.7 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_110_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75007
+ A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A1_M1013_g N_A_110_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1013_d N_A1_M1017_g N_A_110_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75006.2
+ A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_A2_M1007_g N_A_110_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75005.7 A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1007_d N_A2_M1010_g N_A_110_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1021 N_Y_M1021_d N_A2_M1021_g N_A_110_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1027 N_Y_M1021_d N_A2_M1027_g N_A_110_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1029 N_VPWR_M1029_d N_A1_M1029_g N_A_110_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.14 PD=1.32 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1029_d N_B1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75003.7 SB=75003.6
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75003.1 A=0.15
+ P=2.3 MULT=1
MM1011 N_VPWR_M1003_d N_B1_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5 SB=75002.7
+ A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.9 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1000_d N_C1_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.4 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_C1_M1024_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.8 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1024_d N_C1_M1030_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.2 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_B1_M1023_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1 AD=0.675
+ AS=0.135 PD=3.35 PS=1.27 NRD=76.8103 NRS=0 M=1 R=6.66667 SA=75006.6 SB=75000.6
+ A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__o211ai_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o41ai_1.spice.SKY130_FD_SC_HD__O41AI_1.pxi
* Created: Thu Aug 27 14:42:06 2020
* 
x_PM_SKY130_FD_SC_HD__O41AI_1%B1 N_B1_M1008_g N_B1_M1006_g B1 N_B1_c_58_n
+ PM_SKY130_FD_SC_HD__O41AI_1%B1
x_PM_SKY130_FD_SC_HD__O41AI_1%A4 N_A4_M1003_g N_A4_M1007_g A4 A4 A4 A4
+ N_A4_c_84_n A4 PM_SKY130_FD_SC_HD__O41AI_1%A4
x_PM_SKY130_FD_SC_HD__O41AI_1%A3 N_A3_c_119_n N_A3_M1001_g N_A3_M1005_g A3 A3 A3
+ A3 N_A3_c_121_n A3 PM_SKY130_FD_SC_HD__O41AI_1%A3
x_PM_SKY130_FD_SC_HD__O41AI_1%A2 N_A2_M1000_g N_A2_M1002_g N_A2_c_158_n
+ N_A2_c_159_n A2 A2 A2 N_A2_c_160_n A2 PM_SKY130_FD_SC_HD__O41AI_1%A2
x_PM_SKY130_FD_SC_HD__O41AI_1%A1 N_A1_M1009_g N_A1_M1004_g A1 N_A1_c_200_n
+ N_A1_c_201_n PM_SKY130_FD_SC_HD__O41AI_1%A1
x_PM_SKY130_FD_SC_HD__O41AI_1%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_c_226_n
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n VPWR N_VPWR_c_230_n
+ N_VPWR_c_225_n PM_SKY130_FD_SC_HD__O41AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O41AI_1%Y N_Y_M1008_s N_Y_M1006_d N_Y_c_268_n N_Y_c_269_n
+ N_Y_c_264_n Y Y Y N_Y_c_266_n N_Y_c_281_n PM_SKY130_FD_SC_HD__O41AI_1%Y
x_PM_SKY130_FD_SC_HD__O41AI_1%A_109_47# N_A_109_47#_M1008_d N_A_109_47#_M1001_d
+ N_A_109_47#_M1009_d N_A_109_47#_c_310_n N_A_109_47#_c_305_n
+ N_A_109_47#_c_306_n N_A_109_47#_c_318_n N_A_109_47#_c_307_n
+ N_A_109_47#_c_308_n N_A_109_47#_c_312_n N_A_109_47#_c_309_n
+ PM_SKY130_FD_SC_HD__O41AI_1%A_109_47#
x_PM_SKY130_FD_SC_HD__O41AI_1%VGND N_VGND_M1007_d N_VGND_M1000_d N_VGND_c_363_n
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n
+ VGND N_VGND_c_369_n N_VGND_c_370_n PM_SKY130_FD_SC_HD__O41AI_1%VGND
cc_1 VNB N_B1_M1008_g 0.0258462f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB B1 0.00739817f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_B1_c_58_n 0.0363687f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A4_M1003_g 5.5096e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_5 VNB N_A4_M1007_g 0.0202342f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_6 VNB N_A4_c_84_n 0.0448336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A3_c_119_n 0.0162239f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.015
cc_8 VNB A3 0.0036865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A3_c_121_n 0.0191057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A2_c_158_n 0.00317632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_159_n 0.0201408f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_12 VNB N_A2_c_160_n 0.0169356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A1 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_200_n 0.0271099f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_15 VNB N_A1_c_201_n 0.0223997f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_16 VNB N_VPWR_c_225_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_264_n 0.00930481f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_18 VNB Y 0.00878064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_266_n 0.0191417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_109_47#_c_305_n 0.00712135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_109_47#_c_306_n 0.00136544f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_22 VNB N_A_109_47#_c_307_n 0.0164571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_109_47#_c_308_n 0.0183265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_109_47#_c_309_n 0.00740981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_363_n 0.00179054f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB N_VGND_c_364_n 0.0045551f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_27 VNB N_VGND_c_365_n 0.0338183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_366_n 0.00353557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_367_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_368_n 0.00477499f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_369_n 0.0224886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_370_n 0.187786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_B1_M1006_g 0.0268384f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_34 VPB N_B1_c_58_n 0.00817555f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_35 VPB N_A4_M1003_g 0.0232068f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_36 VPB A4 0.00243409f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_37 VPB N_A3_M1005_g 0.0201605f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_38 VPB A3 0.00246507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A3_c_121_n 0.00462864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A2_M1002_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_41 VPB N_A2_c_158_n 0.00176078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A2_c_159_n 0.00501495f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_43 VPB A2 0.0013088f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_44 VPB N_A1_M1004_g 0.0262162f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB A1 0.00713362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A1_c_200_n 0.00473372f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_47 VPB N_VPWR_c_226_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_48 VPB N_VPWR_c_227_n 0.046825f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_49 VPB N_VPWR_c_228_n 0.0155734f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_50 VPB N_VPWR_c_229_n 0.0404601f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_51 VPB N_VPWR_c_230_n 0.0610169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_225_n 0.0498011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB Y 0.0026809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 N_B1_M1006_g N_A4_M1003_g 0.0127862f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_55 N_B1_M1008_g N_A4_M1007_g 0.00938661f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_56 N_B1_c_58_n N_A4_c_84_n 0.0127862f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_57 N_B1_M1006_g N_VPWR_c_227_n 0.00545717f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_58 B1 N_VPWR_c_227_n 0.0194886f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_59 N_B1_c_58_n N_VPWR_c_227_n 0.00562759f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_60 N_B1_M1006_g N_VPWR_c_230_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_61 N_B1_M1006_g N_VPWR_c_225_n 0.0104829f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_62 N_B1_M1006_g N_Y_c_268_n 0.00254657f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_63 N_B1_M1006_g N_Y_c_269_n 0.00918977f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_64 N_B1_M1008_g N_Y_c_264_n 0.00127099f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_65 B1 N_Y_c_264_n 0.0258576f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B1_c_58_n N_Y_c_264_n 0.00706028f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B1_M1008_g Y 0.0221989f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_68 B1 Y 0.0159653f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_69 N_B1_M1008_g N_Y_c_266_n 0.00853413f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_70 N_B1_M1008_g N_A_109_47#_c_310_n 0.00138815f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_71 N_B1_M1008_g N_A_109_47#_c_306_n 4.80492e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_72 N_B1_M1008_g N_A_109_47#_c_312_n 0.00313805f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_73 N_B1_M1008_g N_VGND_c_365_n 0.00424416f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_74 N_B1_M1008_g N_VGND_c_370_n 0.00755765f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_75 N_A4_M1007_g N_A3_c_119_n 0.0260468f $X=1.245 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_76 N_A4_M1003_g N_A3_M1005_g 0.016935f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_77 A4 N_A3_M1005_g 0.00362562f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_78 A4 A3 0.0979774f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A4_c_84_n A3 0.00130936f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A4_M1003_g N_A3_c_121_n 4.00465e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A4_M1007_g N_A3_c_121_n 0.0200183f $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_82 A4 N_A3_c_121_n 2.62319e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A4_M1003_g N_VPWR_c_230_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_84 A4 N_VPWR_c_230_n 0.0122963f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A4_M1003_g N_VPWR_c_225_n 0.0104274f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_86 A4 N_VPWR_c_225_n 0.0109874f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A4_M1003_g N_Y_c_268_n 0.00317169f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A4_M1003_g N_Y_c_269_n 0.0127924f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A4_M1007_g Y 0.00216425f $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_90 A4 Y 0.0256632f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_91 N_A4_c_84_n Y 0.00484198f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A4_M1007_g N_Y_c_281_n 3.51083e-19 $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_93 A4 A_193_297# 0.0257016f $X=1.07 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_94 N_A4_M1007_g N_A_109_47#_c_305_n 0.00999717f $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_95 A4 N_A_109_47#_c_305_n 0.0153079f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A4_c_84_n N_A_109_47#_c_305_n 0.00113821f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_97 A4 N_A_109_47#_c_306_n 0.0112664f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_98 N_A4_c_84_n N_A_109_47#_c_306_n 0.00499404f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A4_M1007_g N_A_109_47#_c_318_n 4.93858e-19 $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A4_c_84_n N_A_109_47#_c_312_n 0.00439247f $X=1.245 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A4_M1007_g N_VGND_c_363_n 0.0090609f $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_102 N_A4_M1007_g N_VGND_c_365_n 0.00350562f $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A4_M1007_g N_VGND_c_370_n 0.00488574f $X=1.245 $Y=0.56 $X2=0 $Y2=0
cc_104 N_A3_M1005_g N_A2_M1002_g 0.06212f $X=1.665 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A3_M1005_g N_A2_c_158_n 2.61427e-19 $X=1.665 $Y=1.985 $X2=0 $Y2=0
cc_106 A3 N_A2_c_158_n 0.027631f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A3_c_121_n N_A2_c_158_n 7.79211e-19 $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_108 A3 N_A2_c_159_n 0.00423262f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_109 N_A3_c_121_n N_A2_c_159_n 0.0219893f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A3_M1005_g A2 8.09612e-19 $X=1.665 $Y=1.985 $X2=0 $Y2=0
cc_111 A3 A2 0.0405154f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_112 N_A3_c_119_n N_A2_c_160_n 0.0124239f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A3_M1005_g N_VPWR_c_230_n 0.0037962f $X=1.665 $Y=1.985 $X2=0 $Y2=0
cc_114 A3 N_VPWR_c_230_n 0.0105675f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A3_M1005_g N_VPWR_c_225_n 0.00606999f $X=1.665 $Y=1.985 $X2=0 $Y2=0
cc_116 A3 N_VPWR_c_225_n 0.0108043f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_117 A3 A_193_297# 0.00907589f $X=1.53 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_118 A3 A_348_297# 0.00774476f $X=1.53 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_119 N_A3_c_119_n N_A_109_47#_c_305_n 0.00845282f $X=1.665 $Y=0.995 $X2=0
+ $Y2=0
cc_120 A3 N_A_109_47#_c_305_n 0.0163508f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A3_c_121_n N_A_109_47#_c_305_n 0.001478f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A3_c_119_n N_A_109_47#_c_318_n 0.0066297f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A3_c_119_n N_A_109_47#_c_309_n 0.00109929f $X=1.665 $Y=0.995 $X2=0
+ $Y2=0
cc_124 A3 N_A_109_47#_c_309_n 0.0104896f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_125 N_A3_c_121_n N_A_109_47#_c_309_n 0.00153445f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A3_c_119_n N_VGND_c_363_n 0.00151363f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A3_c_119_n N_VGND_c_367_n 0.00424416f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A3_c_119_n N_VGND_c_370_n 0.00579048f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_M1002_g N_A1_M1004_g 0.0406049f $X=2.085 $Y=1.985 $X2=0 $Y2=0
cc_130 A2 N_A1_M1004_g 0.00556866f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_131 N_A2_c_158_n A1 0.021657f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A2_c_159_n A1 8.41439e-19 $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A2_c_158_n N_A1_c_200_n 0.00636329f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A2_c_159_n N_A1_c_200_n 0.0220307f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A2_c_160_n N_A1_c_201_n 0.0238041f $X=2.155 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A2_M1002_g N_VPWR_c_229_n 0.00230591f $X=2.085 $Y=1.985 $X2=0 $Y2=0
cc_137 A2 N_VPWR_c_229_n 0.0432714f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_138 N_A2_M1002_g N_VPWR_c_230_n 0.0037962f $X=2.085 $Y=1.985 $X2=0 $Y2=0
cc_139 A2 N_VPWR_c_230_n 0.0121189f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_140 N_A2_M1002_g N_VPWR_c_225_n 0.00558949f $X=2.085 $Y=1.985 $X2=0 $Y2=0
cc_141 A2 N_VPWR_c_225_n 0.0115295f $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_142 A2 A_432_297# 0.0107881f $X=1.99 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_143 N_A2_c_160_n N_A_109_47#_c_318_n 0.00674362f $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A2_c_158_n N_A_109_47#_c_307_n 0.0227435f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A2_c_159_n N_A_109_47#_c_307_n 0.00344866f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A2_c_160_n N_A_109_47#_c_307_n 0.00889201f $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A2_c_160_n N_A_109_47#_c_308_n 5.98596e-19 $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A2_c_158_n N_A_109_47#_c_309_n 0.00337155f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_149 A2 N_A_109_47#_c_309_n 3.90715e-19 $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_150 N_A2_c_160_n N_A_109_47#_c_309_n 0.00109929f $X=2.155 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A2_c_160_n N_VGND_c_364_n 0.00332976f $X=2.155 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_160_n N_VGND_c_367_n 0.00424416f $X=2.155 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A2_c_160_n N_VGND_c_370_n 0.00602715f $X=2.155 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_M1004_g N_VPWR_c_229_n 0.0206173f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_155 A1 N_VPWR_c_229_n 0.0245544f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_200_n N_VPWR_c_229_n 0.00308771f $X=2.665 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_M1004_g N_VPWR_c_230_n 0.0046653f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A1_M1004_g N_VPWR_c_225_n 0.00818715f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A1_c_201_n N_A_109_47#_c_318_n 5.74964e-19 $X=2.655 $Y=0.995 $X2=0
+ $Y2=0
cc_160 A1 N_A_109_47#_c_307_n 0.0368327f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A1_c_200_n N_A_109_47#_c_307_n 0.00358305f $X=2.665 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A1_c_201_n N_A_109_47#_c_307_n 0.010165f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_201_n N_A_109_47#_c_308_n 0.00674362f $X=2.655 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A1_c_201_n N_VGND_c_364_n 0.00291323f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_201_n N_VGND_c_369_n 0.00424416f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_201_n N_VGND_c_370_n 0.0070266f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_167 N_VPWR_c_225_n N_Y_M1006_d 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_c_230_n N_Y_c_269_n 0.0189039f $X=2.63 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_225_n N_Y_c_269_n 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_170 N_VPWR_c_227_n N_Y_c_264_n 7.91944e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_171 N_VPWR_c_227_n Y 0.00222406f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_172 N_VPWR_c_225_n A_193_297# 0.0133331f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_173 N_VPWR_c_225_n A_348_297# 0.00818446f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_174 N_VPWR_c_225_n A_432_297# 0.0091721f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_175 N_Y_c_281_n N_A_109_47#_M1008_d 0.00532792f $X=0.695 $Y=0.905 $X2=-0.19
+ $Y2=-0.24
cc_176 N_Y_c_266_n N_A_109_47#_c_310_n 0.00517226f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_177 N_Y_c_281_n N_A_109_47#_c_306_n 0.0154231f $X=0.695 $Y=0.905 $X2=0 $Y2=0
cc_178 N_Y_c_266_n N_A_109_47#_c_312_n 0.0134111f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_179 Y N_VGND_c_365_n 0.00210502f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_180 N_Y_c_266_n N_VGND_c_365_n 0.0216897f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_181 N_Y_c_281_n N_VGND_c_365_n 0.00267765f $X=0.695 $Y=0.905 $X2=0 $Y2=0
cc_182 N_Y_M1008_s N_VGND_c_370_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_183 Y N_VGND_c_370_n 0.00424379f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_184 N_Y_c_266_n N_VGND_c_370_n 0.0127966f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_185 N_Y_c_281_n N_VGND_c_370_n 0.00475098f $X=0.695 $Y=0.905 $X2=0 $Y2=0
cc_186 N_A_109_47#_c_305_n N_VGND_M1007_d 0.00162006f $X=1.71 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_109_47#_c_307_n N_VGND_M1000_d 0.00245086f $X=2.63 $Y=0.82 $X2=0
+ $Y2=0
cc_188 N_A_109_47#_c_305_n N_VGND_c_363_n 0.0143302f $X=1.71 $Y=0.82 $X2=0 $Y2=0
cc_189 N_A_109_47#_c_307_n N_VGND_c_364_n 0.018519f $X=2.63 $Y=0.82 $X2=0 $Y2=0
cc_190 N_A_109_47#_c_305_n N_VGND_c_365_n 0.00193763f $X=1.71 $Y=0.82 $X2=0
+ $Y2=0
cc_191 N_A_109_47#_c_312_n N_VGND_c_365_n 0.0222091f $X=0.955 $Y=0.38 $X2=0
+ $Y2=0
cc_192 N_A_109_47#_c_305_n N_VGND_c_367_n 0.00193763f $X=1.71 $Y=0.82 $X2=0
+ $Y2=0
cc_193 N_A_109_47#_c_318_n N_VGND_c_367_n 0.0188551f $X=1.875 $Y=0.38 $X2=0
+ $Y2=0
cc_194 N_A_109_47#_c_307_n N_VGND_c_367_n 0.00193763f $X=2.63 $Y=0.82 $X2=0
+ $Y2=0
cc_195 N_A_109_47#_c_307_n N_VGND_c_369_n 0.00193763f $X=2.63 $Y=0.82 $X2=0
+ $Y2=0
cc_196 N_A_109_47#_c_308_n N_VGND_c_369_n 0.0209479f $X=2.795 $Y=0.38 $X2=0
+ $Y2=0
cc_197 N_A_109_47#_M1008_d N_VGND_c_370_n 0.00689388f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_198 N_A_109_47#_M1001_d N_VGND_c_370_n 0.00215201f $X=1.74 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_109_47#_M1009_d N_VGND_c_370_n 0.00225715f $X=2.66 $Y=0.235 $X2=0
+ $Y2=0
cc_200 N_A_109_47#_c_305_n N_VGND_c_370_n 0.00860816f $X=1.71 $Y=0.82 $X2=0
+ $Y2=0
cc_201 N_A_109_47#_c_318_n N_VGND_c_370_n 0.0122069f $X=1.875 $Y=0.38 $X2=0
+ $Y2=0
cc_202 N_A_109_47#_c_307_n N_VGND_c_370_n 0.00859465f $X=2.63 $Y=0.82 $X2=0
+ $Y2=0
cc_203 N_A_109_47#_c_308_n N_VGND_c_370_n 0.0124119f $X=2.795 $Y=0.38 $X2=0
+ $Y2=0
cc_204 N_A_109_47#_c_312_n N_VGND_c_370_n 0.0125064f $X=0.955 $Y=0.38 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__inv_1.pxi.spice
* Created: Tue Sep  1 19:09:55 2020
* 
x_PM_SKY130_FD_SC_HD__INV_1%A N_A_c_24_n N_A_M1000_g N_A_M1001_g A N_A_c_26_n
+ PM_SKY130_FD_SC_HD__INV_1%A
x_PM_SKY130_FD_SC_HD__INV_1%VPWR N_VPWR_M1001_s N_VPWR_c_47_n N_VPWR_c_48_n
+ N_VPWR_c_49_n VPWR N_VPWR_c_50_n N_VPWR_c_46_n PM_SKY130_FD_SC_HD__INV_1%VPWR
x_PM_SKY130_FD_SC_HD__INV_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_60_n N_Y_c_63_n
+ N_Y_c_61_n Y Y Y PM_SKY130_FD_SC_HD__INV_1%Y
x_PM_SKY130_FD_SC_HD__INV_1%VGND N_VGND_M1000_s N_VGND_c_79_n N_VGND_c_80_n
+ N_VGND_c_81_n VGND N_VGND_c_82_n N_VGND_c_83_n PM_SKY130_FD_SC_HD__INV_1%VGND
cc_1 VNB N_A_c_24_n 0.0246111f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=0.995
cc_2 VNB A 0.00854082f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.105
cc_3 VNB N_A_c_26_n 0.0402191f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.16
cc_4 VNB N_VPWR_c_46_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_Y_c_60_n 0.0182459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_Y_c_61_n 0.00657112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB Y 0.0207596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_VGND_c_79_n 0.0308334f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.985
cc_9 VNB N_VGND_c_80_n 0.0123263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_81_n 0.00442067f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_11 VNB N_VGND_c_82_n 0.025344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_83_n 0.123366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VPB N_A_M1001_g 0.0293457f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.985
cc_14 VPB A 3.35665e-19 $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.105
cc_15 VPB N_A_c_26_n 0.0109207f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_16 VPB N_VPWR_c_47_n 0.00491148f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.985
cc_17 VPB N_VPWR_c_48_n 0.0129628f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_18 VPB N_VPWR_c_49_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_19 VPB N_VPWR_c_50_n 0.025344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_46_n 0.063167f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_21 VPB N_Y_c_63_n 0.0317948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_22 VPB Y 0.00883839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB Y 0.00657112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 N_A_M1001_g N_VPWR_c_47_n 0.00444548f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_25 A N_VPWR_c_47_n 0.0158179f $X=0.36 $Y=1.105 $X2=0 $Y2=0
cc_26 N_A_c_26_n N_VPWR_c_47_n 0.00486071f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_27 N_A_M1001_g N_VPWR_c_50_n 0.00541359f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_28 N_A_M1001_g N_VPWR_c_46_n 0.0117186f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_29 N_A_c_24_n N_Y_c_60_n 0.00534153f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_30 N_A_M1001_g N_Y_c_63_n 0.00918977f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_31 N_A_c_24_n N_Y_c_61_n 0.00256049f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_32 N_A_c_24_n Y 0.0207536f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_33 A Y 0.0183958f $X=0.36 $Y=1.105 $X2=0 $Y2=0
cc_34 N_A_M1001_g Y 0.002888f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_35 N_A_c_24_n N_VGND_c_79_n 0.00494327f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_36 A N_VGND_c_79_n 0.0188164f $X=0.36 $Y=1.105 $X2=0 $Y2=0
cc_37 N_A_c_26_n N_VGND_c_79_n 0.00585411f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_38 N_A_c_24_n N_VGND_c_82_n 0.00541359f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_39 N_A_c_24_n N_VGND_c_83_n 0.0117186f $X=0.675 $Y=0.995 $X2=0 $Y2=0
cc_40 N_VPWR_c_46_n N_Y_M1001_d 0.00209319f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_41 N_VPWR_c_50_n N_Y_c_63_n 0.0210382f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_42 N_VPWR_c_46_n N_Y_c_63_n 0.0124268f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_43 Y N_VGND_c_79_n 0.00108376f $X=0.82 $Y=1.105 $X2=0 $Y2=0
cc_44 N_Y_c_60_n N_VGND_c_82_n 0.0210225f $X=0.885 $Y=0.4 $X2=0 $Y2=0
cc_45 N_Y_M1000_d N_VGND_c_83_n 0.00209319f $X=0.75 $Y=0.235 $X2=0 $Y2=0
cc_46 N_Y_c_60_n N_VGND_c_83_n 0.0124193f $X=0.885 $Y=0.4 $X2=0 $Y2=0

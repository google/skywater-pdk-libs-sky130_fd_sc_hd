* File: sky130_fd_sc_hd__o22ai_2.spice.SKY130_FD_SC_HD__O22AI_2.pxi
* Created: Thu Aug 27 14:37:59 2020
* 
x_PM_SKY130_FD_SC_HD__O22AI_2%B1 N_B1_c_69_n N_B1_M1004_g N_B1_M1001_g
+ N_B1_c_70_n N_B1_M1007_g N_B1_M1015_g B1 N_B1_c_71_n N_B1_c_72_n
+ PM_SKY130_FD_SC_HD__O22AI_2%B1
x_PM_SKY130_FD_SC_HD__O22AI_2%B2 N_B2_c_110_n N_B2_M1002_g N_B2_M1010_g
+ N_B2_c_111_n N_B2_M1006_g N_B2_M1012_g B2 N_B2_c_112_n N_B2_c_113_n
+ PM_SKY130_FD_SC_HD__O22AI_2%B2
x_PM_SKY130_FD_SC_HD__O22AI_2%A2 N_A2_c_158_n N_A2_M1008_g N_A2_M1000_g
+ N_A2_c_159_n N_A2_M1014_g N_A2_M1003_g A2 N_A2_c_161_n
+ PM_SKY130_FD_SC_HD__O22AI_2%A2
x_PM_SKY130_FD_SC_HD__O22AI_2%A1 N_A1_c_210_n N_A1_M1009_g N_A1_M1005_g
+ N_A1_c_211_n N_A1_M1011_g N_A1_M1013_g A1 N_A1_c_213_n
+ PM_SKY130_FD_SC_HD__O22AI_2%A1
x_PM_SKY130_FD_SC_HD__O22AI_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1015_s
+ N_A_27_297#_M1012_d N_A_27_297#_c_252_n N_A_27_297#_c_269_p
+ N_A_27_297#_c_253_n N_A_27_297#_c_254_n N_A_27_297#_c_267_p
+ N_A_27_297#_c_263_n N_A_27_297#_c_284_p PM_SKY130_FD_SC_HD__O22AI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__O22AI_2%VPWR N_VPWR_M1001_d N_VPWR_M1005_s N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n VPWR N_VPWR_c_293_n
+ N_VPWR_c_294_n N_VPWR_c_288_n N_VPWR_c_296_n PM_SKY130_FD_SC_HD__O22AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O22AI_2%Y N_Y_M1004_s N_Y_M1002_d N_Y_M1010_s N_Y_M1000_s
+ N_Y_c_343_n N_Y_c_348_n N_Y_c_344_n N_Y_c_345_n N_Y_c_346_n N_Y_c_349_n
+ N_Y_c_350_n Y N_Y_c_352_n Y PM_SKY130_FD_SC_HD__O22AI_2%Y
x_PM_SKY130_FD_SC_HD__O22AI_2%A_475_297# N_A_475_297#_M1000_d
+ N_A_475_297#_M1003_d N_A_475_297#_M1013_d N_A_475_297#_c_431_n
+ N_A_475_297#_c_421_n N_A_475_297#_c_432_n N_A_475_297#_c_418_n
+ N_A_475_297#_c_440_n N_A_475_297#_c_419_n N_A_475_297#_c_420_n
+ N_A_475_297#_c_444_n PM_SKY130_FD_SC_HD__O22AI_2%A_475_297#
x_PM_SKY130_FD_SC_HD__O22AI_2%A_27_47# N_A_27_47#_M1004_d N_A_27_47#_M1007_d
+ N_A_27_47#_M1006_s N_A_27_47#_M1014_s N_A_27_47#_M1011_d N_A_27_47#_c_454_n
+ N_A_27_47#_c_455_n N_A_27_47#_c_464_n N_A_27_47#_c_471_n N_A_27_47#_c_469_n
+ N_A_27_47#_c_456_n N_A_27_47#_c_457_n N_A_27_47#_c_481_n N_A_27_47#_c_458_n
+ N_A_27_47#_c_459_n N_A_27_47#_c_460_n PM_SKY130_FD_SC_HD__O22AI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O22AI_2%VGND N_VGND_M1008_d N_VGND_M1009_s N_VGND_c_534_n
+ N_VGND_c_535_n N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n
+ VGND N_VGND_c_540_n N_VGND_c_541_n PM_SKY130_FD_SC_HD__O22AI_2%VGND
cc_1 VNB N_B1_c_69_n 0.0213689f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_B1_c_70_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_B1_c_71_n 0.0119843f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_4 VNB N_B1_c_72_n 0.0430453f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_5 VNB N_B2_c_110_n 0.0159993f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B2_c_111_n 0.0193754f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_7 VNB N_B2_c_112_n 0.0404324f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_8 VNB N_B2_c_113_n 0.00331652f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_9 VNB N_A2_c_158_n 0.0194756f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_A2_c_159_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_11 VNB A2 0.0029367f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_12 VNB N_A2_c_161_n 0.0390646f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_13 VNB N_A1_c_210_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_14 VNB N_A1_c_211_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_15 VNB A1 0.0116392f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_16 VNB N_A1_c_213_n 0.0426809f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_17 VNB N_VPWR_c_288_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_343_n 0.00315786f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_19 VNB N_Y_c_344_n 0.00219468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_345_n 0.00350868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_346_n 0.0021905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB Y 0.0102314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_454_n 0.0075557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_455_n 0.0210433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_456_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_457_n 0.00144154f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.18
cc_27 VNB N_A_27_47#_c_458_n 0.0143561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_459_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_460_n 0.00384439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_534_n 0.00413609f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.56
cc_31 VNB N_VGND_c_535_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_32 VNB N_VGND_c_536_n 0.0702879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_537_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_34 VNB N_VGND_c_538_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_35 VNB N_VGND_c_539_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=1.16
cc_36 VNB N_VGND_c_540_n 0.0216806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_541_n 0.244474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_B1_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_39 VPB N_B1_M1015_g 0.0185038f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_40 VPB N_B1_c_72_n 0.00740766f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_41 VPB N_B2_M1010_g 0.018814f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_42 VPB N_B2_M1012_g 0.0222273f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_43 VPB N_B2_c_112_n 0.00688651f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_44 VPB N_A2_M1000_g 0.022323f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_45 VPB N_A2_M1003_g 0.018815f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_46 VPB N_A2_c_161_n 0.00689f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_47 VPB N_A1_M1005_g 0.0185038f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_48 VPB N_A1_M1013_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_49 VPB N_A1_c_213_n 0.00740766f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_50 VPB N_A_27_297#_c_252_n 0.00369371f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_51 VPB N_A_27_297#_c_253_n 0.00237544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_254_n 0.00362963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_289_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_54 VPB N_VPWR_c_290_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_55 VPB N_VPWR_c_291_n 0.0689564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_292_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_57 VPB N_VPWR_c_293_n 0.0180608f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_58 VPB N_VPWR_c_294_n 0.0218794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_288_n 0.0634318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_296_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_Y_c_348_n 0.00871165f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_62 VPB N_Y_c_349_n 0.00238006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_Y_c_350_n 0.0023869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB Y 0.0153605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_Y_c_352_n 0.00300151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_475_297#_c_418_n 0.0036062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_475_297#_c_419_n 0.00232133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_475_297#_c_420_n 0.0044132f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.16
cc_69 N_B1_c_70_n N_B2_c_110_n 0.0197588f $X=0.91 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_70 N_B1_M1015_g N_B2_M1010_g 0.0197588f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_71 N_B1_c_71_n N_B2_c_112_n 2.74289e-19 $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B1_c_72_n N_B2_c_112_n 0.0197588f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B1_c_71_n N_B2_c_113_n 0.0176626f $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_74 N_B1_c_72_n N_B2_c_113_n 7.87227e-19 $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B1_c_71_n N_A_27_297#_c_252_n 0.0172172f $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B1_c_72_n N_A_27_297#_c_252_n 0.00220041f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B1_M1001_g N_A_27_297#_c_253_n 0.013451f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B1_M1015_g N_A_27_297#_c_253_n 0.0131689f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B1_c_71_n N_A_27_297#_c_253_n 0.0409752f $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B1_c_72_n N_A_27_297#_c_253_n 0.00234772f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B1_M1001_g N_VPWR_c_289_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_82 N_B1_M1015_g N_VPWR_c_289_n 0.00302074f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_83 N_B1_M1015_g N_VPWR_c_291_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_84 N_B1_M1001_g N_VPWR_c_293_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_85 N_B1_M1001_g N_VPWR_c_288_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_86 N_B1_M1015_g N_VPWR_c_288_n 0.010464f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_87 N_B1_c_69_n N_Y_c_344_n 0.00387612f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B1_c_70_n N_Y_c_344_n 0.00289474f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_c_71_n N_Y_c_344_n 0.0328342f $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B1_c_72_n N_Y_c_344_n 0.00224214f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B1_c_70_n N_Y_c_345_n 0.00762805f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B1_c_70_n N_Y_c_346_n 2.32132e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_93 N_B1_c_69_n N_A_27_47#_c_455_n 4.6346e-19 $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B1_c_71_n N_A_27_47#_c_455_n 0.0137204f $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B1_c_72_n N_A_27_47#_c_455_n 0.00125096f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B1_c_69_n N_A_27_47#_c_464_n 0.00957565f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B1_c_70_n N_A_27_47#_c_464_n 0.0083291f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B1_c_71_n N_A_27_47#_c_464_n 0.00351846f $X=0.82 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B1_c_69_n N_VGND_c_536_n 0.00368123f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B1_c_70_n N_VGND_c_536_n 0.00368123f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_c_69_n N_VGND_c_541_n 0.00621922f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_70_n N_VGND_c_541_n 0.00527354f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B2_c_112_n N_A2_c_161_n 0.00421158f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B2_M1010_g N_A_27_297#_c_254_n 2.57315e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B2_c_113_n N_A_27_297#_c_254_n 0.00733304f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B2_M1010_g N_A_27_297#_c_263_n 0.0121306f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B2_M1012_g N_A_27_297#_c_263_n 0.00984328f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B2_M1010_g N_VPWR_c_291_n 0.00357877f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B2_M1012_g N_VPWR_c_291_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B2_M1010_g N_VPWR_c_288_n 0.00525237f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_111 N_B2_M1012_g N_VPWR_c_288_n 0.00655123f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B2_c_111_n N_Y_c_343_n 0.00964175f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B2_c_112_n N_Y_c_343_n 0.00247123f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B2_c_110_n N_Y_c_344_n 2.32132e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B2_c_110_n N_Y_c_345_n 0.00762314f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B2_c_113_n N_Y_c_345_n 0.0560266f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B2_c_110_n N_Y_c_346_n 0.00289348f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B2_c_111_n N_Y_c_346_n 0.00498062f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B2_c_112_n N_Y_c_346_n 0.00224075f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B2_M1010_g N_Y_c_349_n 5.90444e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B2_c_112_n N_Y_c_349_n 0.00222181f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B2_c_113_n N_Y_c_349_n 0.0204933f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_123 N_B2_c_111_n Y 0.00285931f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B2_M1012_g Y 0.00382312f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_125 N_B2_c_112_n Y 0.00599474f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B2_c_113_n Y 0.0163414f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B2_M1012_g N_Y_c_352_n 0.0135164f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B2_c_112_n N_Y_c_352_n 0.00238426f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B2_c_113_n N_Y_c_352_n 0.018326f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B2_c_110_n N_A_27_47#_c_464_n 0.0083291f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B2_c_111_n N_A_27_47#_c_464_n 0.0083291f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B2_c_111_n N_A_27_47#_c_469_n 0.00392418f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B2_c_111_n N_A_27_47#_c_457_n 5.22916e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B2_c_110_n N_VGND_c_536_n 0.00368123f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B2_c_111_n N_VGND_c_536_n 0.00368123f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B2_c_110_n N_VGND_c_541_n 0.00527354f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B2_c_111_n N_VGND_c_541_n 0.00657241f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A2_c_159_n N_A1_c_210_n 0.0150658f $X=3.15 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_139 N_A2_M1003_g N_A1_M1005_g 0.0150658f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_140 A2 A1 0.0176337f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A2_c_161_n A1 0.00106946f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_142 A2 N_A1_c_213_n 2.068e-19 $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A2_c_161_n N_A1_c_213_n 0.0150658f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_M1000_g N_VPWR_c_291_n 0.00357877f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A2_M1003_g N_VPWR_c_291_n 0.00357877f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A2_M1000_g N_VPWR_c_288_n 0.00655123f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A2_M1003_g N_VPWR_c_288_n 0.00525237f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A2_c_158_n N_Y_c_343_n 0.00101579f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_M1000_g N_Y_c_348_n 0.0135226f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_150 A2 N_Y_c_348_n 0.0183006f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A2_c_161_n N_Y_c_348_n 0.00238134f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A2_M1003_g N_Y_c_350_n 5.90444e-19 $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_153 A2 N_Y_c_350_n 0.0203891f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A2_c_161_n N_Y_c_350_n 0.00222344f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_158_n Y 0.00272643f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_M1000_g Y 0.00364546f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_157 A2 Y 0.0135933f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A2_c_161_n Y 0.00434681f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_M1000_g N_A_475_297#_c_421_n 0.00984328f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A2_M1003_g N_A_475_297#_c_421_n 0.0121306f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A2_M1003_g N_A_475_297#_c_418_n 2.57315e-19 $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A2_c_158_n N_A_27_47#_c_471_n 0.00200126f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_158_n N_A_27_47#_c_469_n 0.00611259f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_159_n N_A_27_47#_c_469_n 4.56713e-19 $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_158_n N_A_27_47#_c_456_n 0.0089828f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A2_c_159_n N_A_27_47#_c_456_n 0.00865686f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_167 A2 N_A_27_47#_c_456_n 0.0364556f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A2_c_161_n N_A_27_47#_c_456_n 0.00222133f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A2_c_158_n N_A_27_47#_c_457_n 0.00389014f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_170 A2 N_A_27_47#_c_457_n 0.0099728f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A2_c_161_n N_A_27_47#_c_457_n 0.00255298f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_c_158_n N_A_27_47#_c_481_n 5.23325e-19 $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_159_n N_A_27_47#_c_481_n 0.00632392f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_c_159_n N_A_27_47#_c_460_n 0.00112787f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_175 A2 N_A_27_47#_c_460_n 0.00230276f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A2_c_158_n N_VGND_c_534_n 0.00268723f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A2_c_159_n N_VGND_c_534_n 0.00146448f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A2_c_158_n N_VGND_c_536_n 0.00426197f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A2_c_159_n N_VGND_c_538_n 0.00423334f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_158_n N_VGND_c_541_n 0.00708259f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A2_c_159_n N_VGND_c_541_n 0.0057435f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_M1005_g N_VPWR_c_290_n 0.00302074f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A1_M1013_g N_VPWR_c_290_n 0.00302074f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A1_M1005_g N_VPWR_c_291_n 0.00585385f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A1_M1013_g N_VPWR_c_294_n 0.00585385f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A1_M1005_g N_VPWR_c_288_n 0.010464f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A1_M1013_g N_VPWR_c_288_n 0.0115008f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_188 A1 N_A_475_297#_c_418_n 0.00771248f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_189 N_A1_M1005_g N_A_475_297#_c_419_n 0.0131689f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A1_M1013_g N_A_475_297#_c_419_n 0.013451f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_191 A1 N_A_475_297#_c_419_n 0.0417028f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_192 N_A1_c_213_n N_A_475_297#_c_419_n 0.00234772f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_193 A1 N_A_475_297#_c_420_n 0.00736234f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_194 N_A1_c_213_n N_A_475_297#_c_420_n 0.00220041f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A1_c_210_n N_A_27_47#_c_481_n 0.00630972f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_211_n N_A_27_47#_c_481_n 5.22228e-19 $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_210_n N_A_27_47#_c_458_n 0.00870364f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_211_n N_A_27_47#_c_458_n 0.00999903f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_199 A1 N_A_27_47#_c_458_n 0.0467034f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_200 N_A1_c_213_n N_A_27_47#_c_458_n 0.00478065f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A1_c_210_n N_A_27_47#_c_459_n 5.22228e-19 $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A1_c_211_n N_A_27_47#_c_459_n 0.00630972f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_210_n N_A_27_47#_c_460_n 0.00112787f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_204 A1 N_A_27_47#_c_460_n 0.0108485f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_205 N_A1_c_210_n N_VGND_c_535_n 0.00146448f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A1_c_211_n N_VGND_c_535_n 0.00268723f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_c_210_n N_VGND_c_538_n 0.00423334f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A1_c_211_n N_VGND_c_540_n 0.00423334f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_210_n N_VGND_c_541_n 0.0057435f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_211_n N_VGND_c_541_n 0.00678032f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_27_297#_c_253_n N_VPWR_M1001_d 0.00165831f $X=0.995 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_212 N_A_27_297#_c_253_n N_VPWR_c_289_n 0.0126919f $X=0.995 $Y=1.54 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_267_p N_VPWR_c_291_n 0.0143053f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_214 N_A_27_297#_c_263_n N_VPWR_c_291_n 0.0489446f $X=1.835 $Y=2.38 $X2=0
+ $Y2=0
cc_215 N_A_27_297#_c_269_p N_VPWR_c_293_n 0.0161885f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_216 N_A_27_297#_M1001_s N_VPWR_c_288_n 0.00315976f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_217 N_A_27_297#_M1015_s N_VPWR_c_288_n 0.00246446f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_218 N_A_27_297#_M1012_d N_VPWR_c_288_n 0.00295147f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_219 N_A_27_297#_c_269_p N_VPWR_c_288_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_220 N_A_27_297#_c_267_p N_VPWR_c_288_n 0.00962794f $X=1.12 $Y=2.295 $X2=0
+ $Y2=0
cc_221 N_A_27_297#_c_263_n N_VPWR_c_288_n 0.0300869f $X=1.835 $Y=2.38 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_c_263_n N_Y_M1010_s 0.00312348f $X=1.835 $Y=2.38 $X2=0 $Y2=0
cc_223 N_A_27_297#_c_253_n N_Y_c_345_n 3.18413e-19 $X=0.995 $Y=1.54 $X2=0 $Y2=0
cc_224 N_A_27_297#_c_254_n N_Y_c_345_n 0.0060312f $X=1.12 $Y=1.625 $X2=0 $Y2=0
cc_225 N_A_27_297#_c_254_n N_Y_c_349_n 0.00271526f $X=1.12 $Y=1.625 $X2=0 $Y2=0
cc_226 N_A_27_297#_c_263_n N_Y_c_349_n 0.0118865f $X=1.835 $Y=2.38 $X2=0 $Y2=0
cc_227 N_A_27_297#_M1012_d Y 5.28596e-19 $X=1.825 $Y=1.485 $X2=0 $Y2=0
cc_228 N_A_27_297#_M1012_d N_Y_c_352_n 0.00322004f $X=1.825 $Y=1.485 $X2=0 $Y2=0
cc_229 N_A_27_297#_c_263_n N_Y_c_352_n 0.00322336f $X=1.835 $Y=2.38 $X2=0 $Y2=0
cc_230 N_A_27_297#_c_284_p N_Y_c_352_n 0.016478f $X=1.96 $Y=1.96 $X2=0 $Y2=0
cc_231 N_A_27_297#_c_284_p N_A_475_297#_c_431_n 0.0246907f $X=1.96 $Y=1.96 $X2=0
+ $Y2=0
cc_232 N_A_27_297#_c_263_n N_A_475_297#_c_432_n 0.00981548f $X=1.835 $Y=2.38
+ $X2=0 $Y2=0
cc_233 N_A_27_297#_c_252_n N_A_27_47#_c_455_n 0.00204459f $X=0.277 $Y=1.625
+ $X2=0 $Y2=0
cc_234 N_VPWR_c_288_n N_Y_M1010_s 0.00216833f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_288_n N_Y_M1000_s 0.00216833f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_c_288_n N_A_475_297#_M1000_d 0.00295147f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_237 N_VPWR_c_288_n N_A_475_297#_M1003_d 0.00246446f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_288_n N_A_475_297#_M1013_d 0.00315976f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_291_n N_A_475_297#_c_421_n 0.0330174f $X=3.655 $Y=2.72 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_288_n N_A_475_297#_c_421_n 0.0204627f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_291_n N_A_475_297#_c_432_n 0.0159273f $X=3.655 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_288_n N_A_475_297#_c_432_n 0.00962421f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_291_n N_A_475_297#_c_440_n 0.0143053f $X=3.655 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_288_n N_A_475_297#_c_440_n 0.00962794f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_M1005_s N_A_475_297#_c_419_n 0.00165831f $X=3.645 $Y=1.485 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_290_n N_A_475_297#_c_419_n 0.0126919f $X=3.78 $Y=1.96 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_294_n N_A_475_297#_c_444_n 0.0161885f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_288_n N_A_475_297#_c_444_n 0.00974347f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_249 N_Y_c_348_n N_A_475_297#_M1000_d 0.00372729f $X=2.815 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_250 N_Y_c_348_n N_A_475_297#_c_431_n 0.016478f $X=2.815 $Y=1.535 $X2=0 $Y2=0
cc_251 N_Y_M1000_s N_A_475_297#_c_421_n 0.00312348f $X=2.805 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_Y_c_348_n N_A_475_297#_c_421_n 0.00322336f $X=2.815 $Y=1.535 $X2=0
+ $Y2=0
cc_253 N_Y_c_350_n N_A_475_297#_c_421_n 0.0118865f $X=2.94 $Y=1.62 $X2=0 $Y2=0
cc_254 N_Y_c_350_n N_A_475_297#_c_418_n 0.00271526f $X=2.94 $Y=1.62 $X2=0 $Y2=0
cc_255 N_Y_c_345_n N_A_27_47#_M1007_d 0.00191752f $X=1.375 $Y=0.775 $X2=0 $Y2=0
cc_256 N_Y_c_343_n N_A_27_47#_M1006_s 0.0101638f $X=2.095 $Y=0.815 $X2=0 $Y2=0
cc_257 N_Y_c_344_n N_A_27_47#_c_455_n 0.0112529f $X=0.865 $Y=0.775 $X2=0 $Y2=0
cc_258 N_Y_M1004_s N_A_27_47#_c_464_n 0.00318958f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_259 N_Y_M1002_d N_A_27_47#_c_464_n 0.00318958f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_260 N_Y_c_343_n N_A_27_47#_c_464_n 0.0296942f $X=2.095 $Y=0.815 $X2=0 $Y2=0
cc_261 N_Y_c_344_n N_A_27_47#_c_464_n 0.015032f $X=0.865 $Y=0.775 $X2=0 $Y2=0
cc_262 N_Y_c_345_n N_A_27_47#_c_464_n 0.0187207f $X=1.375 $Y=0.775 $X2=0 $Y2=0
cc_263 N_Y_c_346_n N_A_27_47#_c_464_n 0.015032f $X=1.705 $Y=0.775 $X2=0 $Y2=0
cc_264 N_Y_c_343_n N_A_27_47#_c_457_n 0.0162997f $X=2.095 $Y=0.815 $X2=0 $Y2=0
cc_265 N_Y_c_348_n N_A_27_47#_c_457_n 0.00169049f $X=2.815 $Y=1.535 $X2=0 $Y2=0
cc_266 N_Y_M1004_s N_VGND_c_541_n 0.00220248f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_267 N_Y_M1002_d N_VGND_c_541_n 0.00220248f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_268 N_A_475_297#_c_420_n N_A_27_47#_c_458_n 0.0067876f $X=4.202 $Y=1.625
+ $X2=0 $Y2=0
cc_269 N_A_475_297#_c_418_n N_A_27_47#_c_460_n 0.00658191f $X=3.36 $Y=1.625
+ $X2=0 $Y2=0
cc_270 N_A_27_47#_c_456_n N_VGND_M1008_d 0.00162089f $X=3.195 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_271 N_A_27_47#_c_458_n N_VGND_M1009_s 0.00162089f $X=4.035 $Y=0.815 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_456_n N_VGND_c_534_n 0.0122559f $X=3.195 $Y=0.815 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_458_n N_VGND_c_535_n 0.0122559f $X=4.035 $Y=0.815 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_454_n N_VGND_c_536_n 0.0143679f $X=0.227 $Y=0.475 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_464_n N_VGND_c_536_n 0.0927884f $X=2.51 $Y=0.39 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_471_n N_VGND_c_536_n 0.00744914f $X=2.595 $Y=0.475 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_456_n N_VGND_c_536_n 0.00205414f $X=3.195 $Y=0.815 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_456_n N_VGND_c_538_n 0.00198695f $X=3.195 $Y=0.815 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_481_n N_VGND_c_538_n 0.0188551f $X=3.36 $Y=0.39 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_458_n N_VGND_c_538_n 0.00198695f $X=4.035 $Y=0.815 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_458_n N_VGND_c_540_n 0.00198695f $X=4.035 $Y=0.815 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_459_n N_VGND_c_540_n 0.0209752f $X=4.2 $Y=0.39 $X2=0 $Y2=0
cc_283 N_A_27_47#_M1004_d N_VGND_c_541_n 0.00229179f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_M1007_d N_VGND_c_541_n 0.00218617f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1006_s N_VGND_c_541_n 0.00683271f $X=1.825 $Y=0.235 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1014_s N_VGND_c_541_n 0.00215201f $X=3.225 $Y=0.235 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1011_d N_VGND_c_541_n 0.00209319f $X=4.065 $Y=0.235 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_454_n N_VGND_c_541_n 0.0102867f $X=0.227 $Y=0.475 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_464_n N_VGND_c_541_n 0.0743659f $X=2.51 $Y=0.39 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_471_n N_VGND_c_541_n 0.00617099f $X=2.595 $Y=0.475 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_456_n N_VGND_c_541_n 0.00846581f $X=3.195 $Y=0.815 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_481_n N_VGND_c_541_n 0.0122069f $X=3.36 $Y=0.39 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_458_n N_VGND_c_541_n 0.00835832f $X=4.035 $Y=0.815 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_459_n N_VGND_c_541_n 0.0124119f $X=4.2 $Y=0.39 $X2=0 $Y2=0

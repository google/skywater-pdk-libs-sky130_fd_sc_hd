# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__buf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 1.660000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 0.255000 2.445000 0.735000 ;
        RECT 2.275000 0.735000 6.645000 0.905000 ;
        RECT 2.275000 1.445000 6.645000 1.615000 ;
        RECT 2.275000 1.615000 2.445000 2.465000 ;
        RECT 3.115000 0.255000 3.285000 0.735000 ;
        RECT 3.115000 1.615000 3.285000 2.465000 ;
        RECT 3.955000 0.255000 4.125000 0.735000 ;
        RECT 3.955000 1.615000 4.125000 2.465000 ;
        RECT 4.710000 0.905000 6.645000 1.445000 ;
        RECT 4.795000 0.255000 4.965000 0.735000 ;
        RECT 4.795000 1.615000 4.965000 2.465000 ;
        RECT 5.635000 0.255000 5.805000 0.735000 ;
        RECT 5.635000 1.615000 5.805000 2.465000 ;
        RECT 6.475000 0.255000 6.645000 0.735000 ;
        RECT 6.475000 1.615000 6.645000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.565000 ;
      RECT 0.175000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  1.445000 2.015000 1.615000 ;
      RECT 0.515000  1.615000 0.845000 2.465000 ;
      RECT 0.595000  0.255000 0.765000 0.735000 ;
      RECT 0.595000  0.735000 2.015000 0.905000 ;
      RECT 0.935000  0.085000 1.265000 0.565000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  1.615000 1.685000 2.465000 ;
      RECT 1.435000  0.260000 1.605000 0.735000 ;
      RECT 1.775000  0.085000 2.105000 0.565000 ;
      RECT 1.840000  0.905000 2.015000 1.075000 ;
      RECT 1.840000  1.075000 4.465000 1.245000 ;
      RECT 1.840000  1.245000 2.015000 1.445000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.615000  0.085000 2.945000 0.565000 ;
      RECT 2.615000  1.835000 2.945000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.565000 ;
      RECT 3.455000  1.835000 3.785000 2.635000 ;
      RECT 4.295000  0.085000 4.625000 0.565000 ;
      RECT 4.295000  1.835000 4.625000 2.635000 ;
      RECT 5.135000  0.085000 5.465000 0.565000 ;
      RECT 5.135000  1.835000 5.465000 2.635000 ;
      RECT 5.975000  0.085000 6.305000 0.565000 ;
      RECT 5.975000  1.835000 6.305000 2.635000 ;
      RECT 6.815000  0.085000 7.145000 0.885000 ;
      RECT 6.815000  1.485000 7.145000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_12
END LIBRARY

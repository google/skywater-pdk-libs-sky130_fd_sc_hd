* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 VGND CLK a_643_369# VNB nshort w=420000u l=150000u
+  ad=1.2937e+12p pd=1.426e+07u as=1.092e+11p ps=1.36e+06u
M1001 a_27_369# a_319_21# a_181_47# VPB phighvt w=640000u l=150000u
+  ad=3.328e+11p pd=3.6e+06u as=2.82e+11p ps=3.18e+06u
M1002 VPWR a_2227_47# Q VPB phighvt w=1e+06u l=150000u
+  ad=1.8638e+12p pd=1.809e+07u as=3.15e+11p ps=2.63e+06u
M1003 a_193_369# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1004 Q a_2227_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_181_47# D a_193_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1129_21# a_997_413# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.428e+11p pd=1.52e+06u as=0p ps=0u
M1007 VPWR a_1781_295# a_1723_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1008 a_997_413# a_809_369# a_181_47# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1009 a_1347_47# a_997_413# a_1129_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u
M1010 VGND a_1597_329# a_2227_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 a_1781_295# a_1597_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1012 a_1525_329# a_997_413# VPWR VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1013 a_181_47# SCE a_109_47# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=8.82e+10p ps=1.26e+06u
M1014 VGND SCE a_319_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1015 a_1514_47# a_997_413# VGND VNB nshort w=640000u l=150000u
+  ad=4.768e+11p pd=2.77e+06u as=0p ps=0u
M1016 a_1781_295# a_1597_329# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1017 a_1597_329# a_643_369# a_1525_329# VPB phighvt w=840000u l=150000u
+  ad=4.158e+11p pd=4e+06u as=0p ps=0u
M1018 VPWR SCD a_27_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_265_47# D a_181_47# VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1020 a_997_413# a_643_369# a_181_47# VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1021 a_1087_47# a_809_369# a_997_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1022 VGND a_1129_21# a_1087_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1597_329# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1597_329# a_2227_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1025 VPWR SCE a_319_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1026 Q a_2227_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.0475e+11p pd=1.93e+06u as=0p ps=0u
M1027 a_809_369# a_643_369# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1028 VPWR SET_B a_1129_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_319_21# a_265_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1815_47# a_643_369# a_1597_329# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.482e+11p ps=2.2e+06u
M1031 a_1723_413# a_809_369# a_1597_329# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1887_47# a_1781_295# a_1815_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1033 VPWR CLK a_643_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1034 a_1081_413# a_643_369# a_997_413# VPB phighvt w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1035 a_809_369# a_643_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1036 VPWR a_1129_21# a_1081_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_109_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND SET_B a_1887_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_2227_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SET_B a_1347_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1597_329# a_809_369# a_1514_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

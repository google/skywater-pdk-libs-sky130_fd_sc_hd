* File: sky130_fd_sc_hd__o31a_4.pex.spice
* Created: Thu Aug 27 14:40:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O31A_4%A_102_21# 1 2 3 12 16 20 24 28 32 36 40 42 46
+ 55 59 60 63 65 67 71 72 74 75 79
c124 74 0 1.68728e-19 $X=3.925 $Y=2.02
c125 65 0 1.24132e-19 $X=3.045 $Y=0.76
c126 59 0 1.49044e-19 $X=2.525 $Y=1.815
r127 75 77 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.455 $Y2=1.16
r128 68 72 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.97
+ $X2=2.525 $Y2=1.97
r129 67 74 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=1.97
+ $X2=3.925 $Y2=1.97
r130 67 68 63.7727 $w=1.98e-07 $l=1.15e-06 $layer=LI1_cond $X=3.76 $Y=1.97
+ $X2=2.61 $Y2=1.97
r131 63 65 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.61 $Y=0.76
+ $X2=3.045 $Y2=0.76
r132 60 72 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.525 $Y=2.07
+ $X2=2.525 $Y2=1.97
r133 60 62 6.1 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.07 $X2=2.525
+ $Y2=2.155
r134 57 72 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.525 $Y=1.87
+ $X2=2.525 $Y2=1.97
r135 57 59 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.525 $Y=1.87
+ $X2=2.525 $Y2=1.815
r136 56 71 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.525 $Y=1.29
+ $X2=2.525 $Y2=1.172
r137 56 59 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.525 $Y=1.29
+ $X2=2.525 $Y2=1.815
r138 55 71 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.525 $Y=1.055
+ $X2=2.525 $Y2=1.172
r139 54 63 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.525 $Y=0.885
+ $X2=2.61 $Y2=0.76
r140 54 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.525 $Y=0.885
+ $X2=2.525 $Y2=1.055
r141 53 79 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.785 $Y=1.16
+ $X2=1.875 $Y2=1.16
r142 53 77 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=1.785 $Y=1.16
+ $X2=1.455 $Y2=1.16
r143 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=1.16 $X2=1.785 $Y2=1.16
r144 49 75 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=1.105 $Y=1.16
+ $X2=1.38 $Y2=1.16
r145 48 52 33.3473 $w=2.33e-07 $l=6.8e-07 $layer=LI1_cond $X=1.105 $Y=1.172
+ $X2=1.785 $Y2=1.172
r146 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.16 $X2=1.105 $Y2=1.16
r147 46 71 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=1.172
+ $X2=2.525 $Y2=1.172
r148 46 52 32.1213 $w=2.33e-07 $l=6.55e-07 $layer=LI1_cond $X=2.44 $Y=1.172
+ $X2=1.785 $Y2=1.172
r149 43 45 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.585 $Y=1.16
+ $X2=1.005 $Y2=1.16
r150 42 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.08 $Y=1.16
+ $X2=1.105 $Y2=1.16
r151 42 45 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.08 $Y=1.16
+ $X2=1.005 $Y2=1.16
r152 38 79 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.875 $Y=1.295
+ $X2=1.875 $Y2=1.16
r153 38 40 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.875 $Y=1.295
+ $X2=1.875 $Y2=1.985
r154 34 79 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.875 $Y=1.025
+ $X2=1.875 $Y2=1.16
r155 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.875 $Y=1.025
+ $X2=1.875 $Y2=0.56
r156 30 77 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.455 $Y=1.295
+ $X2=1.455 $Y2=1.16
r157 30 32 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.455 $Y=1.295
+ $X2=1.455 $Y2=1.985
r158 26 77 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.455 $Y=1.025
+ $X2=1.455 $Y2=1.16
r159 26 28 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.455 $Y=1.025
+ $X2=1.455 $Y2=0.56
r160 22 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.005 $Y=1.295
+ $X2=1.005 $Y2=1.16
r161 22 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.005 $Y=1.295
+ $X2=1.005 $Y2=1.985
r162 18 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.005 $Y=1.025
+ $X2=1.005 $Y2=1.16
r163 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.005 $Y=1.025
+ $X2=1.005 $Y2=0.56
r164 14 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.585 $Y=1.295
+ $X2=0.585 $Y2=1.16
r165 14 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.585 $Y=1.295
+ $X2=0.585 $Y2=1.985
r166 10 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.585 $Y=1.025
+ $X2=0.585 $Y2=1.16
r167 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.585 $Y=1.025
+ $X2=0.585 $Y2=0.56
r168 3 74 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.79
+ $Y=1.485 $X2=3.925 $Y2=2.02
r169 2 62 600 $w=1.7e-07 $l=7.43472e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.485 $X2=2.525 $Y2=2.155
r170 2 59 600 $w=1.7e-07 $l=4.00062e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.485 $X2=2.525 $Y2=1.815
r171 1 65 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.91
+ $Y=0.235 $X2=3.045 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%B1 3 5 6 9 13 17 19 20 21 29 30
c66 30 0 2.33724e-19 $X=3.255 $Y=1.16
c67 29 0 2.66215e-20 $X=3.125 $Y=1.16
r68 32 40 1.96777 $w=3e-07 $l=1.85e-07 $layer=LI1_cond $X=3.15 $Y=1.205
+ $X2=2.965 $Y2=1.205
r69 28 30 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=3.125 $Y=1.16
+ $X2=3.255 $Y2=1.16
r70 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.16 $X2=3.125 $Y2=1.16
r71 26 28 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.835 $Y=1.16
+ $X2=3.125 $Y2=1.16
r72 25 26 22.2174 $w=2.7e-07 $l=1e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=2.835 $Y2=1.16
r73 21 32 10.7561 $w=2.98e-07 $l=2.8e-07 $layer=LI1_cond $X=3.43 $Y=1.205
+ $X2=3.15 $Y2=1.205
r74 20 40 10.1228 $w=3.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=1.53
+ $X2=2.965 $Y2=1.205
r75 19 40 0.467207 $w=3.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.965 $Y=1.19
+ $X2=2.965 $Y2=1.205
r76 19 29 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=2.965 $Y=1.19
+ $X2=2.965 $Y2=1.16
r77 15 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.255 $Y=1.025
+ $X2=3.255 $Y2=1.16
r78 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.255 $Y=1.025
+ $X2=3.255 $Y2=0.56
r79 11 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.835 $Y=1.025
+ $X2=2.835 $Y2=1.16
r80 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.835 $Y=1.025
+ $X2=2.835 $Y2=0.56
r81 7 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.735 $Y=1.295
+ $X2=2.735 $Y2=1.16
r82 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.735 $Y=1.295
+ $X2=2.735 $Y2=1.985
r83 5 25 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.66 $Y=1.16 $X2=2.735
+ $Y2=1.16
r84 5 6 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.66 $Y=1.16 $X2=2.37
+ $Y2=1.16
r85 1 6 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.37 $Y2=1.16
r86 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%A3 3 7 11 15 17 24
c45 24 0 3.82163e-21 $X=4.135 $Y=1.16
c46 17 0 2.0012e-19 $X=3.91 $Y=1.19
c47 3 0 1.24132e-19 $X=3.715 $Y=0.56
r48 22 24 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.135 $Y2=1.16
r49 19 22 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=3.715 $Y=1.16
+ $X2=3.93 $Y2=1.16
r50 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.16 $X2=3.93 $Y2=1.16
r51 13 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.135 $Y=1.295
+ $X2=4.135 $Y2=1.16
r52 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.135 $Y=1.295
+ $X2=4.135 $Y2=1.985
r53 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.135 $Y=1.025
+ $X2=4.135 $Y2=1.16
r54 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.135 $Y=1.025
+ $X2=4.135 $Y2=0.56
r55 5 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.715 $Y=1.295
+ $X2=3.715 $Y2=1.16
r56 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.715 $Y=1.295
+ $X2=3.715 $Y2=1.985
r57 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.715 $Y=1.025
+ $X2=3.715 $Y2=1.16
r58 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.715 $Y=1.025
+ $X2=3.715 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%A2 1 3 6 10 14 18 19 20 21 23 34 37 41 46 56
c89 46 0 5.351e-20 $X=4.825 $Y=1.36
c90 34 0 1.58619e-19 $X=4.555 $Y=1.16
c91 6 0 1.94136e-19 $X=4.555 $Y=1.985
r92 37 40 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.905 $Y=1.16
+ $X2=5.905 $Y2=1.295
r93 37 39 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.905 $Y=1.16
+ $X2=5.905 $Y2=1.025
r94 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.905
+ $Y=1.16 $X2=5.905 $Y2=1.16
r95 35 41 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=4.555 $Y=1.207
+ $X2=4.68 $Y2=1.207
r96 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.555
+ $Y=1.16 $X2=4.555 $Y2=1.16
r97 23 38 5.65587 $w=6.43e-07 $l=3.05e-07 $layer=LI1_cond $X=6.21 $Y=1.377
+ $X2=5.905 $Y2=1.377
r98 21 38 2.8743 $w=6.43e-07 $l=1.55e-07 $layer=LI1_cond $X=5.75 $Y=1.377
+ $X2=5.905 $Y2=1.377
r99 21 56 9.4295 $w=6.43e-07 $l=1.1e-07 $layer=LI1_cond $X=5.75 $Y=1.377
+ $X2=5.64 $Y2=1.377
r100 20 46 5.04691 $w=2.88e-07 $l=1.27e-07 $layer=LI1_cond $X=4.825 $Y=1.487
+ $X2=4.825 $Y2=1.36
r101 19 46 3.50264 $w=2.9e-07 $l=1.53e-07 $layer=LI1_cond $X=4.825 $Y=1.207
+ $X2=4.825 $Y2=1.36
r102 19 41 3.31949 $w=3.05e-07 $l=1.45e-07 $layer=LI1_cond $X=4.825 $Y=1.207
+ $X2=4.68 $Y2=1.207
r103 18 35 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=4.37 $Y=1.207
+ $X2=4.555 $Y2=1.207
r104 17 20 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.97 $Y=1.615
+ $X2=4.825 $Y2=1.615
r105 17 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.97 $Y=1.615
+ $X2=5.64 $Y2=1.615
r106 14 40 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.815 $Y=1.985
+ $X2=5.815 $Y2=1.295
r107 10 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.815 $Y=0.56
+ $X2=5.815 $Y2=1.025
r108 4 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.555 $Y=1.325
+ $X2=4.555 $Y2=1.16
r109 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.555 $Y=1.325
+ $X2=4.555 $Y2=1.985
r110 1 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.555 $Y=0.995
+ $X2=4.555 $Y2=1.16
r111 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.555 $Y=0.995
+ $X2=4.555 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%A1 3 7 11 15 17 24
c52 17 0 1.92011e-19 $X=5.29 $Y=1.19
c53 15 0 5.351e-20 $X=5.395 $Y=1.985
c54 7 0 1.26697e-19 $X=4.975 $Y=1.985
r55 22 24 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.305 $Y=1.16
+ $X2=5.395 $Y2=1.16
r56 19 22 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=4.975 $Y=1.16
+ $X2=5.305 $Y2=1.16
r57 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.305
+ $Y=1.16 $X2=5.305 $Y2=1.16
r58 13 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.395 $Y=1.295
+ $X2=5.395 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.395 $Y=1.295
+ $X2=5.395 $Y2=1.985
r60 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.395 $Y=1.025
+ $X2=5.395 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.395 $Y=1.025
+ $X2=5.395 $Y2=0.56
r62 5 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.975 $Y=1.295
+ $X2=4.975 $Y2=1.16
r63 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.975 $Y=1.295
+ $X2=4.975 $Y2=1.985
r64 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.975 $Y=1.025
+ $X2=4.975 $Y2=1.16
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.975 $Y=1.025
+ $X2=4.975 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%VPWR 1 2 3 4 5 16 18 22 26 32 36 38 40 45 50
+ 55 65 66 72 75 78 81 86
c113 65 0 1.97766e-19 $X=6.21 $Y=2.72
r114 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r115 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r116 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r117 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 69 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r119 66 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.29 $Y2=2.72
r120 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r121 63 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=2.72
+ $X2=5.185 $Y2=2.72
r122 63 65 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.35 $Y=2.72
+ $X2=6.21 $Y2=2.72
r123 62 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r124 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r125 59 62 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r126 59 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r127 58 61 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 56 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=2.72
+ $X2=2.945 $Y2=2.72
r130 56 58 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.11 $Y=2.72
+ $X2=3.45 $Y2=2.72
r131 55 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=2.72
+ $X2=5.185 $Y2=2.72
r132 55 61 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.02 $Y=2.72
+ $X2=4.83 $Y2=2.72
r133 54 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r134 54 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r135 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 51 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.085 $Y2=2.72
r137 51 53 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.53 $Y2=2.72
r138 50 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.945 $Y2=2.72
r139 50 53 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.53 $Y2=2.72
r140 49 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 49 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r142 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r143 46 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.23 $Y2=2.72
r144 46 48 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.61 $Y2=2.72
r145 45 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=2.72
+ $X2=2.085 $Y2=2.72
r146 45 48 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.92 $Y=2.72
+ $X2=1.61 $Y2=2.72
r147 44 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 44 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r149 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r150 41 69 5.73314 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=0.255 $Y2=2.72
r151 41 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=0.69 $Y2=2.72
r152 40 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.23 $Y2=2.72
r153 40 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 38 86 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 34 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.185 $Y=2.635
+ $X2=5.185 $Y2=2.72
r156 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.185 $Y=2.635
+ $X2=5.185 $Y2=2.36
r157 30 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2.72
r158 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2.36
r159 26 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.085 $Y=1.68
+ $X2=2.085 $Y2=2.36
r160 24 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=2.635
+ $X2=2.085 $Y2=2.72
r161 24 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.085 $Y=2.635
+ $X2=2.085 $Y2=2.36
r162 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.72
r163 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.02
r164 16 69 2.85533 $w=4.25e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.297 $Y=2.635
+ $X2=0.255 $Y2=2.72
r165 16 18 17.2189 $w=4.23e-07 $l=6.35e-07 $layer=LI1_cond $X=0.297 $Y=2.635
+ $X2=0.297 $Y2=2
r166 5 36 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=5.05
+ $Y=1.485 $X2=5.185 $Y2=2.36
r167 4 32 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=1.485 $X2=2.945 $Y2=2.36
r168 3 29 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.485 $X2=2.085 $Y2=2.36
r169 3 26 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.485 $X2=2.085 $Y2=1.68
r170 2 22 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.485 $X2=1.23 $Y2=2.02
r171 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.25
+ $Y=1.485 $X2=0.375 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%X 1 2 3 4 15 17 19 21 27 30 31 32 33 44
r48 44 45 0.893119 $w=6.83e-07 $l=5e-08 $layer=LI1_cond $X=0.49 $Y=0.72 $X2=0.49
+ $Y2=0.77
r49 33 55 0.571596 $w=6.83e-07 $l=3.2e-08 $layer=LI1_cond $X=0.49 $Y=1.53
+ $X2=0.49 $Y2=1.562
r50 32 33 6.07321 $w=6.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.49 $Y=1.19
+ $X2=0.49 $Y2=1.53
r51 31 32 6.07321 $w=6.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.49 $Y=0.85
+ $X2=0.49 $Y2=1.19
r52 31 45 1.42899 $w=6.83e-07 $l=8e-08 $layer=LI1_cond $X=0.49 $Y=0.85 $X2=0.49
+ $Y2=0.77
r53 25 27 8.99263 $w=1.83e-07 $l=1.5e-07 $layer=LI1_cond $X=1.657 $Y=1.665
+ $X2=1.657 $Y2=1.815
r54 22 55 7.95557 $w=2.05e-07 $l=4.05e-07 $layer=LI1_cond $X=0.895 $Y=1.562
+ $X2=0.49 $Y2=1.562
r55 21 25 6.83983 $w=2.05e-07 $l=1.41722e-07 $layer=LI1_cond $X=1.565 $Y=1.562
+ $X2=1.657 $Y2=1.665
r56 21 22 36.2483 $w=2.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.562
+ $X2=0.895 $Y2=1.562
r57 20 45 7.21702 $w=2.3e-07 $l=4.05e-07 $layer=LI1_cond $X=0.895 $Y=0.77
+ $X2=0.49 $Y2=0.77
r58 19 30 3.19058 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=1.565 $Y=0.77 $X2=1.665
+ $Y2=0.77
r59 19 20 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=0.77
+ $X2=0.895 $Y2=0.77
r60 15 55 8.07599 $w=6.83e-07 $l=3.44674e-07 $layer=LI1_cond $X=0.787 $Y=1.665
+ $X2=0.49 $Y2=1.562
r61 15 17 8.0403 $w=2.13e-07 $l=1.5e-07 $layer=LI1_cond $X=0.787 $Y=1.665
+ $X2=0.787 $Y2=1.815
r62 4 27 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.485 $X2=1.665 $Y2=1.815
r63 3 17 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=0.66
+ $Y=1.485 $X2=0.795 $Y2=1.815
r64 2 30 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.235 $X2=1.665 $Y2=0.72
r65 1 44 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.235 $X2=0.795 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%A_672_297# 1 2 3 10 15 16 22 23 26
c60 22 0 1.97766e-19 $X=6.21 $Y=2.21
c61 10 0 1.85708e-19 $X=4.26 $Y=1.615
r62 23 30 3.6988 $w=5.93e-07 $l=1.85e-07 $layer=LI1_cond $X=6.21 $Y=2.167
+ $X2=6.025 $Y2=2.167
r63 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.21
+ $X2=6.21 $Y2=2.21
r64 19 26 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=4.385 $Y=2.21
+ $X2=4.385 $Y2=1.815
r65 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.21
+ $X2=4.37 $Y2=2.21
r66 16 18 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=2.21
+ $X2=4.37 $Y2=2.21
r67 15 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.065 $Y=2.21
+ $X2=6.21 $Y2=2.21
r68 15 16 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=6.065 $Y=2.21
+ $X2=4.515 $Y2=2.21
r69 14 26 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.385 $Y=1.7
+ $X2=4.385 $Y2=1.815
r70 10 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.26 $Y=1.615
+ $X2=4.385 $Y2=1.7
r71 10 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.26 $Y=1.615
+ $X2=3.505 $Y2=1.615
r72 3 30 600 $w=1.7e-07 $l=7.34405e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.485 $X2=6.025 $Y2=2.155
r73 2 26 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=4.21
+ $Y=1.485 $X2=4.345 $Y2=1.815
r74 1 12 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.485 $X2=3.505 $Y2=1.615
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%A_926_297# 1 2 9 14 16
c34 14 0 2.55158e-20 $X=4.765 $Y=2.035
r35 10 14 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.85 $Y=1.97 $X2=4.765
+ $Y2=1.97
r36 9 16 3.40825 $w=2e-07 $l=1e-07 $layer=LI1_cond $X=5.52 $Y=1.97 $X2=5.62
+ $Y2=1.97
r37 9 10 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=5.52 $Y=1.97 $X2=4.85
+ $Y2=1.97
r38 2 16 600 $w=1.7e-07 $l=6.138e-07 $layer=licon1_PDIFF $count=1 $X=5.47
+ $Y=1.485 $X2=5.605 $Y2=2.035
r39 1 14 600 $w=1.7e-07 $l=6.138e-07 $layer=licon1_PDIFF $count=1 $X=4.63
+ $Y=1.485 $X2=4.765 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 46 48 53 58 66 76 77 83 86 89 92 97
r111 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r112 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r113 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r114 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r115 80 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r116 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r117 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r118 74 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r119 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r120 71 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=4.765
+ $Y2=0
r121 71 73 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=5.29
+ $Y2=0
r122 70 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r123 70 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r124 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r125 67 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.925
+ $Y2=0
r126 67 69 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.37
+ $Y2=0
r127 66 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.765
+ $Y2=0
r128 66 69 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.37
+ $Y2=0
r129 65 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r130 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r131 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r132 62 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r133 61 64 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r134 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r135 59 86 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.092
+ $Y2=0
r136 59 61 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.53
+ $Y2=0
r137 58 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.925
+ $Y2=0
r138 58 64 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.45
+ $Y2=0
r139 57 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r140 57 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r141 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r142 54 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.23
+ $Y2=0
r143 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.395 $Y=0
+ $X2=1.61 $Y2=0
r144 53 86 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.935 $Y=0
+ $X2=2.092 $Y2=0
r145 53 56 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.935 $Y=0
+ $X2=1.61 $Y2=0
r146 52 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r147 52 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r148 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r149 49 80 5.73314 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r150 49 51 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.69
+ $Y2=0
r151 48 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.23
+ $Y2=0
r152 48 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=0.69 $Y2=0
r153 46 97 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0 $X2=0.23
+ $Y2=0
r154 44 73 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.29
+ $Y2=0
r155 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.605
+ $Y2=0
r156 43 76 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.77 $Y=0 $X2=6.21
+ $Y2=0
r157 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.77 $Y=0 $X2=5.605
+ $Y2=0
r158 39 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=0.085
+ $X2=5.605 $Y2=0
r159 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.605 $Y=0.085
+ $X2=5.605 $Y2=0.36
r160 35 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=0.085
+ $X2=4.765 $Y2=0
r161 35 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.765 $Y=0.085
+ $X2=4.765 $Y2=0.36
r162 31 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r163 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.36
r164 27 86 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.092 $Y=0.085
+ $X2=2.092 $Y2=0
r165 27 29 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=2.092 $Y=0.085
+ $X2=2.092 $Y2=0.38
r166 23 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r167 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.36
r168 19 80 2.85533 $w=4.25e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.297 $Y=0.085
+ $X2=0.255 $Y2=0
r169 19 21 7.99931 $w=4.23e-07 $l=2.95e-07 $layer=LI1_cond $X=0.297 $Y=0.085
+ $X2=0.297 $Y2=0.38
r170 6 41 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.235 $X2=5.605 $Y2=0.36
r171 5 37 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.235 $X2=4.765 $Y2=0.36
r172 4 33 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.79
+ $Y=0.235 $X2=3.925 $Y2=0.36
r173 3 29 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.95
+ $Y=0.235 $X2=2.085 $Y2=0.38
r174 2 25 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.23 $Y2=0.36
r175 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.25
+ $Y=0.235 $X2=0.375 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_4%A_496_47# 1 2 3 4 5 16 24 25 26 29 31 34 36
+ 37 39
r70 35 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=0.76
+ $X2=5.185 $Y2=0.76
r71 34 39 5.55394 $w=4.13e-07 $l=2e-07 $layer=LI1_cond $X=6.147 $Y=0.76
+ $X2=6.147 $Y2=0.56
r72 34 35 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.94 $Y=0.76
+ $X2=5.27 $Y2=0.76
r73 31 37 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=0.635
+ $X2=5.185 $Y2=0.76
r74 31 33 5.38235 $w=1.7e-07 $l=7.5e-08 $layer=LI1_cond $X=5.185 $Y=0.635
+ $X2=5.185 $Y2=0.56
r75 30 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.43 $Y=0.76
+ $X2=4.345 $Y2=0.76
r76 29 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=0.76 $X2=5.185
+ $Y2=0.76
r77 29 30 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.1 $Y=0.76 $X2=4.43
+ $Y2=0.76
r78 26 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.345 $Y=0.635
+ $X2=4.345 $Y2=0.76
r79 26 28 5.38235 $w=1.7e-07 $l=7.5e-08 $layer=LI1_cond $X=4.345 $Y=0.635
+ $X2=4.345 $Y2=0.56
r80 24 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=0.76
+ $X2=4.345 $Y2=0.76
r81 24 25 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=4.26 $Y=0.76
+ $X2=3.57 $Y2=0.76
r82 21 25 6.98266 $w=2.5e-07 $l=1.65831e-07 $layer=LI1_cond $X=3.475 $Y=0.635
+ $X2=3.57 $Y2=0.76
r83 21 23 4.37799 $w=1.88e-07 $l=7.5e-08 $layer=LI1_cond $X=3.475 $Y=0.635
+ $X2=3.475 $Y2=0.56
r84 20 23 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=3.475 $Y=0.465
+ $X2=3.475 $Y2=0.56
r85 16 20 6.83868 $w=2.1e-07 $l=1.44914e-07 $layer=LI1_cond $X=3.38 $Y=0.36
+ $X2=3.475 $Y2=0.465
r86 16 18 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.38 $Y=0.36
+ $X2=2.625 $Y2=0.36
r87 5 39 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.235 $X2=6.025 $Y2=0.56
r88 4 33 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.235 $X2=5.185 $Y2=0.56
r89 3 28 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.21
+ $Y=0.235 $X2=4.345 $Y2=0.56
r90 2 23 182 $w=1.7e-07 $l=3.90832e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.235 $X2=3.475 $Y2=0.56
r91 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.625 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__o22ai_1.spice
* Created: Thu Aug 27 14:37:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o22ai_1.pex.spice"
.subckt sky130_fd_sc_hd__o22ai_1  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_27_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.169 PD=0.935 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_B2_M1005_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.092625 PD=1.005 PS=0.935 NRD=11.076 NRS=1.836 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_27_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.115375 PD=0.92 PS=1.005 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_47#_M1002_d N_A1_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 A_109_297# N_B1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.1125
+ AS=0.26 PD=1.225 PS=2.52 NRD=11.3078 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1003_d N_B2_M1003_g A_109_297# VPB PHIGHVT L=0.15 W=1 AD=0.2325
+ AS=0.1125 PD=1.465 PS=1.225 NRD=0 NRS=11.3078 M=1 R=6.66667 SA=75000.6
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 A_307_297# N_A2_M1000_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.2325 PD=1.21 PS=1.465 NRD=9.8303 NRS=37.4103 M=1 R=6.66667 SA=75001.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_307_297# VPB PHIGHVT L=0.15 W=1 AD=0.27
+ AS=0.105 PD=2.54 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__o22ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a31oi_4.spice.SKY130_FD_SC_HD__A31OI_4.pxi
* Created: Thu Aug 27 14:05:11 2020
* 
x_PM_SKY130_FD_SC_HD__A31OI_4%A3 N_A3_c_86_n N_A3_M1012_g N_A3_M1002_g
+ N_A3_c_87_n N_A3_M1015_g N_A3_M1005_g N_A3_c_88_n N_A3_M1019_g N_A3_M1020_g
+ N_A3_c_89_n N_A3_M1030_g N_A3_M1028_g A3 A3 A3 A3 N_A3_c_90_n
+ PM_SKY130_FD_SC_HD__A31OI_4%A3
x_PM_SKY130_FD_SC_HD__A31OI_4%A2 N_A2_c_155_n N_A2_M1016_g N_A2_M1000_g
+ N_A2_c_156_n N_A2_M1022_g N_A2_M1006_g N_A2_c_157_n N_A2_M1026_g N_A2_M1024_g
+ N_A2_c_158_n N_A2_M1027_g N_A2_M1029_g A2 A2 A2 A2 N_A2_c_160_n
+ PM_SKY130_FD_SC_HD__A31OI_4%A2
x_PM_SKY130_FD_SC_HD__A31OI_4%A1 N_A1_M1004_g N_A1_M1009_g N_A1_c_226_n
+ N_A1_M1010_g N_A1_M1021_g N_A1_c_227_n N_A1_M1013_g N_A1_M1031_g N_A1_c_228_n
+ N_A1_M1017_g N_A1_c_229_n N_A1_M1023_g A1 A1 A1 A1 N_A1_c_231_n
+ PM_SKY130_FD_SC_HD__A31OI_4%A1
x_PM_SKY130_FD_SC_HD__A31OI_4%B1 N_B1_c_296_n N_B1_M1008_g N_B1_M1001_g
+ N_B1_c_297_n N_B1_M1011_g N_B1_M1003_g N_B1_c_298_n N_B1_M1014_g N_B1_M1007_g
+ N_B1_c_299_n N_B1_M1018_g N_B1_M1025_g B1 B1 B1 N_B1_c_300_n N_B1_c_301_n
+ PM_SKY130_FD_SC_HD__A31OI_4%B1
x_PM_SKY130_FD_SC_HD__A31OI_4%A_27_297# N_A_27_297#_M1002_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1028_s N_A_27_297#_M1006_s N_A_27_297#_M1029_s
+ N_A_27_297#_M1009_d N_A_27_297#_M1031_d N_A_27_297#_M1003_s
+ N_A_27_297#_M1025_s N_A_27_297#_c_435_p N_A_27_297#_c_372_n
+ N_A_27_297#_c_376_n N_A_27_297#_c_432_p N_A_27_297#_c_378_n
+ N_A_27_297#_c_433_p N_A_27_297#_c_384_n N_A_27_297#_c_434_p
+ N_A_27_297#_c_388_n N_A_27_297#_c_396_n N_A_27_297#_c_397_n
+ N_A_27_297#_c_436_p N_A_27_297#_c_401_n N_A_27_297#_c_411_n
+ N_A_27_297#_c_412_n N_A_27_297#_c_417_n N_A_27_297#_c_439_p
+ N_A_27_297#_c_382_n N_A_27_297#_c_392_n N_A_27_297#_c_393_n
+ N_A_27_297#_c_395_n N_A_27_297#_c_405_n PM_SKY130_FD_SC_HD__A31OI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A31OI_4%VPWR N_VPWR_M1002_d N_VPWR_M1020_d N_VPWR_M1000_d
+ N_VPWR_M1024_d N_VPWR_M1004_s N_VPWR_M1021_s N_VPWR_c_465_n N_VPWR_c_466_n
+ N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n
+ N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n
+ N_VPWR_c_477_n VPWR N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n
+ N_VPWR_c_464_n N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n
+ PM_SKY130_FD_SC_HD__A31OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A31OI_4%Y N_Y_M1010_s N_Y_M1013_s N_Y_M1023_s N_Y_M1011_s
+ N_Y_M1018_s N_Y_M1001_d N_Y_M1007_d N_Y_c_581_n N_Y_c_595_n N_Y_c_631_p
+ N_Y_c_600_n N_Y_c_633_p N_Y_c_603_n Y Y Y Y N_Y_c_605_n Y Y N_Y_c_612_n
+ PM_SKY130_FD_SC_HD__A31OI_4%Y
x_PM_SKY130_FD_SC_HD__A31OI_4%A_27_47# N_A_27_47#_M1012_d N_A_27_47#_M1015_d
+ N_A_27_47#_M1030_d N_A_27_47#_M1022_s N_A_27_47#_M1027_s N_A_27_47#_c_676_p
+ N_A_27_47#_c_651_n N_A_27_47#_c_655_n N_A_27_47#_c_679_p N_A_27_47#_c_657_n
+ N_A_27_47#_c_682_p N_A_27_47#_c_650_n N_A_27_47#_c_661_n N_A_27_47#_c_669_n
+ PM_SKY130_FD_SC_HD__A31OI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__A31OI_4%VGND N_VGND_M1012_s N_VGND_M1019_s N_VGND_M1008_d
+ N_VGND_M1014_d N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n
+ VGND N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n
+ N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n
+ N_VGND_c_713_n PM_SKY130_FD_SC_HD__A31OI_4%VGND
x_PM_SKY130_FD_SC_HD__A31OI_4%A_445_47# N_A_445_47#_M1016_d N_A_445_47#_M1026_d
+ N_A_445_47#_M1010_d N_A_445_47#_M1017_d N_A_445_47#_c_812_n
+ PM_SKY130_FD_SC_HD__A31OI_4%A_445_47#
cc_1 VNB N_A3_c_86_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A3_c_87_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A3_c_88_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A3_c_89_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A3_c_90_n 0.0941763f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_6 VNB N_A2_c_155_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_7 VNB N_A2_c_156_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_8 VNB N_A2_c_157_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_9 VNB N_A2_c_158_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_10 VNB A2 0.00622401f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_11 VNB N_A2_c_160_n 0.0612088f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_12 VNB N_A1_c_226_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_13 VNB N_A1_c_227_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_14 VNB N_A1_c_228_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_15 VNB N_A1_c_229_n 0.0168748f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_16 VNB A1 0.00159174f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_17 VNB N_A1_c_231_n 0.093262f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_18 VNB N_B1_c_296_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_19 VNB N_B1_c_297_n 0.0157748f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_20 VNB N_B1_c_298_n 0.0157484f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_21 VNB N_B1_c_299_n 0.0212813f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_22 VNB N_B1_c_300_n 0.00205078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B1_c_301_n 0.0770291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_464_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_581_n 0.00209549f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_26 VNB Y 0.00103535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_650_n 0.00297253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_700_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_29 VNB N_VGND_c_701_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_30 VNB N_VGND_c_702_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_31 VNB N_VGND_c_703_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_32 VNB N_VGND_c_704_n 0.0151407f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_33 VNB N_VGND_c_705_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_706_n 0.102905f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_35 VNB N_VGND_c_707_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.16
cc_36 VNB N_VGND_c_708_n 0.0170455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_709_n 0.376687f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.16
cc_38 VNB N_VGND_c_710_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.16
cc_39 VNB N_VGND_c_711_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_712_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_713_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_445_47#_c_812_n 0.00657894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_A3_M1002_g 0.025757f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_A3_M1005_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_45 VPB N_A3_M1020_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_46 VPB N_A3_M1028_g 0.0186099f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_47 VPB N_A3_c_90_n 0.0202265f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_48 VPB N_A2_M1000_g 0.0186099f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_49 VPB N_A2_M1006_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_50 VPB N_A2_M1024_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_51 VPB N_A2_M1029_g 0.0188354f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_52 VPB A2 0.00216413f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_53 VPB N_A2_c_160_n 0.0100219f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_54 VPB N_A1_M1004_g 0.017785f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_55 VPB N_A1_M1009_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A1_M1021_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A1_M1031_g 0.0214914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A1_c_231_n 0.03603f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_59 VPB N_B1_M1001_g 0.0223275f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_60 VPB N_B1_M1003_g 0.0171325f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_61 VPB N_B1_M1007_g 0.0177777f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_62 VPB N_B1_M1025_g 0.0253019f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_63 VPB N_B1_c_300_n 0.00239848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_B1_c_301_n 0.0138634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_465_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_466_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_67 VPB N_VPWR_c_467_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_68 VPB N_VPWR_c_468_n 3.05427e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_469_n 0.0131279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_470_n 3.05427e-19 $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_71 VPB N_VPWR_c_471_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_72 VPB N_VPWR_c_472_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_73 VPB N_VPWR_c_473_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_74 VPB N_VPWR_c_474_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_75 VPB N_VPWR_c_475_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_476_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_477_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_78 VPB N_VPWR_c_478_n 0.0159043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_479_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_480_n 0.0675386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_464_n 0.0480238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_482_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_483_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_484_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB Y 9.69295e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 N_A3_c_89_n N_A2_c_155_n 0.022884f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_87 N_A3_M1028_g N_A2_M1000_g 0.022884f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_88 A3 A2 0.0258519f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A3_c_90_n A2 0.00289706f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_90 A3 N_A2_c_160_n 2.92893e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_91 N_A3_c_90_n N_A2_c_160_n 0.022884f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A3_M1002_g N_A_27_297#_c_372_n 0.015361f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A3_M1005_g N_A_27_297#_c_372_n 0.0141087f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_94 A3 N_A_27_297#_c_372_n 0.0409723f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A3_c_90_n N_A_27_297#_c_372_n 0.00201785f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_96 A3 N_A_27_297#_c_376_n 0.0137245f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A3_c_90_n N_A_27_297#_c_376_n 0.00393893f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A3_M1020_g N_A_27_297#_c_378_n 0.0141528f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A3_M1028_g N_A_27_297#_c_378_n 0.0162466f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_100 A3 N_A_27_297#_c_378_n 0.0340973f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A3_c_90_n N_A_27_297#_c_378_n 0.00201785f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_102 A3 N_A_27_297#_c_382_n 0.0134105f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A3_c_90_n N_A_27_297#_c_382_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A3_M1002_g N_VPWR_c_465_n 0.012183f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A3_M1005_g N_VPWR_c_465_n 0.0102874f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A3_M1020_g N_VPWR_c_465_n 6.0901e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A3_M1005_g N_VPWR_c_466_n 6.0901e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A3_M1020_g N_VPWR_c_466_n 0.0102874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A3_M1028_g N_VPWR_c_466_n 0.0102874f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A3_M1028_g N_VPWR_c_467_n 6.0901e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A3_M1005_g N_VPWR_c_472_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A3_M1020_g N_VPWR_c_472_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A3_M1028_g N_VPWR_c_474_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A3_M1002_g N_VPWR_c_478_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A3_M1002_g N_VPWR_c_464_n 0.008846f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A3_M1005_g N_VPWR_c_464_n 0.00789179f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A3_M1020_g N_VPWR_c_464_n 0.00789179f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A3_M1028_g N_VPWR_c_464_n 0.007919f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A3_c_86_n N_A_27_47#_c_651_n 0.0127817f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A3_c_87_n N_A_27_47#_c_651_n 0.0115294f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_121 A3 N_A_27_47#_c_651_n 0.0375135f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A3_c_90_n N_A_27_47#_c_651_n 0.0019918f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_123 A3 N_A_27_47#_c_655_n 0.0123848f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A3_c_90_n N_A_27_47#_c_655_n 0.00386661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A3_c_88_n N_A_27_47#_c_657_n 0.0115735f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A3_c_89_n N_A_27_47#_c_657_n 0.0136104f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_127 A3 N_A_27_47#_c_657_n 0.0312246f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A3_c_90_n N_A_27_47#_c_657_n 0.0019918f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_129 A3 N_A_27_47#_c_661_n 0.0121035f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A3_c_90_n N_A_27_47#_c_661_n 0.00205824f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A3_c_86_n N_VGND_c_700_n 0.00834749f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A3_c_87_n N_VGND_c_700_n 0.00664421f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A3_c_88_n N_VGND_c_700_n 5.08801e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A3_c_87_n N_VGND_c_701_n 5.08801e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A3_c_88_n N_VGND_c_701_n 0.00664421f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A3_c_89_n N_VGND_c_701_n 0.00784221f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A3_c_86_n N_VGND_c_704_n 0.00339367f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A3_c_87_n N_VGND_c_705_n 0.00339367f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A3_c_88_n N_VGND_c_705_n 0.00339367f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A3_c_89_n N_VGND_c_706_n 0.00339367f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A3_c_86_n N_VGND_c_709_n 0.00489827f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A3_c_87_n N_VGND_c_709_n 0.00394406f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A3_c_88_n N_VGND_c_709_n 0.00394406f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A3_c_89_n N_VGND_c_709_n 0.00397127f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A2_M1029_g N_A1_M1004_g 0.0200133f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_146 A2 A1 0.0203714f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A2_c_160_n A1 3.47199e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_148 A2 N_A1_c_231_n 0.00284587f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A2_c_160_n N_A1_c_231_n 0.0200133f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_M1000_g N_A_27_297#_c_384_n 0.0141087f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_M1006_g N_A_27_297#_c_384_n 0.0141528f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_152 A2 N_A_27_297#_c_384_n 0.0411779f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A2_c_160_n N_A_27_297#_c_384_n 0.00201785f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_M1024_g N_A_27_297#_c_388_n 0.0141528f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A2_M1029_g N_A_27_297#_c_388_n 0.0142272f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_156 A2 N_A_27_297#_c_388_n 0.0411779f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A2_c_160_n N_A_27_297#_c_388_n 0.00201785f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_158 A2 N_A_27_297#_c_392_n 0.007488f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_159 A2 N_A_27_297#_c_393_n 0.0134105f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A2_c_160_n N_A_27_297#_c_393_n 0.00209661f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_161 A2 N_A_27_297#_c_395_n 9.86189e-19 $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A2_M1000_g N_VPWR_c_466_n 6.0901e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_VPWR_c_467_n 0.0102874f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_M1006_g N_VPWR_c_467_n 0.0102874f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A2_M1024_g N_VPWR_c_467_n 6.0901e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A2_M1006_g N_VPWR_c_468_n 6.0901e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A2_M1024_g N_VPWR_c_468_n 0.0102874f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A2_M1029_g N_VPWR_c_468_n 0.0103558f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A2_M1029_g N_VPWR_c_469_n 0.0046653f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A2_M1029_g N_VPWR_c_470_n 6.15726e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A2_M1000_g N_VPWR_c_474_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A2_M1006_g N_VPWR_c_476_n 0.0046653f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_M1024_g N_VPWR_c_476_n 0.0046653f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A2_M1000_g N_VPWR_c_464_n 0.007919f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A2_M1006_g N_VPWR_c_464_n 0.00789179f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A2_M1024_g N_VPWR_c_464_n 0.00789179f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1029_g N_VPWR_c_464_n 0.00796757f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_c_155_n N_A_27_47#_c_650_n 0.011544f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A2_c_156_n N_A_27_47#_c_650_n 0.00847802f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_157_n N_A_27_47#_c_650_n 0.00847802f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A2_c_158_n N_A_27_47#_c_650_n 0.00847802f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_182 A2 N_A_27_47#_c_650_n 0.0872482f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_183 N_A2_c_160_n N_A_27_47#_c_650_n 0.00597539f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_184 A2 N_A_27_47#_c_669_n 0.00680018f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_185 N_A2_c_155_n N_VGND_c_701_n 0.00116167f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A2_c_155_n N_VGND_c_706_n 0.00413298f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A2_c_156_n N_VGND_c_706_n 0.00366111f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A2_c_157_n N_VGND_c_706_n 0.00366111f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A2_c_158_n N_VGND_c_706_n 0.00366111f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_c_155_n N_VGND_c_709_n 0.00570263f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_c_156_n N_VGND_c_709_n 0.00524008f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_157_n N_VGND_c_709_n 0.00524008f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_158_n N_VGND_c_709_n 0.00661716f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_155_n N_A_445_47#_c_812_n 0.00245853f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_156_n N_A_445_47#_c_812_n 0.00789149f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_157_n N_A_445_47#_c_812_n 0.00789149f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_158_n N_A_445_47#_c_812_n 0.00999448f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_229_n N_B1_c_296_n 0.025737f $X=5.61 $Y=1.01 $X2=-0.19 $Y2=-0.24
cc_199 N_A1_M1031_g N_B1_c_300_n 6.01317e-19 $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A1_c_229_n N_B1_c_300_n 4.75953e-19 $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_201 A1 N_B1_c_300_n 0.0203741f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A1_c_231_n N_B1_c_300_n 0.0143656f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_203 N_A1_c_229_n N_B1_c_301_n 0.0215549f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_204 N_A1_M1004_g N_A_27_297#_c_396_n 0.00687412f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A1_M1004_g N_A_27_297#_c_397_n 0.0156314f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A1_M1009_g N_A_27_297#_c_397_n 0.0141528f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_207 A1 N_A_27_297#_c_397_n 0.0355255f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A1_c_231_n N_A_27_297#_c_397_n 0.00209089f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_209 N_A1_M1021_g N_A_27_297#_c_401_n 0.0144059f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A1_M1031_g N_A_27_297#_c_401_n 0.0145014f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_211 A1 N_A_27_297#_c_401_n 0.0546968f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_212 N_A1_c_231_n N_A_27_297#_c_401_n 0.00679219f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_213 A1 N_A_27_297#_c_405_n 0.0134105f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_214 N_A1_c_231_n N_A_27_297#_c_405_n 0.00247295f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_215 N_A1_M1004_g N_VPWR_c_468_n 5.98943e-19 $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A1_M1004_g N_VPWR_c_469_n 0.0046653f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A1_M1004_g N_VPWR_c_470_n 0.0106094f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A1_M1009_g N_VPWR_c_470_n 0.0102874f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A1_M1021_g N_VPWR_c_470_n 6.0901e-19 $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A1_M1009_g N_VPWR_c_471_n 5.08801e-19 $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A1_M1021_g N_VPWR_c_471_n 0.00704125f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A1_M1031_g N_VPWR_c_471_n 0.00873912f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A1_M1009_g N_VPWR_c_479_n 0.0046653f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A1_M1021_g N_VPWR_c_479_n 0.0046653f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A1_M1031_g N_VPWR_c_480_n 0.0046653f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A1_M1004_g N_VPWR_c_464_n 0.00796757f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A1_M1009_g N_VPWR_c_464_n 0.00789179f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A1_M1021_g N_VPWR_c_464_n 0.00789179f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A1_M1031_g N_VPWR_c_464_n 0.00921786f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_c_226_n N_Y_c_581_n 0.00847802f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A1_c_227_n N_Y_c_581_n 0.00847802f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A1_c_228_n N_Y_c_581_n 0.00847802f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A1_c_229_n N_Y_c_581_n 0.0132923f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_234 A1 N_Y_c_581_n 0.0859922f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_235 N_A1_c_231_n N_Y_c_581_n 0.0132757f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_236 N_A1_c_231_n N_A_27_47#_c_650_n 4.06203e-19 $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_237 N_A1_c_229_n N_VGND_c_702_n 0.0018398f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_238 N_A1_c_226_n N_VGND_c_706_n 0.00366111f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A1_c_227_n N_VGND_c_706_n 0.00366111f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A1_c_228_n N_VGND_c_706_n 0.00366111f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A1_c_229_n N_VGND_c_706_n 0.00413298f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_242 N_A1_c_226_n N_VGND_c_709_n 0.00661716f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A1_c_227_n N_VGND_c_709_n 0.00524008f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A1_c_228_n N_VGND_c_709_n 0.00524008f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A1_c_229_n N_VGND_c_709_n 0.00574665f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_246 N_A1_c_226_n N_A_445_47#_c_812_n 0.00999448f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A1_c_227_n N_A_445_47#_c_812_n 0.00789149f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A1_c_228_n N_A_445_47#_c_812_n 0.00789149f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A1_c_229_n N_A_445_47#_c_812_n 0.00363095f $X=5.61 $Y=1.01 $X2=0 $Y2=0
cc_250 A1 N_A_445_47#_c_812_n 0.00478545f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_251 N_A1_c_231_n N_A_445_47#_c_812_n 0.0043895f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_252 N_B1_c_300_n N_A_27_297#_M1031_d 0.00733107f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_253 N_B1_c_300_n N_A_27_297#_M1003_s 0.00219451f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_M1001_g N_A_27_297#_c_401_n 0.00158952f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B1_c_300_n N_A_27_297#_c_401_n 0.00868456f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_M1001_g N_A_27_297#_c_411_n 0.0122312f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B1_M1001_g N_A_27_297#_c_412_n 0.013681f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B1_M1003_g N_A_27_297#_c_412_n 0.00789149f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_259 N_B1_M1007_g N_A_27_297#_c_412_n 0.00789149f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B1_M1025_g N_A_27_297#_c_412_n 0.011511f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B1_c_300_n N_A_27_297#_c_412_n 0.00998857f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_262 N_B1_M1001_g N_A_27_297#_c_417_n 9.23417e-19 $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_263 N_B1_M1001_g N_VPWR_c_480_n 0.00366111f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B1_M1003_g N_VPWR_c_480_n 0.00366111f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B1_M1007_g N_VPWR_c_480_n 0.00366111f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B1_M1025_g N_VPWR_c_480_n 0.00366111f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_267 N_B1_M1001_g N_VPWR_c_464_n 0.00665614f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B1_M1003_g N_VPWR_c_464_n 0.00524008f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B1_M1007_g N_VPWR_c_464_n 0.00524008f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B1_M1025_g N_VPWR_c_464_n 0.0062471f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B1_c_300_n N_Y_M1001_d 0.00219451f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_296_n N_Y_c_581_n 0.00957617f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_273 N_B1_c_297_n N_Y_c_581_n 0.0115735f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B1_c_300_n N_Y_c_581_n 0.0554268f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_275 N_B1_c_301_n N_Y_c_581_n 0.0031865f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B1_M1001_g N_Y_c_595_n 0.004739f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B1_M1003_g N_Y_c_595_n 0.00901269f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1007_g N_Y_c_595_n 0.0113392f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_c_300_n N_Y_c_595_n 0.0291039f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B1_c_301_n N_Y_c_595_n 8.8259e-19 $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_281 N_B1_c_298_n N_Y_c_600_n 0.0142049f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B1_c_300_n N_Y_c_600_n 0.00603295f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_283 N_B1_c_301_n N_Y_c_600_n 3.8744e-19 $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_284 N_B1_c_300_n N_Y_c_603_n 0.0127201f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B1_c_301_n N_Y_c_603_n 0.00205824f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B1_M1025_g N_Y_c_605_n 0.0022776f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_287 N_B1_c_298_n Y 0.00439308f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B1_M1007_g Y 0.00819555f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_289 N_B1_c_299_n Y 0.0093788f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B1_M1025_g Y 0.0153087f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_291 N_B1_c_300_n Y 0.0455217f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_301_n Y 0.0271196f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_293 N_B1_c_299_n N_Y_c_612_n 0.0160497f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B1_c_301_n N_Y_c_612_n 3.61072e-19 $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_295 N_B1_c_296_n N_VGND_c_702_n 0.0093418f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B1_c_297_n N_VGND_c_702_n 0.00664421f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B1_c_298_n N_VGND_c_702_n 5.08801e-19 $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_298 N_B1_c_297_n N_VGND_c_703_n 5.08801e-19 $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_298_n N_VGND_c_703_n 0.00664421f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B1_c_299_n N_VGND_c_703_n 0.00834749f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B1_c_296_n N_VGND_c_706_n 0.00339367f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B1_c_297_n N_VGND_c_707_n 0.00339367f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B1_c_298_n N_VGND_c_707_n 0.00339367f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B1_c_299_n N_VGND_c_708_n 0.00339367f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B1_c_296_n N_VGND_c_709_n 0.00401529f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B1_c_297_n N_VGND_c_709_n 0.00394406f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_c_298_n N_VGND_c_709_n 0.00394406f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_308 N_B1_c_299_n N_VGND_c_709_n 0.00495108f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B1_c_296_n N_A_445_47#_c_812_n 4.913e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A_27_297#_c_372_n N_VPWR_M1002_d 0.00342716f $X=1.015 $Y=1.58 $X2=0.47
+ $Y2=0.995
cc_311 N_A_27_297#_c_378_n N_VPWR_M1020_d 0.00342716f $X=1.855 $Y=1.58 $X2=0.47
+ $Y2=0.56
cc_312 N_A_27_297#_c_384_n N_VPWR_M1000_d 0.00342716f $X=2.695 $Y=1.58 $X2=0.47
+ $Y2=0.56
cc_313 N_A_27_297#_c_388_n N_VPWR_M1024_d 0.00342716f $X=3.535 $Y=1.58 $X2=0.47
+ $Y2=1.325
cc_314 N_A_27_297#_c_397_n N_VPWR_M1004_s 0.0034223f $X=4.395 $Y=1.58 $X2=0.47
+ $Y2=1.985
cc_315 N_A_27_297#_c_401_n N_VPWR_M1021_s 0.00452688f $X=5.235 $Y=1.58 $X2=0.47
+ $Y2=1.985
cc_316 N_A_27_297#_c_372_n N_VPWR_c_465_n 0.0127176f $X=1.015 $Y=1.58 $X2=0
+ $Y2=0
cc_317 N_A_27_297#_c_378_n N_VPWR_c_466_n 0.0127176f $X=1.855 $Y=1.58 $X2=1.73
+ $Y2=1.325
cc_318 N_A_27_297#_c_384_n N_VPWR_c_467_n 0.0127176f $X=2.695 $Y=1.58 $X2=0.15
+ $Y2=1.105
cc_319 N_A_27_297#_c_388_n N_VPWR_c_468_n 0.0127176f $X=3.535 $Y=1.58 $X2=0
+ $Y2=0
cc_320 N_A_27_297#_c_396_n N_VPWR_c_469_n 0.0116048f $X=3.62 $Y=1.96 $X2=0 $Y2=0
cc_321 N_A_27_297#_c_396_n N_VPWR_c_470_n 0.0372674f $X=3.62 $Y=1.96 $X2=0.285
+ $Y2=1.16
cc_322 N_A_27_297#_c_397_n N_VPWR_c_470_n 0.0127176f $X=4.395 $Y=1.58 $X2=0.285
+ $Y2=1.16
cc_323 N_A_27_297#_c_401_n N_VPWR_c_471_n 0.00643049f $X=5.235 $Y=1.58 $X2=1.31
+ $Y2=1.16
cc_324 N_A_27_297#_c_432_p N_VPWR_c_472_n 0.0113958f $X=1.1 $Y=1.96 $X2=1.395
+ $Y2=1.16
cc_325 N_A_27_297#_c_433_p N_VPWR_c_474_n 0.0113958f $X=1.94 $Y=1.96 $X2=0.235
+ $Y2=1.16
cc_326 N_A_27_297#_c_434_p N_VPWR_c_476_n 0.0113958f $X=2.78 $Y=1.96 $X2=0 $Y2=0
cc_327 N_A_27_297#_c_435_p N_VPWR_c_478_n 0.0116048f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_328 N_A_27_297#_c_436_p N_VPWR_c_479_n 0.0113958f $X=4.48 $Y=1.96 $X2=0 $Y2=0
cc_329 N_A_27_297#_c_412_n N_VPWR_c_480_n 0.0906729f $X=7.415 $Y=2.34 $X2=0
+ $Y2=0
cc_330 N_A_27_297#_c_417_n N_VPWR_c_480_n 0.0117106f $X=5.405 $Y=2.34 $X2=0
+ $Y2=0
cc_331 N_A_27_297#_c_439_p N_VPWR_c_480_n 0.0137847f $X=7.54 $Y=2.255 $X2=0
+ $Y2=0
cc_332 N_A_27_297#_M1002_s N_VPWR_c_464_n 0.00525232f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_333 N_A_27_297#_M1005_s N_VPWR_c_464_n 0.00562358f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_334 N_A_27_297#_M1028_s N_VPWR_c_464_n 0.00562358f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_335 N_A_27_297#_M1006_s N_VPWR_c_464_n 0.00562358f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_336 N_A_27_297#_M1029_s N_VPWR_c_464_n 0.00647849f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_337 N_A_27_297#_M1009_d N_VPWR_c_464_n 0.00562358f $X=4.345 $Y=1.485 $X2=0
+ $Y2=0
cc_338 N_A_27_297#_M1031_d N_VPWR_c_464_n 0.00799453f $X=5.185 $Y=1.485 $X2=0
+ $Y2=0
cc_339 N_A_27_297#_M1003_s N_VPWR_c_464_n 0.00217615f $X=6.525 $Y=1.485 $X2=0
+ $Y2=0
cc_340 N_A_27_297#_M1025_s N_VPWR_c_464_n 0.00330547f $X=7.365 $Y=1.485 $X2=0
+ $Y2=0
cc_341 N_A_27_297#_c_435_p N_VPWR_c_464_n 0.00646998f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_342 N_A_27_297#_c_432_p N_VPWR_c_464_n 0.00646998f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_343 N_A_27_297#_c_433_p N_VPWR_c_464_n 0.00646998f $X=1.94 $Y=1.96 $X2=0
+ $Y2=0
cc_344 N_A_27_297#_c_434_p N_VPWR_c_464_n 0.00646998f $X=2.78 $Y=1.96 $X2=0
+ $Y2=0
cc_345 N_A_27_297#_c_396_n N_VPWR_c_464_n 0.00646998f $X=3.62 $Y=1.96 $X2=0
+ $Y2=0
cc_346 N_A_27_297#_c_436_p N_VPWR_c_464_n 0.00646998f $X=4.48 $Y=1.96 $X2=0
+ $Y2=0
cc_347 N_A_27_297#_c_412_n N_VPWR_c_464_n 0.0700398f $X=7.415 $Y=2.34 $X2=0
+ $Y2=0
cc_348 N_A_27_297#_c_417_n N_VPWR_c_464_n 0.006547f $X=5.405 $Y=2.34 $X2=0 $Y2=0
cc_349 N_A_27_297#_c_439_p N_VPWR_c_464_n 0.00943767f $X=7.54 $Y=2.255 $X2=0
+ $Y2=0
cc_350 N_A_27_297#_c_412_n N_Y_M1001_d 0.00325828f $X=7.415 $Y=2.34 $X2=0.47
+ $Y2=1.985
cc_351 N_A_27_297#_c_412_n N_Y_M1007_d 0.00324473f $X=7.415 $Y=2.34 $X2=0 $Y2=0
cc_352 N_A_27_297#_M1003_s N_Y_c_595_n 0.00357959f $X=6.525 $Y=1.485 $X2=0.61
+ $Y2=1.105
cc_353 N_A_27_297#_c_411_n N_Y_c_595_n 0.00441371f $X=5.32 $Y=1.8 $X2=0.61
+ $Y2=1.105
cc_354 N_A_27_297#_c_412_n N_Y_c_595_n 0.0455049f $X=7.415 $Y=2.34 $X2=0.61
+ $Y2=1.105
cc_355 N_A_27_297#_c_412_n N_Y_c_605_n 0.0107229f $X=7.415 $Y=2.34 $X2=1.395
+ $Y2=1.16
cc_356 N_VPWR_c_464_n N_Y_M1001_d 0.00219239f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_357 N_VPWR_c_464_n N_Y_M1007_d 0.00219239f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_358 N_Y_c_581_n N_A_27_47#_c_650_n 0.0145425f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_359 N_Y_c_581_n N_VGND_M1008_d 0.00312394f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_360 N_Y_c_600_n N_VGND_M1014_d 0.00179449f $X=7.045 $Y=0.72 $X2=0 $Y2=0
cc_361 Y N_VGND_M1014_d 0.00123872f $X=7.155 $Y=0.85 $X2=0 $Y2=0
cc_362 N_Y_c_612_n N_VGND_M1014_d 0.00144537f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_363 N_Y_c_581_n N_VGND_c_702_n 0.0159625f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_364 N_Y_c_600_n N_VGND_c_703_n 0.0159297f $X=7.045 $Y=0.72 $X2=0 $Y2=0
cc_365 N_Y_c_581_n N_VGND_c_706_n 0.00775032f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_366 N_Y_c_581_n N_VGND_c_707_n 0.00244309f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_367 N_Y_c_631_p N_VGND_c_707_n 0.0112274f $X=6.66 $Y=0.42 $X2=0 $Y2=0
cc_368 N_Y_c_600_n N_VGND_c_707_n 0.00244309f $X=7.045 $Y=0.72 $X2=0 $Y2=0
cc_369 N_Y_c_633_p N_VGND_c_708_n 0.0111381f $X=7.5 $Y=0.42 $X2=0 $Y2=0
cc_370 N_Y_c_612_n N_VGND_c_708_n 0.00247038f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_371 N_Y_M1010_s N_VGND_c_709_n 0.00212464f $X=4.015 $Y=0.235 $X2=0 $Y2=0
cc_372 N_Y_M1013_s N_VGND_c_709_n 0.00219239f $X=4.845 $Y=0.235 $X2=0 $Y2=0
cc_373 N_Y_M1023_s N_VGND_c_709_n 0.00315309f $X=5.685 $Y=0.235 $X2=0 $Y2=0
cc_374 N_Y_M1011_s N_VGND_c_709_n 0.00249348f $X=6.525 $Y=0.235 $X2=0 $Y2=0
cc_375 N_Y_M1018_s N_VGND_c_709_n 0.00623102f $X=7.365 $Y=0.235 $X2=0 $Y2=0
cc_376 N_Y_c_581_n N_VGND_c_709_n 0.0218108f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_377 N_Y_c_631_p N_VGND_c_709_n 0.00643448f $X=6.66 $Y=0.42 $X2=0 $Y2=0
cc_378 N_Y_c_600_n N_VGND_c_709_n 0.00563684f $X=7.045 $Y=0.72 $X2=0 $Y2=0
cc_379 N_Y_c_633_p N_VGND_c_709_n 0.00637602f $X=7.5 $Y=0.42 $X2=0 $Y2=0
cc_380 N_Y_c_612_n N_VGND_c_709_n 0.00426801f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_381 N_Y_c_581_n N_A_445_47#_M1010_d 0.00312766f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_382 N_Y_c_581_n N_A_445_47#_M1017_d 0.00409876f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_383 N_Y_M1010_s N_A_445_47#_c_812_n 0.00476093f $X=4.015 $Y=0.235 $X2=0 $Y2=0
cc_384 N_Y_M1013_s N_A_445_47#_c_812_n 0.00315945f $X=4.845 $Y=0.235 $X2=0 $Y2=0
cc_385 N_Y_c_581_n N_A_445_47#_c_812_n 0.0797583f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_651_n N_VGND_M1012_s 0.00312394f $X=1.015 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_387 N_A_27_47#_c_657_n N_VGND_M1019_s 0.00312394f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_651_n N_VGND_c_700_n 0.0159625f $X=1.015 $Y=0.72 $X2=0 $Y2=0
cc_389 N_A_27_47#_c_657_n N_VGND_c_701_n 0.0159625f $X=1.855 $Y=0.72 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_676_p N_VGND_c_704_n 0.01143f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_391 N_A_27_47#_c_651_n N_VGND_c_704_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_651_n N_VGND_c_705_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_679_p N_VGND_c_705_n 0.0112274f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_657_n N_VGND_c_705_n 0.00244309f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_657_n N_VGND_c_706_n 0.00244309f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_682_p N_VGND_c_706_n 0.0112274f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_397 N_A_27_47#_c_650_n N_VGND_c_706_n 0.00245287f $X=3.62 $Y=0.72 $X2=0 $Y2=0
cc_398 N_A_27_47#_M1012_d N_VGND_c_709_n 0.00368727f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_M1015_d N_VGND_c_709_n 0.00249348f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_M1030_d N_VGND_c_709_n 0.00249348f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_M1022_s N_VGND_c_709_n 0.00219239f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_M1027_s N_VGND_c_709_n 0.00212464f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_676_p N_VGND_c_709_n 0.00643448f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_651_n N_VGND_c_709_n 0.00984256f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_679_p N_VGND_c_709_n 0.00643448f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_406 N_A_27_47#_c_657_n N_VGND_c_709_n 0.00984256f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_682_p N_VGND_c_709_n 0.00643448f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_408 N_A_27_47#_c_650_n N_VGND_c_709_n 0.00707809f $X=3.62 $Y=0.72 $X2=0 $Y2=0
cc_409 N_A_27_47#_c_650_n N_A_445_47#_M1016_d 0.00312766f $X=3.62 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_410 N_A_27_47#_c_650_n N_A_445_47#_M1026_d 0.00312766f $X=3.62 $Y=0.72 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_M1022_s N_A_445_47#_c_812_n 0.00315945f $X=2.645 $Y=0.235
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_M1027_s N_A_445_47#_c_812_n 0.00498385f $X=3.485 $Y=0.235
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_650_n N_A_445_47#_c_812_n 0.0797583f $X=3.62 $Y=0.72 $X2=0
+ $Y2=0
cc_414 N_VGND_c_709_n N_A_445_47#_M1016_d 0.00217615f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_415 N_VGND_c_709_n N_A_445_47#_M1026_d 0.00217615f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_709_n N_A_445_47#_M1010_d 0.00217615f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_709_n N_A_445_47#_M1017_d 0.00217615f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_702_n N_A_445_47#_c_812_n 0.00545039f $X=6.24 $Y=0.38 $X2=0
+ $Y2=0
cc_419 N_VGND_c_706_n N_A_445_47#_c_812_n 0.151358f $X=6.075 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_709_n N_A_445_47#_c_812_n 0.117456f $X=7.59 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.420000 1.020000 8.195000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.027500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 0.635000 8.195000 0.850000 ;
        RECT 4.870000 0.850000 5.250000 1.445000 ;
        RECT 4.870000 1.445000 7.720000 1.615000 ;
        RECT 4.870000 1.615000 5.200000 2.125000 ;
        RECT 5.710000 1.615000 6.040000 2.125000 ;
        RECT 6.550000 1.615000 6.880000 2.125000 ;
        RECT 7.390000 1.615000 7.720000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.695000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.695000 0.995000 ;
      RECT 0.500000  0.995000 4.700000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.035000  0.255000 1.205000 0.655000 ;
      RECT 1.035000  0.655000 4.700000 0.825000 ;
      RECT 1.075000  1.555000 4.700000 1.725000 ;
      RECT 1.075000  1.725000 1.285000 2.465000 ;
      RECT 1.375000  0.085000 1.705000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.875000  0.255000 2.045000 0.655000 ;
      RECT 1.955000  1.725000 2.125000 2.465000 ;
      RECT 2.215000  0.085000 2.545000 0.485000 ;
      RECT 2.295000  1.895000 2.625000 2.635000 ;
      RECT 2.715000  0.255000 2.885000 0.655000 ;
      RECT 2.795000  1.725000 2.965000 2.465000 ;
      RECT 3.055000  0.085000 3.385000 0.485000 ;
      RECT 3.135000  1.895000 3.465000 2.635000 ;
      RECT 3.555000  0.255000 3.725000 0.655000 ;
      RECT 3.635000  1.725000 3.805000 2.465000 ;
      RECT 3.895000  0.085000 4.235000 0.485000 ;
      RECT 3.975000  1.895000 4.305000 2.635000 ;
      RECT 4.405000  0.255000 8.195000 0.465000 ;
      RECT 4.405000  0.465000 4.700000 0.655000 ;
      RECT 4.475000  1.725000 4.700000 2.295000 ;
      RECT 4.475000  2.295000 8.195000 2.465000 ;
      RECT 5.370000  1.785000 5.540000 2.295000 ;
      RECT 6.210000  1.785000 6.380000 2.295000 ;
      RECT 7.050000  1.785000 7.220000 2.295000 ;
      RECT 7.890000  1.445000 8.195000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_8
END LIBRARY

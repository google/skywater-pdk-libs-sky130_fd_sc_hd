* File: sky130_fd_sc_hd__o311ai_0.pex.spice
* Created: Tue Sep  1 19:24:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311AI_0%A1 3 7 9 10 11 23
r27 20 23 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.405 $Y=1.16
+ $X2=0.615 $Y2=1.16
r28 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.16 $X2=0.405 $Y2=1.16
r29 10 11 6.50157 $w=6.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.432 $Y=1.19
+ $X2=0.432 $Y2=1.53
r30 10 21 0.573668 $w=6.38e-07 $l=3e-08 $layer=LI1_cond $X=0.432 $Y=1.19
+ $X2=0.432 $Y2=1.16
r31 9 21 5.9279 $w=6.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.432 $Y=0.85
+ $X2=0.432 $Y2=1.16
r32 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.325
+ $X2=0.615 $Y2=1.16
r33 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.615 $Y=1.325
+ $X2=0.615 $Y2=2.165
r34 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=1.16
r35 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%A2 3 7 9 10 11 12 18 19
c39 7 0 1.55302e-19 $X=1.035 $Y=2.165
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r41 11 12 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.105 $Y=1.87
+ $X2=1.105 $Y2=2.21
r42 10 11 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.105 $Y=1.53
+ $X2=1.105 $Y2=1.87
r43 9 10 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.105 $Y=1.19
+ $X2=1.105 $Y2=1.53
r44 9 19 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=1.105 $Y=1.19 $X2=1.105
+ $Y2=1.16
r45 5 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.325
+ $X2=1.035 $Y2=1.16
r46 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.035 $Y=1.325
+ $X2=1.035 $Y2=2.165
r47 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=0.995
+ $X2=1.035 $Y2=1.16
r48 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.035 $Y=0.995
+ $X2=1.035 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%A3 3 7 9 12
r31 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.16
+ $X2=1.515 $Y2=1.325
r32 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.16
+ $X2=1.515 $Y2=0.995
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=1.16 $X2=1.515 $Y2=1.16
r34 9 13 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=1.16
+ $X2=1.515 $Y2=1.16
r35 7 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.455 $Y=2.165
+ $X2=1.455 $Y2=1.325
r36 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.455 $Y=0.445
+ $X2=1.455 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%B1 3 7 9 12
r36 12 15 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.16
+ $X2=2.135 $Y2=1.325
r37 12 14 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.16
+ $X2=2.135 $Y2=0.995
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.16 $X2=2.115 $Y2=1.16
r39 7 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.215 $Y=0.445
+ $X2=2.215 $Y2=0.995
r40 3 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.055 $Y=2.165
+ $X2=2.055 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%C1 3 7 9 10 16
r26 13 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.575 $Y=1.16
+ $X2=2.915 $Y2=1.16
r27 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.16 $X2=2.915 $Y2=1.16
r28 9 10 11.7134 $w=3.03e-07 $l=3.1e-07 $layer=LI1_cond $X=2.982 $Y=0.85
+ $X2=2.982 $Y2=1.16
r29 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.325
+ $X2=2.575 $Y2=1.16
r30 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.575 $Y=1.325
+ $X2=2.575 $Y2=2.165
r31 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=1.16
r32 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%VPWR 1 2 7 9 13 16 17 18 28 29
r37 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r40 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 23 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 22 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r45 20 32 8.12166 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=0.78 $Y=2.72 $X2=0.39
+ $Y2=2.72
r46 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=2.72 $X2=1.15
+ $Y2=2.72
r47 18 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 16 25 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.15 $Y=2.72 $X2=2.07
+ $Y2=2.72
r49 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=2.72
+ $X2=2.315 $Y2=2.72
r50 15 28 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.48 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.72
+ $X2=2.315 $Y2=2.72
r52 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=2.635
+ $X2=2.315 $Y2=2.72
r53 11 13 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=2.315 $Y=2.635
+ $X2=2.315 $Y2=1.995
r54 7 32 2.64475 $w=6.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.432 $Y=2.635
+ $X2=0.39 $Y2=2.72
r55 7 9 11.0142 $w=6.93e-07 $l=6.4e-07 $layer=LI1_cond $X=0.432 $Y=2.635
+ $X2=0.432 $Y2=1.995
r56 2 13 300 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=2 $X=2.13
+ $Y=1.845 $X2=2.315 $Y2=1.995
r57 1 9 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.26
+ $Y=1.845 $X2=0.405 $Y2=1.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%Y 1 2 3 10 12 13 14 15 16 17 18 19 20
c47 10 0 1.55302e-19 $X=1.98 $Y=1.58
r48 48 50 4.23692 $w=3.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.66 $Y=0.425
+ $X2=2.785 $Y2=0.425
r49 20 58 5.3022 $w=4.83e-07 $l=2.15e-07 $layer=LI1_cond $X=2.892 $Y=2.21
+ $X2=2.892 $Y2=1.995
r50 19 58 3.08268 $w=4.83e-07 $l=1.25e-07 $layer=LI1_cond $X=2.892 $Y=1.87
+ $X2=2.892 $Y2=1.995
r51 19 54 5.05559 $w=4.83e-07 $l=2.05e-07 $layer=LI1_cond $X=2.892 $Y=1.87
+ $X2=2.892 $Y2=1.665
r52 18 50 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=2.99 $Y=0.425
+ $X2=2.785 $Y2=0.425
r53 17 41 2.73602 $w=3.5e-07 $l=2.77262e-07 $layer=LI1_cond $X=2.79 $Y=1.58
+ $X2=2.552 $Y2=1.495
r54 17 54 2.73602 $w=3.5e-07 $l=1.38109e-07 $layer=LI1_cond $X=2.79 $Y=1.58
+ $X2=2.892 $Y2=1.665
r55 17 41 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.552 $Y=1.47
+ $X2=2.552 $Y2=1.495
r56 16 17 15.0086 $w=2.13e-07 $l=2.8e-07 $layer=LI1_cond $X=2.552 $Y=1.19
+ $X2=2.552 $Y2=1.47
r57 15 16 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.552 $Y=0.85
+ $X2=2.552 $Y2=1.19
r58 14 48 2.82669 $w=3.4e-07 $l=1.08e-07 $layer=LI1_cond $X=2.552 $Y=0.425
+ $X2=2.66 $Y2=0.425
r59 14 15 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=2.552 $Y=0.595
+ $X2=2.552 $Y2=0.85
r60 13 36 4.67558 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.705 $Y=2.21
+ $X2=1.705 $Y2=1.995
r61 12 36 2.71836 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=1.87
+ $X2=1.705 $Y2=1.995
r62 11 12 4.45811 $w=5.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.87
r63 10 17 19.7147 $w=2.88e-07 $l=4.65e-07 $layer=LI1_cond $X=1.98 $Y=1.58
+ $X2=2.445 $Y2=1.58
r64 10 11 9.64472 $w=1.7e-07 $l=3.14643e-07 $layer=LI1_cond $X=1.98 $Y=1.58
+ $X2=1.705 $Y2=1.665
r65 3 58 300 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=2 $X=2.65
+ $Y=1.845 $X2=2.815 $Y2=1.995
r66 2 36 300 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.845 $X2=1.755 $Y2=1.995
r67 1 50 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.65
+ $Y=0.235 $X2=2.785 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%VGND 1 2 7 9 11 15 17 24 25 31
r43 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r44 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r45 22 25 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r46 22 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r47 21 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r48 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r49 19 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.245
+ $Y2=0
r50 19 21 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.61
+ $Y2=0
r51 17 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r52 17 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r53 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r54 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.36
r55 12 28 6.29768 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.285
+ $Y2=0
r56 11 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=1.245
+ $Y2=0
r57 11 12 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.57
+ $Y2=0
r58 7 28 2.80634 $w=4.85e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.327 $Y=0.085
+ $X2=0.285 $Y2=0
r59 7 9 8.87811 $w=4.83e-07 $l=3.6e-07 $layer=LI1_cond $X=0.327 $Y=0.085
+ $X2=0.327 $Y2=0.445
r60 2 15 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.235 $X2=1.245 $Y2=0.36
r61 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.26
+ $Y=0.235 $X2=0.405 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_0%A_138_47# 1 2 9 11 12 15
r26 13 15 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.665 $Y=0.655
+ $X2=1.665 $Y2=0.445
r27 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=0.74
+ $X2=1.665 $Y2=0.655
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.58 $Y=0.74
+ $X2=0.91 $Y2=0.74
r29 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.825 $Y=0.655
+ $X2=0.91 $Y2=0.74
r30 7 9 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.825 $Y=0.655
+ $X2=0.825 $Y2=0.445
r31 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.235 $X2=1.665 $Y2=0.445
r32 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.235 $X2=0.825 $Y2=0.445
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.915000 0.275000 13.255000 0.825000 ;
        RECT 12.915000 1.495000 13.255000 2.450000 ;
        RECT 13.070000 0.825000 13.255000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.500000 0.255000 11.830000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.345000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.765000 0.825000 1.675000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.550000 1.075000 0.840000 1.120000 ;
        RECT 0.550000 1.120000 2.675000 1.260000 ;
        RECT 0.550000 1.260000 0.840000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.015000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.885000 1.415000  9.110000 1.525000 ;
        RECT 8.885000 1.525000 10.075000 1.725000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.115000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.825000 1.415000 9.115000 1.460000 ;
        RECT 8.825000 1.600000 9.115000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.590000 ;
        RECT 2.905000 1.590000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.340000 0.085000 ;
        RECT  0.085000  0.085000  0.480000 0.595000 ;
        RECT  1.825000  0.085000  2.005000 0.545000 ;
        RECT  2.690000  0.085000  3.030000 0.555000 ;
        RECT  3.630000  0.085000  3.940000 0.545000 ;
        RECT  5.610000  0.085000  6.095000 0.465000 ;
        RECT  6.735000  0.085000  7.630000 0.805000 ;
        RECT 10.220000  0.085000 10.390000 0.545000 ;
        RECT 11.120000  0.085000 11.330000 0.885000 ;
        RECT 12.540000  0.085000 12.745000 0.825000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 13.340000 2.805000 ;
        RECT  0.515000 2.195000  0.765000 2.635000 ;
        RECT  2.690000 2.140000  3.030000 2.635000 ;
        RECT  3.595000 2.275000  3.925000 2.635000 ;
        RECT  5.945000 2.275000  6.275000 2.635000 ;
        RECT  7.005000 2.125000  7.960000 2.635000 ;
        RECT  9.195000 2.235000  9.525000 2.635000 ;
        RECT 10.135000 2.235000 10.465000 2.635000 ;
        RECT 11.120000 1.485000 11.330000 2.635000 ;
        RECT 12.575000 1.575000 12.745000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 1.845000  1.105000 2.025000 ;
      RECT  0.085000 2.025000  0.345000 2.465000 ;
      RECT  0.875000 0.280000  1.655000 0.560000 ;
      RECT  0.935000 2.025000  1.105000 2.255000 ;
      RECT  0.935000 2.255000  2.045000 2.465000 ;
      RECT  1.295000 1.870000  1.695000 2.075000 ;
      RECT  1.380000 0.560000  1.655000 0.590000 ;
      RECT  1.380000 0.590000  1.660000 0.600000 ;
      RECT  1.395000 0.600000  1.660000 0.605000 ;
      RECT  1.405000 0.605000  1.660000 0.610000 ;
      RECT  1.420000 0.610000  1.660000 0.615000 ;
      RECT  1.430000 0.615000  1.670000 0.620000 ;
      RECT  1.440000 0.620000  1.670000 0.630000 ;
      RECT  1.445000 0.630000  1.670000 0.635000 ;
      RECT  1.460000 0.635000  1.670000 0.645000 ;
      RECT  1.475000 0.645000  1.670000 0.655000 ;
      RECT  1.475000 0.655000  1.695000 0.665000 ;
      RECT  1.495000 0.665000  1.695000 0.705000 ;
      RECT  1.505000 0.705000  1.695000 1.870000 ;
      RECT  1.865000 0.715000  2.515000 0.905000 ;
      RECT  1.865000 0.905000  2.200000 1.770000 ;
      RECT  1.865000 1.770000  2.520000 2.085000 ;
      RECT  2.260000 0.255000  2.515000 0.715000 ;
      RECT  2.270000 2.085000  2.520000 2.465000 ;
      RECT  3.255000 1.775000  3.995000 1.955000 ;
      RECT  3.255000 1.955000  3.425000 2.325000 ;
      RECT  3.270000 0.255000  3.455000 0.715000 ;
      RECT  3.270000 0.715000  3.995000 0.885000 ;
      RECT  3.735000 0.885000  3.995000 1.775000 ;
      RECT  4.095000 2.135000  4.440000 2.465000 ;
      RECT  4.110000 0.255000  4.335000 0.585000 ;
      RECT  4.165000 0.585000  4.335000 1.090000 ;
      RECT  4.165000 1.090000  4.490000 1.420000 ;
      RECT  4.165000 1.420000  4.440000 2.135000 ;
      RECT  4.505000 0.255000  4.830000 0.920000 ;
      RECT  4.610000 1.590000  4.915000 1.615000 ;
      RECT  4.610000 1.615000  4.830000 2.465000 ;
      RECT  4.660000 0.920000  4.830000 1.445000 ;
      RECT  4.660000 1.445000  4.915000 1.590000 ;
      RECT  5.000000 0.255000  5.440000 1.225000 ;
      RECT  5.000000 1.225000  7.660000 1.275000 ;
      RECT  5.030000 2.135000  5.755000 2.465000 ;
      RECT  5.085000 1.275000  6.435000 1.395000 ;
      RECT  5.205000 1.575000  5.415000 1.955000 ;
      RECT  5.585000 1.395000  5.755000 2.135000 ;
      RECT  5.610000 0.635000  6.535000 0.805000 ;
      RECT  5.610000 0.805000  5.975000 1.015000 ;
      RECT  5.925000 1.575000  6.095000 1.935000 ;
      RECT  5.925000 1.935000  6.765000 2.105000 ;
      RECT  6.250000 0.975000  7.660000 1.225000 ;
      RECT  6.275000 0.255000  6.535000 0.635000 ;
      RECT  6.550000 2.105000  6.765000 2.450000 ;
      RECT  7.190000 1.495000  8.005000 1.955000 ;
      RECT  7.300000 1.275000  7.660000 1.325000 ;
      RECT  7.835000 0.695000  9.040000 0.895000 ;
      RECT  7.835000 0.895000  8.005000 1.495000 ;
      RECT  8.130000 2.125000  8.935000 2.460000 ;
      RECT  8.365000 1.075000  8.595000 1.905000 ;
      RECT  8.410000 0.275000  9.825000 0.445000 ;
      RECT  8.765000 1.895000 10.465000 2.065000 ;
      RECT  8.765000 2.065000  8.935000 2.125000 ;
      RECT  8.810000 0.895000  9.040000 1.245000 ;
      RECT  9.290000 0.855000  9.465000 1.185000 ;
      RECT  9.290000 1.185000 10.895000 1.355000 ;
      RECT  9.655000 0.445000  9.825000 0.845000 ;
      RECT  9.655000 0.845000 10.545000 1.015000 ;
      RECT  9.695000 2.065000  9.910000 2.450000 ;
      RECT 10.245000 1.525000 10.465000 1.895000 ;
      RECT 10.560000 0.255000 10.895000 0.540000 ;
      RECT 10.635000 1.355000 10.895000 2.465000 ;
      RECT 10.715000 0.540000 10.895000 1.185000 ;
      RECT 12.060000 0.255000 12.270000 0.995000 ;
      RECT 12.060000 0.995000 12.900000 1.325000 ;
      RECT 12.060000 1.325000 12.270000 2.465000 ;
    LAYER mcon ;
      RECT 1.525000 1.445000 1.695000 1.615000 ;
      RECT 3.825000 1.785000 3.995000 1.955000 ;
      RECT 4.285000 1.105000 4.455000 1.275000 ;
      RECT 4.745000 1.445000 4.915000 1.615000 ;
      RECT 5.205000 1.785000 5.375000 1.955000 ;
      RECT 7.505000 1.785000 7.675000 1.955000 ;
      RECT 8.425000 1.105000 8.595000 1.275000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.735000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.655000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.445000 1.755000 7.735000 1.800000 ;
      RECT 7.445000 1.940000 7.735000 1.985000 ;
      RECT 8.365000 1.075000 8.655000 1.120000 ;
      RECT 8.365000 1.260000 8.655000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfsbp_1

* File: sky130_fd_sc_hd__and3_4.pex.spice
* Created: Tue Sep  1 18:57:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND3_4%A 3 6 8 9 10 11 12 19 20 21 23
c33 20 0 1.08553e-20 $X=0.79 $Y=1.16
r34 19 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.79 $Y=1.16
+ $X2=0.79 $Y2=1.325
r35 19 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.79 $Y=1.16
+ $X2=0.79 $Y2=0.995
r36 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.79
+ $Y=1.16 $X2=0.79 $Y2=1.16
r37 12 20 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=1.167 $X2=0.79
+ $Y2=1.167
r38 12 28 10.8563 $w=3.43e-07 $l=3.25e-07 $layer=LI1_cond $X=0.69 $Y=1.167
+ $X2=0.365 $Y2=1.167
r39 10 11 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.24 $Y=1.87
+ $X2=0.24 $Y2=2.21
r40 9 10 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.24 $Y=1.53 $X2=0.24
+ $Y2=1.87
r41 9 23 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.53 $X2=0.24
+ $Y2=1.34
r42 8 23 4.08986 $w=2.5e-07 $l=1.73e-07 $layer=LI1_cond $X=0.24 $Y=1.167
+ $X2=0.24 $Y2=1.34
r43 8 28 2.9551 $w=3.45e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=1.167
+ $X2=0.365 $Y2=1.167
r44 6 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.85 $Y=1.985
+ $X2=0.85 $Y2=1.325
r45 3 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.85 $Y=0.56 $X2=0.85
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_4%B 3 6 8 9 13 15
c35 8 0 6.96876e-20 $X=1.065 $Y=0.765
c36 6 0 1.08553e-20 $X=1.395 $Y=1.985
r37 13 16 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.302 $Y=1.16
+ $X2=1.302 $Y2=1.325
r38 13 15 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.302 $Y=1.16
+ $X2=1.302 $Y2=0.995
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r40 9 14 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=1.21 $Y=1.19 $X2=1.21
+ $Y2=1.16
r41 8 14 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=1.21 $Y=0.85 $X2=1.21
+ $Y2=1.16
r42 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.395 $Y=1.985
+ $X2=1.395 $Y2=1.325
r43 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.395 $Y=0.56
+ $X2=1.395 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_4%C 3 6 8 11 12 13
c40 13 0 1.63729e-19 $X=1.815 $Y=0.995
c41 11 0 1.91186e-19 $X=1.815 $Y=1.16
c42 6 0 6.96876e-20 $X=1.825 $Y=1.985
r43 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=1.815 $Y2=1.325
r44 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=1.815 $Y2=0.995
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.16 $X2=1.815 $Y2=1.16
r46 8 12 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.61 $Y=1.16
+ $X2=1.815 $Y2=1.16
r47 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.825 $Y=1.985
+ $X2=1.825 $Y2=1.325
r48 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.755 $Y=0.56
+ $X2=1.755 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_4%A_94_47# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 40 42 43 44 48 50 52 55 57 63 67 71 72 76 83
c136 55 0 1.91186e-19 $X=2.175 $Y=1.02
c137 44 0 1.63729e-19 $X=1.535 $Y=0.47
r138 80 81 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.76 $Y=1.16
+ $X2=3.19 $Y2=1.16
r139 72 74 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=1.63 $Y=0.47
+ $X2=1.63 $Y2=0.71
r140 67 69 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=0.632 $Y=0.38
+ $X2=0.632 $Y2=0.47
r141 64 83 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.44 $Y=1.16
+ $X2=3.62 $Y2=1.16
r142 64 81 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.44 $Y=1.16
+ $X2=3.19 $Y2=1.16
r143 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r144 61 80 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.42 $Y=1.16
+ $X2=2.76 $Y2=1.16
r145 61 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.42 $Y=1.16 $X2=2.33
+ $Y2=1.16
r146 60 63 35.0893 $w=3.33e-07 $l=1.02e-06 $layer=LI1_cond $X=2.42 $Y=1.187
+ $X2=3.44 $Y2=1.187
r147 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.42
+ $Y=1.16 $X2=2.42 $Y2=1.16
r148 58 76 0.271299 $w=3.35e-07 $l=1.05e-07 $layer=LI1_cond $X=2.28 $Y=1.187
+ $X2=2.175 $Y2=1.187
r149 58 60 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=2.28 $Y=1.187
+ $X2=2.42 $Y2=1.187
r150 56 76 7.47207 $w=2.1e-07 $l=1.68e-07 $layer=LI1_cond $X=2.175 $Y=1.355
+ $X2=2.175 $Y2=1.187
r151 56 57 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=2.175 $Y=1.355
+ $X2=2.175 $Y2=1.58
r152 55 76 7.47207 $w=2.1e-07 $l=1.67e-07 $layer=LI1_cond $X=2.175 $Y=1.02
+ $X2=2.175 $Y2=1.187
r153 54 55 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.175 $Y=0.805
+ $X2=2.175 $Y2=1.02
r154 53 74 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=0.71
+ $X2=1.63 $Y2=0.71
r155 52 54 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=2.07 $Y=0.71
+ $X2=2.175 $Y2=0.805
r156 52 53 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=2.07 $Y=0.71
+ $X2=1.725 $Y2=0.71
r157 51 71 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.61
+ $Y2=1.665
r158 50 57 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.07 $Y=1.665
+ $X2=2.175 $Y2=1.58
r159 50 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.07 $Y=1.665
+ $X2=1.7 $Y2=1.665
r160 46 71 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.75
+ $X2=1.61 $Y2=1.665
r161 46 48 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=1.61 $Y=1.75
+ $X2=1.61 $Y2=1.96
r162 45 69 4.05585 $w=1.9e-07 $l=1.68e-07 $layer=LI1_cond $X=0.8 $Y=0.47
+ $X2=0.632 $Y2=0.47
r163 44 72 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.535 $Y=0.47
+ $X2=1.63 $Y2=0.47
r164 44 45 42.9043 $w=1.88e-07 $l=7.35e-07 $layer=LI1_cond $X=1.535 $Y=0.47
+ $X2=0.8 $Y2=0.47
r165 42 71 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.52 $Y=1.665 $X2=1.61
+ $Y2=1.665
r166 42 43 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=0.725 $Y2=1.665
r167 38 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.635 $Y=1.75
+ $X2=0.725 $Y2=1.665
r168 38 40 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.635 $Y=1.75
+ $X2=0.635 $Y2=1.96
r169 34 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.62 $Y=1.325
+ $X2=3.62 $Y2=1.16
r170 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.62 $Y=1.325
+ $X2=3.62 $Y2=1.985
r171 31 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.62 $Y2=1.16
r172 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.62 $Y2=0.56
r173 27 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.325
+ $X2=3.19 $Y2=1.16
r174 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.19 $Y=1.325
+ $X2=3.19 $Y2=1.985
r175 24 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=0.995
+ $X2=3.19 $Y2=1.16
r176 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.19 $Y=0.995
+ $X2=3.19 $Y2=0.56
r177 20 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.325
+ $X2=2.76 $Y2=1.16
r178 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.76 $Y=1.325
+ $X2=2.76 $Y2=1.985
r179 17 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=0.995
+ $X2=2.76 $Y2=1.16
r180 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.76 $Y=0.995
+ $X2=2.76 $Y2=0.56
r181 13 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.325
+ $X2=2.33 $Y2=1.16
r182 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.33 $Y=1.325
+ $X2=2.33 $Y2=1.985
r183 10 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=0.995
+ $X2=2.33 $Y2=1.16
r184 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.33 $Y=0.995
+ $X2=2.33 $Y2=0.56
r185 3 48 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=1.485 $X2=1.61 $Y2=1.96
r186 2 40 300 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=2 $X=0.47
+ $Y=1.485 $X2=0.635 $Y2=1.96
r187 1 67 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=0.47
+ $Y=0.235 $X2=0.635 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_4%VPWR 1 2 3 4 15 19 23 25 27 29 31 36 41 46 52
+ 55 58 62
r63 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r65 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 50 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 50 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 47 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=2.975 $Y2=2.72
r71 47 49 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 46 61 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.67 $Y=2.72
+ $X2=3.905 $Y2=2.72
r73 46 49 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.67 $Y=2.72
+ $X2=3.45 $Y2=2.72
r74 45 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 45 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=2.72
+ $X2=2.075 $Y2=2.72
r78 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.24 $Y=2.72
+ $X2=2.53 $Y2=2.72
r79 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.975 $Y2=2.72
r80 41 44 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.53 $Y2=2.72
r81 40 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r82 40 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r84 37 52 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=1.12 $Y2=2.72
r85 37 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=1.61 $Y2=2.72
r86 36 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=2.075 $Y2=2.72
r87 36 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=1.61
+ $Y2=2.72
r88 34 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 31 52 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.12 $Y2=2.72
r91 31 33 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.69 $Y2=2.72
r92 29 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r93 25 61 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.835 $Y=2.635
+ $X2=3.905 $Y2=2.72
r94 25 27 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.835 $Y=2.635
+ $X2=3.835 $Y2=2.02
r95 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.72
r96 21 23 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.02
r97 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=2.635
+ $X2=2.075 $Y2=2.72
r98 17 19 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.075 $Y=2.635
+ $X2=2.075 $Y2=2.02
r99 13 52 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r100 13 15 16.3464 $w=4.48e-07 $l=6.15e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.02
r101 4 27 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=3.695
+ $Y=1.485 $X2=3.835 $Y2=2.02
r102 3 23 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=2.835
+ $Y=1.485 $X2=2.975 $Y2=2.02
r103 2 19 300 $w=1.7e-07 $l=6.1632e-07 $layer=licon1_PDIFF $count=2 $X=1.9
+ $Y=1.485 $X2=2.075 $Y2=2.02
r104 1 15 300 $w=1.7e-07 $l=6.29206e-07 $layer=licon1_PDIFF $count=2 $X=0.925
+ $Y=1.485 $X2=1.13 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_4%X 1 2 3 4 15 17 19 20 23 27 29 31 36 38 40 42
+ 45 47
r56 45 47 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=3.915 $Y=0.845
+ $X2=3.915 $Y2=0.85
r57 42 45 3.11269 $w=2.8e-07 $l=1.15e-07 $layer=LI1_cond $X=3.915 $Y=0.73
+ $X2=3.915 $Y2=0.845
r58 42 47 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=3.915 $Y=0.89
+ $X2=3.915 $Y2=0.85
r59 41 42 26.5473 $w=2.78e-07 $l=6.45e-07 $layer=LI1_cond $X=3.915 $Y=1.535
+ $X2=3.915 $Y2=0.89
r60 34 36 4.38803 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.545 $Y=0.68
+ $X2=2.64 $Y2=0.68
r61 32 40 4.43576 $w=2.27e-07 $l=9.5e-08 $layer=LI1_cond $X=3.5 $Y=1.65
+ $X2=3.405 $Y2=1.65
r62 31 41 6.90206 $w=2.3e-07 $l=1.88944e-07 $layer=LI1_cond $X=3.775 $Y=1.65
+ $X2=3.915 $Y2=1.535
r63 31 32 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.775 $Y=1.65
+ $X2=3.5 $Y2=1.65
r64 30 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.5 $Y=0.73 $X2=3.405
+ $Y2=0.73
r65 29 42 3.78936 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.775 $Y=0.73
+ $X2=3.915 $Y2=0.73
r66 29 30 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.775 $Y=0.73
+ $X2=3.5 $Y2=0.73
r67 25 40 1.99853 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=1.65
r68 25 27 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=1.96
r69 21 38 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.405 $Y=0.615
+ $X2=3.405 $Y2=0.73
r70 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.405 $Y=0.615
+ $X2=3.405 $Y2=0.42
r71 19 40 4.43576 $w=2.27e-07 $l=9.64883e-08 $layer=LI1_cond $X=3.31 $Y=1.647
+ $X2=3.405 $Y2=1.65
r72 19 20 34.3172 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=3.31 $Y=1.647
+ $X2=2.64 $Y2=1.647
r73 17 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.31 $Y=0.73
+ $X2=3.405 $Y2=0.73
r74 17 36 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.31 $Y=0.73
+ $X2=2.64 $Y2=0.73
r75 13 20 6.87974 $w=2.25e-07 $l=1.5331e-07 $layer=LI1_cond $X=2.545 $Y=1.76
+ $X2=2.64 $Y2=1.647
r76 13 15 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=2.545 $Y=1.76
+ $X2=2.545 $Y2=1.96
r77 4 40 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.485 $X2=3.405 $Y2=1.62
r78 4 27 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=1.485 $X2=3.405 $Y2=1.96
r79 3 15 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=2.405
+ $Y=1.485 $X2=2.545 $Y2=1.96
r80 2 38 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.235 $X2=3.405 $Y2=0.76
r81 2 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.235 $X2=3.405 $Y2=0.42
r82 1 34 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=2.405
+ $Y=0.235 $X2=2.545 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_4%VGND 1 2 3 12 16 18 20 22 24 32 37 43 46 50
r68 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r69 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r70 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r71 41 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r72 41 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r73 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r74 38 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=2.975
+ $Y2=0
r75 38 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.45
+ $Y2=0
r76 37 49 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.905
+ $Y2=0
r77 37 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.45
+ $Y2=0
r78 36 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r79 36 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r80 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r81 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.07
+ $Y2=0
r82 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.53
+ $Y2=0
r83 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.975
+ $Y2=0
r84 32 35 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.53
+ $Y2=0
r85 31 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r86 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r87 26 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r88 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.07
+ $Y2=0
r89 24 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.61
+ $Y2=0
r90 22 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r91 22 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r92 18 49 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.905 $Y2=0
r93 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0.36
r94 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=0.085
+ $X2=2.975 $Y2=0
r95 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.975 $Y=0.085
+ $X2=2.975 $Y2=0.36
r96 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0
r97 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0.36
r98 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.835 $Y2=0.36
r99 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.235 $X2=2.975 $Y2=0.36
r100 1 12 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.235 $X2=2.07 $Y2=0.36
.ends


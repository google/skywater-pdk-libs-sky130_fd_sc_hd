# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.510000 1.560000 12.780000 2.465000 ;
        RECT 12.520000 0.255000 12.780000 0.760000 ;
        RECT 12.600000 0.760000 12.780000 1.560000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.880000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  1.875000  0.085000  2.205000 0.560000 ;
        RECT  2.395000  0.085000  2.725000 0.825000 ;
        RECT  4.445000  0.085000  4.775000 0.540000 ;
        RECT  6.915000  0.085000  7.245000 0.545000 ;
        RECT  9.085000  0.085000  9.255000 0.525000 ;
        RECT 10.720000  0.085000 10.890000 0.545000 ;
        RECT 12.010000  0.085000 12.340000 0.465000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 12.880000 2.805000 ;
        RECT  0.530000 2.135000  0.860000 2.635000 ;
        RECT  2.320000 2.040000  2.490000 2.635000 ;
        RECT  4.300000 2.275000  4.630000 2.635000 ;
        RECT  6.410000 2.355000  6.740000 2.635000 ;
        RECT  7.375000 2.175000  7.745000 2.635000 ;
        RECT  9.360000 2.195000  9.610000 2.635000 ;
        RECT 10.120000 2.255000 10.450000 2.635000 ;
        RECT 10.720000 1.495000 10.970000 2.635000 ;
        RECT 12.010000 1.875000 12.340000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.090000 1.795000  0.865000 1.965000 ;
      RECT  0.090000 1.965000  0.345000 2.465000 ;
      RECT  0.095000 0.345000  0.345000 0.635000 ;
      RECT  0.095000 0.635000  0.835000 0.805000 ;
      RECT  0.660000 0.805000  0.835000 0.995000 ;
      RECT  0.660000 0.995000  0.975000 1.325000 ;
      RECT  0.660000 1.325000  0.865000 1.795000 ;
      RECT  1.015000 0.345000  1.315000 0.675000 ;
      RECT  1.035000 1.730000  1.315000 1.900000 ;
      RECT  1.035000 1.900000  1.205000 2.465000 ;
      RECT  1.145000 0.675000  1.315000 1.730000 ;
      RECT  1.535000 0.395000  1.705000 0.730000 ;
      RECT  1.535000 0.730000  2.225000 0.900000 ;
      RECT  1.900000 2.055000  2.150000 2.400000 ;
      RECT  1.980000 1.260000  2.470000 1.455000 ;
      RECT  1.980000 1.455000  2.150000 2.055000 ;
      RECT  2.055000 0.900000  2.225000 0.995000 ;
      RECT  2.055000 0.995000  3.085000 1.185000 ;
      RECT  2.055000 1.185000  2.470000 1.260000 ;
      RECT  2.915000 0.255000  3.850000 0.425000 ;
      RECT  2.915000 0.425000  3.085000 0.995000 ;
      RECT  3.255000 0.675000  3.425000 1.015000 ;
      RECT  3.255000 1.015000  3.460000 1.185000 ;
      RECT  3.290000 1.185000  3.460000 1.935000 ;
      RECT  3.290000 1.935000  5.075000 2.105000 ;
      RECT  3.460000 2.105000  3.630000 2.465000 ;
      RECT  3.680000 0.425000  3.850000 1.685000 ;
      RECT  4.565000 0.715000  5.145000 0.895000 ;
      RECT  4.565000 0.895000  4.735000 1.935000 ;
      RECT  4.905000 1.065000  5.075000 1.395000 ;
      RECT  4.905000 2.105000  5.075000 2.185000 ;
      RECT  4.905000 2.185000  5.275000 2.435000 ;
      RECT  4.975000 0.335000  5.315000 0.505000 ;
      RECT  4.975000 0.505000  5.145000 0.715000 ;
      RECT  5.245000 1.575000  5.495000 1.955000 ;
      RECT  5.325000 0.705000  5.975000 1.035000 ;
      RECT  5.325000 1.035000  5.495000 1.575000 ;
      RECT  5.470000 2.135000  5.835000 2.465000 ;
      RECT  5.485000 0.305000  6.335000 0.475000 ;
      RECT  5.665000 1.215000  7.375000 1.385000 ;
      RECT  5.665000 1.385000  5.835000 2.135000 ;
      RECT  6.005000 1.935000  7.165000 2.105000 ;
      RECT  6.005000 2.105000  6.175000 2.375000 ;
      RECT  6.165000 0.475000  6.335000 1.215000 ;
      RECT  6.285000 1.595000  7.715000 1.765000 ;
      RECT  6.995000 2.105000  7.165000 2.375000 ;
      RECT  7.205000 1.005000  7.375000 1.215000 ;
      RECT  7.455000 0.275000  7.785000 0.445000 ;
      RECT  7.455000 0.445000  7.715000 0.835000 ;
      RECT  7.455000 1.765000  7.715000 1.835000 ;
      RECT  7.455000 1.835000  8.140000 2.005000 ;
      RECT  7.545000 0.835000  7.715000 1.595000 ;
      RECT  7.885000 0.705000  8.095000 1.495000 ;
      RECT  7.885000 1.495000  8.520000 1.655000 ;
      RECT  7.885000 1.655000  8.870000 1.665000 ;
      RECT  7.970000 2.005000  8.140000 2.465000 ;
      RECT  8.005000 0.255000  8.915000 0.535000 ;
      RECT  8.310000 1.665000  8.870000 1.935000 ;
      RECT  8.310000 1.935000  8.840000 1.955000 ;
      RECT  8.320000 2.125000  9.190000 2.465000 ;
      RECT  8.405000 0.920000  8.575000 1.325000 ;
      RECT  8.745000 0.535000  8.915000 1.315000 ;
      RECT  8.745000 1.315000  9.210000 1.485000 ;
      RECT  9.015000 2.035000  9.210000 2.115000 ;
      RECT  9.015000 2.115000  9.190000 2.125000 ;
      RECT  9.040000 1.485000  9.210000 1.575000 ;
      RECT  9.040000 1.575000 10.205000 1.745000 ;
      RECT  9.040000 1.745000  9.210000 2.035000 ;
      RECT  9.125000 0.695000  9.655000 0.865000 ;
      RECT  9.125000 0.865000  9.295000 1.145000 ;
      RECT  9.485000 0.295000 10.515000 0.465000 ;
      RECT  9.485000 0.465000  9.655000 0.695000 ;
      RECT  9.780000 1.915000 10.545000 2.085000 ;
      RECT  9.780000 2.085000  9.950000 2.375000 ;
      RECT 10.345000 0.465000 10.515000 0.995000 ;
      RECT 10.345000 0.995000 11.020000 1.295000 ;
      RECT 10.375000 1.295000 11.020000 1.325000 ;
      RECT 10.375000 1.325000 10.545000 1.915000 ;
      RECT 11.650000 1.535000 12.325000 1.705000 ;
      RECT 11.650000 1.705000 11.830000 2.465000 ;
      RECT 11.660000 0.255000 11.830000 0.635000 ;
      RECT 11.660000 0.635000 12.325000 0.805000 ;
      RECT 12.155000 0.805000 12.325000 1.060000 ;
      RECT 12.155000 1.060000 12.430000 1.390000 ;
      RECT 12.155000 1.390000 12.325000 1.535000 ;
    LAYER mcon ;
      RECT 0.805000 1.105000 0.975000 1.275000 ;
      RECT 1.035000 1.785000 1.205000 1.955000 ;
      RECT 4.905000 1.105000 5.075000 1.275000 ;
      RECT 5.325000 1.785000 5.495000 1.955000 ;
      RECT 8.405000 1.105000 8.575000 1.275000 ;
      RECT 8.445000 1.785000 8.615000 1.955000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrbp_1
END LIBRARY

* File: sky130_fd_sc_hd__a222oi_1.spice.SKY130_FD_SC_HD__A222OI_1.pxi
* Created: Thu Aug 27 14:02:19 2020
* 
x_PM_SKY130_FD_SC_HD__A222OI_1%C1 N_C1_M1011_g N_C1_M1009_g C1 N_C1_c_63_n
+ N_C1_c_64_n N_C1_c_65_n C1 PM_SKY130_FD_SC_HD__A222OI_1%C1
x_PM_SKY130_FD_SC_HD__A222OI_1%C2 N_C2_M1004_g N_C2_M1001_g C2 N_C2_c_94_n
+ N_C2_c_95_n PM_SKY130_FD_SC_HD__A222OI_1%C2
x_PM_SKY130_FD_SC_HD__A222OI_1%B2 N_B2_M1003_g N_B2_M1008_g B2 N_B2_c_128_n
+ N_B2_c_129_n PM_SKY130_FD_SC_HD__A222OI_1%B2
x_PM_SKY130_FD_SC_HD__A222OI_1%B1 N_B1_M1005_g N_B1_M1007_g B1 N_B1_c_163_n
+ N_B1_c_164_n PM_SKY130_FD_SC_HD__A222OI_1%B1
x_PM_SKY130_FD_SC_HD__A222OI_1%A1 N_A1_M1006_g N_A1_M1002_g A1 N_A1_c_196_n
+ N_A1_c_197_n PM_SKY130_FD_SC_HD__A222OI_1%A1
x_PM_SKY130_FD_SC_HD__A222OI_1%A2 N_A2_M1010_g N_A2_M1000_g A2 N_A2_c_228_n
+ N_A2_c_229_n PM_SKY130_FD_SC_HD__A222OI_1%A2
x_PM_SKY130_FD_SC_HD__A222OI_1%Y N_Y_M1011_s N_Y_M1005_d N_Y_M1009_s N_Y_M1001_d
+ N_Y_c_252_n N_Y_c_255_n N_Y_c_265_n N_Y_c_253_n N_Y_c_270_n N_Y_c_256_n
+ N_Y_c_287_n N_Y_c_290_n N_Y_c_257_n N_Y_c_258_n N_Y_c_259_n N_Y_c_312_p Y Y
+ PM_SKY130_FD_SC_HD__A222OI_1%Y
x_PM_SKY130_FD_SC_HD__A222OI_1%A_109_297# N_A_109_297#_M1009_d
+ N_A_109_297#_M1008_d N_A_109_297#_c_346_p N_A_109_297#_c_330_n
+ N_A_109_297#_c_331_n N_A_109_297#_c_344_p
+ PM_SKY130_FD_SC_HD__A222OI_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A222OI_1%A_311_297# N_A_311_297#_M1008_s
+ N_A_311_297#_M1007_d N_A_311_297#_M1000_d N_A_311_297#_c_356_n
+ N_A_311_297#_c_368_n N_A_311_297#_c_364_n N_A_311_297#_c_365_n
+ N_A_311_297#_c_357_n N_A_311_297#_c_366_n N_A_311_297#_c_374_n
+ N_A_311_297#_c_358_n N_A_311_297#_c_379_n N_A_311_297#_c_359_n
+ PM_SKY130_FD_SC_HD__A222OI_1%A_311_297#
x_PM_SKY130_FD_SC_HD__A222OI_1%VPWR N_VPWR_M1002_d N_VPWR_c_405_n N_VPWR_c_419_n
+ N_VPWR_c_406_n N_VPWR_c_407_n VPWR N_VPWR_c_408_n N_VPWR_c_404_n VPWR
+ PM_SKY130_FD_SC_HD__A222OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A222OI_1%VGND N_VGND_M1004_d N_VGND_M1010_d N_VGND_c_451_n
+ N_VGND_c_452_n VGND N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n
+ N_VGND_c_456_n VGND PM_SKY130_FD_SC_HD__A222OI_1%VGND
cc_1 VNB N_C1_c_63_n 0.0330844f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_2 VNB N_C1_c_64_n 0.0141583f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_3 VNB N_C1_c_65_n 0.0228156f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1
cc_4 VNB C2 0.0050758f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_5 VNB N_C2_c_94_n 0.0217917f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_6 VNB N_C2_c_95_n 0.0192453f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1
cc_7 VNB B2 0.00422551f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_8 VNB N_B2_c_128_n 0.0239373f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_9 VNB N_B2_c_129_n 0.0200757f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1
cc_10 VNB B1 0.00334856f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_11 VNB N_B1_c_163_n 0.0202448f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_12 VNB N_B1_c_164_n 0.0172355f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1
cc_13 VNB A1 0.00693299f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_14 VNB N_A1_c_196_n 0.0202476f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_15 VNB N_A1_c_197_n 0.0184496f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1
cc_16 VNB A2 0.0150009f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=1.09
cc_17 VNB N_A2_c_228_n 0.0234535f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.165
cc_18 VNB N_A2_c_229_n 0.0231349f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1
cc_19 VNB N_Y_c_252_n 0.0153416f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.157
cc_20 VNB N_Y_c_253_n 0.00745159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.0100708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_404_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_451_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_452_n 0.0267372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_453_n 0.0454414f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.157
cc_26 VNB N_VGND_c_454_n 0.0237516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_455_n 0.0178414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_456_n 0.199562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_C1_M1009_g 0.0258556f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_30 VPB N_C1_c_63_n 0.00957375f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_31 VPB N_C1_c_64_n 8.68599e-19 $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_32 VPB N_C2_M1001_g 0.0223758f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB C2 0.00107657f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_34 VPB N_C2_c_94_n 0.00473711f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_35 VPB N_B2_M1008_g 0.0226665f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB B2 3.33593e-19 $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_37 VPB N_B2_c_128_n 0.00649153f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_38 VPB N_B1_M1007_g 0.0189004f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB B1 0.00187612f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_40 VPB N_B1_c_163_n 0.0047554f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_41 VPB N_A1_M1002_g 0.0195444f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_42 VPB A1 0.00161044f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_43 VPB N_A1_c_196_n 0.00475837f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_44 VPB N_A2_M1000_g 0.02655f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB A2 0.00169445f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=1.09
cc_46 VPB N_A2_c_228_n 0.00454717f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_47 VPB N_Y_c_255_n 0.00964646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_Y_c_256_n 0.00476645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_257_n 0.00841329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_258_n 0.0214669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_Y_c_259_n 0.00787519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB Y 0.00277209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_109_297#_c_330_n 0.0111892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_311_297#_c_356_n 0.00430192f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.165
cc_55 VPB N_A_311_297#_c_357_n 0.0198658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_311_297#_c_358_n 0.0116537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_311_297#_c_359_n 0.00859245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_405_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_406_n 0.0705502f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.165
cc_60 VPB N_VPWR_c_407_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1
cc_61 VPB N_VPWR_c_408_n 0.0193344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_404_n 0.0469289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 N_C1_M1009_g N_C2_M1001_g 0.027761f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_64 N_C1_c_63_n C2 0.00104617f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_65 N_C1_c_64_n C2 0.0258586f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_66 N_C1_c_63_n N_C2_c_94_n 0.038913f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_67 N_C1_c_64_n N_C2_c_94_n 3.60288e-19 $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_68 N_C1_c_65_n N_C2_c_95_n 0.038913f $X=0.325 $Y=1 $X2=0 $Y2=0
cc_69 N_C1_c_65_n N_Y_c_252_n 0.00677814f $X=0.325 $Y=1 $X2=0 $Y2=0
cc_70 N_C1_M1009_g N_Y_c_255_n 0.00205643f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_71 N_C1_c_63_n N_Y_c_255_n 0.00669979f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_72 N_C1_c_64_n N_Y_c_255_n 0.0243799f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_73 N_C1_c_64_n N_Y_c_265_n 0.00794644f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_74 N_C1_c_65_n N_Y_c_265_n 0.00784669f $X=0.325 $Y=1 $X2=0 $Y2=0
cc_75 N_C1_c_63_n N_Y_c_253_n 0.00648158f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_76 N_C1_c_64_n N_Y_c_253_n 0.0227068f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_77 N_C1_c_65_n N_Y_c_253_n 8.84837e-19 $X=0.325 $Y=1 $X2=0 $Y2=0
cc_78 N_C1_M1009_g N_Y_c_270_n 0.00990148f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_79 N_C1_c_64_n N_Y_c_270_n 0.00794644f $X=0.38 $Y=1.165 $X2=0 $Y2=0
cc_80 N_C1_M1009_g N_Y_c_257_n 0.00313853f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_81 N_C1_M1009_g N_A_109_297#_c_331_n 0.00327186f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_82 N_C1_M1009_g N_VPWR_c_406_n 0.00510626f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_83 N_C1_M1009_g N_VPWR_c_404_n 0.00968865f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_84 N_C1_c_65_n N_VGND_c_454_n 0.00414303f $X=0.325 $Y=1 $X2=0 $Y2=0
cc_85 N_C1_c_65_n N_VGND_c_455_n 0.00186996f $X=0.325 $Y=1 $X2=0 $Y2=0
cc_86 N_C1_c_65_n N_VGND_c_456_n 0.00654541f $X=0.325 $Y=1 $X2=0 $Y2=0
cc_87 N_C2_c_94_n N_B2_c_128_n 0.00407805f $X=0.89 $Y=1.165 $X2=0 $Y2=0
cc_88 N_C2_c_95_n N_Y_c_252_n 0.00148545f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_89 C2 N_Y_c_265_n 0.0222407f $X=0.82 $Y=1.09 $X2=0 $Y2=0
cc_90 N_C2_c_94_n N_Y_c_265_n 0.00276586f $X=0.89 $Y=1.165 $X2=0 $Y2=0
cc_91 N_C2_c_95_n N_Y_c_265_n 0.0132688f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_92 N_C2_M1001_g N_Y_c_270_n 0.0101695f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 C2 N_Y_c_270_n 0.0167953f $X=0.82 $Y=1.09 $X2=0 $Y2=0
cc_94 N_C2_c_94_n N_Y_c_270_n 0.00145711f $X=0.89 $Y=1.165 $X2=0 $Y2=0
cc_95 N_C2_M1001_g N_Y_c_256_n 0.00485099f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_96 C2 N_Y_c_259_n 0.00508029f $X=0.82 $Y=1.09 $X2=0 $Y2=0
cc_97 N_C2_c_94_n N_Y_c_259_n 2.1076e-19 $X=0.89 $Y=1.165 $X2=0 $Y2=0
cc_98 C2 Y 0.0256311f $X=0.82 $Y=1.09 $X2=0 $Y2=0
cc_99 N_C2_c_94_n Y 0.00150745f $X=0.89 $Y=1.165 $X2=0 $Y2=0
cc_100 N_C2_c_95_n Y 0.00537776f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_101 N_C2_M1001_g N_A_109_297#_c_330_n 0.0114517f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_102 N_C2_M1001_g N_A_109_297#_c_331_n 0.00710241f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_C2_M1001_g N_A_311_297#_c_356_n 0.00282221f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_C2_M1001_g N_VPWR_c_406_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_105 N_C2_M1001_g N_VPWR_c_404_n 0.00662944f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 N_C2_c_95_n N_VGND_c_454_n 0.00340533f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_107 N_C2_c_95_n N_VGND_c_455_n 0.0106756f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_108 N_C2_c_95_n N_VGND_c_456_n 0.00385622f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_109 N_B2_M1008_g N_B1_M1007_g 0.043499f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_110 B2 B1 0.0258384f $X=1.755 $Y=1.09 $X2=0 $Y2=0
cc_111 N_B2_c_128_n B1 0.00106525f $X=1.82 $Y=1.165 $X2=0 $Y2=0
cc_112 B2 N_B1_c_163_n 3.80173e-19 $X=1.755 $Y=1.09 $X2=0 $Y2=0
cc_113 N_B2_c_128_n N_B1_c_163_n 0.0390259f $X=1.82 $Y=1.165 $X2=0 $Y2=0
cc_114 N_B2_c_129_n N_B1_c_164_n 0.0390259f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_115 N_B2_M1008_g N_Y_c_256_n 0.00456908f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_116 B2 N_Y_c_287_n 0.0191329f $X=1.755 $Y=1.09 $X2=0 $Y2=0
cc_117 N_B2_c_128_n N_Y_c_287_n 0.00342142f $X=1.82 $Y=1.165 $X2=0 $Y2=0
cc_118 N_B2_c_129_n N_Y_c_287_n 0.0135459f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_119 N_B2_c_129_n N_Y_c_290_n 0.00169984f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_120 N_B2_M1008_g N_Y_c_259_n 0.00630435f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_121 B2 Y 0.024609f $X=1.755 $Y=1.09 $X2=0 $Y2=0
cc_122 N_B2_c_128_n Y 0.00138609f $X=1.82 $Y=1.165 $X2=0 $Y2=0
cc_123 N_B2_c_129_n Y 0.00546293f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_124 N_B2_M1008_g N_A_109_297#_c_330_n 0.0104925f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_125 N_B2_M1008_g N_A_311_297#_c_356_n 0.00164765f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_126 B2 N_A_311_297#_c_356_n 0.0050766f $X=1.755 $Y=1.09 $X2=0 $Y2=0
cc_127 N_B2_c_128_n N_A_311_297#_c_356_n 0.00262732f $X=1.82 $Y=1.165 $X2=0
+ $Y2=0
cc_128 N_B2_M1008_g N_A_311_297#_c_364_n 7.59208e-19 $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_B2_M1008_g N_A_311_297#_c_365_n 8.95701e-19 $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_B2_M1008_g N_A_311_297#_c_366_n 0.0141455f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_131 B2 N_A_311_297#_c_366_n 0.00537711f $X=1.755 $Y=1.09 $X2=0 $Y2=0
cc_132 N_B2_M1008_g N_VPWR_c_406_n 0.00357877f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_133 N_B2_M1008_g N_VPWR_c_404_n 0.00662944f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_134 N_B2_c_129_n N_VGND_c_453_n 0.00426565f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_135 N_B2_c_129_n N_VGND_c_455_n 0.0125724f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_136 N_B2_c_129_n N_VGND_c_456_n 0.00714369f $X=1.81 $Y=1 $X2=0 $Y2=0
cc_137 N_B1_M1007_g N_A1_M1002_g 0.0148938f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_138 B1 A1 0.0258687f $X=2.225 $Y=1.09 $X2=0 $Y2=0
cc_139 N_B1_c_163_n A1 0.00180205f $X=2.31 $Y=1.165 $X2=0 $Y2=0
cc_140 B1 N_A1_c_196_n 3.82001e-19 $X=2.225 $Y=1.09 $X2=0 $Y2=0
cc_141 N_B1_c_163_n N_A1_c_196_n 0.0203108f $X=2.31 $Y=1.165 $X2=0 $Y2=0
cc_142 N_B1_c_164_n N_A1_c_197_n 0.010879f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_143 B1 N_Y_c_287_n 0.0183236f $X=2.225 $Y=1.09 $X2=0 $Y2=0
cc_144 N_B1_c_163_n N_Y_c_287_n 7.30673e-19 $X=2.31 $Y=1.165 $X2=0 $Y2=0
cc_145 N_B1_c_164_n N_Y_c_287_n 0.00917045f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_146 N_B1_c_164_n N_Y_c_290_n 0.00572028f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_147 N_B1_M1007_g N_A_311_297#_c_368_n 0.0113592f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_148 B1 N_A_311_297#_c_368_n 0.00842948f $X=2.225 $Y=1.09 $X2=0 $Y2=0
cc_149 N_B1_M1007_g N_A_311_297#_c_364_n 0.00398048f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_150 B1 N_A_311_297#_c_364_n 0.0046921f $X=2.225 $Y=1.09 $X2=0 $Y2=0
cc_151 N_B1_c_163_n N_A_311_297#_c_364_n 2.94234e-19 $X=2.31 $Y=1.165 $X2=0
+ $Y2=0
cc_152 N_B1_M1007_g N_A_311_297#_c_365_n 0.0062068f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B1_M1007_g N_A_311_297#_c_374_n 0.00242223f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_B1_M1007_g N_VPWR_c_406_n 0.00541359f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B1_M1007_g N_VPWR_c_404_n 0.00967871f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B1_c_164_n N_VGND_c_453_n 0.00423984f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_157 N_B1_c_164_n N_VGND_c_456_n 0.00584475f $X=2.31 $Y=1 $X2=0 $Y2=0
cc_158 N_A1_M1002_g N_A2_M1000_g 0.0232602f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_159 A1 A2 0.0260296f $X=2.705 $Y=1.09 $X2=0 $Y2=0
cc_160 N_A1_c_196_n A2 0.00180897f $X=2.79 $Y=1.165 $X2=0 $Y2=0
cc_161 A1 N_A2_c_228_n 3.78749e-19 $X=2.705 $Y=1.09 $X2=0 $Y2=0
cc_162 N_A1_c_196_n N_A2_c_228_n 0.0203289f $X=2.79 $Y=1.165 $X2=0 $Y2=0
cc_163 N_A1_c_197_n N_A2_c_229_n 0.0332815f $X=2.79 $Y=1 $X2=0 $Y2=0
cc_164 N_A1_M1002_g N_A_311_297#_c_364_n 0.00271412f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_165 A1 N_A_311_297#_c_364_n 0.00382056f $X=2.705 $Y=1.09 $X2=0 $Y2=0
cc_166 N_A1_M1002_g N_A_311_297#_c_374_n 0.00313631f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A1_M1002_g N_A_311_297#_c_358_n 2.06999e-19 $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A1_M1002_g N_A_311_297#_c_379_n 0.0101953f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_169 A1 N_A_311_297#_c_379_n 0.0153323f $X=2.705 $Y=1.09 $X2=0 $Y2=0
cc_170 N_A1_c_196_n N_A_311_297#_c_379_n 7.14516e-19 $X=2.79 $Y=1.165 $X2=0
+ $Y2=0
cc_171 N_A1_M1002_g N_VPWR_c_405_n 0.00277568f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A1_M1002_g N_VPWR_c_419_n 0.00287535f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A1_M1002_g N_VPWR_c_406_n 0.00510626f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A1_M1002_g N_VPWR_c_404_n 0.00877947f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A1_c_197_n N_VGND_c_452_n 0.00286189f $X=2.79 $Y=1 $X2=0 $Y2=0
cc_176 N_A1_c_197_n N_VGND_c_453_n 0.00585385f $X=2.79 $Y=1 $X2=0 $Y2=0
cc_177 N_A1_c_197_n N_VGND_c_456_n 0.0110778f $X=2.79 $Y=1 $X2=0 $Y2=0
cc_178 N_A2_M1000_g N_A_311_297#_c_358_n 0.00555699f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A2_c_228_n N_A_311_297#_c_358_n 0.00257612f $X=3.27 $Y=1.165 $X2=0
+ $Y2=0
cc_180 N_A2_M1000_g N_A_311_297#_c_379_n 0.00843175f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_181 A2 N_A_311_297#_c_379_n 0.0217171f $X=3.215 $Y=1.07 $X2=0 $Y2=0
cc_182 N_A2_M1000_g N_A_311_297#_c_359_n 0.00343123f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A2_M1000_g N_VPWR_c_405_n 0.00423848f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A2_M1000_g N_VPWR_c_408_n 0.00541359f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A2_M1000_g N_VPWR_c_404_n 0.0107463f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_186 A2 N_VGND_c_452_n 0.0114486f $X=3.215 $Y=1.07 $X2=0 $Y2=0
cc_187 N_A2_c_228_n N_VGND_c_452_n 0.00259233f $X=3.27 $Y=1.165 $X2=0 $Y2=0
cc_188 N_A2_c_229_n N_VGND_c_452_n 0.0176141f $X=3.27 $Y=1 $X2=0 $Y2=0
cc_189 N_A2_c_229_n N_VGND_c_453_n 0.0046653f $X=3.27 $Y=1 $X2=0 $Y2=0
cc_190 N_A2_c_229_n N_VGND_c_456_n 0.00814192f $X=3.27 $Y=1 $X2=0 $Y2=0
cc_191 N_Y_c_270_n N_A_109_297#_M1009_d 0.00655095f $X=1.015 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_192 N_Y_M1001_d N_A_109_297#_c_330_n 0.00629265f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_193 N_Y_c_270_n N_A_109_297#_c_330_n 0.00277132f $X=1.015 $Y=1.585 $X2=0
+ $Y2=0
cc_194 N_Y_c_259_n N_A_109_297#_c_330_n 0.01373f $X=1.1 $Y=1.665 $X2=0 $Y2=0
cc_195 N_Y_c_270_n N_A_109_297#_c_331_n 0.0142964f $X=1.015 $Y=1.585 $X2=0 $Y2=0
cc_196 N_Y_c_259_n N_A_311_297#_c_366_n 0.0048154f $X=1.1 $Y=1.665 $X2=0 $Y2=0
cc_197 N_Y_c_257_n N_VPWR_c_406_n 0.0208882f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_198 N_Y_M1009_s N_VPWR_c_404_n 0.00209319f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_199 N_Y_M1001_d N_VPWR_c_404_n 0.00210147f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_200 N_Y_c_257_n N_VPWR_c_404_n 0.0123452f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_201 N_Y_c_265_n A_109_47# 0.00535658f $X=1.255 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_202 N_Y_c_265_n N_VGND_M1004_d 0.0122978f $X=1.255 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_203 N_Y_c_287_n N_VGND_M1004_d 0.012968f $X=2.315 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_204 N_Y_c_312_p N_VGND_M1004_d 0.00456789f $X=1.367 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_205 Y N_VGND_M1004_d 0.00234717f $X=1.255 $Y=1.09 $X2=-0.19 $Y2=-0.24
cc_206 N_Y_c_287_n N_VGND_c_453_n 0.0105145f $X=2.315 $Y=0.73 $X2=0 $Y2=0
cc_207 N_Y_c_290_n N_VGND_c_453_n 0.0152618f $X=2.48 $Y=0.38 $X2=0 $Y2=0
cc_208 N_Y_c_252_n N_VGND_c_454_n 0.0207701f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_209 N_Y_c_265_n N_VGND_c_454_n 0.0065519f $X=1.255 $Y=0.73 $X2=0 $Y2=0
cc_210 N_Y_c_252_n N_VGND_c_455_n 0.00755777f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_211 N_Y_c_265_n N_VGND_c_455_n 0.0231635f $X=1.255 $Y=0.73 $X2=0 $Y2=0
cc_212 N_Y_c_287_n N_VGND_c_455_n 0.00901698f $X=2.315 $Y=0.73 $X2=0 $Y2=0
cc_213 N_Y_c_312_p N_VGND_c_455_n 0.0179745f $X=1.367 $Y=0.73 $X2=0 $Y2=0
cc_214 N_Y_M1011_s N_VGND_c_456_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_215 N_Y_M1005_d N_VGND_c_456_n 0.00300852f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_216 N_Y_c_252_n N_VGND_c_456_n 0.0123637f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_217 N_Y_c_265_n N_VGND_c_456_n 0.0131351f $X=1.255 $Y=0.73 $X2=0 $Y2=0
cc_218 N_Y_c_287_n N_VGND_c_456_n 0.0190645f $X=2.315 $Y=0.73 $X2=0 $Y2=0
cc_219 N_Y_c_290_n N_VGND_c_456_n 0.0121726f $X=2.48 $Y=0.38 $X2=0 $Y2=0
cc_220 N_Y_c_312_p N_VGND_c_456_n 0.00114853f $X=1.367 $Y=0.73 $X2=0 $Y2=0
cc_221 N_Y_c_287_n A_393_47# 0.00535658f $X=2.315 $Y=0.73 $X2=-0.19 $Y2=-0.24
cc_222 N_A_109_297#_c_330_n N_A_311_297#_M1008_s 0.00545924f $X=2.015 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_223 N_A_109_297#_c_330_n N_A_311_297#_c_356_n 0.0115135f $X=2.015 $Y=2.38
+ $X2=0 $Y2=0
cc_224 N_A_109_297#_c_331_n N_A_311_297#_c_356_n 0.00343074f $X=0.68 $Y=1.96
+ $X2=0 $Y2=0
cc_225 N_A_109_297#_M1008_d N_A_311_297#_c_368_n 0.00710142f $X=1.965 $Y=1.485
+ $X2=0 $Y2=0
cc_226 N_A_109_297#_c_344_p N_A_311_297#_c_368_n 0.00768758f $X=2.1 $Y=2.3 $X2=0
+ $Y2=0
cc_227 N_A_109_297#_c_330_n N_A_311_297#_c_366_n 0.00466557f $X=2.015 $Y=2.38
+ $X2=0 $Y2=0
cc_228 N_A_109_297#_c_346_p N_VPWR_c_406_n 0.0113535f $X=0.68 $Y=2.295 $X2=0
+ $Y2=0
cc_229 N_A_109_297#_c_330_n N_VPWR_c_406_n 0.0729478f $X=2.015 $Y=2.38 $X2=0
+ $Y2=0
cc_230 N_A_109_297#_c_331_n N_VPWR_c_406_n 9.40997e-19 $X=0.68 $Y=1.96 $X2=0
+ $Y2=0
cc_231 N_A_109_297#_c_344_p N_VPWR_c_406_n 0.0108432f $X=2.1 $Y=2.3 $X2=0 $Y2=0
cc_232 N_A_109_297#_M1009_d N_VPWR_c_404_n 0.00233719f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_109_297#_M1008_d N_VPWR_c_404_n 0.00384769f $X=1.965 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_A_109_297#_c_346_p N_VPWR_c_404_n 0.0065228f $X=0.68 $Y=2.295 $X2=0
+ $Y2=0
cc_235 N_A_109_297#_c_330_n N_VPWR_c_404_n 0.0450487f $X=2.015 $Y=2.38 $X2=0
+ $Y2=0
cc_236 N_A_109_297#_c_331_n N_VPWR_c_404_n 0.0020407f $X=0.68 $Y=1.96 $X2=0
+ $Y2=0
cc_237 N_A_109_297#_c_344_p N_VPWR_c_404_n 0.0063548f $X=2.1 $Y=2.3 $X2=0 $Y2=0
cc_238 N_A_311_297#_c_379_n N_VPWR_M1002_d 0.00904351f $X=3.22 $Y=1.617
+ $X2=-0.19 $Y2=1.305
cc_239 N_A_311_297#_c_359_n N_VPWR_c_405_n 0.0123166f $X=3.42 $Y=2.34 $X2=0
+ $Y2=0
cc_240 N_A_311_297#_c_379_n N_VPWR_c_419_n 0.0149709f $X=3.22 $Y=1.617 $X2=0
+ $Y2=0
cc_241 N_A_311_297#_c_374_n N_VPWR_c_406_n 0.018754f $X=2.52 $Y=2.34 $X2=0 $Y2=0
cc_242 N_A_311_297#_c_359_n N_VPWR_c_408_n 0.0216052f $X=3.42 $Y=2.34 $X2=0
+ $Y2=0
cc_243 N_A_311_297#_M1008_s N_VPWR_c_404_n 0.00210147f $X=1.555 $Y=1.485 $X2=0
+ $Y2=0
cc_244 N_A_311_297#_M1007_d N_VPWR_c_404_n 0.00215201f $X=2.385 $Y=1.485 $X2=0
+ $Y2=0
cc_245 N_A_311_297#_M1000_d N_VPWR_c_404_n 0.00209319f $X=3.285 $Y=1.485 $X2=0
+ $Y2=0
cc_246 N_A_311_297#_c_374_n N_VPWR_c_404_n 0.0121401f $X=2.52 $Y=2.34 $X2=0
+ $Y2=0
cc_247 N_A_311_297#_c_359_n N_VPWR_c_404_n 0.0127303f $X=3.42 $Y=2.34 $X2=0
+ $Y2=0
cc_248 A_109_47# N_VGND_c_456_n 0.00248276f $X=0.545 $Y=0.235 $X2=0.26 $Y2=2.255
cc_249 N_VGND_c_456_n A_393_47# 0.00248276f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_250 N_VGND_c_456_n A_561_47# 0.014106f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

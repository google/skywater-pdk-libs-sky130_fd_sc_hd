* File: sky130_fd_sc_hd__probe_p_8.pxi.spice
* Created: Tue Sep  1 19:29:25 2020
* 
x_PM_SKY130_FD_SC_HD__PROBE_P_8%A N_A_M1007_g N_A_M1002_g N_A_M1012_g
+ N_A_M1004_g N_A_c_120_n N_A_M1021_g N_A_M1013_g A A A
+ PM_SKY130_FD_SC_HD__PROBE_P_8%A
x_PM_SKY130_FD_SC_HD__PROBE_P_8%A_27_47# N_A_27_47#_M1007_d N_A_27_47#_M1012_d
+ N_A_27_47#_M1002_s N_A_27_47#_M1004_s N_A_27_47#_M1000_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1003_g N_A_27_47#_M1005_g N_A_27_47#_M1009_g N_A_27_47#_M1006_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1008_g N_A_27_47#_M1014_g N_A_27_47#_M1011_g
+ N_A_27_47#_M1016_g N_A_27_47#_M1015_g N_A_27_47#_M1017_g N_A_27_47#_M1019_g
+ N_A_27_47#_M1018_g N_A_27_47#_M1020_g N_A_27_47#_c_227_n N_A_27_47#_c_464_p
+ N_A_27_47#_c_210_n N_A_27_47#_c_211_n N_A_27_47#_c_228_n N_A_27_47#_c_229_n
+ N_A_27_47#_c_249_n N_A_27_47#_c_398_p N_A_27_47#_c_212_n N_A_27_47#_c_213_n
+ N_A_27_47#_c_214_n N_A_27_47#_c_215_n N_A_27_47#_c_231_n N_A_27_47#_c_216_n
+ N_A_27_47#_c_217_n N_A_27_47#_c_218_n PM_SKY130_FD_SC_HD__PROBE_P_8%A_27_47#
x_PM_SKY130_FD_SC_HD__PROBE_P_8%VPWR N_VPWR_M1002_d N_VPWR_M1013_d
+ N_VPWR_M1005_d N_VPWR_M1008_d N_VPWR_M1015_d N_VPWR_M1020_d N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n
+ N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n
+ N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n VPWR VPWR
+ N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_490_n N_VPWR_c_509_n N_VPWR_c_510_n
+ PM_SKY130_FD_SC_HD__PROBE_P_8%VPWR
x_PM_SKY130_FD_SC_HD__PROBE_P_8%noxref_6 N_noxref_6_M1000_d N_noxref_6_M1009_d
+ N_noxref_6_M1014_d N_noxref_6_M1017_d N_noxref_6_M1001_s N_noxref_6_M1006_s
+ N_noxref_6_M1011_s N_noxref_6_M1019_s N_noxref_6_c_646_n N_noxref_6_c_648_n
+ N_noxref_6_c_608_n N_noxref_6_c_609_n N_noxref_6_c_620_n N_noxref_6_c_621_n
+ N_noxref_6_c_667_n N_noxref_6_c_669_n N_noxref_6_c_610_n N_noxref_6_c_622_n
+ N_noxref_6_c_679_n N_noxref_6_c_681_n N_noxref_6_c_611_n N_noxref_6_c_623_n
+ N_noxref_6_c_612_n N_noxref_6_c_846_p N_noxref_6_c_794_n N_noxref_6_c_613_n
+ N_noxref_6_c_624_n N_noxref_6_c_614_n N_noxref_6_c_625_n N_noxref_6_c_615_n
+ N_noxref_6_c_626_n N_noxref_6_c_627_n N_noxref_6_c_616_n N_noxref_6_c_617_n
+ N_noxref_6_c_630_n N_noxref_6_c_618_n N_noxref_6_c_640_n N_noxref_6_c_632_n
+ N_noxref_6_R23_noxref_pos N_noxref_6_c_619_n
+ PM_SKY130_FD_SC_HD__PROBE_P_8%noxref_6
x_PM_SKY130_FD_SC_HD__PROBE_P_8%VGND N_VGND_M1007_s N_VGND_M1021_s
+ N_VGND_M1003_s N_VGND_M1010_s N_VGND_M1016_s N_VGND_M1018_s N_VGND_c_870_n
+ N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n N_VGND_c_875_n
+ N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n N_VGND_c_880_n
+ N_VGND_c_881_n N_VGND_c_882_n VGND VGND N_VGND_c_883_n VGND N_VGND_c_884_n
+ N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n
+ PM_SKY130_FD_SC_HD__PROBE_P_8%VGND
x_PM_SKY130_FD_SC_HD__PROBE_P_8%X X N_X_R23_noxref_neg
+ PM_SKY130_FD_SC_HD__PROBE_P_8%X
cc_1 VNB N_A_M1007_g 0.0228678f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1012_g 0.0170552f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_A_M1004_g 4.49778e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_4 VNB N_A_c_120_n 0.067134f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_5 VNB N_A_M1021_g 0.0169759f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_6 VNB N_A_M1013_g 4.42879e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_7 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_8 VNB N_A_27_47#_M1000_g 0.016824f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_9 VNB N_A_27_47#_M1001_g 4.20085e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_10 VNB N_A_27_47#_M1003_g 0.0164556f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_11 VNB N_A_27_47#_M1005_g 4.04623e-19 $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_12 VNB N_A_27_47#_M1009_g 0.0164701f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_13 VNB N_A_27_47#_M1006_g 4.04623e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_14 VNB N_A_27_47#_M1010_g 0.0164701f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_15 VNB N_A_27_47#_M1008_g 4.04623e-19 $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_16 VNB N_A_27_47#_M1014_g 0.0164484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_M1011_g 3.90963e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_M1016_g 0.0164123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_M1015_g 3.77304e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_M1017_g 0.016313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_M1019_g 3.7605e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_M1018_g 0.0233974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1020_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_210_n 0.00292127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_211_n 0.00183779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_212_n 9.42264e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_213_n 0.00900752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_214_n 0.00262633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_215_n 0.00211055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_216_n 0.00127298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_217_n 0.00132922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_218_n 0.150406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_490_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_noxref_6_c_608_n 0.00223004f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_35 VNB N_noxref_6_c_609_n 0.00111804f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_36 VNB N_noxref_6_c_610_n 0.00223004f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.175
cc_37 VNB N_noxref_6_c_611_n 0.00247147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_noxref_6_c_612_n 0.00113458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_noxref_6_c_613_n 9.73172e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_noxref_6_c_614_n 9.73172e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_noxref_6_c_615_n 2.04274e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_noxref_6_c_616_n 0.00951408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_noxref_6_c_617_n 0.00496574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_noxref_6_c_618_n 0.00128099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_noxref_6_c_619_n 0.00960561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_870_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.295
cc_47 VNB N_VGND_c_871_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_48 VNB N_VGND_c_872_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_873_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_50 VNB N_VGND_c_874_n 0.0112357f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_51 VNB N_VGND_c_875_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_52 VNB N_VGND_c_876_n 0.0309017f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_53 VNB N_VGND_c_877_n 0.0112511f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.175
cc_54 VNB N_VGND_c_878_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_879_n 0.0118636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_880_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_881_n 0.0112357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_882_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_883_n 0.0152765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_884_n 0.011863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_885_n 0.0172587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_886_n 0.292703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_887_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_888_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_889_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VPB N_A_M1002_g 0.0266267f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_A_M1004_g 0.0191647f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_A_c_120_n 0.00598216f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_69 VPB N_A_M1013_g 0.0191158f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_70 VPB N_A_27_47#_M1001_g 0.0189935f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_71 VPB N_A_27_47#_M1005_g 0.0182326f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_72 VPB N_A_27_47#_M1006_g 0.0182471f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_73 VPB N_A_27_47#_M1008_g 0.0182471f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_74 VPB N_A_27_47#_M1011_g 0.0181617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_M1015_g 0.0180762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_M1019_g 0.0180222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_M1020_g 0.0264665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_227_n 0.0331497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_228_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_229_n 0.0106324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_214_n 0.00763528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_231_n 0.00297261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_491_n 0.00410835f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.295
cc_84 VPB N_VPWR_c_492_n 0.00354062f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_85 VPB N_VPWR_c_493_n 3.15634e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_494_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.16
cc_87 VPB N_VPWR_c_495_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_88 VPB N_VPWR_c_496_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_89 VPB N_VPWR_c_497_n 0.0444458f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_90 VPB N_VPWR_c_498_n 0.0178658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_499_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_500_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_501_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_502_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_503_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_504_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_505_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_506_n 0.0124659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_507_n 0.0172587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_490_n 0.0596433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_509_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_510_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_noxref_6_c_620_n 0.0024098f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_104 VPB N_noxref_6_c_621_n 0.00138209f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_105 VPB N_noxref_6_c_622_n 0.0024098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_noxref_6_c_623_n 0.0025638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_noxref_6_c_624_n 0.00105115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_noxref_6_c_625_n 0.00105115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_noxref_6_c_626_n 0.00163765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_noxref_6_c_627_n 0.00180391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_noxref_6_c_616_n 0.00135411f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_noxref_6_c_617_n 0.00345636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_noxref_6_c_630_n 0.00420815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_noxref_6_c_618_n 9.71416e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_noxref_6_c_632_n 7.55234e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_noxref_6_c_619_n 0.0102093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 N_A_M1021_g N_A_27_47#_M1000_g 0.0260955f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_118 N_A_M1013_g N_A_27_47#_M1001_g 0.0260955f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1002_g N_A_27_47#_c_227_n 0.0106215f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_M1004_g N_A_27_47#_c_227_n 7.66249e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_M1007_g N_A_27_47#_c_210_n 0.0126041f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A_M1012_g N_A_27_47#_c_210_n 0.0114493f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_123 N_A_c_120_n N_A_27_47#_c_210_n 0.00322376f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_124 A N_A_27_47#_c_210_n 0.0473007f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_125 N_A_c_120_n N_A_27_47#_c_211_n 0.00413894f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_126 A N_A_27_47#_c_211_n 0.0138086f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A_M1002_g N_A_27_47#_c_228_n 0.0107189f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_M1004_g N_A_27_47#_c_228_n 0.0107189f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_c_120_n N_A_27_47#_c_228_n 0.00198252f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_130 A N_A_27_47#_c_228_n 0.0578998f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A_M1002_g N_A_27_47#_c_229_n 0.00168781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_c_120_n N_A_27_47#_c_229_n 0.00600433f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_133 A N_A_27_47#_c_229_n 0.0231044f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_M1002_g N_A_27_47#_c_249_n 7.67038e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1004_g N_A_27_47#_c_249_n 0.0107272f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1013_g N_A_27_47#_c_249_n 0.0106426f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1021_g N_A_27_47#_c_212_n 0.012104f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_138 A N_A_27_47#_c_212_n 0.00392548f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A_M1021_g N_A_27_47#_c_213_n 0.004229f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_c_120_n N_A_27_47#_c_214_n 0.00450613f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_141 A N_A_27_47#_c_214_n 0.00222755f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_142 N_A_M1004_g N_A_27_47#_c_231_n 0.00139111f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_c_120_n N_A_27_47#_c_231_n 0.00198252f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_144 N_A_M1013_g N_A_27_47#_c_231_n 0.0125562f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_c_120_n N_A_27_47#_c_216_n 0.00213376f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_146 A N_A_27_47#_c_216_n 0.0138019f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A_c_120_n N_A_27_47#_c_217_n 0.00167713f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_148 A N_A_27_47#_c_217_n 0.0141757f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A_c_120_n N_A_27_47#_c_218_n 0.0260955f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_150 N_A_M1002_g N_VPWR_c_491_n 0.00268723f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1004_g N_VPWR_c_491_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1013_g N_VPWR_c_492_n 0.00191527f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_VPWR_c_498_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_M1004_g N_VPWR_c_500_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1013_g N_VPWR_c_500_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1002_g N_VPWR_c_490_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1004_g N_VPWR_c_490_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_M1013_g N_VPWR_c_490_n 0.00927191f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1012_g N_noxref_6_c_618_n 4.18822e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_M1004_g N_noxref_6_c_618_n 5.21833e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_c_120_n N_noxref_6_c_618_n 0.00382357f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_162 N_A_M1021_g N_noxref_6_c_618_n 0.00242414f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A_M1013_g N_noxref_6_c_618_n 0.00515026f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_164 A N_noxref_6_c_618_n 0.00108623f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A_M1012_g N_noxref_6_c_640_n 2.58214e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A_M1004_g N_noxref_6_c_640_n 3.20593e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_c_120_n N_noxref_6_c_640_n 0.00531804f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_168 N_A_M1021_g N_noxref_6_c_640_n 0.00612881f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A_M1013_g N_noxref_6_c_640_n 0.00240196f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_170 A N_noxref_6_c_640_n 0.00120253f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A_M1007_g N_VGND_c_870_n 0.0094499f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A_M1012_g N_VGND_c_870_n 0.00772492f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A_M1021_g N_VGND_c_870_n 5.9099e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A_M1012_g N_VGND_c_871_n 5.9433e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_M1021_g N_VGND_c_871_n 0.00761022f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_M1012_g N_VGND_c_877_n 0.00350562f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_M1021_g N_VGND_c_877_n 0.00350562f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_M1007_g N_VGND_c_883_n 0.00350562f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A_M1007_g N_VGND_c_886_n 0.00517665f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_M1012_g N_VGND_c_886_n 0.00418574f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_M1021_g N_VGND_c_886_n 0.00412878f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_M1013_g X 0.00156409f $X=1.31 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_183 N_A_27_47#_c_228_n N_VPWR_M1002_d 0.00185611f $X=0.935 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_184 N_A_27_47#_c_231_n N_VPWR_M1013_d 0.00281475f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_228_n N_VPWR_c_491_n 0.0104788f $X=0.935 $Y=1.53 $X2=0 $Y2=0
cc_186 N_A_27_47#_M1001_g N_VPWR_c_492_n 0.0020122f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_249_n N_VPWR_c_492_n 0.0299702f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_215_n N_VPWR_c_492_n 2.25712e-19 $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_231_n N_VPWR_c_492_n 0.0103872f $X=1.507 $Y=1.53 $X2=0 $Y2=0
cc_190 N_A_27_47#_M1001_g N_VPWR_c_493_n 9.17051e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1005_g N_VPWR_c_493_n 0.0108489f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_27_47#_M1006_g N_VPWR_c_493_n 0.0106635f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_27_47#_M1008_g N_VPWR_c_493_n 8.84103e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1006_g N_VPWR_c_494_n 8.84103e-19 $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1008_g N_VPWR_c_494_n 0.0106635f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1011_g N_VPWR_c_494_n 0.0106635f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_27_47#_M1015_g N_VPWR_c_494_n 8.84103e-19 $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_M1011_g N_VPWR_c_495_n 0.0046653f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1015_g N_VPWR_c_495_n 0.0046653f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_27_47#_M1011_g N_VPWR_c_496_n 8.84103e-19 $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_M1015_g N_VPWR_c_496_n 0.0106635f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1019_g N_VPWR_c_496_n 0.0106995f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_27_47#_M1020_g N_VPWR_c_496_n 8.84564e-19 $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_M1019_g N_VPWR_c_497_n 8.09564e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1020_g N_VPWR_c_497_n 0.0157572f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_227_n N_VPWR_c_498_n 0.0210382f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_249_n N_VPWR_c_500_n 0.0189039f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1001_g N_VPWR_c_502_n 0.00585385f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1005_g N_VPWR_c_502_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1006_g N_VPWR_c_504_n 0.0046653f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_27_47#_M1008_g N_VPWR_c_504_n 0.0046653f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_27_47#_M1019_g N_VPWR_c_506_n 0.0046653f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_27_47#_M1020_g N_VPWR_c_506_n 0.0046653f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_27_47#_M1002_s N_VPWR_c_490_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1004_s N_VPWR_c_490_n 0.00215201f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_M1001_g N_VPWR_c_490_n 0.00984197f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_M1005_g N_VPWR_c_490_n 0.00731944f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_M1006_g N_VPWR_c_490_n 0.00731944f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_M1008_g N_VPWR_c_490_n 0.00731944f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1011_g N_VPWR_c_490_n 0.00731944f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_M1015_g N_VPWR_c_490_n 0.00731944f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_M1019_g N_VPWR_c_490_n 0.00785732f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_M1020_g N_VPWR_c_490_n 0.00796766f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_227_n N_VPWR_c_490_n 0.0124268f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_249_n N_VPWR_c_490_n 0.0122217f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_226 N_A_27_47#_M1000_g N_noxref_6_c_646_n 0.00121957f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_M1003_g N_noxref_6_c_646_n 0.00121957f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1001_g N_noxref_6_c_648_n 0.00205258f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1005_g N_noxref_6_c_648_n 0.00195397f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_249_n N_noxref_6_c_648_n 0.00454491f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1003_g N_noxref_6_c_608_n 0.0105482f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1009_g N_noxref_6_c_608_n 0.0109265f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_215_n N_noxref_6_c_608_n 0.0490878f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_218_n N_noxref_6_c_608_n 0.00202003f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_M1000_g N_noxref_6_c_609_n 0.0011364f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_212_n N_noxref_6_c_609_n 0.00844934f $X=1.42 $Y=0.82 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_215_n N_noxref_6_c_609_n 0.0137623f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_218_n N_noxref_6_c_609_n 0.00208213f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1005_g N_noxref_6_c_620_n 0.0122351f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1006_g N_noxref_6_c_620_n 0.0125142f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_215_n N_noxref_6_c_620_n 0.0428422f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_218_n N_noxref_6_c_620_n 0.00197712f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_M1001_g N_noxref_6_c_621_n 0.0010746f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_215_n N_noxref_6_c_621_n 0.0120817f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_231_n N_noxref_6_c_621_n 0.00870005f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_218_n N_noxref_6_c_621_n 0.00205043f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_M1009_g N_noxref_6_c_667_n 0.00121957f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1010_g N_noxref_6_c_667_n 0.00121957f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1006_g N_noxref_6_c_669_n 0.00195397f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1008_g N_noxref_6_c_669_n 0.00195397f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1010_g N_noxref_6_c_610_n 0.0109707f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1014_g N_noxref_6_c_610_n 0.0109707f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_215_n N_noxref_6_c_610_n 0.0488959f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_218_n N_noxref_6_c_610_n 0.00202003f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1008_g N_noxref_6_c_622_n 0.0125584f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1011_g N_noxref_6_c_622_n 0.0125584f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_215_n N_noxref_6_c_622_n 0.0425781f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_218_n N_noxref_6_c_622_n 0.00197712f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1014_g N_noxref_6_c_679_n 0.00121957f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1016_g N_noxref_6_c_679_n 0.00121957f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1011_g N_noxref_6_c_681_n 0.00195397f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1015_g N_noxref_6_c_681_n 0.00195397f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1016_g N_noxref_6_c_611_n 0.0109265f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1017_g N_noxref_6_c_611_n 0.00870955f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_215_n N_noxref_6_c_611_n 0.0238195f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_218_n N_noxref_6_c_611_n 0.00204324f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_M1015_g N_noxref_6_c_623_n 0.0125584f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1019_g N_noxref_6_c_623_n 0.0109215f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_215_n N_noxref_6_c_623_n 0.0204251f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_218_n N_noxref_6_c_623_n 0.001731f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1016_g N_noxref_6_c_612_n 5.83668e-19 $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1017_g N_noxref_6_c_612_n 0.00306769f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1018_g N_noxref_6_c_612_n 0.00307239f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_218_n N_noxref_6_c_612_n 0.00498725f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_215_n N_noxref_6_c_613_n 0.0137623f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_218_n N_noxref_6_c_613_n 0.00208213f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_215_n N_noxref_6_c_624_n 0.0120817f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_218_n N_noxref_6_c_624_n 0.00205043f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_215_n N_noxref_6_c_614_n 0.0131988f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_218_n N_noxref_6_c_614_n 0.00193766f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_215_n N_noxref_6_c_625_n 0.0113996f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_218_n N_noxref_6_c_625_n 0.00166072f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1017_g N_noxref_6_c_615_n 0.00272967f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_M1018_g N_noxref_6_c_615_n 0.00114299f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1015_g N_noxref_6_c_626_n 8.35458e-19 $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1019_g N_noxref_6_c_626_n 0.00740053f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1020_g N_noxref_6_c_626_n 0.0052532f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_215_n N_noxref_6_c_626_n 0.00732938f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_218_n N_noxref_6_c_626_n 0.0114051f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1019_g N_noxref_6_c_627_n 2.22048e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_215_n N_noxref_6_c_627_n 0.00392059f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_218_n N_noxref_6_c_627_n 0.00299048f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1019_g N_noxref_6_c_616_n 0.00352352f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_218_n N_noxref_6_c_616_n 0.00556094f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1020_g N_noxref_6_c_617_n 0.00666556f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_218_n N_noxref_6_c_617_n 0.0169938f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1011_g N_noxref_6_c_630_n 8.61503e-19 $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1015_g N_noxref_6_c_630_n 0.00294243f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_215_n N_noxref_6_c_630_n 0.0182206f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_218_n N_noxref_6_c_630_n 0.0107749f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1000_g N_noxref_6_c_618_n 0.00299603f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1001_g N_noxref_6_c_618_n 0.00345649f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_M1003_g N_noxref_6_c_618_n 0.00216773f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_M1005_g N_noxref_6_c_618_n 0.00223217f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1009_g N_noxref_6_c_618_n 0.00216955f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1006_g N_noxref_6_c_618_n 0.00222181f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1010_g N_noxref_6_c_618_n 0.00216955f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_M1008_g N_noxref_6_c_618_n 0.00221025f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1014_g N_noxref_6_c_618_n 0.00215562f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1011_g N_noxref_6_c_618_n 0.00208137f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_M1016_g N_noxref_6_c_618_n 0.00181943f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_M1015_g N_noxref_6_c_618_n 0.00145196f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_M1017_g N_noxref_6_c_618_n 8.42392e-19 $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1019_g N_noxref_6_c_618_n 0.00147202f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_249_n N_noxref_6_c_618_n 0.0014224f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_398_p N_noxref_6_c_618_n 3.55572e-19 $X=1.1 $Y=0.56 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_212_n N_noxref_6_c_618_n 0.00308681f $X=1.42 $Y=0.82 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_213_n N_noxref_6_c_618_n 0.00258043f $X=1.507 $Y=1.075 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_214_n N_noxref_6_c_618_n 0.0030166f $X=1.507 $Y=1.445 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_215_n N_noxref_6_c_618_n 0.00890046f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_231_n N_noxref_6_c_618_n 0.00400474f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_217_n N_noxref_6_c_618_n 3.47197e-19 $X=1.507 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_218_n N_noxref_6_c_618_n 0.00244823f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1000_g N_noxref_6_c_640_n 0.00178028f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1003_g N_noxref_6_c_640_n 0.00176611f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_M1009_g N_noxref_6_c_640_n 0.00176611f $X=2.57 $Y=0.56 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_M1010_g N_noxref_6_c_640_n 0.00176611f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_M1014_g N_noxref_6_c_640_n 0.00176611f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_M1016_g N_noxref_6_c_640_n 0.00176611f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_M1017_g N_noxref_6_c_640_n 0.00568178f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_M1019_g N_noxref_6_c_640_n 0.00745955f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_227_n N_noxref_6_c_640_n 6.11998e-19 $X=0.26 $Y=1.63 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_249_n N_noxref_6_c_640_n 0.00615941f $X=1.1 $Y=1.63 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_398_p N_noxref_6_c_640_n 0.00120869f $X=1.1 $Y=0.56 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_212_n N_noxref_6_c_640_n 0.0035243f $X=1.42 $Y=0.82 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_231_n N_noxref_6_c_640_n 0.00375854f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_218_n N_noxref_6_c_640_n 7.93234e-19 $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_M1008_g N_noxref_6_c_632_n 3.07854e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_M1011_g N_noxref_6_c_632_n 0.00154019f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1019_g N_noxref_6_c_632_n 4.86156e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_215_n N_noxref_6_c_632_n 0.00312295f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_218_n N_noxref_6_c_632_n 0.00421165f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_M1008_g N_noxref_6_c_619_n 4.89114e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_M1014_g N_noxref_6_c_619_n 0.00138846f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_M1011_g N_noxref_6_c_619_n 0.00230703f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_M1016_g N_noxref_6_c_619_n 0.00355547f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_M1015_g N_noxref_6_c_619_n 0.00372276f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_M1017_g N_noxref_6_c_619_n 2.43988e-19 $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_M1019_g N_noxref_6_c_619_n 7.37946e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_215_n N_noxref_6_c_619_n 0.00349157f $X=3.88 $Y=1.16 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_218_n N_noxref_6_c_619_n 0.00327537f $X=4.67 $Y=1.16 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_210_n N_VGND_M1007_s 0.00162006f $X=1.015 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_353 N_A_27_47#_c_212_n N_VGND_M1021_s 0.00281281f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_210_n N_VGND_c_870_n 0.016419f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_355 N_A_27_47#_M1000_g N_VGND_c_871_n 0.00788658f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_27_47#_M1003_g N_VGND_c_871_n 5.81128e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_212_n N_VGND_c_871_n 0.0182088f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_215_n N_VGND_c_871_n 0.00255027f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A_27_47#_M1000_g N_VGND_c_872_n 5.81128e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_27_47#_M1003_g N_VGND_c_872_n 0.00760925f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_27_47#_M1009_g N_VGND_c_872_n 0.00760925f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_27_47#_M1010_g N_VGND_c_872_n 5.81128e-19 $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_27_47#_M1009_g N_VGND_c_873_n 5.81128e-19 $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_27_47#_M1010_g N_VGND_c_873_n 0.00760925f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_27_47#_M1014_g N_VGND_c_873_n 0.00760925f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A_27_47#_M1016_g N_VGND_c_873_n 5.81128e-19 $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A_27_47#_M1014_g N_VGND_c_874_n 0.00350562f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_27_47#_M1016_g N_VGND_c_874_n 0.00350562f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_369 N_A_27_47#_M1014_g N_VGND_c_875_n 5.81128e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_27_47#_M1016_g N_VGND_c_875_n 0.00760925f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_27_47#_M1017_g N_VGND_c_875_n 0.00760925f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_27_47#_M1018_g N_VGND_c_875_n 5.81128e-19 $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A_27_47#_M1017_g N_VGND_c_876_n 7.31324e-19 $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A_27_47#_M1018_g N_VGND_c_876_n 0.0121041f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_375 N_A_27_47#_c_210_n N_VGND_c_877_n 0.00193763f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_398_p N_VGND_c_877_n 0.0110017f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A_27_47#_c_212_n N_VGND_c_877_n 0.00249618f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_378 N_A_27_47#_M1000_g N_VGND_c_879_n 0.0046653f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_379 N_A_27_47#_M1003_g N_VGND_c_879_n 0.00350562f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_380 N_A_27_47#_M1009_g N_VGND_c_881_n 0.00350562f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_381 N_A_27_47#_M1010_g N_VGND_c_881_n 0.00350562f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_382 N_A_27_47#_c_464_p N_VGND_c_883_n 0.0115672f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_210_n N_VGND_c_883_n 0.00193763f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1017_g N_VGND_c_884_n 0.0035053f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A_27_47#_M1018_g N_VGND_c_884_n 0.0046653f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_386 N_A_27_47#_M1007_d N_VGND_c_886_n 0.00377256f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_M1012_d N_VGND_c_886_n 0.00266498f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1000_g N_VGND_c_886_n 0.00729505f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_389 N_A_27_47#_M1003_g N_VGND_c_886_n 0.00396954f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_390 N_A_27_47#_M1009_g N_VGND_c_886_n 0.00396954f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_391 N_A_27_47#_M1010_g N_VGND_c_886_n 0.00396954f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_392 N_A_27_47#_M1014_g N_VGND_c_886_n 0.00372552f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_393 N_A_27_47#_M1016_g N_VGND_c_886_n 0.00364147f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_394 N_A_27_47#_M1017_g N_VGND_c_886_n 0.00414969f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_395 N_A_27_47#_M1018_g N_VGND_c_886_n 0.00796766f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_396 N_A_27_47#_c_464_p N_VGND_c_886_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_397 N_A_27_47#_c_210_n N_VGND_c_886_n 0.00895872f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_398_p N_VGND_c_886_n 0.00644569f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_399 N_A_27_47#_c_212_n N_VGND_c_886_n 0.00479056f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_400 N_A_27_47#_M1001_g X 0.00204351f $X=1.73 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_401 N_A_27_47#_M1005_g X 0.00166552f $X=2.15 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_402 N_A_27_47#_M1006_g X 0.00166552f $X=2.57 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_403 N_A_27_47#_M1008_g X 0.00166552f $X=2.99 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_404 N_A_27_47#_M1011_g X 0.00166552f $X=3.41 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_405 N_A_27_47#_M1015_g X 0.00166552f $X=3.83 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_406 N_A_27_47#_M1019_g X 0.00399484f $X=4.25 $Y=1.985 $X2=-0.19 $Y2=-0.24
cc_407 N_A_27_47#_c_249_n X 0.00390964f $X=1.1 $Y=1.63 $X2=-0.19 $Y2=-0.24
cc_408 N_VPWR_c_490_n N_noxref_6_M1001_s 0.00498929f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_490_n N_noxref_6_M1006_s 0.00498929f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_490_n N_noxref_6_M1011_s 0.00498929f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_490_n N_noxref_6_M1019_s 0.00570907f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_492_n N_noxref_6_c_648_n 0.00932276f $X=1.52 $Y=2 $X2=0 $Y2=0
cc_413 N_VPWR_c_493_n N_noxref_6_c_648_n 0.0299716f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_414 N_VPWR_c_502_n N_noxref_6_c_648_n 0.0113958f $X=2.195 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_c_490_n N_noxref_6_c_648_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_M1005_d N_noxref_6_c_620_n 0.00138461f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_493_n N_noxref_6_c_620_n 0.0179526f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_418 N_VPWR_c_493_n N_noxref_6_c_669_n 0.0299716f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_419 N_VPWR_c_494_n N_noxref_6_c_669_n 0.0299716f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_420 N_VPWR_c_504_n N_noxref_6_c_669_n 0.0113958f $X=3.035 $Y=2.72 $X2=0 $Y2=0
cc_421 N_VPWR_c_490_n N_noxref_6_c_669_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_M1008_d N_noxref_6_c_622_n 0.00138461f $X=3.065 $Y=1.485 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_494_n N_noxref_6_c_622_n 0.0179526f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_424 N_VPWR_c_494_n N_noxref_6_c_681_n 0.0299716f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_425 N_VPWR_c_495_n N_noxref_6_c_681_n 0.0113958f $X=3.875 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_c_496_n N_noxref_6_c_681_n 0.0299716f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_427 N_VPWR_c_490_n N_noxref_6_c_681_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_M1015_d N_noxref_6_c_623_n 0.00138461f $X=3.905 $Y=1.485 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_496_n N_noxref_6_c_623_n 0.0179676f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_430 N_VPWR_c_506_n N_noxref_6_c_794_n 0.0113958f $X=4.715 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_c_490_n N_noxref_6_c_794_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_432 N_VPWR_c_497_n N_noxref_6_c_616_n 0.00227769f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_433 N_VPWR_c_497_n N_noxref_6_c_617_n 0.0107017f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_434 N_VPWR_M1013_d N_noxref_6_c_618_n 0.00108834f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_VPWR_M1015_d N_noxref_6_c_618_n 0.00247526f $X=3.905 $Y=1.485 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_492_n N_noxref_6_c_618_n 0.00251602f $X=1.52 $Y=2 $X2=0 $Y2=0
cc_437 N_VPWR_c_493_n N_noxref_6_c_618_n 0.00486812f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_438 N_VPWR_c_494_n N_noxref_6_c_618_n 0.00477242f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_439 N_VPWR_c_496_n N_noxref_6_c_618_n 0.00424153f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_440 N_VPWR_c_490_n N_noxref_6_c_618_n 0.0466821f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_441 N_VPWR_c_491_n N_noxref_6_c_640_n 2.61592e-19 $X=0.68 $Y=2 $X2=0 $Y2=0
cc_442 N_VPWR_c_492_n N_noxref_6_c_640_n 3.05197e-19 $X=1.52 $Y=2 $X2=0 $Y2=0
cc_443 N_VPWR_c_493_n N_noxref_6_c_640_n 2.12444e-19 $X=2.36 $Y=2 $X2=0 $Y2=0
cc_444 N_VPWR_c_494_n N_noxref_6_c_640_n 2.12444e-19 $X=3.2 $Y=2 $X2=0 $Y2=0
cc_445 N_VPWR_c_497_n N_VGND_c_876_n 0.00516367f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_446 N_VPWR_M1013_d X 0.00158966f $X=1.385 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_447 N_VPWR_c_491_n X 5.01252e-19 $X=0.68 $Y=2 $X2=-0.19 $Y2=-0.24
cc_448 N_VPWR_c_492_n X 0.00312271f $X=1.52 $Y=2 $X2=-0.19 $Y2=-0.24
cc_449 N_VPWR_c_493_n X 0.00514275f $X=2.36 $Y=2 $X2=-0.19 $Y2=-0.24
cc_450 N_VPWR_c_494_n X 0.00514275f $X=3.2 $Y=2 $X2=-0.19 $Y2=-0.24
cc_451 N_VPWR_c_496_n X 0.00487846f $X=4.04 $Y=2 $X2=-0.19 $Y2=-0.24
cc_452 N_VPWR_c_490_n X 0.0376037f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_453 N_noxref_6_c_618_n N_VGND_M1021_s 0.00306096f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_454 N_noxref_6_c_608_n N_VGND_M1003_s 0.0011982f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_455 N_noxref_6_c_618_n N_VGND_M1003_s 0.00306096f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_456 N_noxref_6_c_610_n N_VGND_M1010_s 0.0011982f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_457 N_noxref_6_c_618_n N_VGND_M1010_s 0.00306096f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_458 N_noxref_6_c_611_n N_VGND_M1016_s 0.0011982f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_459 N_noxref_6_c_618_n N_VGND_M1016_s 0.00339068f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_460 N_noxref_6_c_646_n N_VGND_c_871_n 0.0117314f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_461 N_noxref_6_c_618_n N_VGND_c_871_n 0.00256166f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_462 N_noxref_6_c_640_n N_VGND_c_871_n 0.00553005f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_463 N_noxref_6_c_646_n N_VGND_c_872_n 0.0117314f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_464 N_noxref_6_c_608_n N_VGND_c_872_n 0.0221953f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_465 N_noxref_6_c_667_n N_VGND_c_872_n 0.0117314f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_466 N_noxref_6_c_618_n N_VGND_c_872_n 0.00255021f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_467 N_noxref_6_c_640_n N_VGND_c_872_n 0.00544447f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_468 N_noxref_6_c_667_n N_VGND_c_873_n 0.0117314f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_469 N_noxref_6_c_610_n N_VGND_c_873_n 0.0221953f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_470 N_noxref_6_c_679_n N_VGND_c_873_n 0.0117314f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_471 N_noxref_6_c_618_n N_VGND_c_873_n 0.00255021f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_472 N_noxref_6_c_640_n N_VGND_c_873_n 0.00544447f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_473 N_noxref_6_c_610_n N_VGND_c_874_n 0.00290993f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_474 N_noxref_6_c_679_n N_VGND_c_874_n 0.0113595f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_475 N_noxref_6_c_611_n N_VGND_c_874_n 0.00290993f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_476 N_noxref_6_c_679_n N_VGND_c_875_n 0.0117314f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_477 N_noxref_6_c_611_n N_VGND_c_875_n 0.0221755f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_478 N_noxref_6_c_618_n N_VGND_c_875_n 0.0021616f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_479 N_noxref_6_c_640_n N_VGND_c_875_n 0.00543815f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_480 N_noxref_6_c_616_n N_VGND_c_876_n 0.00222764f $X=4.765 $Y=1.19 $X2=0
+ $Y2=0
cc_481 N_noxref_6_c_617_n N_VGND_c_876_n 0.0107205f $X=4.765 $Y=1.19 $X2=0 $Y2=0
cc_482 N_noxref_6_c_618_n N_VGND_c_876_n 6.42778e-19 $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_483 N_noxref_6_c_640_n N_VGND_c_876_n 4.2528e-19 $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_484 N_noxref_6_c_646_n N_VGND_c_879_n 0.0113595f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_485 N_noxref_6_c_608_n N_VGND_c_879_n 0.00290993f $X=2.695 $Y=0.82 $X2=0
+ $Y2=0
cc_486 N_noxref_6_c_608_n N_VGND_c_881_n 0.00290993f $X=2.695 $Y=0.82 $X2=0
+ $Y2=0
cc_487 N_noxref_6_c_667_n N_VGND_c_881_n 0.0113595f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_488 N_noxref_6_c_610_n N_VGND_c_881_n 0.00290993f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_489 N_noxref_6_c_611_n N_VGND_c_884_n 0.00144667f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_490 N_noxref_6_c_846_p N_VGND_c_884_n 0.0113958f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_491 N_noxref_6_c_615_n N_VGND_c_884_n 8.77886e-19 $X=4.417 $Y=0.82 $X2=0
+ $Y2=0
cc_492 N_noxref_6_M1000_d N_VGND_c_886_n 0.00363964f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_noxref_6_M1009_d N_VGND_c_886_n 0.00231603f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_494 N_noxref_6_M1014_d N_VGND_c_886_n 0.00181772f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_495 N_noxref_6_M1017_d N_VGND_c_886_n 0.00418582f $X=4.325 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_noxref_6_c_646_n N_VGND_c_886_n 0.0064623f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_497 N_noxref_6_c_608_n N_VGND_c_886_n 0.00887359f $X=2.695 $Y=0.82 $X2=0
+ $Y2=0
cc_498 N_noxref_6_c_667_n N_VGND_c_886_n 0.0064623f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_499 N_noxref_6_c_610_n N_VGND_c_886_n 0.00887359f $X=3.535 $Y=0.82 $X2=0
+ $Y2=0
cc_500 N_noxref_6_c_679_n N_VGND_c_886_n 0.0064623f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_501 N_noxref_6_c_611_n N_VGND_c_886_n 0.00685389f $X=4.29 $Y=0.82 $X2=0 $Y2=0
cc_502 N_noxref_6_c_846_p N_VGND_c_886_n 0.00646998f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_503 N_noxref_6_c_615_n N_VGND_c_886_n 0.00218249f $X=4.417 $Y=0.82 $X2=0
+ $Y2=0
cc_504 N_noxref_6_c_618_n N_VGND_c_886_n 0.0513297f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_505 N_noxref_6_c_640_n N_VGND_c_886_n 0.0522017f $X=3.56 $Y=1.27 $X2=0 $Y2=0
cc_506 N_noxref_6_c_632_n N_VGND_c_886_n 0.0119334f $X=3.985 $Y=1.19 $X2=0 $Y2=0
cc_507 N_noxref_6_M1001_s X 0.00158966f $X=1.805 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_508 N_noxref_6_M1006_s X 0.00158966f $X=2.645 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_509 N_noxref_6_M1011_s X 0.00158966f $X=3.485 $Y=1.485 $X2=-0.19 $Y2=-0.24
cc_510 N_noxref_6_c_648_n X 0.00304954f $X=1.94 $Y=1.755 $X2=-0.19 $Y2=-0.24
cc_511 N_noxref_6_c_669_n X 0.0029886f $X=2.78 $Y=1.755 $X2=-0.19 $Y2=-0.24
cc_512 N_noxref_6_c_681_n X 0.0029886f $X=3.62 $Y=1.755 $X2=-0.19 $Y2=-0.24
cc_513 N_noxref_6_c_794_n X 0.0011968f $X=4.46 $Y=1.755 $X2=-0.19 $Y2=-0.24

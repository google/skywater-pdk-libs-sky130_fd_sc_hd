* NGSPICE file created from sky130_fd_sc_hd__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_285_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=3.575e+11p ps=3.7e+06u
M1001 VGND A2 a_285_47# VNB nshort w=650000u l=150000u
+  ad=6.5975e+11p pd=5.93e+06u as=0p ps=0u
M1002 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.19e+12p pd=1.038e+07u as=5.5e+11p ps=5.1e+06u
M1003 a_114_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u
M1004 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A1 a_114_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1011 Y B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__dfstp_1.spice.SKY130_FD_SC_HD__DFSTP_1.pxi
* Created: Thu Aug 27 14:15:15 2020
* 
x_PM_SKY130_FD_SC_HD__DFSTP_1%CLK N_CLK_c_220_n N_CLK_c_215_n N_CLK_M1028_g
+ N_CLK_c_221_n N_CLK_M1014_g N_CLK_c_216_n N_CLK_c_222_n CLK CLK N_CLK_c_218_n
+ N_CLK_c_219_n PM_SKY130_FD_SC_HD__DFSTP_1%CLK
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_27_47# N_A_27_47#_M1028_s N_A_27_47#_M1014_s
+ N_A_27_47#_M1016_g N_A_27_47#_M1000_g N_A_27_47#_c_260_n N_A_27_47#_M1024_g
+ N_A_27_47#_M1031_g N_A_27_47#_M1026_g N_A_27_47#_M1011_g N_A_27_47#_c_517_p
+ N_A_27_47#_c_261_n N_A_27_47#_c_262_n N_A_27_47#_c_276_n N_A_27_47#_c_388_p
+ N_A_27_47#_c_263_n N_A_27_47#_c_264_n N_A_27_47#_c_265_n N_A_27_47#_c_266_n
+ N_A_27_47#_c_267_n N_A_27_47#_c_268_n N_A_27_47#_c_280_n N_A_27_47#_c_269_n
+ N_A_27_47#_c_270_n N_A_27_47#_c_281_n N_A_27_47#_c_282_n N_A_27_47#_c_283_n
+ N_A_27_47#_c_284_n N_A_27_47#_c_285_n N_A_27_47#_c_271_n N_A_27_47#_c_287_n
+ N_A_27_47#_c_288_n N_A_27_47#_c_289_n N_A_27_47#_c_290_n N_A_27_47#_c_272_n
+ PM_SKY130_FD_SC_HD__DFSTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DFSTP_1%D N_D_M1005_g N_D_M1022_g D D N_D_c_535_n
+ N_D_c_536_n PM_SKY130_FD_SC_HD__DFSTP_1%D
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_193_47# N_A_193_47#_M1016_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1006_g N_A_193_47#_c_573_n N_A_193_47#_c_574_n
+ N_A_193_47#_M1015_g N_A_193_47#_c_576_n N_A_193_47#_M1009_g
+ N_A_193_47#_c_578_n N_A_193_47#_M1008_g N_A_193_47#_c_579_n
+ N_A_193_47#_c_580_n N_A_193_47#_c_581_n N_A_193_47#_c_582_n
+ N_A_193_47#_c_583_n N_A_193_47#_c_584_n N_A_193_47#_c_585_n
+ N_A_193_47#_c_586_n N_A_193_47#_c_587_n N_A_193_47#_c_588_n
+ N_A_193_47#_c_589_n N_A_193_47#_c_590_n PM_SKY130_FD_SC_HD__DFSTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_652_21# N_A_652_21#_M1003_d N_A_652_21#_M1023_d
+ N_A_652_21#_M1021_g N_A_652_21#_M1004_g N_A_652_21#_c_774_n
+ N_A_652_21#_c_858_p N_A_652_21#_c_775_n N_A_652_21#_c_769_n
+ N_A_652_21#_c_770_n N_A_652_21#_c_777_n N_A_652_21#_c_778_n
+ N_A_652_21#_c_779_n N_A_652_21#_c_771_n PM_SKY130_FD_SC_HD__DFSTP_1%A_652_21#
x_PM_SKY130_FD_SC_HD__DFSTP_1%SET_B N_SET_B_c_883_n N_SET_B_M1023_g
+ N_SET_B_M1002_g N_SET_B_M1001_g N_SET_B_M1018_g N_SET_B_c_887_n
+ N_SET_B_c_897_n N_SET_B_c_888_n N_SET_B_c_889_n SET_B N_SET_B_c_891_n
+ N_SET_B_c_892_n N_SET_B_c_959_p N_SET_B_c_893_n
+ PM_SKY130_FD_SC_HD__DFSTP_1%SET_B
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_476_47# N_A_476_47#_M1024_d N_A_476_47#_M1006_d
+ N_A_476_47#_c_1018_n N_A_476_47#_M1003_g N_A_476_47#_c_1019_n
+ N_A_476_47#_M1017_g N_A_476_47#_c_1020_n N_A_476_47#_M1013_g
+ N_A_476_47#_c_1021_n N_A_476_47#_M1019_g N_A_476_47#_c_1022_n
+ N_A_476_47#_c_1045_n N_A_476_47#_c_1051_n N_A_476_47#_c_1030_n
+ N_A_476_47#_c_1023_n N_A_476_47#_c_1024_n N_A_476_47#_c_1025_n
+ N_A_476_47#_c_1026_n N_A_476_47#_c_1027_n
+ PM_SKY130_FD_SC_HD__DFSTP_1%A_476_47#
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_1182_261# N_A_1182_261#_M1007_d
+ N_A_1182_261#_M1010_d N_A_1182_261#_M1027_g N_A_1182_261#_M1012_g
+ N_A_1182_261#_c_1177_n N_A_1182_261#_c_1182_n N_A_1182_261#_c_1183_n
+ N_A_1182_261#_c_1214_p N_A_1182_261#_c_1178_n N_A_1182_261#_c_1179_n
+ N_A_1182_261#_c_1185_n N_A_1182_261#_c_1186_n
+ PM_SKY130_FD_SC_HD__DFSTP_1%A_1182_261#
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_1032_413# N_A_1032_413#_M1009_d
+ N_A_1032_413#_M1026_d N_A_1032_413#_M1018_s N_A_1032_413#_M1007_g
+ N_A_1032_413#_M1010_g N_A_1032_413#_c_1257_n N_A_1032_413#_M1030_g
+ N_A_1032_413#_M1029_g N_A_1032_413#_c_1259_n N_A_1032_413#_c_1278_n
+ N_A_1032_413#_c_1270_n N_A_1032_413#_c_1287_n N_A_1032_413#_c_1260_n
+ N_A_1032_413#_c_1261_n N_A_1032_413#_c_1272_n N_A_1032_413#_c_1262_n
+ N_A_1032_413#_c_1273_n N_A_1032_413#_c_1274_n N_A_1032_413#_c_1362_n
+ N_A_1032_413#_c_1263_n N_A_1032_413#_c_1264_n N_A_1032_413#_c_1265_n
+ PM_SKY130_FD_SC_HD__DFSTP_1%A_1032_413#
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_1602_47# N_A_1602_47#_M1030_s
+ N_A_1602_47#_M1029_s N_A_1602_47#_M1020_g N_A_1602_47#_M1025_g
+ N_A_1602_47#_c_1420_n N_A_1602_47#_c_1421_n N_A_1602_47#_c_1422_n
+ N_A_1602_47#_c_1428_n N_A_1602_47#_c_1429_n N_A_1602_47#_c_1423_n
+ N_A_1602_47#_c_1424_n PM_SKY130_FD_SC_HD__DFSTP_1%A_1602_47#
x_PM_SKY130_FD_SC_HD__DFSTP_1%VPWR N_VPWR_M1014_d N_VPWR_M1022_s N_VPWR_M1004_d
+ N_VPWR_M1017_d N_VPWR_M1027_d N_VPWR_M1018_d N_VPWR_M1029_d N_VPWR_c_1477_n
+ N_VPWR_c_1478_n N_VPWR_c_1479_n N_VPWR_c_1480_n N_VPWR_c_1481_n
+ N_VPWR_c_1482_n VPWR VPWR N_VPWR_c_1483_n N_VPWR_c_1484_n N_VPWR_c_1485_n
+ N_VPWR_c_1486_n N_VPWR_c_1487_n N_VPWR_c_1488_n N_VPWR_c_1489_n
+ N_VPWR_c_1476_n N_VPWR_c_1491_n N_VPWR_c_1492_n N_VPWR_c_1493_n
+ N_VPWR_c_1494_n N_VPWR_c_1495_n N_VPWR_c_1496_n N_VPWR_c_1497_n
+ PM_SKY130_FD_SC_HD__DFSTP_1%VPWR
x_PM_SKY130_FD_SC_HD__DFSTP_1%A_381_47# N_A_381_47#_M1005_d N_A_381_47#_M1022_d
+ N_A_381_47#_c_1641_n N_A_381_47#_c_1646_n N_A_381_47#_c_1642_n
+ N_A_381_47#_c_1648_n N_A_381_47#_c_1644_n N_A_381_47#_c_1650_n
+ N_A_381_47#_c_1651_n PM_SKY130_FD_SC_HD__DFSTP_1%A_381_47#
x_PM_SKY130_FD_SC_HD__DFSTP_1%Q N_Q_M1020_d N_Q_M1025_d N_Q_c_1707_n
+ N_Q_c_1710_n N_Q_c_1708_n Q Q Q PM_SKY130_FD_SC_HD__DFSTP_1%Q
x_PM_SKY130_FD_SC_HD__DFSTP_1%VGND N_VGND_M1028_d N_VGND_M1005_s N_VGND_M1021_d
+ N_VGND_M1019_s N_VGND_M1001_d N_VGND_M1030_d N_VGND_c_1723_n N_VGND_c_1724_n
+ N_VGND_c_1725_n N_VGND_c_1726_n N_VGND_c_1727_n N_VGND_c_1728_n VGND VGND
+ N_VGND_c_1729_n N_VGND_c_1730_n N_VGND_c_1731_n N_VGND_c_1732_n
+ N_VGND_c_1733_n N_VGND_c_1734_n N_VGND_c_1735_n N_VGND_c_1736_n
+ N_VGND_c_1737_n N_VGND_c_1738_n N_VGND_c_1739_n N_VGND_c_1740_n
+ N_VGND_c_1741_n PM_SKY130_FD_SC_HD__DFSTP_1%VGND
cc_1 VNB N_CLK_c_215_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_216_n 0.0229857f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK 0.0187424f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_CLK_c_218_n 0.01953f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_CLK_c_219_n 0.0141141f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1016_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_260_n 0.0180458f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_8 VNB N_A_27_47#_c_261_n 0.00174761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_262_n 0.00643757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_263_n 0.00246672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_264_n 0.004477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_265_n 0.0327379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_266_n 0.00635368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_267_n 0.00811013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_268_n 0.00156998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_269_n 0.00506957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_270_n 0.0255871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_271_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_272_n 0.0159476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_M1005_g 0.0205663f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_21 VNB N_D_c_535_n 0.0258802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_D_c_536_n 0.00442451f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_23 VNB N_A_193_47#_c_573_n 0.0133397f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_24 VNB N_A_193_47#_c_574_n 0.00435992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_M1015_g 0.0199596f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_26 VNB N_A_193_47#_c_576_n 0.00878847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_M1009_g 0.0339128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_578_n 0.00977928f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_29 VNB N_A_193_47#_c_579_n 0.0187369f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_30 VNB N_A_193_47#_c_580_n 0.0191962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_581_n 0.00569477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_582_n 0.0012554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_583_n 0.0157358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_584_n 0.00235584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_585_n 0.00199889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_586_n 0.00146001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_587_n 0.00222242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_588_n 0.0249277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_589_n 0.00499852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_590_n 0.0161628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_652_21#_M1021_g 0.0422385f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_42 VNB N_A_652_21#_c_769_n 0.00136482f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_652_21#_c_770_n 0.00318738f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_44 VNB N_A_652_21#_c_771_n 0.00545975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_SET_B_c_883_n 0.0308821f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_46 VNB N_SET_B_M1023_g 0.00706345f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_47 VNB N_SET_B_M1002_g 0.0179723f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_48 VNB N_SET_B_M1001_g 0.0186416f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_49 VNB N_SET_B_c_887_n 0.00770175f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_50 VNB N_SET_B_c_888_n 0.0255769f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_51 VNB N_SET_B_c_889_n 0.00449682f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_52 VNB SET_B 0.00658023f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_53 VNB N_SET_B_c_891_n 0.0134128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_892_n 0.0020958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_893_n 0.0030779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_476_47#_c_1018_n 0.017726f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_57 VNB N_A_476_47#_c_1019_n 0.0138425f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_58 VNB N_A_476_47#_c_1020_n 0.0553275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_476_47#_c_1021_n 0.0177765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_476_47#_c_1022_n 0.00507008f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_61 VNB N_A_476_47#_c_1023_n 0.0043153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_476_47#_c_1024_n 0.00446117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_476_47#_c_1025_n 0.00392752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_476_47#_c_1026_n 0.00107462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_476_47#_c_1027_n 0.0145875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1182_261#_M1012_g 0.0377839f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_67 VNB N_A_1182_261#_c_1177_n 0.00810921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1182_261#_c_1178_n 0.00703862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1182_261#_c_1179_n 0.00490354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1032_413#_M1007_g 0.0319034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1032_413#_c_1257_n 0.03953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1032_413#_M1030_g 0.0411298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1032_413#_c_1259_n 0.00547482f $X=-0.19 $Y=-0.24 $X2=0.265
+ $Y2=1.19
cc_74 VNB N_A_1032_413#_c_1260_n 0.00479234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1032_413#_c_1261_n 0.00125329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1032_413#_c_1262_n 0.00913165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1032_413#_c_1263_n 7.5989e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1032_413#_c_1264_n 0.0124184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1032_413#_c_1265_n 0.00481971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1602_47#_c_1420_n 0.00302836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1602_47#_c_1421_n 0.0043507f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_82 VNB N_A_1602_47#_c_1422_n 0.0228329f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_83 VNB N_A_1602_47#_c_1423_n 7.97391e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1602_47#_c_1424_n 0.0197447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VPWR_c_1476_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_381_47#_c_1641_n 0.00882858f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_87 VNB N_A_381_47#_c_1642_n 0.00229891f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_88 VNB N_Q_c_1707_n 0.00479254f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_89 VNB N_Q_c_1708_n 0.0232324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB Q 0.0154962f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_91 VNB N_VGND_c_1723_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1724_n 0.00492922f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_93 VNB N_VGND_c_1725_n 0.00404464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1726_n 0.0198618f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_95 VNB N_VGND_c_1727_n 0.00985311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1728_n 0.00262294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1729_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1730_n 0.0164349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1731_n 0.0451324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1732_n 0.0303862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1733_n 0.0272431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1734_n 0.47633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1735_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1736_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1737_n 0.0056662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1738_n 0.00612673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1739_n 0.0408815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1740_n 0.0122102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1741_n 0.00427022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VPB N_CLK_c_220_n 0.0118724f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_111 VPB N_CLK_c_221_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_112 VPB N_CLK_c_222_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_113 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_114 VPB N_CLK_c_218_n 0.0100888f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_115 VPB N_A_27_47#_M1000_g 0.0364742f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_116 VPB N_A_27_47#_M1031_g 0.021588f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_117 VPB N_A_27_47#_M1026_g 0.0205628f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_118 VPB N_A_27_47#_c_276_n 0.00121034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_263_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_264_n 0.00245106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_266_n 0.00547613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_280_n 0.00355155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_281_n 0.0141666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_282_n 0.00241912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_47#_c_283_n 0.011654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_27_47#_c_284_n 0.0016702f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_285_n 0.00390757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_271_n 0.0115872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_287_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_288_n 0.00575159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_289_n 0.0281846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_290_n 0.00634002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_D_M1022_g 0.0293669f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_134 VPB N_D_c_535_n 0.00538482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_D_c_536_n 0.00459652f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_136 VPB N_A_193_47#_M1006_g 0.0466922f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_137 VPB N_A_193_47#_c_573_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_138 VPB N_A_193_47#_c_574_n 0.00328709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_193_47#_c_578_n 0.0116784f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_140 VPB N_A_193_47#_M1008_g 0.0394871f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_141 VPB N_A_193_47#_c_579_n 0.0122605f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_142 VPB N_A_193_47#_c_587_n 0.00217849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_193_47#_c_590_n 0.0183602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_652_21#_M1021_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_145 VPB N_A_652_21#_M1004_g 0.0208799f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_146 VPB N_A_652_21#_c_774_n 0.00189033f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_147 VPB N_A_652_21#_c_775_n 0.00247793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_652_21#_c_770_n 0.0027381f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_149 VPB N_A_652_21#_c_777_n 0.00460198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_652_21#_c_778_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_151 VPB N_A_652_21#_c_779_n 0.00112185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_SET_B_M1023_g 0.0474843f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_153 VPB N_SET_B_M1018_g 0.038305f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_154 VPB N_SET_B_c_887_n 0.0123607f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_155 VPB N_SET_B_c_897_n 0.00992356f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_156 VPB N_A_476_47#_M1017_g 0.0334449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_476_47#_M1013_g 0.0324152f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_158 VPB N_A_476_47#_c_1030_n 0.0121057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_476_47#_c_1024_n 0.00542515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_476_47#_c_1025_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_476_47#_c_1026_n 0.00262972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_476_47#_c_1027_n 0.0308068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_1182_261#_M1027_g 0.0268094f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_164 VPB N_A_1182_261#_c_1177_n 0.0277544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1182_261#_c_1182_n 0.0164657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1182_261#_c_1183_n 0.0160465f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_167 VPB N_A_1182_261#_c_1178_n 0.00309392f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1182_261#_c_1185_n 0.018178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_1182_261#_c_1186_n 0.008614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1032_413#_M1010_g 0.0263696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_1032_413#_c_1257_n 0.029899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1032_413#_M1029_g 0.0408779f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_173 VPB N_A_1032_413#_c_1259_n 0.00428118f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.19
cc_174 VPB N_A_1032_413#_c_1270_n 0.00422026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1032_413#_c_1260_n 0.00190145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1032_413#_c_1272_n 0.0150397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1032_413#_c_1273_n 0.0037282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1032_413#_c_1274_n 2.86428e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1032_413#_c_1263_n 2.77041e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1032_413#_c_1264_n 0.00840405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_1032_413#_c_1265_n 0.0046931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1602_47#_M1025_g 0.0226675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1602_47#_c_1421_n 0.0044838f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_184 VPB N_A_1602_47#_c_1422_n 0.00502506f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_185 VPB N_A_1602_47#_c_1428_n 0.00606637f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.19
cc_186 VPB N_A_1602_47#_c_1429_n 0.00377036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1477_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_188 VPB N_VPWR_c_1478_n 0.00578936f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_189 VPB N_VPWR_c_1479_n 0.0114969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1480_n 3.97306e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1481_n 0.00366994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1482_n 0.00289339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1483_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1484_n 0.0163072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1485_n 0.0416374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1486_n 0.0313047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1487_n 0.01851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1488_n 0.0303512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1489_n 0.0277678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1476_n 0.0824326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1491_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1492_n 0.00507833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1493_n 0.0091704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1494_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1495_n 0.011387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1496_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1497_n 0.00427244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_381_47#_c_1641_n 0.00799498f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_209 VPB N_A_381_47#_c_1644_n 0.00185682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_Q_c_1710_n 0.00479254f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_211 VPB N_Q_c_1708_n 0.0150909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB Q 0.0208614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 N_CLK_c_215_n N_A_27_47#_M1016_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_214 CLK N_A_27_47#_M1016_g 3.09846e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_215 N_CLK_c_219_n N_A_27_47#_M1016_g 0.00508029f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_216 N_CLK_c_222_n N_A_27_47#_M1000_g 0.0276478f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_217 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_218 N_CLK_c_218_n N_A_27_47#_M1000_g 0.00530924f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_219 N_CLK_c_215_n N_A_27_47#_c_261_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_220 N_CLK_c_216_n N_A_27_47#_c_261_n 0.00787672f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_221 CLK N_A_27_47#_c_261_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_222 N_CLK_c_216_n N_A_27_47#_c_262_n 0.0059979f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_223 CLK N_A_27_47#_c_262_n 0.014414f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_224 N_CLK_c_218_n N_A_27_47#_c_262_n 3.2891e-19 $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_225 N_CLK_c_221_n N_A_27_47#_c_276_n 0.0128144f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_226 N_CLK_c_222_n N_A_27_47#_c_276_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_227 CLK N_A_27_47#_c_276_n 0.00728212f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_228 N_CLK_c_216_n N_A_27_47#_c_263_n 0.00189711f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_229 N_CLK_c_222_n N_A_27_47#_c_263_n 0.00440146f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_230 CLK N_A_27_47#_c_263_n 0.0517133f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_231 N_CLK_c_218_n N_A_27_47#_c_263_n 9.99252e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_232 N_CLK_c_219_n N_A_27_47#_c_263_n 0.00246929f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_233 N_CLK_c_221_n N_A_27_47#_c_280_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_234 N_CLK_c_222_n N_A_27_47#_c_280_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_235 CLK N_A_27_47#_c_280_n 0.0153363f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_236 N_CLK_c_218_n N_A_27_47#_c_280_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_237 N_CLK_c_221_n N_A_27_47#_c_282_n 0.00103212f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_238 CLK N_A_27_47#_c_271_n 0.00161876f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_239 N_CLK_c_218_n N_A_27_47#_c_271_n 0.0169694f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_240 N_CLK_c_221_n N_VPWR_c_1477_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_241 N_CLK_c_221_n N_VPWR_c_1483_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_221_n N_VPWR_c_1476_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_243 N_CLK_c_215_n N_VGND_c_1723_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_244 N_CLK_c_215_n N_VGND_c_1729_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_245 N_CLK_c_216_n N_VGND_c_1729_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_246 N_CLK_c_215_n N_VGND_c_1734_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_260_n N_D_M1005_g 0.0210908f $X=2.305 $Y=0.705 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_264_n N_D_M1005_g 0.00120175f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_288_n N_D_M1022_g 7.92917e-19 $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_264_n N_D_c_535_n 0.00106119f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_265_n N_D_c_535_n 0.00155965f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_264_n N_D_c_536_n 0.0453933f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_265_n N_D_c_536_n 2.37218e-19 $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_281_n N_D_c_536_n 0.00575757f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_288_n N_D_c_536_n 0.00408526f $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_281_n N_A_193_47#_M1000_d 6.81311e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1031_g N_A_193_47#_M1006_g 0.0190899f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_264_n N_A_193_47#_M1006_g 0.00534395f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_281_n N_A_193_47#_M1006_g 0.00702647f $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_284_n N_A_193_47#_M1006_g 5.24592e-19 $X=2.7 $Y=1.87 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_287_n N_A_193_47#_M1006_g 0.0174486f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_288_n N_A_193_47#_M1006_g 0.0104483f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_264_n N_A_193_47#_c_573_n 0.010154f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_283_n N_A_193_47#_c_573_n 3.83457e-19 $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_287_n N_A_193_47#_c_573_n 0.0212221f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_288_n N_A_193_47#_c_573_n 0.00654686f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_264_n N_A_193_47#_c_574_n 0.00204176f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_265_n N_A_193_47#_c_574_n 0.0232669f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_260_n N_A_193_47#_M1015_g 0.0128107f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_264_n N_A_193_47#_M1015_g 4.45841e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_265_n N_A_193_47#_M1015_g 0.0214266f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_266_n N_A_193_47#_M1009_g 0.00410946f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_c_267_n N_A_193_47#_M1009_g 0.011907f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_269_n N_A_193_47#_M1009_g 0.00270619f $X=5.985 $Y=0.81 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_270_n N_A_193_47#_M1009_g 0.020941f $X=5.985 $Y=0.93 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_272_n N_A_193_47#_M1009_g 0.0125268f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_267_n N_A_193_47#_c_578_n 2.6295e-19 $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1026_g N_A_193_47#_M1008_g 0.0175641f $X=5.085 $Y=2.275 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_266_n N_A_193_47#_M1008_g 0.00215568f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_280 N_A_27_47#_c_285_n N_A_193_47#_M1008_g 0.00442284f $X=5.335 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_289_n N_A_193_47#_M1008_g 0.0159766f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_290_n N_A_193_47#_M1008_g 0.00180554f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_266_n N_A_193_47#_c_579_n 0.0035853f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_267_n N_A_193_47#_c_579_n 0.00337501f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_285_n N_A_193_47#_c_579_n 8.69467e-19 $X=5.335 $Y=1.87 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_289_n N_A_193_47#_c_579_n 0.0106619f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_290_n N_A_193_47#_c_579_n 0.00101144f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_264_n N_A_193_47#_c_580_n 0.0173333f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_265_n N_A_193_47#_c_580_n 0.0059767f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1016_g N_A_193_47#_c_581_n 0.00654297f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_261_n N_A_193_47#_c_581_n 0.00215348f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_263_n N_A_193_47#_c_581_n 0.00507209f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_c_264_n N_A_193_47#_c_582_n 0.00934078f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_266_n N_A_193_47#_c_583_n 0.0118781f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_267_n N_A_193_47#_c_583_n 0.00166232f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_289_n N_A_193_47#_c_583_n 9.1133e-19 $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_290_n N_A_193_47#_c_583_n 0.00282033f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_283_n N_A_193_47#_c_584_n 0.0952174f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_264_n N_A_193_47#_c_585_n 4.74166e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_266_n N_A_193_47#_c_586_n 0.00254764f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_301 N_A_27_47#_c_267_n N_A_193_47#_c_586_n 0.00143429f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_285_n N_A_193_47#_c_586_n 0.0144457f $X=5.335 $Y=1.87 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_290_n N_A_193_47#_c_586_n 0.00167414f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_266_n N_A_193_47#_c_587_n 0.0285066f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_267_n N_A_193_47#_c_587_n 0.0123872f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_285_n N_A_193_47#_c_587_n 6.9568e-19 $X=5.335 $Y=1.87 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_289_n N_A_193_47#_c_587_n 6.19272e-19 $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_290_n N_A_193_47#_c_587_n 0.0119993f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_264_n N_A_193_47#_c_588_n 0.00674133f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_260_n N_A_193_47#_c_589_n 5.14023e-19 $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_264_n N_A_193_47#_c_589_n 0.0210004f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_265_n N_A_193_47#_c_589_n 0.00154674f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_287_n N_A_193_47#_c_589_n 3.18577e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_288_n N_A_193_47#_c_589_n 0.00339609f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_M1016_g N_A_193_47#_c_590_n 0.0272829f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_261_n N_A_193_47#_c_590_n 0.011891f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_388_p N_A_193_47#_c_590_n 0.00826851f $X=0.725 $Y=1.795
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_c_263_n N_A_193_47#_c_590_n 0.0701354f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_281_n N_A_193_47#_c_590_n 0.0247331f $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_282_n N_A_193_47#_c_590_n 0.00185693f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_264_n N_A_652_21#_M1021_g 5.35023e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_283_n N_A_652_21#_M1004_g 0.00197541f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_283_n N_A_652_21#_c_774_n 0.0147195f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_M1026_g N_A_652_21#_c_775_n 6.97636e-19 $X=5.085 $Y=2.275
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_283_n N_A_652_21#_c_775_n 0.022507f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_285_n N_A_652_21#_c_775_n 9.07105e-19 $X=5.335 $Y=1.87 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_290_n N_A_652_21#_c_775_n 0.00938889f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_266_n N_A_652_21#_c_770_n 0.0421767f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_283_n N_A_652_21#_c_770_n 0.00751374f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_289_n N_A_652_21#_c_770_n 2.32128e-19 $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_290_n N_A_652_21#_c_770_n 0.0137093f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_283_n N_A_652_21#_c_777_n 0.0157473f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_M1031_g N_A_652_21#_c_778_n 0.0161874f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_283_n N_A_652_21#_c_778_n 0.00193898f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_287_n N_A_652_21#_c_778_n 0.00927772f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_283_n N_A_652_21#_c_779_n 0.00782494f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_266_n N_A_652_21#_c_771_n 0.0133315f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_268_n N_A_652_21#_c_771_n 0.0121229f $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_283_n N_SET_B_M1023_g 0.00205491f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_266_n N_SET_B_c_891_n 0.00399047f $X=4.985 $Y=1.655 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_267_n N_SET_B_c_891_n 0.0293235f $X=5.82 $Y=0.81 $X2=0 $Y2=0
cc_342 N_A_27_47#_c_268_n N_SET_B_c_891_n 0.00574094f $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_269_n N_SET_B_c_891_n 0.0167082f $X=5.985 $Y=0.81 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_266_n N_A_476_47#_c_1019_n 2.85114e-19 $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_283_n N_A_476_47#_M1017_g 0.00187886f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_266_n N_A_476_47#_c_1020_n 0.00470216f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_267_n N_A_476_47#_c_1020_n 0.00749989f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_268_n N_A_476_47#_c_1020_n 0.00602324f $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_289_n N_A_476_47#_c_1020_n 0.00228641f $X=5.175 $Y=1.74
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_283_n N_A_476_47#_M1013_g 0.00241494f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_289_n N_A_476_47#_M1013_g 0.0565606f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_290_n N_A_476_47#_M1013_g 0.00171839f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_267_n N_A_476_47#_c_1021_n 0.00413822f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_M1031_g N_A_476_47#_c_1045_n 0.00904177f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_281_n N_A_476_47#_c_1045_n 2.09728e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_283_n N_A_476_47#_c_1045_n 0.00506942f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_284_n N_A_476_47#_c_1045_n 0.00303545f $X=2.7 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_287_n N_A_476_47#_c_1045_n 0.00186639f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_288_n N_A_476_47#_c_1045_n 0.0152514f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_264_n N_A_476_47#_c_1051_n 0.00676006f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_265_n N_A_476_47#_c_1051_n 9.25786e-19 $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_M1031_g N_A_476_47#_c_1030_n 0.00650943f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_264_n N_A_476_47#_c_1030_n 0.00666284f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_283_n N_A_476_47#_c_1030_n 0.013911f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_284_n N_A_476_47#_c_1030_n 0.00149623f $X=2.7 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_287_n N_A_476_47#_c_1030_n 0.00203066f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_c_288_n N_A_476_47#_c_1030_n 0.0282877f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_283_n N_A_476_47#_c_1024_n 0.00472657f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_264_n N_A_476_47#_c_1025_n 0.00728915f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_283_n N_A_476_47#_c_1025_n 0.00456576f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_283_n N_A_476_47#_c_1026_n 0.00248872f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_266_n N_A_476_47#_c_1027_n 0.00628168f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_283_n N_A_476_47#_c_1027_n 0.00148193f $X=5.19 $Y=1.87 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_269_n N_A_1182_261#_M1012_g 8.41348e-19 $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_272_n N_A_1182_261#_M1012_g 0.0628006f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_269_n N_A_1182_261#_c_1177_n 3.76765e-19 $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_270_n N_A_1182_261#_c_1177_n 0.0136804f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_M1026_g N_A_1032_413#_c_1278_n 0.00503271f $X=5.085 $Y=2.275
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_283_n N_A_1032_413#_c_1278_n 2.55921e-19 $X=5.19 $Y=1.87
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_285_n N_A_1032_413#_c_1278_n 0.00456317f $X=5.335 $Y=1.87
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_289_n N_A_1032_413#_c_1278_n 9.00165e-19 $X=5.175 $Y=1.74
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_290_n N_A_1032_413#_c_1278_n 0.0149056f $X=5.175 $Y=1.74
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_266_n N_A_1032_413#_c_1270_n 0.00537793f $X=4.985 $Y=1.655
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_285_n N_A_1032_413#_c_1270_n 0.00798359f $X=5.335 $Y=1.87
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_c_289_n N_A_1032_413#_c_1270_n 4.1977e-19 $X=5.175 $Y=1.74
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_290_n N_A_1032_413#_c_1270_n 0.0211007f $X=5.175 $Y=1.74
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_267_n N_A_1032_413#_c_1287_n 0.00680222f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_269_n N_A_1032_413#_c_1287_n 0.0126727f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_270_n N_A_1032_413#_c_1287_n 5.72459e-19 $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_272_n N_A_1032_413#_c_1287_n 0.00790984f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_267_n N_A_1032_413#_c_1260_n 0.00194166f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_269_n N_A_1032_413#_c_1260_n 0.0183126f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_c_270_n N_A_1032_413#_c_1260_n 0.00282863f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_267_n N_A_1032_413#_c_1261_n 0.00583458f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_269_n N_A_1032_413#_c_1262_n 0.0218685f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_270_n N_A_1032_413#_c_1262_n 0.00156489f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_272_n N_A_1032_413#_c_1262_n 0.00248854f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_M1026_g N_A_1032_413#_c_1274_n 0.0010081f $X=5.085 $Y=2.275
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_388_p N_VPWR_M1014_d 6.91013e-19 $X=0.725 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_400 N_A_27_47#_c_282_n N_VPWR_M1014_d 0.00195102f $X=0.84 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_401 N_A_27_47#_M1000_g N_VPWR_c_1477_n 0.00827983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_276_n N_VPWR_c_1477_n 0.00355272f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_388_p N_VPWR_c_1477_n 0.0133497f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_280_n N_VPWR_c_1477_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_405 N_A_27_47#_c_282_n N_VPWR_c_1477_n 0.00347913f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_M1000_g N_VPWR_c_1478_n 0.00190407f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_281_n N_VPWR_c_1478_n 0.00166908f $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_M1026_g N_VPWR_c_1480_n 0.00190036f $X=5.085 $Y=2.275 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_283_n N_VPWR_c_1480_n 0.001212f $X=5.19 $Y=1.87 $X2=0 $Y2=0
cc_410 N_A_27_47#_c_276_n N_VPWR_c_1483_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_411 N_A_27_47#_c_280_n N_VPWR_c_1483_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_412 N_A_27_47#_M1000_g N_VPWR_c_1484_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_M1031_g N_VPWR_c_1485_n 0.00367119f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_M1026_g N_VPWR_c_1486_n 0.00427125f $X=5.085 $Y=2.275 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_290_n N_VPWR_c_1486_n 0.0032218f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_M1000_g N_VPWR_c_1476_n 0.00536257f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_M1031_g N_VPWR_c_1476_n 0.00562272f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_M1026_g N_VPWR_c_1476_n 0.00582964f $X=5.085 $Y=2.275 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_276_n N_VPWR_c_1476_n 0.00396423f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_280_n N_VPWR_c_1476_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_281_n N_VPWR_c_1476_n 0.0735427f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_422 N_A_27_47#_c_282_n N_VPWR_c_1476_n 0.0144757f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_423 N_A_27_47#_c_283_n N_VPWR_c_1476_n 0.112922f $X=5.19 $Y=1.87 $X2=0 $Y2=0
cc_424 N_A_27_47#_c_284_n N_VPWR_c_1476_n 0.0160117f $X=2.7 $Y=1.87 $X2=0 $Y2=0
cc_425 N_A_27_47#_c_285_n N_VPWR_c_1476_n 0.016077f $X=5.335 $Y=1.87 $X2=0 $Y2=0
cc_426 N_A_27_47#_c_288_n N_VPWR_c_1476_n 3.19863e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_290_n N_VPWR_c_1476_n 0.00251853f $X=5.175 $Y=1.74 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_283_n N_VPWR_c_1493_n 0.0014214f $X=5.19 $Y=1.87 $X2=0 $Y2=0
cc_429 N_A_27_47#_c_281_n N_A_381_47#_M1022_d 8.84929e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_260_n N_A_381_47#_c_1646_n 0.00225228f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_264_n N_A_381_47#_c_1646_n 0.00713576f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_281_n N_A_381_47#_c_1648_n 0.019313f $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_281_n N_A_381_47#_c_1644_n 0.0157335f $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_260_n N_A_381_47#_c_1650_n 0.00399753f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_281_n N_A_381_47#_c_1651_n 0.0109514f $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_284_n N_A_381_47#_c_1651_n 0.00154103f $X=2.7 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_288_n N_A_381_47#_c_1651_n 0.00827849f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_261_n N_VGND_M1028_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_439 N_A_27_47#_M1016_g N_VGND_c_1723_n 0.0078844f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_c_261_n N_VGND_c_1723_n 0.0170164f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_441 N_A_27_47#_c_271_n N_VGND_c_1723_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_M1016_g N_VGND_c_1724_n 0.00296522f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_260_n N_VGND_c_1724_n 0.00120909f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_267_n N_VGND_c_1727_n 3.70426e-19 $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_268_n N_VGND_c_1727_n 0.0129707f $X=5.07 $Y=0.81 $X2=0 $Y2=0
cc_446 N_A_27_47#_c_517_p N_VGND_c_1729_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_261_n N_VGND_c_1729_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_M1016_g N_VGND_c_1730_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_260_n N_VGND_c_1731_n 0.00556304f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_264_n N_VGND_c_1731_n 0.00113905f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_265_n N_VGND_c_1731_n 2.48118e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_M1028_s N_VGND_c_1734_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1016_g N_VGND_c_1734_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_260_n N_VGND_c_1734_n 0.00678262f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_517_p N_VGND_c_1734_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_261_n N_VGND_c_1734_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_264_n N_VGND_c_1734_n 0.00122477f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_267_n N_VGND_c_1734_n 0.00610914f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_268_n N_VGND_c_1734_n 4.92512e-19 $X=5.07 $Y=0.81 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_272_n N_VGND_c_1734_n 0.00522127f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_267_n N_VGND_c_1739_n 0.00797153f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_272_n N_VGND_c_1739_n 0.00368123f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_463 N_D_M1022_g N_A_193_47#_c_574_n 0.0303627f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_464 N_D_c_535_n N_A_193_47#_c_574_n 0.00467503f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_465 N_D_c_536_n N_A_193_47#_c_574_n 0.00330794f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_466 N_D_M1005_g N_A_193_47#_c_580_n 0.00395556f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_467 N_D_c_535_n N_A_193_47#_c_580_n 8.88354e-19 $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_468 N_D_c_536_n N_A_193_47#_c_580_n 0.0127149f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_469 N_D_M1005_g N_A_193_47#_c_590_n 0.00372305f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_470 N_D_M1022_g N_A_193_47#_c_590_n 0.00471318f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_471 N_D_M1022_g N_VPWR_c_1478_n 0.0116766f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_472 N_D_M1022_g N_VPWR_c_1485_n 0.0035268f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_473 N_D_M1022_g N_VPWR_c_1476_n 0.00402871f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_474 N_D_M1005_g N_A_381_47#_c_1641_n 0.00557005f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_475 N_D_M1022_g N_A_381_47#_c_1641_n 0.0115166f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_476 N_D_c_535_n N_A_381_47#_c_1641_n 0.00753248f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_477 N_D_c_536_n N_A_381_47#_c_1641_n 0.0473419f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_478 N_D_M1005_g N_A_381_47#_c_1646_n 0.0126635f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_479 N_D_c_535_n N_A_381_47#_c_1646_n 0.0014463f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_480 N_D_c_536_n N_A_381_47#_c_1646_n 0.0217898f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_481 N_D_M1022_g N_A_381_47#_c_1648_n 0.011823f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_482 N_D_c_536_n N_A_381_47#_c_1648_n 0.0109323f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_483 N_D_c_536_n N_A_381_47#_c_1651_n 0.0137404f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_484 N_D_M1005_g N_VGND_c_1724_n 0.00942273f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_485 N_D_M1005_g N_VGND_c_1731_n 0.00339367f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_486 N_D_M1005_g N_VGND_c_1734_n 0.00393034f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_487 N_A_193_47#_M1015_g N_A_652_21#_M1021_g 0.0245694f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_488 N_A_193_47#_c_576_n N_A_652_21#_M1021_g 0.0105189f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_489 N_A_193_47#_c_583_n N_A_652_21#_M1021_g 7.74803e-19 $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_490 N_A_193_47#_c_585_n N_A_652_21#_M1021_g 0.00642269f $X=3.015 $Y=0.85
+ $X2=0 $Y2=0
cc_491 N_A_193_47#_c_588_n N_A_652_21#_M1021_g 0.0200662f $X=2.915 $Y=0.93 $X2=0
+ $Y2=0
cc_492 N_A_193_47#_c_589_n N_A_652_21#_M1021_g 0.00189958f $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_493 N_A_193_47#_c_583_n N_A_652_21#_c_774_n 5.47854e-19 $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_494 N_A_193_47#_c_583_n N_A_652_21#_c_775_n 0.00115455f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_495 N_A_193_47#_c_583_n N_A_652_21#_c_770_n 0.0150994f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_496 N_A_193_47#_c_583_n N_A_652_21#_c_777_n 8.37667e-19 $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_497 N_A_193_47#_c_583_n N_A_652_21#_c_771_n 0.00658398f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_498 N_A_193_47#_c_583_n N_SET_B_c_883_n 0.00386718f $X=5.19 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_499 N_A_193_47#_c_583_n N_SET_B_M1023_g 0.00121673f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_500 N_A_193_47#_c_583_n SET_B 0.00617024f $X=5.19 $Y=1.19 $X2=0 $Y2=0
cc_501 N_A_193_47#_M1009_g N_SET_B_c_891_n 0.00472752f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_502 N_A_193_47#_c_579_n N_SET_B_c_891_n 6.41485e-19 $X=5.49 $Y=1.26 $X2=0
+ $Y2=0
cc_503 N_A_193_47#_c_583_n N_SET_B_c_891_n 0.0876451f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_504 N_A_193_47#_c_586_n N_SET_B_c_891_n 0.02693f $X=5.335 $Y=1.19 $X2=0 $Y2=0
cc_505 N_A_193_47#_c_587_n N_SET_B_c_891_n 0.00112669f $X=5.335 $Y=1.19 $X2=0
+ $Y2=0
cc_506 N_A_193_47#_c_583_n N_SET_B_c_892_n 0.026499f $X=5.19 $Y=1.19 $X2=0 $Y2=0
cc_507 N_A_193_47#_c_583_n N_A_476_47#_c_1019_n 0.00253485f $X=5.19 $Y=1.19
+ $X2=0 $Y2=0
cc_508 N_A_193_47#_c_579_n N_A_476_47#_c_1020_n 0.00775418f $X=5.49 $Y=1.26
+ $X2=0 $Y2=0
cc_509 N_A_193_47#_c_583_n N_A_476_47#_c_1020_n 0.00107838f $X=5.19 $Y=1.19
+ $X2=0 $Y2=0
cc_510 N_A_193_47#_c_587_n N_A_476_47#_c_1020_n 2.11256e-19 $X=5.335 $Y=1.19
+ $X2=0 $Y2=0
cc_511 N_A_193_47#_M1009_g N_A_476_47#_c_1021_n 0.0518139f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_193_47#_M1006_g N_A_476_47#_c_1045_n 0.00285915f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_513 N_A_193_47#_M1015_g N_A_476_47#_c_1051_n 0.00883573f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_514 N_A_193_47#_c_580_n N_A_476_47#_c_1051_n 0.00579266f $X=2.87 $Y=0.85
+ $X2=0 $Y2=0
cc_515 N_A_193_47#_c_585_n N_A_476_47#_c_1051_n 0.00257401f $X=3.015 $Y=0.85
+ $X2=0 $Y2=0
cc_516 N_A_193_47#_c_588_n N_A_476_47#_c_1051_n 5.24878e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_517 N_A_193_47#_c_589_n N_A_476_47#_c_1051_n 0.0194937f $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_518 N_A_193_47#_M1006_g N_A_476_47#_c_1030_n 8.73767e-19 $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_519 N_A_193_47#_c_584_n N_A_476_47#_c_1030_n 3.03433e-19 $X=3.16 $Y=1.19
+ $X2=0 $Y2=0
cc_520 N_A_193_47#_M1015_g N_A_476_47#_c_1023_n 0.00119254f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_c_576_n N_A_476_47#_c_1023_n 8.54957e-19 $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_522 N_A_193_47#_c_583_n N_A_476_47#_c_1023_n 0.0145635f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_523 N_A_193_47#_c_585_n N_A_476_47#_c_1023_n 0.0138897f $X=3.015 $Y=0.85
+ $X2=0 $Y2=0
cc_524 N_A_193_47#_c_588_n N_A_476_47#_c_1023_n 7.78235e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_525 N_A_193_47#_c_589_n N_A_476_47#_c_1023_n 0.0244377f $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_526 N_A_193_47#_c_583_n N_A_476_47#_c_1024_n 0.0232188f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_c_576_n N_A_476_47#_c_1025_n 0.00268952f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_528 N_A_193_47#_c_583_n N_A_476_47#_c_1025_n 0.0109965f $X=5.19 $Y=1.19 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_c_584_n N_A_476_47#_c_1025_n 0.00666557f $X=3.16 $Y=1.19
+ $X2=0 $Y2=0
cc_530 N_A_193_47#_c_588_n N_A_476_47#_c_1025_n 5.70846e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_531 N_A_193_47#_c_589_n N_A_476_47#_c_1025_n 0.0053097f $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_532 N_A_193_47#_c_583_n N_A_476_47#_c_1026_n 0.00996075f $X=5.19 $Y=1.19
+ $X2=0 $Y2=0
cc_533 N_A_193_47#_c_578_n N_A_476_47#_c_1027_n 5.50204e-19 $X=5.625 $Y=1.455
+ $X2=0 $Y2=0
cc_534 N_A_193_47#_c_579_n N_A_476_47#_c_1027_n 0.00447301f $X=5.49 $Y=1.26
+ $X2=0 $Y2=0
cc_535 N_A_193_47#_c_583_n N_A_476_47#_c_1027_n 0.00376918f $X=5.19 $Y=1.19
+ $X2=0 $Y2=0
cc_536 N_A_193_47#_M1009_g N_A_1182_261#_M1012_g 0.00242755f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_c_578_n N_A_1182_261#_c_1177_n 0.0407077f $X=5.625 $Y=1.455
+ $X2=0 $Y2=0
cc_538 N_A_193_47#_M1008_g N_A_1182_261#_c_1182_n 0.0407077f $X=5.625 $Y=2.275
+ $X2=0 $Y2=0
cc_539 N_A_193_47#_M1008_g N_A_1032_413#_c_1278_n 0.00768489f $X=5.625 $Y=2.275
+ $X2=0 $Y2=0
cc_540 N_A_193_47#_c_578_n N_A_1032_413#_c_1270_n 0.00103911f $X=5.625 $Y=1.455
+ $X2=0 $Y2=0
cc_541 N_A_193_47#_M1008_g N_A_1032_413#_c_1270_n 0.0101633f $X=5.625 $Y=2.275
+ $X2=0 $Y2=0
cc_542 N_A_193_47#_c_587_n N_A_1032_413#_c_1270_n 0.00496139f $X=5.335 $Y=1.19
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_c_578_n N_A_1032_413#_c_1261_n 0.00804748f $X=5.625 $Y=1.455
+ $X2=0 $Y2=0
cc_544 N_A_193_47#_c_586_n N_A_1032_413#_c_1261_n 0.00202294f $X=5.335 $Y=1.19
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_587_n N_A_1032_413#_c_1261_n 0.0123091f $X=5.335 $Y=1.19
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_M1008_g N_A_1032_413#_c_1272_n 2.49577e-19 $X=5.625 $Y=2.275
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_M1009_g N_A_1032_413#_c_1262_n 0.00203086f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_M1008_g N_A_1032_413#_c_1274_n 0.0116631f $X=5.625 $Y=2.275
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_590_n N_VPWR_c_1477_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_550 N_A_193_47#_M1006_g N_VPWR_c_1478_n 0.00113058f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_551 N_A_193_47#_c_590_n N_VPWR_c_1478_n 0.0226552f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_552 N_A_193_47#_c_590_n N_VPWR_c_1484_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_553 N_A_193_47#_M1006_g N_VPWR_c_1485_n 0.00541732f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_554 N_A_193_47#_M1008_g N_VPWR_c_1486_n 0.00369426f $X=5.625 $Y=2.275 $X2=0
+ $Y2=0
cc_555 N_A_193_47#_M1006_g N_VPWR_c_1476_n 0.00632491f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_556 N_A_193_47#_M1008_g N_VPWR_c_1476_n 0.00544628f $X=5.625 $Y=2.275 $X2=0
+ $Y2=0
cc_557 N_A_193_47#_c_590_n N_VPWR_c_1476_n 0.00409094f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_558 N_A_193_47#_M1008_g N_VPWR_c_1495_n 0.00197636f $X=5.625 $Y=2.275 $X2=0
+ $Y2=0
cc_559 N_A_193_47#_c_580_n N_A_381_47#_M1005_d 4.25819e-19 $X=2.87 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_560 N_A_193_47#_c_580_n N_A_381_47#_c_1641_n 0.0148354f $X=2.87 $Y=0.85 $X2=0
+ $Y2=0
cc_561 N_A_193_47#_c_581_n N_A_381_47#_c_1641_n 0.00136171f $X=1.3 $Y=0.85 $X2=0
+ $Y2=0
cc_562 N_A_193_47#_c_590_n N_A_381_47#_c_1641_n 0.0675451f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_563 N_A_193_47#_c_580_n N_A_381_47#_c_1646_n 0.0198802f $X=2.87 $Y=0.85 $X2=0
+ $Y2=0
cc_564 N_A_193_47#_c_589_n N_A_381_47#_c_1646_n 0.0019894f $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_565 N_A_193_47#_c_580_n N_A_381_47#_c_1642_n 0.00435863f $X=2.87 $Y=0.85
+ $X2=0 $Y2=0
cc_566 N_A_193_47#_c_581_n N_A_381_47#_c_1642_n 0.00141243f $X=1.3 $Y=0.85 $X2=0
+ $Y2=0
cc_567 N_A_193_47#_c_590_n N_A_381_47#_c_1642_n 0.0138319f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_568 N_A_193_47#_c_590_n N_A_381_47#_c_1644_n 0.0114342f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_569 N_A_193_47#_M1006_g N_A_381_47#_c_1651_n 0.0102511f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_570 N_A_193_47#_c_580_n N_VGND_c_1724_n 0.0012296f $X=2.87 $Y=0.85 $X2=0
+ $Y2=0
cc_571 N_A_193_47#_c_590_n N_VGND_c_1724_n 0.00823827f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_572 N_A_193_47#_c_590_n N_VGND_c_1730_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_573 N_A_193_47#_M1015_g N_VGND_c_1731_n 0.00359964f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_574 N_A_193_47#_M1016_d N_VGND_c_1734_n 0.0033946f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_575 N_A_193_47#_M1015_g N_VGND_c_1734_n 0.00564268f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_576 N_A_193_47#_M1009_g N_VGND_c_1734_n 0.00571363f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_577 N_A_193_47#_c_580_n N_VGND_c_1734_n 0.0731727f $X=2.87 $Y=0.85 $X2=0
+ $Y2=0
cc_578 N_A_193_47#_c_581_n N_VGND_c_1734_n 0.0151433f $X=1.3 $Y=0.85 $X2=0 $Y2=0
cc_579 N_A_193_47#_c_585_n N_VGND_c_1734_n 0.0153531f $X=3.015 $Y=0.85 $X2=0
+ $Y2=0
cc_580 N_A_193_47#_c_590_n N_VGND_c_1734_n 0.00372614f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_581 N_A_193_47#_M1009_g N_VGND_c_1739_n 0.00437852f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_582 N_A_193_47#_c_589_n A_586_47# 0.00109904f $X=2.915 $Y=0.93 $X2=-0.19
+ $Y2=-0.24
cc_583 N_A_652_21#_M1021_g N_SET_B_c_883_n 0.0189903f $X=3.335 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_584 N_A_652_21#_c_770_n N_SET_B_c_883_n 7.68518e-19 $X=4.635 $Y=1.835
+ $X2=-0.19 $Y2=-0.24
cc_585 N_A_652_21#_M1021_g N_SET_B_M1023_g 0.0137896f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_586 N_A_652_21#_M1004_g N_SET_B_M1023_g 0.0113783f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_587 N_A_652_21#_c_774_n N_SET_B_M1023_g 0.0139954f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_588 N_A_652_21#_c_777_n N_SET_B_M1023_g 0.00563707f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_589 N_A_652_21#_c_778_n N_SET_B_M1023_g 0.0201938f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_590 N_A_652_21#_M1021_g N_SET_B_M1002_g 0.0141659f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_591 N_A_652_21#_c_769_n N_SET_B_M1002_g 0.00124922f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_592 N_A_652_21#_c_771_n N_SET_B_M1002_g 3.79959e-19 $X=4.635 $Y=0.895 $X2=0
+ $Y2=0
cc_593 N_A_652_21#_M1021_g SET_B 0.00110794f $X=3.335 $Y=0.445 $X2=0 $Y2=0
cc_594 N_A_652_21#_c_771_n SET_B 0.0144301f $X=4.635 $Y=0.895 $X2=0 $Y2=0
cc_595 N_A_652_21#_c_769_n N_SET_B_c_891_n 9.52814e-19 $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_596 N_A_652_21#_c_771_n N_SET_B_c_891_n 0.0205287f $X=4.635 $Y=0.895 $X2=0
+ $Y2=0
cc_597 N_A_652_21#_c_771_n N_SET_B_c_892_n 0.00258368f $X=4.635 $Y=0.895 $X2=0
+ $Y2=0
cc_598 N_A_652_21#_c_769_n N_A_476_47#_c_1018_n 0.00809901f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_599 N_A_652_21#_c_771_n N_A_476_47#_c_1018_n 4.6818e-19 $X=4.635 $Y=0.895
+ $X2=0 $Y2=0
cc_600 N_A_652_21#_c_770_n N_A_476_47#_c_1019_n 0.00249424f $X=4.635 $Y=1.835
+ $X2=0 $Y2=0
cc_601 N_A_652_21#_c_771_n N_A_476_47#_c_1019_n 0.00354719f $X=4.635 $Y=0.895
+ $X2=0 $Y2=0
cc_602 N_A_652_21#_c_775_n N_A_476_47#_M1017_g 0.0138123f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_603 N_A_652_21#_c_770_n N_A_476_47#_M1017_g 0.00542756f $X=4.635 $Y=1.835
+ $X2=0 $Y2=0
cc_604 N_A_652_21#_c_769_n N_A_476_47#_c_1020_n 0.00253676f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_605 N_A_652_21#_c_770_n N_A_476_47#_c_1020_n 2.30787e-19 $X=4.635 $Y=1.835
+ $X2=0 $Y2=0
cc_606 N_A_652_21#_c_771_n N_A_476_47#_c_1020_n 0.0156344f $X=4.635 $Y=0.895
+ $X2=0 $Y2=0
cc_607 N_A_652_21#_c_775_n N_A_476_47#_M1013_g 0.00928157f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_608 N_A_652_21#_c_770_n N_A_476_47#_M1013_g 0.0054278f $X=4.635 $Y=1.835
+ $X2=0 $Y2=0
cc_609 N_A_652_21#_c_769_n N_A_476_47#_c_1021_n 0.0042575f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_610 N_A_652_21#_c_771_n N_A_476_47#_c_1022_n 0.00182092f $X=4.635 $Y=0.895
+ $X2=0 $Y2=0
cc_611 N_A_652_21#_M1004_g N_A_476_47#_c_1045_n 0.00202046f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_612 N_A_652_21#_M1021_g N_A_476_47#_c_1051_n 0.00854236f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_613 N_A_652_21#_M1021_g N_A_476_47#_c_1030_n 0.015293f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_614 N_A_652_21#_c_777_n N_A_476_47#_c_1030_n 0.0366983f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_615 N_A_652_21#_M1021_g N_A_476_47#_c_1023_n 0.018811f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_616 N_A_652_21#_c_774_n N_A_476_47#_c_1024_n 0.00881126f $X=3.99 $Y=1.96
+ $X2=0 $Y2=0
cc_617 N_A_652_21#_c_779_n N_A_476_47#_c_1024_n 0.00337624f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_618 N_A_652_21#_M1021_g N_A_476_47#_c_1025_n 0.0109017f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_619 N_A_652_21#_c_777_n N_A_476_47#_c_1025_n 0.0171213f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_620 N_A_652_21#_c_778_n N_A_476_47#_c_1025_n 0.0011995f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_621 N_A_652_21#_c_775_n N_A_476_47#_c_1026_n 0.0079382f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_622 N_A_652_21#_c_770_n N_A_476_47#_c_1026_n 0.0231083f $X=4.635 $Y=1.835
+ $X2=0 $Y2=0
cc_623 N_A_652_21#_c_779_n N_A_476_47#_c_1026_n 0.00169427f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_624 N_A_652_21#_c_771_n N_A_476_47#_c_1026_n 0.0037745f $X=4.635 $Y=0.895
+ $X2=0 $Y2=0
cc_625 N_A_652_21#_c_775_n N_A_476_47#_c_1027_n 0.0029883f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_626 N_A_652_21#_c_770_n N_A_476_47#_c_1027_n 0.0136869f $X=4.635 $Y=1.835
+ $X2=0 $Y2=0
cc_627 N_A_652_21#_c_771_n N_A_476_47#_c_1027_n 0.00440033f $X=4.635 $Y=0.895
+ $X2=0 $Y2=0
cc_628 N_A_652_21#_c_774_n N_VPWR_M1004_d 0.00131929f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_629 N_A_652_21#_c_777_n N_VPWR_M1004_d 0.00154452f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_630 N_A_652_21#_c_775_n N_VPWR_M1017_d 0.00161389f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_631 N_A_652_21#_c_774_n N_VPWR_c_1479_n 0.00266175f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_632 N_A_652_21#_c_858_p N_VPWR_c_1479_n 0.0070924f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_633 N_A_652_21#_c_775_n N_VPWR_c_1479_n 0.00248431f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_634 N_A_652_21#_c_775_n N_VPWR_c_1480_n 0.0155298f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_635 N_A_652_21#_M1004_g N_VPWR_c_1485_n 0.00532975f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_636 N_A_652_21#_c_777_n N_VPWR_c_1485_n 0.00105935f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_637 N_A_652_21#_c_775_n N_VPWR_c_1486_n 0.00123954f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_638 N_A_652_21#_M1023_d N_VPWR_c_1476_n 0.00202389f $X=3.94 $Y=2.065 $X2=0
+ $Y2=0
cc_639 N_A_652_21#_M1004_g N_VPWR_c_1476_n 0.0066225f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_640 N_A_652_21#_c_774_n N_VPWR_c_1476_n 0.00255051f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_641 N_A_652_21#_c_858_p N_VPWR_c_1476_n 0.00288476f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_642 N_A_652_21#_c_775_n N_VPWR_c_1476_n 0.0036803f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_643 N_A_652_21#_c_777_n N_VPWR_c_1476_n 0.00138626f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_644 N_A_652_21#_M1004_g N_VPWR_c_1493_n 0.00326498f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_645 N_A_652_21#_c_774_n N_VPWR_c_1493_n 0.0101842f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_646 N_A_652_21#_c_777_n N_VPWR_c_1493_n 0.0109284f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_647 N_A_652_21#_c_778_n N_VPWR_c_1493_n 6.81742e-19 $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_648 N_A_652_21#_M1021_g N_VGND_c_1725_n 0.0040279f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_649 N_A_652_21#_c_769_n N_VGND_c_1726_n 0.0118981f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_650 N_A_652_21#_c_771_n N_VGND_c_1726_n 0.00276209f $X=4.635 $Y=0.895 $X2=0
+ $Y2=0
cc_651 N_A_652_21#_c_769_n N_VGND_c_1727_n 0.0177704f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_652 N_A_652_21#_M1021_g N_VGND_c_1731_n 0.0035977f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_653 N_A_652_21#_M1003_d N_VGND_c_1734_n 0.00186029f $X=4.34 $Y=0.235 $X2=0
+ $Y2=0
cc_654 N_A_652_21#_M1021_g N_VGND_c_1734_n 0.00580574f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_655 N_A_652_21#_c_769_n N_VGND_c_1734_n 0.00426169f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_656 N_A_652_21#_c_771_n N_VGND_c_1734_n 0.002078f $X=4.635 $Y=0.895 $X2=0
+ $Y2=0
cc_657 N_SET_B_M1002_g N_A_476_47#_c_1018_n 0.0270653f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_883_n N_A_476_47#_c_1019_n 0.0146844f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_891_n N_A_476_47#_c_1019_n 8.12862e-19 $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_892_n N_A_476_47#_c_1019_n 7.4235e-19 $X=4.08 $Y=0.85 $X2=0
+ $Y2=0
cc_661 N_SET_B_M1023_g N_A_476_47#_M1017_g 0.0336841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_891_n N_A_476_47#_c_1020_n 0.00259966f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_883_n N_A_476_47#_c_1022_n 0.0270653f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_664 SET_B N_A_476_47#_c_1022_n 0.0021684f $X=3.85 $Y=0.765 $X2=0 $Y2=0
cc_665 N_SET_B_c_891_n N_A_476_47#_c_1022_n 0.00277782f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_892_n N_A_476_47#_c_1022_n 7.4235e-19 $X=4.08 $Y=0.85 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_883_n N_A_476_47#_c_1023_n 0.00218199f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_668 N_SET_B_M1023_g N_A_476_47#_c_1023_n 6.04572e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_669 N_SET_B_M1002_g N_A_476_47#_c_1023_n 0.00184201f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_670 SET_B N_A_476_47#_c_1023_n 0.0243796f $X=3.85 $Y=0.765 $X2=0 $Y2=0
cc_671 N_SET_B_c_892_n N_A_476_47#_c_1023_n 0.00110622f $X=4.08 $Y=0.85 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_883_n N_A_476_47#_c_1024_n 0.00307815f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_673 N_SET_B_M1023_g N_A_476_47#_c_1024_n 0.0103672f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_674 SET_B N_A_476_47#_c_1024_n 0.0263655f $X=3.85 $Y=0.765 $X2=0 $Y2=0
cc_675 N_SET_B_c_891_n N_A_476_47#_c_1024_n 2.2446e-19 $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_892_n N_A_476_47#_c_1024_n 6.51468e-19 $X=4.08 $Y=0.85 $X2=0
+ $Y2=0
cc_677 N_SET_B_M1023_g N_A_476_47#_c_1025_n 5.20457e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_678 N_SET_B_M1023_g N_A_476_47#_c_1026_n 0.00354841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_891_n N_A_476_47#_c_1026_n 0.00236582f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_680 N_SET_B_M1023_g N_A_476_47#_c_1027_n 0.0205296f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_681 N_SET_B_M1001_g N_A_1182_261#_M1012_g 0.0588503f $X=6.785 $Y=0.445 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_887_n N_A_1182_261#_M1012_g 0.0108133f $X=6.915 $Y=1.535 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_889_n N_A_1182_261#_M1012_g 0.00109086f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_684 N_SET_B_M1018_g N_A_1182_261#_c_1182_n 0.00284189f $X=6.925 $Y=2.275
+ $X2=0 $Y2=0
cc_685 N_SET_B_c_897_n N_A_1182_261#_c_1182_n 0.00234806f $X=6.915 $Y=1.685
+ $X2=0 $Y2=0
cc_686 N_SET_B_c_887_n N_A_1182_261#_c_1183_n 0.00234806f $X=6.915 $Y=1.535
+ $X2=0 $Y2=0
cc_687 N_SET_B_c_888_n N_A_1182_261#_c_1178_n 2.40668e-19 $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_889_n N_A_1182_261#_c_1178_n 0.00183264f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_959_p N_A_1182_261#_c_1178_n 0.00159132f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_893_n N_A_1182_261#_c_1178_n 0.00928478f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_691 N_SET_B_M1018_g N_A_1182_261#_c_1185_n 0.00936381f $X=6.925 $Y=2.275
+ $X2=0 $Y2=0
cc_692 N_SET_B_c_897_n N_A_1182_261#_c_1185_n 0.00778928f $X=6.915 $Y=1.685
+ $X2=0 $Y2=0
cc_693 N_SET_B_M1001_g N_A_1032_413#_M1007_g 0.0164397f $X=6.785 $Y=0.445 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_888_n N_A_1032_413#_M1007_g 0.00943035f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_889_n N_A_1032_413#_M1007_g 5.48549e-19 $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_959_p N_A_1032_413#_M1007_g 0.00242743f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_893_n N_A_1032_413#_M1007_g 0.00669129f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_887_n N_A_1032_413#_M1010_g 0.00412516f $X=6.915 $Y=1.535 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_897_n N_A_1032_413#_M1010_g 0.0260901f $X=6.915 $Y=1.685 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_891_n N_A_1032_413#_c_1287_n 0.00655755f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_891_n N_A_1032_413#_c_1260_n 0.0101452f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_891_n N_A_1032_413#_c_1261_n 0.00400607f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_703 N_SET_B_M1018_g N_A_1032_413#_c_1272_n 0.00433068f $X=6.925 $Y=2.275
+ $X2=0 $Y2=0
cc_704 N_SET_B_M1001_g N_A_1032_413#_c_1262_n 0.002614f $X=6.785 $Y=0.445 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_887_n N_A_1032_413#_c_1262_n 0.00101786f $X=6.915 $Y=1.535
+ $X2=0 $Y2=0
cc_706 N_SET_B_c_888_n N_A_1032_413#_c_1262_n 0.00156588f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_889_n N_A_1032_413#_c_1262_n 0.0232334f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_891_n N_A_1032_413#_c_1262_n 0.0182014f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_959_p N_A_1032_413#_c_1262_n 3.21596e-19 $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_887_n N_A_1032_413#_c_1263_n 6.30503e-19 $X=6.915 $Y=1.535
+ $X2=0 $Y2=0
cc_711 N_SET_B_c_959_p N_A_1032_413#_c_1263_n 0.00119139f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_893_n N_A_1032_413#_c_1263_n 0.0126036f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_888_n N_A_1032_413#_c_1264_n 0.0220269f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_893_n N_A_1032_413#_c_1264_n 0.00349124f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_887_n N_A_1032_413#_c_1265_n 0.0102848f $X=6.915 $Y=1.535 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_897_n N_A_1032_413#_c_1265_n 5.5231e-19 $X=6.915 $Y=1.685 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_888_n N_A_1032_413#_c_1265_n 0.00347344f $X=6.845 $Y=0.98 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_889_n N_A_1032_413#_c_1265_n 0.0229298f $X=7.01 $Y=0.9 $X2=0
+ $Y2=0
cc_719 N_SET_B_c_891_n N_A_1032_413#_c_1265_n 0.00944298f $X=7.05 $Y=0.85 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_959_p N_A_1032_413#_c_1265_n 7.31634e-19 $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_721 N_SET_B_c_893_n N_A_1032_413#_c_1265_n 0.00833263f $X=7.195 $Y=0.85 $X2=0
+ $Y2=0
cc_722 N_SET_B_M1023_g N_VPWR_c_1479_n 0.00368415f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_723 N_SET_B_M1023_g N_VPWR_c_1480_n 7.26951e-19 $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_724 N_SET_B_M1018_g N_VPWR_c_1481_n 0.00327827f $X=6.925 $Y=2.275 $X2=0 $Y2=0
cc_725 N_SET_B_M1018_g N_VPWR_c_1487_n 0.00585385f $X=6.925 $Y=2.275 $X2=0 $Y2=0
cc_726 N_SET_B_M1023_g N_VPWR_c_1476_n 0.00406312f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_727 N_SET_B_M1018_g N_VPWR_c_1476_n 0.0121898f $X=6.925 $Y=2.275 $X2=0 $Y2=0
cc_728 N_SET_B_M1023_g N_VPWR_c_1493_n 0.00699603f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_729 N_SET_B_M1018_g N_VPWR_c_1495_n 0.00306764f $X=6.925 $Y=2.275 $X2=0 $Y2=0
cc_730 N_SET_B_c_959_p N_VGND_M1001_d 0.00132095f $X=7.195 $Y=0.85 $X2=0 $Y2=0
cc_731 N_SET_B_c_893_n N_VGND_M1001_d 9.16065e-19 $X=7.195 $Y=0.85 $X2=0 $Y2=0
cc_732 N_SET_B_c_883_n N_VGND_c_1725_n 0.00103531f $X=3.865 $Y=1.145 $X2=0 $Y2=0
cc_733 N_SET_B_M1002_g N_VGND_c_1725_n 0.0134999f $X=3.905 $Y=0.445 $X2=0 $Y2=0
cc_734 SET_B N_VGND_c_1725_n 0.0214436f $X=3.85 $Y=0.765 $X2=0 $Y2=0
cc_735 N_SET_B_c_892_n N_VGND_c_1725_n 0.0023818f $X=4.08 $Y=0.85 $X2=0 $Y2=0
cc_736 N_SET_B_c_891_n N_VGND_c_1727_n 0.00554763f $X=7.05 $Y=0.85 $X2=0 $Y2=0
cc_737 N_SET_B_c_889_n N_VGND_c_1734_n 9.40071e-19 $X=7.01 $Y=0.9 $X2=0 $Y2=0
cc_738 SET_B N_VGND_c_1734_n 0.00108472f $X=3.85 $Y=0.765 $X2=0 $Y2=0
cc_739 N_SET_B_c_891_n N_VGND_c_1734_n 0.136444f $X=7.05 $Y=0.85 $X2=0 $Y2=0
cc_740 N_SET_B_c_892_n N_VGND_c_1734_n 0.0148244f $X=4.08 $Y=0.85 $X2=0 $Y2=0
cc_741 N_SET_B_c_959_p N_VGND_c_1734_n 0.0145428f $X=7.195 $Y=0.85 $X2=0 $Y2=0
cc_742 N_SET_B_c_893_n N_VGND_c_1734_n 2.23886e-19 $X=7.195 $Y=0.85 $X2=0 $Y2=0
cc_743 N_SET_B_M1001_g N_VGND_c_1740_n 0.02016f $X=6.785 $Y=0.445 $X2=0 $Y2=0
cc_744 N_SET_B_c_888_n N_VGND_c_1740_n 6.12458e-19 $X=6.845 $Y=0.98 $X2=0 $Y2=0
cc_745 N_SET_B_c_889_n N_VGND_c_1740_n 0.0407925f $X=7.01 $Y=0.9 $X2=0 $Y2=0
cc_746 N_SET_B_c_891_n N_VGND_c_1740_n 0.00168626f $X=7.05 $Y=0.85 $X2=0 $Y2=0
cc_747 N_SET_B_c_959_p N_VGND_c_1740_n 0.00338224f $X=7.195 $Y=0.85 $X2=0 $Y2=0
cc_748 N_A_476_47#_M1013_g N_A_1032_413#_c_1278_n 8.92621e-19 $X=4.705 $Y=2.275
+ $X2=0 $Y2=0
cc_749 N_A_476_47#_M1017_g N_VPWR_c_1479_n 0.00339367f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_750 N_A_476_47#_M1017_g N_VPWR_c_1480_n 0.00730335f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_751 N_A_476_47#_M1013_g N_VPWR_c_1480_n 0.00918253f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_752 N_A_476_47#_c_1045_n N_VPWR_c_1485_n 0.0377433f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_753 N_A_476_47#_M1013_g N_VPWR_c_1486_n 0.00392729f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_754 N_A_476_47#_M1006_d N_VPWR_c_1476_n 0.00173085f $X=2.39 $Y=2.065 $X2=0
+ $Y2=0
cc_755 N_A_476_47#_M1017_g N_VPWR_c_1476_n 0.00379591f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_756 N_A_476_47#_M1013_g N_VPWR_c_1476_n 0.00396629f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_757 N_A_476_47#_c_1045_n N_VPWR_c_1476_n 0.0132511f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_758 N_A_476_47#_M1017_g N_VPWR_c_1493_n 7.14614e-19 $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_759 N_A_476_47#_c_1045_n N_A_381_47#_c_1651_n 0.0102747f $X=3.02 $Y=2.335
+ $X2=0 $Y2=0
cc_760 N_A_476_47#_c_1045_n A_562_413# 0.00859792f $X=3.02 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_761 N_A_476_47#_c_1030_n A_562_413# 0.00578953f $X=3.105 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_762 N_A_476_47#_c_1018_n N_VGND_c_1725_n 0.00301834f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_763 N_A_476_47#_c_1018_n N_VGND_c_1726_n 0.00541969f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_764 N_A_476_47#_c_1020_n N_VGND_c_1726_n 0.0011731f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_765 N_A_476_47#_c_1018_n N_VGND_c_1727_n 0.00362321f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_766 N_A_476_47#_c_1020_n N_VGND_c_1727_n 0.00665809f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_767 N_A_476_47#_c_1021_n N_VGND_c_1727_n 0.00456783f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_768 N_A_476_47#_c_1051_n N_VGND_c_1731_n 0.055608f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_769 N_A_476_47#_M1024_d N_VGND_c_1734_n 0.00275359f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_770 N_A_476_47#_c_1018_n N_VGND_c_1734_n 0.00742824f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_771 N_A_476_47#_c_1020_n N_VGND_c_1734_n 3.98471e-19 $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_772 N_A_476_47#_c_1021_n N_VGND_c_1734_n 0.00674913f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_773 N_A_476_47#_c_1051_n N_VGND_c_1734_n 0.0218827f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_774 N_A_476_47#_c_1021_n N_VGND_c_1739_n 0.00437852f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_775 N_A_476_47#_c_1051_n A_586_47# 0.00568226f $X=3.27 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_776 N_A_1182_261#_c_1178_n N_A_1032_413#_M1007_g 0.00942388f $X=7.755
+ $Y=1.575 $X2=0 $Y2=0
cc_777 N_A_1182_261#_c_1178_n N_A_1032_413#_M1010_g 0.00513051f $X=7.755
+ $Y=1.575 $X2=0 $Y2=0
cc_778 N_A_1182_261#_c_1185_n N_A_1032_413#_M1010_g 0.0144865f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_779 N_A_1182_261#_c_1178_n N_A_1032_413#_c_1257_n 0.0232556f $X=7.755
+ $Y=1.575 $X2=0 $Y2=0
cc_780 N_A_1182_261#_c_1179_n N_A_1032_413#_c_1257_n 0.0033418f $X=7.755
+ $Y=0.515 $X2=0 $Y2=0
cc_781 N_A_1182_261#_c_1186_n N_A_1032_413#_c_1257_n 0.00452123f $X=7.755
+ $Y=1.67 $X2=0 $Y2=0
cc_782 N_A_1182_261#_c_1178_n N_A_1032_413#_M1030_g 0.00180277f $X=7.755
+ $Y=1.575 $X2=0 $Y2=0
cc_783 N_A_1182_261#_c_1179_n N_A_1032_413#_M1030_g 6.69263e-19 $X=7.755
+ $Y=0.515 $X2=0 $Y2=0
cc_784 N_A_1182_261#_c_1214_p N_A_1032_413#_M1029_g 0.00122441f $X=7.615 $Y=1.87
+ $X2=0 $Y2=0
cc_785 N_A_1182_261#_c_1178_n N_A_1032_413#_M1029_g 6.46443e-19 $X=7.755
+ $Y=1.575 $X2=0 $Y2=0
cc_786 N_A_1182_261#_c_1186_n N_A_1032_413#_M1029_g 9.16556e-19 $X=7.755 $Y=1.67
+ $X2=0 $Y2=0
cc_787 N_A_1182_261#_c_1177_n N_A_1032_413#_c_1270_n 0.00400855f $X=6.405
+ $Y=1.38 $X2=0 $Y2=0
cc_788 N_A_1182_261#_c_1185_n N_A_1032_413#_c_1270_n 0.0133834f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_789 N_A_1182_261#_M1012_g N_A_1032_413#_c_1287_n 0.00585858f $X=6.405
+ $Y=0.445 $X2=0 $Y2=0
cc_790 N_A_1182_261#_c_1177_n N_A_1032_413#_c_1260_n 0.0136825f $X=6.405 $Y=1.38
+ $X2=0 $Y2=0
cc_791 N_A_1182_261#_c_1185_n N_A_1032_413#_c_1260_n 0.026737f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_792 N_A_1182_261#_M1027_g N_A_1032_413#_c_1272_n 0.0119267f $X=5.985 $Y=2.275
+ $X2=0 $Y2=0
cc_793 N_A_1182_261#_c_1182_n N_A_1032_413#_c_1272_n 0.00460004f $X=6.07
+ $Y=1.825 $X2=0 $Y2=0
cc_794 N_A_1182_261#_c_1185_n N_A_1032_413#_c_1272_n 0.0654175f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_795 N_A_1182_261#_M1012_g N_A_1032_413#_c_1262_n 0.014625f $X=6.405 $Y=0.445
+ $X2=0 $Y2=0
cc_796 N_A_1182_261#_M1027_g N_A_1032_413#_c_1273_n 0.00296198f $X=5.985
+ $Y=2.275 $X2=0 $Y2=0
cc_797 N_A_1182_261#_M1027_g N_A_1032_413#_c_1274_n 0.00444241f $X=5.985
+ $Y=2.275 $X2=0 $Y2=0
cc_798 N_A_1182_261#_c_1182_n N_A_1032_413#_c_1274_n 0.00400855f $X=6.07
+ $Y=1.825 $X2=0 $Y2=0
cc_799 N_A_1182_261#_M1012_g N_A_1032_413#_c_1362_n 0.00335259f $X=6.405
+ $Y=0.445 $X2=0 $Y2=0
cc_800 N_A_1182_261#_c_1177_n N_A_1032_413#_c_1362_n 0.00418281f $X=6.405
+ $Y=1.38 $X2=0 $Y2=0
cc_801 N_A_1182_261#_c_1185_n N_A_1032_413#_c_1362_n 0.0136304f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_802 N_A_1182_261#_c_1178_n N_A_1032_413#_c_1263_n 0.0172431f $X=7.755
+ $Y=1.575 $X2=0 $Y2=0
cc_803 N_A_1182_261#_c_1185_n N_A_1032_413#_c_1264_n 0.0032134f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_804 N_A_1182_261#_c_1185_n N_A_1032_413#_c_1265_n 0.0723173f $X=7.53 $Y=1.67
+ $X2=0 $Y2=0
cc_805 N_A_1182_261#_c_1178_n N_A_1602_47#_c_1420_n 0.0219446f $X=7.755 $Y=1.575
+ $X2=0 $Y2=0
cc_806 N_A_1182_261#_c_1179_n N_A_1602_47#_c_1420_n 0.0234463f $X=7.755 $Y=0.515
+ $X2=0 $Y2=0
cc_807 N_A_1182_261#_c_1214_p N_A_1602_47#_c_1428_n 0.0257383f $X=7.615 $Y=1.87
+ $X2=0 $Y2=0
cc_808 N_A_1182_261#_c_1214_p N_A_1602_47#_c_1429_n 0.00670342f $X=7.615 $Y=1.87
+ $X2=0 $Y2=0
cc_809 N_A_1182_261#_c_1178_n N_A_1602_47#_c_1429_n 0.0166195f $X=7.755 $Y=1.575
+ $X2=0 $Y2=0
cc_810 N_A_1182_261#_c_1186_n N_A_1602_47#_c_1429_n 0.014454f $X=7.755 $Y=1.67
+ $X2=0 $Y2=0
cc_811 N_A_1182_261#_c_1178_n N_A_1602_47#_c_1423_n 0.0230781f $X=7.755 $Y=1.575
+ $X2=0 $Y2=0
cc_812 N_A_1182_261#_c_1185_n N_VPWR_M1018_d 0.00225674f $X=7.53 $Y=1.67 $X2=0
+ $Y2=0
cc_813 N_A_1182_261#_c_1185_n N_VPWR_c_1481_n 0.0195228f $X=7.53 $Y=1.67 $X2=0
+ $Y2=0
cc_814 N_A_1182_261#_M1027_g N_VPWR_c_1486_n 8.50188e-19 $X=5.985 $Y=2.275 $X2=0
+ $Y2=0
cc_815 N_A_1182_261#_c_1214_p N_VPWR_c_1488_n 0.00727431f $X=7.615 $Y=1.87 $X2=0
+ $Y2=0
cc_816 N_A_1182_261#_M1010_d N_VPWR_c_1476_n 0.00535012f $X=7.48 $Y=1.645 $X2=0
+ $Y2=0
cc_817 N_A_1182_261#_M1027_g N_VPWR_c_1476_n 0.00145798f $X=5.985 $Y=2.275 $X2=0
+ $Y2=0
cc_818 N_A_1182_261#_c_1214_p N_VPWR_c_1476_n 0.00614354f $X=7.615 $Y=1.87 $X2=0
+ $Y2=0
cc_819 N_A_1182_261#_M1027_g N_VPWR_c_1495_n 0.0145664f $X=5.985 $Y=2.275 $X2=0
+ $Y2=0
cc_820 N_A_1182_261#_c_1179_n N_VGND_c_1732_n 0.0131701f $X=7.755 $Y=0.515 $X2=0
+ $Y2=0
cc_821 N_A_1182_261#_M1007_d N_VGND_c_1734_n 0.00391384f $X=7.48 $Y=0.235 $X2=0
+ $Y2=0
cc_822 N_A_1182_261#_M1012_g N_VGND_c_1734_n 0.00501331f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_823 N_A_1182_261#_c_1179_n N_VGND_c_1734_n 0.0114301f $X=7.755 $Y=0.515 $X2=0
+ $Y2=0
cc_824 N_A_1182_261#_M1012_g N_VGND_c_1739_n 0.00367922f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_825 N_A_1182_261#_M1012_g N_VGND_c_1740_n 0.00242905f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_826 N_A_1032_413#_c_1259_n N_A_1602_47#_M1025_g 0.0230602f $X=8.345 $Y=1.26
+ $X2=0 $Y2=0
cc_827 N_A_1032_413#_M1030_g N_A_1602_47#_c_1420_n 0.0175367f $X=8.345 $Y=0.445
+ $X2=0 $Y2=0
cc_828 N_A_1032_413#_M1030_g N_A_1602_47#_c_1421_n 0.0076587f $X=8.345 $Y=0.445
+ $X2=0 $Y2=0
cc_829 N_A_1032_413#_c_1259_n N_A_1602_47#_c_1421_n 0.0103507f $X=8.345 $Y=1.26
+ $X2=0 $Y2=0
cc_830 N_A_1032_413#_M1030_g N_A_1602_47#_c_1422_n 0.0214041f $X=8.345 $Y=0.445
+ $X2=0 $Y2=0
cc_831 N_A_1032_413#_M1010_g N_A_1602_47#_c_1428_n 0.00145954f $X=7.405 $Y=2.065
+ $X2=0 $Y2=0
cc_832 N_A_1032_413#_c_1257_n N_A_1602_47#_c_1428_n 0.00240579f $X=8.27 $Y=1.26
+ $X2=0 $Y2=0
cc_833 N_A_1032_413#_M1029_g N_A_1602_47#_c_1428_n 0.0057641f $X=8.345 $Y=2.165
+ $X2=0 $Y2=0
cc_834 N_A_1032_413#_M1010_g N_A_1602_47#_c_1429_n 6.55852e-19 $X=7.405 $Y=2.065
+ $X2=0 $Y2=0
cc_835 N_A_1032_413#_c_1257_n N_A_1602_47#_c_1429_n 0.00670725f $X=8.27 $Y=1.26
+ $X2=0 $Y2=0
cc_836 N_A_1032_413#_M1029_g N_A_1602_47#_c_1429_n 0.0165499f $X=8.345 $Y=2.165
+ $X2=0 $Y2=0
cc_837 N_A_1032_413#_c_1259_n N_A_1602_47#_c_1429_n 0.00186719f $X=8.345 $Y=1.26
+ $X2=0 $Y2=0
cc_838 N_A_1032_413#_c_1257_n N_A_1602_47#_c_1423_n 0.0115739f $X=8.27 $Y=1.26
+ $X2=0 $Y2=0
cc_839 N_A_1032_413#_M1030_g N_A_1602_47#_c_1423_n 0.00213726f $X=8.345 $Y=0.445
+ $X2=0 $Y2=0
cc_840 N_A_1032_413#_c_1259_n N_A_1602_47#_c_1423_n 6.49734e-19 $X=8.345 $Y=1.26
+ $X2=0 $Y2=0
cc_841 N_A_1032_413#_M1030_g N_A_1602_47#_c_1424_n 0.0197757f $X=8.345 $Y=0.445
+ $X2=0 $Y2=0
cc_842 N_A_1032_413#_c_1272_n N_VPWR_M1027_d 0.00216018f $X=6.56 $Y=2 $X2=0
+ $Y2=0
cc_843 N_A_1032_413#_c_1278_n N_VPWR_c_1480_n 0.00537013f $X=5.59 $Y=2.29 $X2=0
+ $Y2=0
cc_844 N_A_1032_413#_M1010_g N_VPWR_c_1481_n 0.0153912f $X=7.405 $Y=2.065 $X2=0
+ $Y2=0
cc_845 N_A_1032_413#_c_1272_n N_VPWR_c_1481_n 0.00850121f $X=6.56 $Y=2 $X2=0
+ $Y2=0
cc_846 N_A_1032_413#_M1029_g N_VPWR_c_1482_n 0.00609621f $X=8.345 $Y=2.165 $X2=0
+ $Y2=0
cc_847 N_A_1032_413#_c_1278_n N_VPWR_c_1486_n 0.0200526f $X=5.59 $Y=2.29 $X2=0
+ $Y2=0
cc_848 N_A_1032_413#_c_1272_n N_VPWR_c_1486_n 0.00267646f $X=6.56 $Y=2 $X2=0
+ $Y2=0
cc_849 N_A_1032_413#_c_1274_n N_VPWR_c_1486_n 0.00720374f $X=5.675 $Y=2 $X2=0
+ $Y2=0
cc_850 N_A_1032_413#_c_1272_n N_VPWR_c_1487_n 0.0036467f $X=6.56 $Y=2 $X2=0
+ $Y2=0
cc_851 N_A_1032_413#_c_1273_n N_VPWR_c_1487_n 0.0101929f $X=6.715 $Y=2.21 $X2=0
+ $Y2=0
cc_852 N_A_1032_413#_M1010_g N_VPWR_c_1488_n 0.0046653f $X=7.405 $Y=2.065 $X2=0
+ $Y2=0
cc_853 N_A_1032_413#_M1029_g N_VPWR_c_1488_n 0.00542953f $X=8.345 $Y=2.165 $X2=0
+ $Y2=0
cc_854 N_A_1032_413#_M1026_d N_VPWR_c_1476_n 0.00263666f $X=5.16 $Y=2.065 $X2=0
+ $Y2=0
cc_855 N_A_1032_413#_M1018_s N_VPWR_c_1476_n 0.00394021f $X=6.59 $Y=2.065 $X2=0
+ $Y2=0
cc_856 N_A_1032_413#_M1010_g N_VPWR_c_1476_n 0.00934473f $X=7.405 $Y=2.065 $X2=0
+ $Y2=0
cc_857 N_A_1032_413#_M1029_g N_VPWR_c_1476_n 0.0110121f $X=8.345 $Y=2.165 $X2=0
+ $Y2=0
cc_858 N_A_1032_413#_c_1278_n N_VPWR_c_1476_n 0.00937878f $X=5.59 $Y=2.29 $X2=0
+ $Y2=0
cc_859 N_A_1032_413#_c_1272_n N_VPWR_c_1476_n 0.0124969f $X=6.56 $Y=2 $X2=0
+ $Y2=0
cc_860 N_A_1032_413#_c_1273_n N_VPWR_c_1476_n 0.0086238f $X=6.715 $Y=2.21 $X2=0
+ $Y2=0
cc_861 N_A_1032_413#_c_1274_n N_VPWR_c_1476_n 0.00578252f $X=5.675 $Y=2 $X2=0
+ $Y2=0
cc_862 N_A_1032_413#_c_1272_n N_VPWR_c_1495_n 0.0270337f $X=6.56 $Y=2 $X2=0
+ $Y2=0
cc_863 N_A_1032_413#_c_1273_n N_VPWR_c_1495_n 0.00887045f $X=6.715 $Y=2.21 $X2=0
+ $Y2=0
cc_864 N_A_1032_413#_c_1274_n N_VPWR_c_1495_n 0.0115187f $X=5.675 $Y=2 $X2=0
+ $Y2=0
cc_865 N_A_1032_413#_c_1272_n A_1140_413# 0.00166681f $X=6.56 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_866 N_A_1032_413#_c_1274_n A_1140_413# 0.00336335f $X=5.675 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_867 N_A_1032_413#_M1030_g N_VGND_c_1728_n 0.00587725f $X=8.345 $Y=0.445 $X2=0
+ $Y2=0
cc_868 N_A_1032_413#_M1007_g N_VGND_c_1732_n 0.00505556f $X=7.405 $Y=0.505 $X2=0
+ $Y2=0
cc_869 N_A_1032_413#_M1030_g N_VGND_c_1732_n 0.00544863f $X=8.345 $Y=0.445 $X2=0
+ $Y2=0
cc_870 N_A_1032_413#_M1009_d N_VGND_c_1734_n 0.00218745f $X=5.64 $Y=0.235 $X2=0
+ $Y2=0
cc_871 N_A_1032_413#_M1007_g N_VGND_c_1734_n 0.00991048f $X=7.405 $Y=0.505 $X2=0
+ $Y2=0
cc_872 N_A_1032_413#_M1030_g N_VGND_c_1734_n 0.0111099f $X=8.345 $Y=0.445 $X2=0
+ $Y2=0
cc_873 N_A_1032_413#_c_1287_n N_VGND_c_1734_n 0.0135115f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_874 N_A_1032_413#_c_1287_n N_VGND_c_1739_n 0.0361566f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_875 N_A_1032_413#_M1007_g N_VGND_c_1740_n 0.0188937f $X=7.405 $Y=0.505 $X2=0
+ $Y2=0
cc_876 N_A_1032_413#_c_1263_n N_VGND_c_1740_n 2.67651e-19 $X=7.325 $Y=1.26 $X2=0
+ $Y2=0
cc_877 N_A_1032_413#_c_1287_n A_1224_47# 0.00244121f $X=6.32 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_878 N_A_1602_47#_c_1428_n N_VPWR_c_1481_n 0.00150514f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_879 N_A_1602_47#_M1025_g N_VPWR_c_1482_n 0.0168002f $X=8.82 $Y=1.985 $X2=0
+ $Y2=0
cc_880 N_A_1602_47#_c_1421_n N_VPWR_c_1482_n 0.00939656f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_881 N_A_1602_47#_c_1422_n N_VPWR_c_1482_n 0.00188681f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_882 N_A_1602_47#_c_1429_n N_VPWR_c_1482_n 0.0431561f $X=8.135 $Y=1.915 $X2=0
+ $Y2=0
cc_883 N_A_1602_47#_c_1428_n N_VPWR_c_1488_n 0.0166647f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_884 N_A_1602_47#_M1025_g N_VPWR_c_1489_n 0.00505556f $X=8.82 $Y=1.985 $X2=0
+ $Y2=0
cc_885 N_A_1602_47#_M1029_s N_VPWR_c_1476_n 0.00211564f $X=8.01 $Y=1.845 $X2=0
+ $Y2=0
cc_886 N_A_1602_47#_M1025_g N_VPWR_c_1476_n 0.00995901f $X=8.82 $Y=1.985 $X2=0
+ $Y2=0
cc_887 N_A_1602_47#_c_1428_n N_VPWR_c_1476_n 0.0121504f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_888 N_A_1602_47#_M1025_g N_Q_c_1708_n 0.0113745f $X=8.82 $Y=1.985 $X2=0 $Y2=0
cc_889 N_A_1602_47#_c_1421_n N_Q_c_1708_n 0.026319f $X=8.765 $Y=1.16 $X2=0 $Y2=0
cc_890 N_A_1602_47#_c_1422_n N_Q_c_1708_n 0.00757092f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_891 N_A_1602_47#_c_1424_n N_Q_c_1708_n 0.00666969f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_892 N_A_1602_47#_c_1420_n N_VGND_c_1728_n 0.0143899f $X=8.135 $Y=0.51 $X2=0
+ $Y2=0
cc_893 N_A_1602_47#_c_1421_n N_VGND_c_1728_n 0.0102661f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_894 N_A_1602_47#_c_1422_n N_VGND_c_1728_n 0.00198004f $X=8.765 $Y=1.16 $X2=0
+ $Y2=0
cc_895 N_A_1602_47#_c_1424_n N_VGND_c_1728_n 0.00905698f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_896 N_A_1602_47#_c_1420_n N_VGND_c_1732_n 0.00973496f $X=8.135 $Y=0.51 $X2=0
+ $Y2=0
cc_897 N_A_1602_47#_c_1424_n N_VGND_c_1733_n 0.00505556f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_898 N_A_1602_47#_M1030_s N_VGND_c_1734_n 0.00359633f $X=8.01 $Y=0.235 $X2=0
+ $Y2=0
cc_899 N_A_1602_47#_c_1420_n N_VGND_c_1734_n 0.00895081f $X=8.135 $Y=0.51 $X2=0
+ $Y2=0
cc_900 N_A_1602_47#_c_1424_n N_VGND_c_1734_n 0.00995901f $X=8.765 $Y=0.995 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1476_n N_A_381_47#_M1022_d 0.00325229f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_902 N_VPWR_M1022_s N_A_381_47#_c_1641_n 0.00237137f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_903 N_VPWR_M1022_s N_A_381_47#_c_1648_n 0.00471078f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1478_n N_A_381_47#_c_1648_n 0.00880041f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1485_n N_A_381_47#_c_1648_n 0.0018545f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1476_n N_A_381_47#_c_1648_n 0.00198108f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_907 N_VPWR_M1022_s N_A_381_47#_c_1644_n 0.00187968f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_908 N_VPWR_c_1478_n N_A_381_47#_c_1644_n 0.0114817f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_909 N_VPWR_c_1484_n N_A_381_47#_c_1644_n 3.86777e-19 $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_910 N_VPWR_c_1476_n N_A_381_47#_c_1644_n 7.1462e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1485_n N_A_381_47#_c_1651_n 0.0115924f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_912 N_VPWR_c_1476_n N_A_381_47#_c_1651_n 0.00307944f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1476_n A_562_413# 0.00355877f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_914 N_VPWR_c_1476_n A_956_413# 0.00279018f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_915 N_VPWR_c_1476_n A_1140_413# 0.00223276f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_916 N_VPWR_c_1476_n N_Q_M1025_d 0.00401809f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_917 N_VPWR_c_1489_n Q 0.00922946f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_918 N_VPWR_c_1476_n Q 0.00900208f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_919 N_A_381_47#_c_1641_n N_VGND_M1005_s 0.00105184f $X=1.515 $Y=1.795 $X2=0
+ $Y2=0
cc_920 N_A_381_47#_c_1646_n N_VGND_M1005_s 0.00264874f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_921 N_A_381_47#_c_1642_n N_VGND_M1005_s 0.0019591f $X=1.6 $Y=0.73 $X2=0 $Y2=0
cc_922 N_A_381_47#_c_1646_n N_VGND_c_1724_n 0.00883988f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_923 N_A_381_47#_c_1642_n N_VGND_c_1724_n 0.0114461f $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_924 N_A_381_47#_c_1642_n N_VGND_c_1730_n 4.97798e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_925 N_A_381_47#_c_1646_n N_VGND_c_1731_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_926 N_A_381_47#_c_1650_n N_VGND_c_1731_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_927 N_A_381_47#_M1005_d N_VGND_c_1734_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_928 N_A_381_47#_c_1646_n N_VGND_c_1734_n 0.00232804f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_929 N_A_381_47#_c_1642_n N_VGND_c_1734_n 8.52239e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_930 N_A_381_47#_c_1650_n N_VGND_c_1734_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_931 Q N_VGND_c_1733_n 0.016502f $X=8.97 $Y=0.425 $X2=0 $Y2=0
cc_932 N_Q_M1020_d N_VGND_c_1734_n 0.00387432f $X=8.895 $Y=0.235 $X2=0 $Y2=0
cc_933 Q N_VGND_c_1734_n 0.00967853f $X=8.97 $Y=0.425 $X2=0 $Y2=0
cc_934 N_VGND_c_1734_n A_586_47# 0.0022723f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_935 N_VGND_c_1734_n A_796_47# 0.0023931f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_936 N_VGND_c_1734_n A_1056_47# 0.00198596f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_937 N_VGND_c_1734_n A_1224_47# 0.00140476f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_938 N_VGND_c_1734_n A_1296_47# 0.0028857f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__xnor2_2.spice.SKY130_FD_SC_HD__XNOR2_2.pxi
* Created: Thu Aug 27 14:49:04 2020
* 
x_PM_SKY130_FD_SC_HD__XNOR2_2%B N_B_c_96_n N_B_M1008_g N_B_M1003_g N_B_c_97_n
+ N_B_M1015_g N_B_M1018_g N_B_c_98_n N_B_M1010_g N_B_M1012_g N_B_c_99_n
+ N_B_M1016_g N_B_M1017_g N_B_c_129_p N_B_c_107_n N_B_c_108_n N_B_c_125_p
+ N_B_c_100_n N_B_c_109_n N_B_c_110_n B N_B_c_101_n N_B_c_102_n
+ PM_SKY130_FD_SC_HD__XNOR2_2%B
x_PM_SKY130_FD_SC_HD__XNOR2_2%A N_A_c_215_n N_A_M1007_g N_A_M1009_g N_A_c_216_n
+ N_A_M1013_g N_A_M1011_g N_A_c_217_n N_A_M1014_g N_A_M1002_g N_A_c_218_n
+ N_A_M1019_g N_A_M1005_g N_A_c_219_n N_A_c_220_n A N_A_c_221_n N_A_c_249_n
+ PM_SKY130_FD_SC_HD__XNOR2_2%A
x_PM_SKY130_FD_SC_HD__XNOR2_2%A_27_297# N_A_27_297#_M1008_s N_A_27_297#_M1003_s
+ N_A_27_297#_M1018_s N_A_27_297#_M1011_d N_A_27_297#_c_310_n
+ N_A_27_297#_M1000_g N_A_27_297#_M1001_g N_A_27_297#_c_311_n
+ N_A_27_297#_M1004_g N_A_27_297#_M1006_g N_A_27_297#_c_312_n
+ N_A_27_297#_c_313_n N_A_27_297#_c_314_n N_A_27_297#_c_338_n
+ N_A_27_297#_c_344_n N_A_27_297#_c_322_n N_A_27_297#_c_363_n
+ N_A_27_297#_c_323_n N_A_27_297#_c_324_n N_A_27_297#_c_315_n
+ N_A_27_297#_c_316_n N_A_27_297#_c_317_n N_A_27_297#_c_326_n
+ N_A_27_297#_c_356_n N_A_27_297#_c_357_n N_A_27_297#_c_318_n
+ PM_SKY130_FD_SC_HD__XNOR2_2%A_27_297#
x_PM_SKY130_FD_SC_HD__XNOR2_2%VPWR N_VPWR_M1003_d N_VPWR_M1009_s N_VPWR_M1002_s
+ N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n
+ N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n
+ VPWR N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_459_n
+ N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_447_n
+ PM_SKY130_FD_SC_HD__XNOR2_2%VPWR
x_PM_SKY130_FD_SC_HD__XNOR2_2%A_474_297# N_A_474_297#_M1002_d
+ N_A_474_297#_M1005_d N_A_474_297#_M1017_s N_A_474_297#_c_554_n
+ N_A_474_297#_c_584_n N_A_474_297#_c_560_n N_A_474_297#_c_562_n
+ N_A_474_297#_c_573_n N_A_474_297#_c_556_n N_A_474_297#_c_558_n
+ PM_SKY130_FD_SC_HD__XNOR2_2%A_474_297#
x_PM_SKY130_FD_SC_HD__XNOR2_2%Y N_Y_M1000_d N_Y_M1004_d N_Y_M1012_d N_Y_M1001_s
+ N_Y_c_612_n N_Y_c_609_n N_Y_c_638_n N_Y_c_610_n N_Y_c_611_n N_Y_c_624_n Y
+ PM_SKY130_FD_SC_HD__XNOR2_2%Y
x_PM_SKY130_FD_SC_HD__XNOR2_2%A_27_47# N_A_27_47#_M1008_d N_A_27_47#_M1015_d
+ N_A_27_47#_M1013_s N_A_27_47#_c_661_n N_A_27_47#_c_670_n N_A_27_47#_c_662_n
+ N_A_27_47#_c_663_n N_A_27_47#_c_664_n PM_SKY130_FD_SC_HD__XNOR2_2%A_27_47#
x_PM_SKY130_FD_SC_HD__XNOR2_2%VGND N_VGND_M1007_d N_VGND_M1014_s N_VGND_M1019_s
+ N_VGND_M1016_d N_VGND_c_703_n N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n
+ N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n
+ N_VGND_c_712_n N_VGND_c_713_n N_VGND_c_714_n VGND N_VGND_c_715_n
+ N_VGND_c_716_n PM_SKY130_FD_SC_HD__XNOR2_2%VGND
x_PM_SKY130_FD_SC_HD__XNOR2_2%A_560_47# N_A_560_47#_M1014_d N_A_560_47#_M1010_s
+ N_A_560_47#_M1000_s N_A_560_47#_c_796_n N_A_560_47#_c_791_n
+ N_A_560_47#_c_792_n N_A_560_47#_c_801_n N_A_560_47#_c_793_n
+ N_A_560_47#_c_794_n N_A_560_47#_c_795_n PM_SKY130_FD_SC_HD__XNOR2_2%A_560_47#
cc_1 VNB N_B_c_96_n 0.0191418f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_B_c_97_n 0.0161688f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_B_c_98_n 0.0163545f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.995
cc_4 VNB N_B_c_99_n 0.0218312f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.995
cc_5 VNB N_B_c_100_n 0.00545644f $X=-0.19 $Y=-0.24 $X2=3.755 $Y2=1.16
cc_6 VNB N_B_c_101_n 0.0345208f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_7 VNB N_B_c_102_n 0.0395067f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=1.16
cc_8 VNB N_A_c_215_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_9 VNB N_A_c_216_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_10 VNB N_A_c_217_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.995
cc_11 VNB N_A_c_218_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.995
cc_12 VNB N_A_c_219_n 0.0510052f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.18
cc_13 VNB N_A_c_220_n 0.0255324f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_14 VNB N_A_c_221_n 0.0269042f $X=-0.19 $Y=-0.24 $X2=0.875 $Y2=1.445
cc_15 VNB N_A_27_297#_c_310_n 0.0214899f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_16 VNB N_A_27_297#_c_311_n 0.0190697f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=1.985
cc_17 VNB N_A_27_297#_c_312_n 0.0205105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_313_n 0.0112022f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_19 VNB N_A_27_297#_c_314_n 0.00562166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_315_n 0.0014749f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_21 VNB N_A_27_297#_c_316_n 0.00418379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_297#_c_317_n 0.00192645f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_297#_c_318_n 0.039041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_447_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_609_n 0.00241737f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.995
cc_26 VNB N_Y_c_610_n 0.0094867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_611_n 0.0433703f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.56
cc_28 VNB N_A_27_47#_c_661_n 0.00961138f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_29 VNB N_A_27_47#_c_662_n 0.00358652f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.995
cc_30 VNB N_A_27_47#_c_663_n 0.00609203f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.56
cc_31 VNB N_A_27_47#_c_664_n 0.00472644f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=1.985
cc_32 VNB N_VGND_c_703_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.995
cc_33 VNB N_VGND_c_704_n 0.00566097f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=1.985
cc_34 VNB N_VGND_c_705_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.56
cc_35 VNB N_VGND_c_706_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=1.985
cc_36 VNB N_VGND_c_707_n 0.036159f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.18
cc_37 VNB N_VGND_c_708_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_38 VNB N_VGND_c_709_n 0.0218603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_710_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0.875 $Y2=1.285
cc_40 VNB N_VGND_c_711_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=3.015 $Y2=1.285
cc_41 VNB N_VGND_c_712_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=3.015 $Y2=1.445
cc_42 VNB N_VGND_c_713_n 0.0174412f $X=-0.19 $Y=-0.24 $X2=3.755 $Y2=1.18
cc_43 VNB N_VGND_c_714_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=3.755 $Y2=1.16
cc_44 VNB N_VGND_c_715_n 0.042967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_716_n 0.309767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_560_47#_c_791_n 0.00248283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_560_47#_c_792_n 0.00289865f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.995
cc_48 VNB N_A_560_47#_c_793_n 0.00243379f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.995
cc_49 VNB N_A_560_47#_c_794_n 0.00224987f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=0.56
cc_50 VNB N_A_560_47#_c_795_n 0.0160859f $X=-0.19 $Y=-0.24 $X2=4.02 $Y2=1.325
cc_51 VPB N_B_M1003_g 0.0218915f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_52 VPB N_B_M1018_g 0.0178886f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_53 VPB N_B_M1012_g 0.0189073f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=1.985
cc_54 VPB N_B_M1017_g 0.0233065f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=1.985
cc_55 VPB N_B_c_107_n 0.0010643f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.445
cc_56 VPB N_B_c_108_n 0.00111437f $X=-0.19 $Y=1.305 $X2=3.015 $Y2=1.445
cc_57 VPB N_B_c_109_n 3.58755e-19 $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.53
cc_58 VPB N_B_c_110_n 0.0187016f $X=-0.19 $Y=1.305 $X2=2.93 $Y2=1.53
cc_59 VPB N_B_c_101_n 0.00477025f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_60 VPB N_B_c_102_n 0.00530143f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=1.16
cc_61 VPB N_A_M1009_g 0.0183682f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_62 VPB N_A_M1011_g 0.025044f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_63 VPB N_A_M1002_g 0.0249968f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=1.985
cc_64 VPB N_A_M1005_g 0.0181328f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=1.985
cc_65 VPB N_A_c_219_n 0.0170727f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.18
cc_66 VPB N_A_c_220_n 0.00394613f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_67 VPB N_A_c_221_n 0.00372033f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.445
cc_68 VPB N_A_27_297#_M1001_g 0.0218604f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=1.325
cc_69 VPB N_A_27_297#_M1006_g 0.0220154f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=1.325
cc_70 VPB N_A_27_297#_c_312_n 0.0206091f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_297#_c_322_n 0.0079379f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.53
cc_72 VPB N_A_27_297#_c_323_n 0.0153085f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_73 VPB N_A_27_297#_c_324_n 0.00177887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_297#_c_315_n 0.00373325f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_75 VPB N_A_27_297#_c_326_n 0.0274163f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.53
cc_76 VPB N_A_27_297#_c_318_n 0.00428376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_448_n 0.00454762f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=1.325
cc_78 VPB N_VPWR_c_449_n 0.00454762f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=0.995
cc_79 VPB N_VPWR_c_450_n 0.00516508f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=1.985
cc_80 VPB N_VPWR_c_451_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.18
cc_81 VPB N_VPWR_c_452_n 0.0131574f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_82 VPB N_VPWR_c_453_n 0.0375473f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.285
cc_83 VPB N_VPWR_c_454_n 0.0379282f $X=-0.19 $Y=1.305 $X2=3.015 $Y2=1.445
cc_84 VPB N_VPWR_c_455_n 0.00478242f $X=-0.19 $Y=1.305 $X2=3.1 $Y2=1.18
cc_85 VPB N_VPWR_c_456_n 0.0167335f $X=-0.19 $Y=1.305 $X2=3.755 $Y2=1.16
cc_86 VPB N_VPWR_c_457_n 0.0151708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_458_n 0.0312617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_459_n 0.0169155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_460_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_461_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_462_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_447_n 0.0506842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_Y_c_612_n 0.0081428f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_94 VPB N_Y_c_611_n 0.0074506f $X=-0.19 $Y=1.305 $X2=4.02 $Y2=0.56
cc_95 VPB Y 0.0171019f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.285
cc_96 N_B_c_97_n N_A_c_215_n 0.0195418f $X=0.905 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_97 N_B_M1018_g N_A_M1009_g 0.0195418f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B_c_110_n N_A_M1009_g 0.010384f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_99 N_B_c_110_n N_A_M1011_g 0.0124706f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_100 N_B_c_108_n N_A_M1002_g 0.0025712f $X=3.015 $Y=1.445 $X2=0 $Y2=0
cc_101 N_B_c_110_n N_A_M1002_g 0.0148082f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_102 N_B_c_98_n N_A_c_218_n 0.0279744f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B_M1012_g N_A_M1005_g 0.0279744f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B_c_108_n N_A_M1005_g 0.00286987f $X=3.015 $Y=1.445 $X2=0 $Y2=0
cc_105 N_B_c_110_n N_A_M1005_g 0.00440759f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_106 N_B_c_110_n N_A_c_219_n 0.0154578f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_107 N_B_c_108_n N_A_c_220_n 0.00389291f $X=3.015 $Y=1.445 $X2=0 $Y2=0
cc_108 N_B_c_125_p N_A_c_220_n 0.00933351f $X=3.1 $Y=1.18 $X2=0 $Y2=0
cc_109 N_B_c_100_n N_A_c_220_n 0.0093613f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B_c_110_n N_A_c_220_n 0.00111167f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_111 N_B_c_102_n N_A_c_220_n 0.0279744f $X=4.02 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B_c_129_p N_A_c_221_n 9.43616e-19 $X=0.79 $Y=1.18 $X2=0 $Y2=0
cc_113 N_B_c_107_n N_A_c_221_n 0.00100797f $X=0.875 $Y=1.445 $X2=0 $Y2=0
cc_114 N_B_c_110_n N_A_c_221_n 0.00214031f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_115 N_B_c_101_n N_A_c_221_n 0.0195418f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B_c_129_p N_A_c_249_n 0.010458f $X=0.79 $Y=1.18 $X2=0 $Y2=0
cc_117 N_B_c_125_p N_A_c_249_n 0.0133646f $X=3.1 $Y=1.18 $X2=0 $Y2=0
cc_118 N_B_c_110_n N_A_c_249_n 0.103577f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_119 N_B_c_101_n N_A_c_249_n 8.44684e-19 $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_c_110_n N_A_27_297#_M1018_s 0.00165831f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_121 N_B_c_110_n N_A_27_297#_M1011_d 0.00308507f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_122 N_B_c_96_n N_A_27_297#_c_312_n 0.0279065f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_129_p N_A_27_297#_c_312_n 0.0165247f $X=0.79 $Y=1.18 $X2=0 $Y2=0
cc_124 N_B_c_107_n N_A_27_297#_c_312_n 0.00583811f $X=0.875 $Y=1.445 $X2=0 $Y2=0
cc_125 N_B_c_109_n N_A_27_297#_c_312_n 0.00396363f $X=0.96 $Y=1.53 $X2=0 $Y2=0
cc_126 N_B_c_96_n N_A_27_297#_c_314_n 0.0152531f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_97_n N_A_27_297#_c_314_n 0.00351551f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B_c_129_p N_A_27_297#_c_314_n 0.0268528f $X=0.79 $Y=1.18 $X2=0 $Y2=0
cc_129 N_B_c_101_n N_A_27_297#_c_314_n 0.00222641f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_M1003_g N_A_27_297#_c_338_n 0.013602f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B_M1018_g N_A_27_297#_c_338_n 0.0104707f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B_c_129_p N_A_27_297#_c_338_n 0.00804975f $X=0.79 $Y=1.18 $X2=0 $Y2=0
cc_133 N_B_c_109_n N_A_27_297#_c_338_n 0.00971246f $X=0.96 $Y=1.53 $X2=0 $Y2=0
cc_134 N_B_c_110_n N_A_27_297#_c_338_n 0.00129352f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_135 N_B_c_101_n N_A_27_297#_c_338_n 0.00165009f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B_c_110_n N_A_27_297#_c_344_n 0.0317352f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_137 N_B_c_100_n N_A_27_297#_c_322_n 0.00559778f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B_c_110_n N_A_27_297#_c_322_n 0.0608669f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_139 N_B_M1012_g N_A_27_297#_c_323_n 0.0118326f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B_M1017_g N_A_27_297#_c_323_n 0.0143203f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B_c_100_n N_A_27_297#_c_323_n 0.0339105f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B_c_102_n N_A_27_297#_c_323_n 0.00293762f $X=4.02 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B_c_100_n N_A_27_297#_c_324_n 0.0142097f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B_c_110_n N_A_27_297#_c_324_n 0.0119195f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_145 N_B_c_102_n N_A_27_297#_c_315_n 0.00519427f $X=4.02 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B_c_100_n N_A_27_297#_c_316_n 0.00519147f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B_c_102_n N_A_27_297#_c_316_n 0.00358725f $X=4.02 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B_c_110_n N_A_27_297#_c_356_n 0.0126919f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_149 N_B_c_110_n N_A_27_297#_c_357_n 0.0165158f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_150 N_B_c_110_n N_VPWR_M1009_s 0.00166235f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_151 N_B_c_110_n N_VPWR_M1002_s 0.00164824f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_152 N_B_M1003_g N_VPWR_c_448_n 0.00302074f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B_M1018_g N_VPWR_c_448_n 0.00157837f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B_M1017_g N_VPWR_c_451_n 0.00214938f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B_M1012_g N_VPWR_c_454_n 0.00359305f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B_M1017_g N_VPWR_c_454_n 0.00357877f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B_M1003_g N_VPWR_c_456_n 0.00441875f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_158 N_B_M1018_g N_VPWR_c_457_n 0.00441875f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B_M1003_g N_VPWR_c_447_n 0.0068285f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B_M1018_g N_VPWR_c_447_n 0.00588739f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B_M1012_g N_VPWR_c_447_n 0.00486683f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_162 N_B_M1017_g N_VPWR_c_447_n 0.00664485f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_163 N_B_c_110_n N_A_474_297#_M1002_d 0.00304026f $X=2.93 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_164 N_B_M1012_g N_A_474_297#_c_554_n 0.0065265f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B_M1017_g N_A_474_297#_c_554_n 0.00872269f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_166 N_B_M1012_g N_A_474_297#_c_556_n 0.00411447f $X=3.565 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_B_M1017_g N_A_474_297#_c_556_n 8.39194e-19 $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_168 N_B_M1012_g N_A_474_297#_c_558_n 0.00590837f $X=3.565 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_B_M1017_g N_A_474_297#_c_558_n 7.98874e-19 $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_170 N_B_M1017_g N_Y_c_612_n 0.0113377f $X=4.02 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B_c_96_n N_A_27_47#_c_661_n 0.00892725f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B_c_97_n N_A_27_47#_c_661_n 0.0109056f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B_c_129_p N_A_27_47#_c_661_n 0.00267312f $X=0.79 $Y=1.18 $X2=0 $Y2=0
cc_174 N_B_c_97_n N_A_27_47#_c_662_n 4.16929e-19 $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B_c_110_n N_A_27_47#_c_662_n 0.00843334f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_176 N_B_c_98_n N_VGND_c_705_n 0.00268723f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B_c_99_n N_VGND_c_706_n 0.00438629f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B_c_96_n N_VGND_c_707_n 0.00357877f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B_c_97_n N_VGND_c_707_n 0.00357877f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B_c_98_n N_VGND_c_713_n 0.00423334f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B_c_99_n N_VGND_c_713_n 0.00423334f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B_c_96_n N_VGND_c_716_n 0.00619348f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B_c_97_n N_VGND_c_716_n 0.00525237f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_98_n N_VGND_c_716_n 0.00583365f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B_c_99_n N_VGND_c_716_n 0.00713252f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B_c_98_n N_A_560_47#_c_796_n 5.22228e-19 $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_c_98_n N_A_560_47#_c_791_n 0.00865686f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B_c_100_n N_A_560_47#_c_791_n 0.0372562f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B_c_125_p N_A_560_47#_c_792_n 0.0147217f $X=3.1 $Y=1.18 $X2=0 $Y2=0
cc_190 N_B_c_110_n N_A_560_47#_c_792_n 0.00574269f $X=2.93 $Y=1.53 $X2=0 $Y2=0
cc_191 N_B_c_98_n N_A_560_47#_c_801_n 0.00630972f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B_c_99_n N_A_560_47#_c_801_n 0.0110139f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B_c_98_n N_A_560_47#_c_793_n 0.00115677f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B_c_99_n N_A_560_47#_c_793_n 0.00140826f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B_c_100_n N_A_560_47#_c_793_n 0.0279387f $X=3.755 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B_c_102_n N_A_560_47#_c_793_n 0.00319915f $X=4.02 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B_c_99_n N_A_560_47#_c_795_n 0.0124093f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_M1009_g N_A_27_297#_c_344_n 0.0104325f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_M1011_g N_A_27_297#_c_344_n 0.0104897f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_M1002_g N_A_27_297#_c_322_n 0.0126468f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_M1005_g N_A_27_297#_c_322_n 0.01158f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_c_220_n N_A_27_297#_c_322_n 2.49536e-19 $X=3.145 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_M1005_g N_A_27_297#_c_363_n 0.00359553f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_M1005_g N_A_27_297#_c_324_n 0.00160334f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_M1002_g N_A_27_297#_c_357_n 0.00445973f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A_M1009_g N_VPWR_c_449_n 0.00157837f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_M1011_g N_VPWR_c_449_n 0.00302074f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_M1002_g N_VPWR_c_450_n 0.00321753f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_M1005_g N_VPWR_c_450_n 0.00321753f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_M1005_g N_VPWR_c_454_n 0.00585385f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_M1009_g N_VPWR_c_457_n 0.00441875f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_M1011_g N_VPWR_c_458_n 0.00441875f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_M1002_g N_VPWR_c_458_n 0.00585385f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_M1009_g N_VPWR_c_447_n 0.00588739f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_M1011_g N_VPWR_c_447_n 0.00718625f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_M1002_g N_VPWR_c_447_n 0.00609727f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_M1005_g N_VPWR_c_447_n 0.00483015f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_M1002_g N_A_474_297#_c_560_n 0.00165616f $X=2.725 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_M1005_g N_A_474_297#_c_560_n 0.00237973f $X=3.145 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_M1002_g N_A_474_297#_c_562_n 0.00183751f $X=2.725 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_M1005_g N_A_474_297#_c_556_n 4.31699e-19 $X=3.145 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_c_215_n N_A_27_47#_c_670_n 0.00255288f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_c_215_n N_A_27_47#_c_662_n 0.00492325f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_c_216_n N_A_27_47#_c_662_n 4.58193e-19 $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_c_249_n N_A_27_47#_c_662_n 0.00191873f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_c_215_n N_A_27_47#_c_663_n 0.00870364f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_216_n N_A_27_47#_c_663_n 0.00995225f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_c_219_n N_A_27_47#_c_663_n 0.00537465f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_c_221_n N_A_27_47#_c_663_n 0.00222133f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_c_249_n N_A_27_47#_c_663_n 0.0627481f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_c_215_n N_A_27_47#_c_664_n 5.22228e-19 $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_216_n N_A_27_47#_c_664_n 0.00630972f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_c_215_n N_VGND_c_703_n 0.00268723f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_c_216_n N_VGND_c_703_n 0.00268723f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_c_216_n N_VGND_c_704_n 0.00298279f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_c_217_n N_VGND_c_704_n 0.00360182f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_c_219_n N_VGND_c_704_n 0.00331219f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_c_249_n N_VGND_c_704_n 0.0136993f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_c_218_n N_VGND_c_705_n 0.00146448f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_c_215_n N_VGND_c_707_n 0.00421816f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_c_216_n N_VGND_c_709_n 0.00423334f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_217_n N_VGND_c_711_n 0.00541359f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_218_n N_VGND_c_711_n 0.00423334f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_215_n N_VGND_c_716_n 0.00575258f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_216_n N_VGND_c_716_n 0.00704237f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_217_n N_VGND_c_716_n 0.0108276f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_c_218_n N_VGND_c_716_n 0.0057435f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_c_217_n N_A_560_47#_c_796_n 0.00539651f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_c_218_n N_A_560_47#_c_796_n 0.00630972f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_218_n N_A_560_47#_c_791_n 0.00865686f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_217_n N_A_560_47#_c_792_n 0.00300399f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_218_n N_A_560_47#_c_792_n 0.00113159f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_c_220_n N_A_560_47#_c_792_n 0.00254391f $X=3.145 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_c_218_n N_A_560_47#_c_801_n 5.21666e-19 $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_27_297#_c_338_n N_VPWR_M1003_d 0.00417282f $X=0.99 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A_27_297#_c_344_n N_VPWR_M1009_s 0.00317395f $X=1.83 $Y=1.875 $X2=0
+ $Y2=0
cc_257 N_A_27_297#_c_322_n N_VPWR_M1002_s 0.00307924f $X=3.31 $Y=1.87 $X2=0
+ $Y2=0
cc_258 N_A_27_297#_c_323_n N_VPWR_M1001_d 0.00464908f $X=4.635 $Y=1.54 $X2=0
+ $Y2=0
cc_259 N_A_27_297#_c_338_n N_VPWR_c_448_n 0.0123469f $X=0.99 $Y=1.875 $X2=0
+ $Y2=0
cc_260 N_A_27_297#_c_344_n N_VPWR_c_449_n 0.0123469f $X=1.83 $Y=1.875 $X2=0
+ $Y2=0
cc_261 N_A_27_297#_c_322_n N_VPWR_c_450_n 0.011057f $X=3.31 $Y=1.87 $X2=0 $Y2=0
cc_262 N_A_27_297#_M1001_g N_VPWR_c_451_n 0.00338128f $X=4.96 $Y=1.985 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_M1006_g N_VPWR_c_453_n 0.00345498f $X=5.38 $Y=1.985 $X2=0
+ $Y2=0
cc_264 N_A_27_297#_c_338_n N_VPWR_c_456_n 0.0020229f $X=0.99 $Y=1.875 $X2=0
+ $Y2=0
cc_265 N_A_27_297#_c_326_n N_VPWR_c_456_n 0.0204751f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_266 N_A_27_297#_c_338_n N_VPWR_c_457_n 0.0020229f $X=0.99 $Y=1.875 $X2=0
+ $Y2=0
cc_267 N_A_27_297#_c_344_n N_VPWR_c_457_n 0.0020229f $X=1.83 $Y=1.875 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_c_356_n N_VPWR_c_457_n 0.0142343f $X=1.115 $Y=1.96 $X2=0
+ $Y2=0
cc_269 N_A_27_297#_c_344_n N_VPWR_c_458_n 0.0020229f $X=1.83 $Y=1.875 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_c_357_n N_VPWR_c_458_n 0.0158369f $X=1.955 $Y=1.96 $X2=0
+ $Y2=0
cc_271 N_A_27_297#_M1001_g N_VPWR_c_459_n 0.00441875f $X=4.96 $Y=1.985 $X2=0
+ $Y2=0
cc_272 N_A_27_297#_M1006_g N_VPWR_c_459_n 0.00585385f $X=5.38 $Y=1.985 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_M1003_s N_VPWR_c_447_n 0.0022569f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_M1018_s N_VPWR_c_447_n 0.0022335f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_M1011_d N_VPWR_c_447_n 0.00240124f $X=1.82 $Y=1.485 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_M1001_g N_VPWR_c_447_n 0.0072312f $X=4.96 $Y=1.985 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_M1006_g N_VPWR_c_447_n 0.0115702f $X=5.38 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_A_27_297#_c_338_n N_VPWR_c_447_n 0.00802398f $X=0.99 $Y=1.875 $X2=0
+ $Y2=0
cc_279 N_A_27_297#_c_344_n N_VPWR_c_447_n 0.00802398f $X=1.83 $Y=1.875 $X2=0
+ $Y2=0
cc_280 N_A_27_297#_c_322_n N_VPWR_c_447_n 0.0117001f $X=3.31 $Y=1.87 $X2=0 $Y2=0
cc_281 N_A_27_297#_c_326_n N_VPWR_c_447_n 0.0120542f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_c_356_n N_VPWR_c_447_n 0.00955092f $X=1.115 $Y=1.96 $X2=0
+ $Y2=0
cc_283 N_A_27_297#_c_357_n N_VPWR_c_447_n 0.00955092f $X=1.955 $Y=1.96 $X2=0
+ $Y2=0
cc_284 N_A_27_297#_c_322_n N_A_474_297#_M1002_d 0.00539951f $X=3.31 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_285 N_A_27_297#_c_322_n N_A_474_297#_M1005_d 0.00236176f $X=3.31 $Y=1.87
+ $X2=0 $Y2=0
cc_286 N_A_27_297#_c_363_n N_A_474_297#_M1005_d 0.00175548f $X=3.395 $Y=1.785
+ $X2=0 $Y2=0
cc_287 N_A_27_297#_c_324_n N_A_474_297#_M1005_d 0.00132259f $X=3.48 $Y=1.54
+ $X2=0 $Y2=0
cc_288 N_A_27_297#_c_323_n N_A_474_297#_M1017_s 0.00276803f $X=4.635 $Y=1.54
+ $X2=0 $Y2=0
cc_289 N_A_27_297#_c_323_n N_A_474_297#_c_554_n 0.00184635f $X=4.635 $Y=1.54
+ $X2=0 $Y2=0
cc_290 N_A_27_297#_c_322_n N_A_474_297#_c_560_n 0.0133232f $X=3.31 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_c_322_n N_A_474_297#_c_562_n 0.00905671f $X=3.31 $Y=1.87
+ $X2=0 $Y2=0
cc_292 N_A_27_297#_c_357_n N_A_474_297#_c_562_n 0.00270019f $X=1.955 $Y=1.96
+ $X2=0 $Y2=0
cc_293 N_A_27_297#_c_322_n N_A_474_297#_c_573_n 0.0139782f $X=3.31 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_c_357_n N_A_474_297#_c_573_n 0.0152341f $X=1.955 $Y=1.96
+ $X2=0 $Y2=0
cc_295 N_A_27_297#_c_322_n N_A_474_297#_c_556_n 0.0045174f $X=3.31 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_27_297#_c_323_n N_A_474_297#_c_556_n 0.00259926f $X=4.635 $Y=1.54
+ $X2=0 $Y2=0
cc_297 N_A_27_297#_c_322_n N_A_474_297#_c_558_n 0.0118411f $X=3.31 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_27_297#_c_323_n N_A_474_297#_c_558_n 0.00109076f $X=4.635 $Y=1.54
+ $X2=0 $Y2=0
cc_299 N_A_27_297#_c_323_n N_Y_M1012_d 0.00233412f $X=4.635 $Y=1.54 $X2=0 $Y2=0
cc_300 N_A_27_297#_M1001_g N_Y_c_612_n 0.0141764f $X=4.96 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_323_n N_Y_c_612_n 0.0594936f $X=4.635 $Y=1.54 $X2=0 $Y2=0
cc_302 N_A_27_297#_c_317_n N_Y_c_612_n 0.0056604f $X=5.13 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_27_297#_c_310_n N_Y_c_609_n 0.0083291f $X=4.96 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_27_297#_c_311_n N_Y_c_609_n 0.0115911f $X=5.38 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_27_297#_c_311_n N_Y_c_611_n 0.0213879f $X=5.38 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_27_297#_c_317_n N_Y_c_611_n 0.0121436f $X=5.13 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A_27_297#_c_323_n N_Y_c_624_n 0.0124408f $X=4.635 $Y=1.54 $X2=0 $Y2=0
cc_308 N_A_27_297#_M1001_g Y 7.03933e-19 $X=4.96 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_27_297#_M1006_g Y 0.0210846f $X=5.38 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_27_297#_c_323_n Y 0.00700876f $X=4.635 $Y=1.54 $X2=0 $Y2=0
cc_311 N_A_27_297#_c_315_n Y 0.00255273f $X=4.72 $Y=1.455 $X2=0 $Y2=0
cc_312 N_A_27_297#_c_317_n Y 0.0181901f $X=5.13 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_27_297#_c_318_n Y 0.00222985f $X=5.38 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_27_297#_c_313_n N_A_27_47#_M1008_d 0.00318623f $X=0.315 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_315 N_A_27_297#_c_314_n N_A_27_47#_M1008_d 3.84519e-19 $X=0.695 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_316 N_A_27_297#_M1008_s N_A_27_47#_c_661_n 0.00305026f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_317 N_A_27_297#_c_313_n N_A_27_47#_c_661_n 0.0165567f $X=0.315 $Y=0.77 $X2=0
+ $Y2=0
cc_318 N_A_27_297#_c_314_n N_A_27_47#_c_661_n 0.0260973f $X=0.695 $Y=0.73 $X2=0
+ $Y2=0
cc_319 N_A_27_297#_c_314_n N_A_27_47#_c_662_n 0.00752753f $X=0.695 $Y=0.73 $X2=0
+ $Y2=0
cc_320 N_A_27_297#_c_310_n N_VGND_c_706_n 0.00252945f $X=4.96 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_27_297#_c_313_n N_VGND_c_707_n 3.97819e-19 $X=0.315 $Y=0.77 $X2=0
+ $Y2=0
cc_322 N_A_27_297#_c_310_n N_VGND_c_715_n 0.00368123f $X=4.96 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_27_297#_c_311_n N_VGND_c_715_n 0.00368123f $X=5.38 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_27_297#_M1008_s N_VGND_c_716_n 0.00216833f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_325 N_A_27_297#_c_310_n N_VGND_c_716_n 0.00657241f $X=4.96 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A_27_297#_c_311_n N_VGND_c_716_n 0.00630397f $X=5.38 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_27_297#_c_313_n N_VGND_c_716_n 0.00112342f $X=0.315 $Y=0.77 $X2=0
+ $Y2=0
cc_328 N_A_27_297#_c_323_n N_A_560_47#_c_793_n 5.77138e-19 $X=4.635 $Y=1.54
+ $X2=0 $Y2=0
cc_329 N_A_27_297#_c_310_n N_A_560_47#_c_794_n 0.00498188f $X=4.96 $Y=0.995
+ $X2=0 $Y2=0
cc_330 N_A_27_297#_c_311_n N_A_560_47#_c_794_n 0.00422352f $X=5.38 $Y=0.995
+ $X2=0 $Y2=0
cc_331 N_A_27_297#_c_318_n N_A_560_47#_c_794_n 0.00224214f $X=5.38 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_27_297#_c_310_n N_A_560_47#_c_795_n 0.00990301f $X=4.96 $Y=0.995
+ $X2=0 $Y2=0
cc_333 N_A_27_297#_c_323_n N_A_560_47#_c_795_n 0.0211811f $X=4.635 $Y=1.54 $X2=0
+ $Y2=0
cc_334 N_A_27_297#_c_316_n N_A_560_47#_c_795_n 0.0141654f $X=4.805 $Y=1.16 $X2=0
+ $Y2=0
cc_335 N_A_27_297#_c_317_n N_A_560_47#_c_795_n 0.0355006f $X=5.13 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_447_n N_A_474_297#_M1002_d 0.00145723f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_337 N_VPWR_c_447_n N_A_474_297#_M1005_d 0.00117976f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_447_n N_A_474_297#_M1017_s 0.00207714f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_454_n N_A_474_297#_c_554_n 0.0309112f $X=4.625 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_447_n N_A_474_297#_c_554_n 0.0178255f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_451_n N_A_474_297#_c_584_n 0.0180653f $X=4.75 $Y=2.3 $X2=0 $Y2=0
cc_342 N_VPWR_c_454_n N_A_474_297#_c_584_n 0.0151213f $X=4.625 $Y=2.72 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_447_n N_A_474_297#_c_584_n 0.00938089f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_344 N_VPWR_M1002_s N_A_474_297#_c_560_n 2.19468e-19 $X=2.8 $Y=1.485 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_450_n N_A_474_297#_c_560_n 0.013287f $X=2.935 $Y=2.3 $X2=0 $Y2=0
cc_346 N_VPWR_c_454_n N_A_474_297#_c_560_n 8.75468e-19 $X=4.625 $Y=2.72 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_458_n N_A_474_297#_c_560_n 5.44986e-19 $X=2.81 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_447_n N_A_474_297#_c_560_n 0.0519243f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_450_n N_A_474_297#_c_562_n 0.00133907f $X=2.935 $Y=2.3 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_458_n N_A_474_297#_c_562_n 4.35969e-19 $X=2.81 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_447_n N_A_474_297#_c_562_n 0.0282617f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_450_n N_A_474_297#_c_573_n 0.00589098f $X=2.935 $Y=2.3 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_458_n N_A_474_297#_c_573_n 0.0151494f $X=2.81 $Y=2.72 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_447_n N_A_474_297#_c_573_n 0.00264208f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_450_n N_A_474_297#_c_556_n 3.05262e-19 $X=2.935 $Y=2.3 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_447_n N_A_474_297#_c_556_n 0.0280917f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_450_n N_A_474_297#_c_558_n 0.0050191f $X=2.935 $Y=2.3 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_454_n N_A_474_297#_c_558_n 0.0182182f $X=4.625 $Y=2.72 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_447_n N_A_474_297#_c_558_n 0.00293817f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_447_n N_Y_M1012_d 0.00244138f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_361 N_VPWR_c_447_n N_Y_M1001_s 0.00333586f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_362 N_VPWR_M1001_d N_Y_c_612_n 0.0051974f $X=4.625 $Y=1.485 $X2=0 $Y2=0
cc_363 N_VPWR_c_451_n N_Y_c_612_n 0.0159284f $X=4.75 $Y=2.3 $X2=0 $Y2=0
cc_364 N_VPWR_c_454_n N_Y_c_612_n 0.0039015f $X=4.625 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_c_459_n N_Y_c_612_n 0.00201582f $X=5.465 $Y=2.72 $X2=0 $Y2=0
cc_366 N_VPWR_c_447_n N_Y_c_612_n 0.012325f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_367 N_VPWR_c_459_n N_Y_c_638_n 0.00424887f $X=5.465 $Y=2.72 $X2=0 $Y2=0
cc_368 N_VPWR_c_447_n N_Y_c_638_n 0.00763999f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_M1006_d Y 0.0031554f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_370 N_VPWR_c_453_n Y 0.0320301f $X=5.59 $Y=1.96 $X2=0 $Y2=0
cc_371 N_A_474_297#_c_554_n N_Y_M1012_d 0.00412801f $X=4.105 $Y=2.38 $X2=0.485
+ $Y2=0.56
cc_372 N_A_474_297#_M1017_s N_Y_c_612_n 0.00500976f $X=4.095 $Y=1.485 $X2=0.905
+ $Y2=1.985
cc_373 N_A_474_297#_c_554_n N_Y_c_612_n 0.00520504f $X=4.105 $Y=2.38 $X2=0.905
+ $Y2=1.985
cc_374 N_A_474_297#_c_584_n N_Y_c_612_n 0.0150265f $X=4.23 $Y=2.3 $X2=0.905
+ $Y2=1.985
cc_375 N_A_474_297#_c_554_n N_Y_c_624_n 0.0116894f $X=4.105 $Y=2.38 $X2=4.02
+ $Y2=1.325
cc_376 N_A_474_297#_c_556_n N_Y_c_624_n 0.00147036f $X=3.47 $Y=2.21 $X2=4.02
+ $Y2=1.325
cc_377 N_Y_c_609_n N_VGND_c_706_n 0.0100248f $X=5.505 $Y=0.39 $X2=0 $Y2=0
cc_378 N_Y_c_609_n N_VGND_c_715_n 0.039179f $X=5.505 $Y=0.39 $X2=0 $Y2=0
cc_379 N_Y_c_610_n N_VGND_c_715_n 0.0207814f $X=5.7 $Y=0.475 $X2=0 $Y2=0
cc_380 N_Y_M1000_d N_VGND_c_716_n 0.0021262f $X=4.625 $Y=0.235 $X2=0 $Y2=0
cc_381 N_Y_M1004_d N_VGND_c_716_n 0.00212536f $X=5.455 $Y=0.235 $X2=0 $Y2=0
cc_382 N_Y_c_609_n N_VGND_c_716_n 0.0316767f $X=5.505 $Y=0.39 $X2=0 $Y2=0
cc_383 N_Y_c_610_n N_VGND_c_716_n 0.0146438f $X=5.7 $Y=0.475 $X2=0 $Y2=0
cc_384 N_Y_c_609_n N_A_560_47#_M1000_s 0.00318958f $X=5.505 $Y=0.39 $X2=0 $Y2=0
cc_385 N_Y_c_609_n N_A_560_47#_c_794_n 0.015032f $X=5.505 $Y=0.39 $X2=0 $Y2=0
cc_386 N_Y_c_611_n N_A_560_47#_c_794_n 0.0112926f $X=5.59 $Y=0.73 $X2=0 $Y2=0
cc_387 Y N_A_560_47#_c_794_n 0.0012404f $X=5.705 $Y=1.445 $X2=0 $Y2=0
cc_388 N_Y_M1000_d N_A_560_47#_c_795_n 0.00319929f $X=4.625 $Y=0.235 $X2=0 $Y2=0
cc_389 N_Y_c_609_n N_A_560_47#_c_795_n 0.0177508f $X=5.505 $Y=0.39 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_663_n N_VGND_M1007_d 0.00162089f $X=1.79 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_391 N_A_27_47#_c_663_n N_VGND_c_703_n 0.0122559f $X=1.79 $Y=0.815 $X2=0 $Y2=0
cc_392 N_A_27_47#_c_663_n N_VGND_c_704_n 0.00976972f $X=1.79 $Y=0.815 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_664_n N_VGND_c_704_n 0.0238522f $X=1.955 $Y=0.39 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_661_n N_VGND_c_707_n 0.052604f $X=1.03 $Y=0.365 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_670_n N_VGND_c_707_n 0.0152108f $X=1.155 $Y=0.475 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_663_n N_VGND_c_707_n 0.00198695f $X=1.79 $Y=0.815 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_663_n N_VGND_c_709_n 0.00198695f $X=1.79 $Y=0.815 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_664_n N_VGND_c_709_n 0.0209479f $X=1.955 $Y=0.39 $X2=0 $Y2=0
cc_399 N_A_27_47#_M1008_d N_VGND_c_716_n 0.00221642f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_M1015_d N_VGND_c_716_n 0.00215206f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_M1013_s N_VGND_c_716_n 0.00225715f $X=1.82 $Y=0.235 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_661_n N_VGND_c_716_n 0.0331327f $X=1.03 $Y=0.365 $X2=0 $Y2=0
cc_403 N_A_27_47#_c_670_n N_VGND_c_716_n 0.00940698f $X=1.155 $Y=0.475 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_663_n N_VGND_c_716_n 0.00835832f $X=1.79 $Y=0.815 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_664_n N_VGND_c_716_n 0.0124119f $X=1.955 $Y=0.39 $X2=0 $Y2=0
cc_406 N_VGND_c_716_n N_A_560_47#_M1014_d 0.00215201f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_407 N_VGND_c_716_n N_A_560_47#_M1010_s 0.00243306f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_716_n N_A_560_47#_M1000_s 0.00220248f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_711_n N_A_560_47#_c_796_n 0.0188551f $X=3.27 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_716_n N_A_560_47#_c_796_n 0.0122069f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_M1019_s N_A_560_47#_c_791_n 0.00162089f $X=3.22 $Y=0.235 $X2=0
+ $Y2=0
cc_412 N_VGND_c_705_n N_A_560_47#_c_791_n 0.0122559f $X=3.355 $Y=0.39 $X2=0
+ $Y2=0
cc_413 N_VGND_c_711_n N_A_560_47#_c_791_n 0.00198695f $X=3.27 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_713_n N_A_560_47#_c_791_n 0.00198695f $X=4.145 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_716_n N_A_560_47#_c_791_n 0.00835832f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_704_n N_A_560_47#_c_792_n 0.00830019f $X=2.515 $Y=0.39 $X2=0
+ $Y2=0
cc_417 N_VGND_c_713_n N_A_560_47#_c_801_n 0.0213082f $X=4.145 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_716_n N_A_560_47#_c_801_n 0.0135533f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_M1016_d N_A_560_47#_c_795_n 0.00315681f $X=4.095 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_VGND_c_706_n N_A_560_47#_c_795_n 0.0127273f $X=4.23 $Y=0.39 $X2=0 $Y2=0
cc_421 N_VGND_c_713_n N_A_560_47#_c_795_n 0.00198695f $X=4.145 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_715_n N_A_560_47#_c_795_n 0.00409419f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_716_n N_A_560_47#_c_795_n 0.012649f $X=5.75 $Y=0 $X2=0 $Y2=0

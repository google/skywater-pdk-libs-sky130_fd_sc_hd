* File: sky130_fd_sc_hd__xnor2_1.spice.pex
* Created: Thu Aug 27 14:48:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XNOR2_1%B 3 7 10 14 16 17 19 20 22 23 28 29 30 32 36
c91 28 0 1.4951e-19 $X=0.51 $Y=1.16
c92 20 0 9.65133e-20 $X=2.23 $Y=1.16
r93 34 36 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.67 $Y=1.53 $X2=0.69
+ $Y2=1.53
r94 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r95 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r96 23 34 4.20453 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.547 $Y=1.53
+ $X2=0.67 $Y2=1.53
r97 23 29 11.134 $w=3.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.547 $Y=1.445
+ $X2=0.547 $Y2=1.16
r98 23 36 2.0877 $w=1.68e-07 $l=3.2e-08 $layer=LI1_cond $X=0.722 $Y=1.53
+ $X2=0.69 $Y2=1.53
r99 22 23 70.0032 $w=1.68e-07 $l=1.073e-06 $layer=LI1_cond $X=1.795 $Y=1.53
+ $X2=0.722 $Y2=1.53
r100 20 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=1.325
r101 20 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=0.995
r102 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.16 $X2=2.23 $Y2=1.16
r103 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.965 $Y=1.16
+ $X2=2.23 $Y2=1.16
r104 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.88 $Y=1.445
+ $X2=1.795 $Y2=1.53
r105 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.88 $Y=1.245
+ $X2=1.965 $Y2=1.16
r106 15 16 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=1.245
+ $X2=1.88 $Y2=1.445
r107 14 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.29 $Y=0.56
+ $X2=2.29 $Y2=0.995
r108 10 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.985
+ $X2=2.17 $Y2=1.325
r109 7 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.57 $Y=0.56
+ $X2=0.57 $Y2=0.995
r110 1 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.325
+ $X2=0.51 $Y2=1.16
r111 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.51 $Y=1.325
+ $X2=0.51 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_1%A 1 3 6 8 10 13 15 22 23
c49 22 0 9.65133e-20 $X=1.435 $Y=1.16
c50 13 0 1.71597e-19 $X=1.81 $Y=1.985
r51 21 23 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.435 $Y=1.16
+ $X2=1.81 $Y2=1.16
r52 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.435
+ $Y=1.16 $X2=1.435 $Y2=1.16
r53 19 21 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.35 $Y=1.16
+ $X2=1.435 $Y2=1.16
r54 17 19 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=1.35 $Y2=1.16
r55 15 22 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=1.435 $Y2=1.175
r56 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.325
+ $X2=1.81 $Y2=1.16
r57 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.81 $Y=1.325
+ $X2=1.81 $Y2=1.985
r58 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=1.16
r59 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=0.56
r60 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.16
r61 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.93 $Y=1.325 $X2=0.93
+ $Y2=1.985
r62 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r63 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.93 $Y=0.995 $X2=0.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_1%A_47_47# 1 2 9 11 13 15 16 17 20 22 25 26 27
+ 30 31 34 37
c105 37 0 1.4951e-19 $X=0.72 $Y=1.87
c106 27 0 1.71597e-19 $X=2.305 $Y=1.5
r107 34 36 16.2536 $w=4.63e-07 $l=4.35e-07 $layer=LI1_cond $X=0.317 $Y=0.39
+ $X2=0.317 $Y2=0.825
r108 31 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=1.325
r109 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.16 $X2=2.71 $Y2=1.16
r110 28 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.71 $Y=1.415
+ $X2=2.71 $Y2=1.16
r111 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.625 $Y=1.5
+ $X2=2.71 $Y2=1.415
r112 26 27 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.625 $Y=1.5
+ $X2=2.305 $Y2=1.5
r113 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=1.585
+ $X2=2.305 $Y2=1.5
r114 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.22 $Y=1.585
+ $X2=2.22 $Y2=1.785
r115 23 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=1.87
+ $X2=0.72 $Y2=1.87
r116 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=1.87
+ $X2=2.22 $Y2=1.785
r117 22 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.135 $Y=1.87
+ $X2=0.885 $Y2=1.87
r118 18 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.955
+ $X2=0.72 $Y2=1.87
r119 18 20 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.955
+ $X2=0.72 $Y2=1.96
r120 16 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=1.87
+ $X2=0.72 $Y2=1.87
r121 16 17 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.555 $Y=1.87
+ $X2=0.255 $Y2=1.87
r122 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.785
+ $X2=0.255 $Y2=1.87
r123 15 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.17 $Y=1.785
+ $X2=0.17 $Y2=0.825
r124 11 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.995
+ $X2=2.71 $Y2=1.16
r125 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.71 $Y=0.995
+ $X2=2.71 $Y2=0.56
r126 9 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.65 $Y=1.985
+ $X2=2.65 $Y2=1.325
r127 2 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.72 $Y2=1.96
r128 1 34 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_1%VPWR 1 2 3 10 12 14 16 18 25 36 42 45
r50 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 40 42 9.09332 $w=6.78e-07 $l=7.5e-08 $layer=LI1_cond $X=1.61 $Y=2.465
+ $X2=1.685 $Y2=2.465
r52 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 38 40 0.175894 $w=6.78e-07 $l=1e-08 $layer=LI1_cond $X=1.6 $Y=2.465 $X2=1.61
+ $Y2=2.465
r54 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 34 38 7.91522 $w=6.78e-07 $l=4.5e-07 $layer=LI1_cond $X=1.15 $Y=2.465
+ $X2=1.6 $Y2=2.465
r56 34 36 9.44511 $w=6.78e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=2.465
+ $X2=1.055 $Y2=2.465
r57 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 29 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 29 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 28 42 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=1.685 $Y2=2.72
r61 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 25 44 4.47956 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=3.017 $Y2=2.72
r63 25 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 23 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.055 $Y2=2.72
r66 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 21 31 4.51997 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r68 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 18 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 14 44 3.03811 $w=3e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.965 $Y=2.635
+ $X2=3.017 $Y2=2.72
r72 14 16 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=2.965 $Y=2.635
+ $X2=2.965 $Y2=2.29
r73 10 31 2.9977 $w=3e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.192 $Y2=2.72
r74 10 12 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.235 $Y2=2.34
r75 3 16 600 $w=1.7e-07 $l=8.882e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=1.485 $X2=2.9 $Y2=2.29
r76 2 38 300 $w=1.7e-07 $l=1.0616e-06 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=1.485 $X2=1.6 $Y2=2.29
r77 1 12 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.3 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_1%Y 1 2 8 10 14 16 18 21 24
r41 21 24 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=1.855 $X2=2.965
+ $Y2=1.855
r42 21 24 1.66364 $w=1.98e-07 $l=3e-08 $layer=LI1_cond $X=2.935 $Y=1.855
+ $X2=2.965 $Y2=1.855
r43 18 20 12.2417 $w=3.18e-07 $l=2.7e-07 $layer=LI1_cond $X=2.975 $Y=0.555
+ $X2=2.975 $Y2=0.825
r44 16 21 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=2.645 $Y=1.855
+ $X2=2.935 $Y2=1.855
r45 12 14 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.44 $Y=2.21
+ $X2=2.56 $Y2=2.21
r46 10 21 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.05 $Y=1.755 $X2=3.05
+ $Y2=1.855
r47 10 20 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.05 $Y=1.755
+ $X2=3.05 $Y2=0.825
r48 8 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=2.125
+ $X2=2.56 $Y2=2.21
r49 7 16 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.56 $Y=1.955
+ $X2=2.645 $Y2=1.855
r50 7 8 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.56 $Y=1.955 $X2=2.56
+ $Y2=2.125
r51 2 12 600 $w=1.7e-07 $l=8.16701e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.44 $Y2=2.21
r52 1 18 182 $w=1.7e-07 $l=3.97995e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.235 $X2=2.96 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_1%VGND 1 2 9 13 16 17 18 24 30 31 34
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r46 31 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r48 28 34 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.07
+ $Y2=0
r49 28 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.99
+ $Y2=0
r50 27 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r51 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r52 24 34 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.07
+ $Y2=0
r53 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=1.61
+ $Y2=0
r54 22 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r55 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r57 16 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.69
+ $Y2=0
r58 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.14
+ $Y2=0
r59 15 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.61
+ $Y2=0
r60 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.14
+ $Y2=0
r61 11 34 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0
r62 11 13 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0.39
r63 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085 $X2=1.14
+ $Y2=0
r64 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.39
r65 2 13 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.08 $Y2=0.39
r66 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_1%A_285_47# 1 2 9 11 12 13
r34 13 15 5.30435 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=2.53 $Y=0.655 $X2=2.53
+ $Y2=0.555
r35 11 13 24.8344 $w=1.96e-07 $l=4.14518e-07 $layer=LI1_cond $X=2.135 $Y=0.82
+ $X2=2.53 $Y2=0.78
r36 11 12 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.135 $Y=0.82
+ $X2=1.725 $Y2=0.82
r37 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.56 $Y=0.735
+ $X2=1.725 $Y2=0.82
r38 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.56 $Y=0.735
+ $X2=1.56 $Y2=0.39
r39 2 15 182 $w=1.7e-07 $l=3.81576e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=2.5 $Y2=0.555
r40 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.425
+ $Y=0.235 $X2=1.56 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__a2bb2oi_2.pxi.spice
* Created: Thu Aug 27 14:03:38 2020
* 
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%B1 N_B1_M1002_g N_B1_M1004_g N_B1_c_84_n
+ N_B1_M1003_g N_B1_M1005_g N_B1_c_85_n N_B1_c_86_n N_B1_c_94_n B1 B1
+ N_B1_c_87_n N_B1_c_88_n N_B1_c_89_n PM_SKY130_FD_SC_HD__A2BB2OI_2%B1
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%B2 N_B2_c_159_n N_B2_M1011_g N_B2_M1007_g
+ N_B2_c_160_n N_B2_M1016_g N_B2_M1008_g B2 N_B2_c_162_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_2%B2
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%A_442_21# N_A_442_21#_M1014_s
+ N_A_442_21#_M1012_d N_A_442_21#_M1010_s N_A_442_21#_c_202_n
+ N_A_442_21#_M1001_g N_A_442_21#_M1000_g N_A_442_21#_c_203_n
+ N_A_442_21#_M1006_g N_A_442_21#_M1015_g N_A_442_21#_c_204_n
+ N_A_442_21#_c_211_n N_A_442_21#_c_220_p N_A_442_21#_c_205_n
+ N_A_442_21#_c_226_p N_A_442_21#_c_279_p N_A_442_21#_c_206_n
+ N_A_442_21#_c_207_n N_A_442_21#_c_208_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_2%A_442_21#
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%A1_N N_A1_N_c_308_n N_A1_N_M1014_g
+ N_A1_N_M1009_g N_A1_N_c_309_n N_A1_N_M1017_g N_A1_N_M1019_g A1_N
+ N_A1_N_c_311_n PM_SKY130_FD_SC_HD__A2BB2OI_2%A1_N
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%A2_N N_A2_N_c_355_n N_A2_N_M1012_g
+ N_A2_N_M1010_g N_A2_N_c_356_n N_A2_N_M1018_g N_A2_N_M1013_g A2_N
+ N_A2_N_c_358_n PM_SKY130_FD_SC_HD__A2BB2OI_2%A2_N
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%A_54_297# N_A_54_297#_M1004_s
+ N_A_54_297#_M1007_s N_A_54_297#_M1005_s N_A_54_297#_M1015_s
+ N_A_54_297#_c_425_p N_A_54_297#_c_399_n N_A_54_297#_c_394_n
+ N_A_54_297#_c_417_p N_A_54_297#_c_403_n N_A_54_297#_c_395_n
+ N_A_54_297#_c_420_p N_A_54_297#_c_412_n N_A_54_297#_c_406_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_2%A_54_297#
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%VPWR N_VPWR_M1004_d N_VPWR_M1008_d
+ N_VPWR_M1009_d N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n
+ VPWR N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_437_n N_VPWR_c_445_n
+ N_VPWR_c_446_n N_VPWR_c_447_n PM_SKY130_FD_SC_HD__A2BB2OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%Y N_Y_M1011_d N_Y_M1001_d N_Y_M1000_d
+ N_Y_c_513_n N_Y_c_522_n N_Y_c_514_n N_Y_c_515_n Y Y Y
+ PM_SKY130_FD_SC_HD__A2BB2OI_2%Y
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%A_662_297# N_A_662_297#_M1009_s
+ N_A_662_297#_M1019_s N_A_662_297#_M1013_d N_A_662_297#_c_567_n
+ N_A_662_297#_c_568_n N_A_662_297#_c_569_n N_A_662_297#_c_591_n
+ N_A_662_297#_c_593_n N_A_662_297#_c_563_n N_A_662_297#_c_564_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_2%A_662_297#
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%VGND N_VGND_M1002_s N_VGND_M1003_s
+ N_VGND_M1006_s N_VGND_M1017_d N_VGND_M1018_s N_VGND_c_597_n N_VGND_c_598_n
+ N_VGND_c_599_n N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n
+ N_VGND_c_604_n N_VGND_c_605_n N_VGND_c_606_n VGND N_VGND_c_607_n
+ N_VGND_c_608_n N_VGND_c_609_n N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_2%VGND
x_PM_SKY130_FD_SC_HD__A2BB2OI_2%A_136_47# N_A_136_47#_M1002_d
+ N_A_136_47#_M1016_s N_A_136_47#_c_681_n N_A_136_47#_c_680_n
+ N_A_136_47#_c_685_n PM_SKY130_FD_SC_HD__A2BB2OI_2%A_136_47#
cc_1 VNB N_B1_c_84_n 0.0162054f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.995
cc_2 VNB N_B1_c_85_n 0.00395886f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_3 VNB N_B1_c_86_n 0.0190084f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_4 VNB N_B1_c_87_n 0.0282041f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_5 VNB N_B1_c_88_n 0.0218917f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_6 VNB N_B1_c_89_n 0.0223869f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.345
cc_7 VNB N_B2_c_159_n 0.0161504f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.995
cc_8 VNB N_B2_c_160_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.995
cc_9 VNB B2 0.00164678f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.445
cc_10 VNB N_B2_c_162_n 0.0308143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_442_21#_c_202_n 0.0159859f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.56
cc_12 VNB N_A_442_21#_c_203_n 0.0187921f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_13 VNB N_A_442_21#_c_204_n 0.00498466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_442_21#_c_205_n 0.00553724f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.325
cc_15 VNB N_A_442_21#_c_206_n 0.00586414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_442_21#_c_207_n 0.0523376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_442_21#_c_208_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_N_c_308_n 0.020695f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.995
cc_19 VNB N_A1_N_c_309_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.995
cc_20 VNB A1_N 0.0092683f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.445
cc_21 VNB N_A1_N_c_311_n 0.0325581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_N_c_355_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.995
cc_23 VNB N_A2_N_c_356_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.995
cc_24 VNB A2_N 0.0312609f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.445
cc_25 VNB N_A2_N_c_358_n 0.0385514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_437_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.345
cc_27 VNB N_Y_c_513_n 0.010208f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.56
cc_28 VNB N_Y_c_514_n 0.00219468f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_29 VNB N_Y_c_515_n 4.05044e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_30 VNB Y 8.57147e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_597_n 0.00650164f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_32 VNB N_VGND_c_598_n 0.00410177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_599_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_600_n 0.00661728f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_35 VNB N_VGND_c_601_n 0.0120081f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=1.16
cc_36 VNB N_VGND_c_602_n 0.00326621f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.53
cc_37 VNB N_VGND_c_603_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.345
cc_38 VNB N_VGND_c_604_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_605_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.345
cc_40 VNB N_VGND_c_606_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0.657 $Y2=1.345
cc_41 VNB N_VGND_c_607_n 0.0359098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_608_n 0.0123263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_609_n 0.28929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_610_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_611_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_612_n 0.0197313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_136_47#_c_680_n 0.00330644f $X=-0.19 $Y=-0.24 $X2=1.865 $Y2=0.56
cc_48 VPB N_B1_M1004_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.985
cc_49 VPB N_B1_M1005_g 0.0172429f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.985
cc_50 VPB N_B1_c_85_n 0.00253424f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_51 VPB N_B1_c_86_n 0.00441099f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_52 VPB N_B1_c_94_n 0.00954818f $X=-0.19 $Y=1.305 $X2=1.7 $Y2=1.53
cc_53 VPB N_B1_c_87_n 0.00483422f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_54 VPB N_B1_c_89_n 0.0233291f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.345
cc_55 VPB N_B2_M1007_g 0.0183442f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.985
cc_56 VPB N_B2_M1008_g 0.0183389f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.985
cc_57 VPB N_B2_c_162_n 0.00405367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_442_21#_M1000_g 0.0187511f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.445
cc_59 VPB N_A_442_21#_M1015_g 0.0213583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_442_21#_c_211_n 0.020341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_442_21#_c_206_n 0.00758654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_442_21#_c_207_n 0.0140332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A1_N_M1009_g 0.0236533f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.985
cc_64 VPB N_A1_N_M1019_g 0.0184042f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.985
cc_65 VPB N_A1_N_c_311_n 0.00426088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A2_N_M1010_g 0.0184042f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.985
cc_67 VPB N_A2_N_M1013_g 0.025194f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.985
cc_68 VPB N_A2_N_c_358_n 0.00479918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_54_297#_c_394_n 0.00692367f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_70 VPB N_A_54_297#_c_395_n 0.00148118f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_71 VPB N_VPWR_c_438_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_439_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.865 $Y2=1.16
cc_73 VPB N_VPWR_c_440_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.7 $Y2=1.53
cc_74 VPB N_VPWR_c_441_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_442_n 0.0485343f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_76 VPB N_VPWR_c_443_n 0.0400401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_437_n 0.0692809f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.345
cc_78 VPB N_VPWR_c_445_n 0.0265498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_446_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_447_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB Y 0.00117056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_662_297#_c_563_n 0.00389675f $X=-0.19 $Y=1.305 $X2=1.7 $Y2=1.53
cc_83 VPB N_A_662_297#_c_564_n 0.00163726f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_84 N_B1_c_88_n N_B2_c_159_n 0.0241679f $X=0.545 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_85 N_B1_M1004_g N_B2_M1007_g 0.0241679f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_86 N_B1_c_94_n N_B2_M1007_g 0.0103235f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_87 N_B1_c_84_n N_B2_c_160_n 0.0269138f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B1_M1005_g N_B2_M1008_g 0.0432836f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B1_c_94_n N_B2_M1008_g 0.0108086f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_90 N_B1_c_85_n B2 0.0134455f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B1_c_86_n B2 2.20976e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B1_c_94_n B2 0.0381541f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_93 N_B1_c_87_n B2 7.56849e-19 $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_c_89_n B2 0.0146287f $X=0.71 $Y=1.345 $X2=0 $Y2=0
cc_95 N_B1_c_85_n N_B2_c_162_n 0.00527477f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B1_c_86_n N_B2_c_162_n 0.022397f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B1_c_94_n N_B2_c_162_n 0.00214031f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_98 N_B1_c_87_n N_B2_c_162_n 0.0241679f $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B1_c_89_n N_B2_c_162_n 0.00505778f $X=0.71 $Y=1.345 $X2=0 $Y2=0
cc_100 N_B1_c_84_n N_A_442_21#_c_202_n 0.0261689f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_M1005_g N_A_442_21#_M1000_g 0.0262864f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_c_94_n N_A_442_21#_M1000_g 0.00148978f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_103 N_B1_c_85_n N_A_442_21#_c_207_n 0.00300327f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B1_c_86_n N_A_442_21#_c_207_n 0.0224305f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B1_c_89_n N_A_54_297#_M1004_s 0.00271859f $X=0.71 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_106 N_B1_c_94_n N_A_54_297#_M1007_s 0.00165831f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_107 N_B1_c_94_n N_A_54_297#_M1005_s 0.00186821f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_108 N_B1_M1004_g N_A_54_297#_c_399_n 0.00956194f $X=0.605 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_B1_c_89_n N_A_54_297#_c_399_n 0.0325821f $X=0.71 $Y=1.345 $X2=0 $Y2=0
cc_110 N_B1_c_87_n N_A_54_297#_c_394_n 3.80105e-19 $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B1_c_89_n N_A_54_297#_c_394_n 0.017911f $X=0.71 $Y=1.345 $X2=0 $Y2=0
cc_112 N_B1_M1005_g N_A_54_297#_c_403_n 0.0095558f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B1_c_86_n N_A_54_297#_c_403_n 2.78509e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_c_94_n N_A_54_297#_c_403_n 0.0357686f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_115 N_B1_c_94_n N_A_54_297#_c_406_n 0.0126919f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_116 N_B1_c_94_n N_VPWR_M1004_d 0.00166235f $X=1.7 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_117 N_B1_c_94_n N_VPWR_M1008_d 0.00165255f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_118 N_B1_M1004_g N_VPWR_c_438_n 0.00302074f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B1_M1005_g N_VPWR_c_440_n 0.00302074f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_M1005_g N_VPWR_c_442_n 0.00585385f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B1_M1004_g N_VPWR_c_437_n 0.00697288f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1005_g N_VPWR_c_437_n 0.00593924f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1004_g N_VPWR_c_445_n 0.00585385f $X=0.605 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_c_84_n N_Y_c_513_n 0.0121351f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B1_c_85_n N_Y_c_513_n 0.0255336f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B1_c_86_n N_Y_c_513_n 0.00296008f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_c_94_n N_Y_c_513_n 0.0071501f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_128 N_B1_c_84_n N_Y_c_522_n 8.6161e-19 $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B1_c_84_n N_Y_c_514_n 3.91234e-19 $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_85_n Y 0.0177855f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B1_c_86_n Y 6.36716e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B1_c_94_n Y 0.00562939f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_133 N_B1_c_87_n N_VGND_c_597_n 0.00176309f $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B1_c_88_n N_VGND_c_597_n 0.00460417f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B1_c_89_n N_VGND_c_597_n 0.0144842f $X=0.71 $Y=1.345 $X2=0 $Y2=0
cc_136 N_B1_c_84_n N_VGND_c_598_n 0.00268723f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_84_n N_VGND_c_607_n 0.00421857f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_88_n N_VGND_c_607_n 0.00539841f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_84_n N_VGND_c_609_n 0.00577981f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_88_n N_VGND_c_609_n 0.0105526f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_c_88_n N_A_136_47#_c_681_n 0.00266812f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_94_n N_A_136_47#_c_680_n 0.00700049f $X=1.7 $Y=1.53 $X2=0 $Y2=0
cc_143 N_B1_c_88_n N_A_136_47#_c_680_n 0.00511819f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B1_c_89_n N_A_136_47#_c_680_n 0.0049108f $X=0.71 $Y=1.345 $X2=0 $Y2=0
cc_145 N_B1_c_84_n N_A_136_47#_c_685_n 0.00302655f $X=1.865 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B2_M1007_g N_A_54_297#_c_399_n 0.00956194f $X=1.025 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_B2_M1008_g N_A_54_297#_c_403_n 0.00956194f $X=1.445 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_B2_M1007_g N_VPWR_c_438_n 0.00157837f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B2_M1007_g N_VPWR_c_439_n 0.00585385f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B2_M1008_g N_VPWR_c_439_n 0.00585385f $X=1.445 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B2_M1008_g N_VPWR_c_440_n 0.00157837f $X=1.445 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B2_M1007_g N_VPWR_c_437_n 0.00591203f $X=1.025 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B2_M1008_g N_VPWR_c_437_n 0.00591203f $X=1.445 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B2_c_160_n N_Y_c_513_n 0.00811447f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_159_n N_Y_c_514_n 0.00381649f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B2_c_160_n N_Y_c_514_n 0.00298551f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_157 B2 N_Y_c_514_n 0.029959f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_158 N_B2_c_162_n N_Y_c_514_n 0.00224214f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B2_c_159_n N_VGND_c_607_n 0.00357877f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_160_n N_VGND_c_607_n 0.00357877f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_159_n N_VGND_c_609_n 0.00525237f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B2_c_160_n N_VGND_c_609_n 0.00525237f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B2_c_159_n N_A_136_47#_c_685_n 0.0105669f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_160_n N_A_136_47#_c_685_n 0.00930415f $X=1.445 $Y=0.995 $X2=0
+ $Y2=0
cc_165 B2 N_A_136_47#_c_685_n 0.00310861f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A_442_21#_c_204_n N_A1_N_c_308_n 0.0108074f $X=3.69 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_442_21#_c_220_p N_A1_N_c_308_n 0.0109565f $X=3.855 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_442_21#_c_206_n N_A1_N_c_308_n 0.00258192f $X=2.915 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_442_21#_c_208_n N_A1_N_c_308_n 0.00113286f $X=3.855 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_170 N_A_442_21#_c_211_n N_A1_N_M1009_g 0.0123532f $X=4.57 $Y=1.53 $X2=0 $Y2=0
cc_171 N_A_442_21#_c_220_p N_A1_N_c_309_n 0.00630972f $X=3.855 $Y=0.39 $X2=0
+ $Y2=0
cc_172 N_A_442_21#_c_205_n N_A1_N_c_309_n 0.00865686f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_173 N_A_442_21#_c_226_p N_A1_N_c_309_n 5.22228e-19 $X=4.695 $Y=0.39 $X2=0
+ $Y2=0
cc_174 N_A_442_21#_c_208_n N_A1_N_c_309_n 0.00113286f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_175 N_A_442_21#_c_211_n N_A1_N_M1019_g 0.0103235f $X=4.57 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A_442_21#_c_204_n A1_N 0.0281469f $X=3.69 $Y=0.815 $X2=0 $Y2=0
cc_177 N_A_442_21#_c_211_n A1_N 0.0649161f $X=4.57 $Y=1.53 $X2=0 $Y2=0
cc_178 N_A_442_21#_c_205_n A1_N 0.0132155f $X=4.53 $Y=0.815 $X2=0 $Y2=0
cc_179 N_A_442_21#_c_206_n A1_N 0.0161058f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_442_21#_c_207_n A1_N 8.32501e-19 $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_442_21#_c_208_n A1_N 0.0265405f $X=3.855 $Y=0.815 $X2=0 $Y2=0
cc_182 N_A_442_21#_c_211_n N_A1_N_c_311_n 0.00214031f $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_A_442_21#_c_206_n N_A1_N_c_311_n 0.00322402f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_442_21#_c_207_n N_A1_N_c_311_n 0.0068545f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_442_21#_c_208_n N_A1_N_c_311_n 0.00230339f $X=3.855 $Y=0.815 $X2=0
+ $Y2=0
cc_186 N_A_442_21#_c_220_p N_A2_N_c_355_n 5.22228e-19 $X=3.855 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_442_21#_c_205_n N_A2_N_c_355_n 0.0103016f $X=4.53 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_442_21#_c_226_p N_A2_N_c_355_n 0.00630972f $X=4.695 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_442_21#_c_211_n N_A2_N_M1010_g 0.0137782f $X=4.57 $Y=1.53 $X2=0 $Y2=0
cc_190 N_A_442_21#_c_205_n N_A2_N_c_356_n 0.00262807f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_191 N_A_442_21#_c_226_p N_A2_N_c_356_n 0.00539651f $X=4.695 $Y=0.39 $X2=0
+ $Y2=0
cc_192 N_A_442_21#_c_211_n N_A2_N_M1013_g 5.91109e-19 $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_193 N_A_442_21#_c_211_n A2_N 0.0282825f $X=4.57 $Y=1.53 $X2=0 $Y2=0
cc_194 N_A_442_21#_c_205_n A2_N 0.0316767f $X=4.53 $Y=0.815 $X2=0 $Y2=0
cc_195 N_A_442_21#_c_211_n N_A2_N_c_358_n 0.00222344f $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_442_21#_c_205_n N_A2_N_c_358_n 0.00230339f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_197 N_A_442_21#_c_206_n N_A_54_297#_M1015_s 0.00296633f $X=2.915 $Y=1.16
+ $X2=0 $Y2=0
cc_198 N_A_442_21#_M1000_g N_A_54_297#_c_395_n 0.0121306f $X=2.285 $Y=1.985
+ $X2=0 $Y2=0
cc_199 N_A_442_21#_M1015_g N_A_54_297#_c_395_n 0.0116622f $X=2.705 $Y=1.985
+ $X2=0 $Y2=0
cc_200 N_A_442_21#_c_206_n N_A_54_297#_c_412_n 0.0120421f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_201 N_A_442_21#_c_207_n N_A_54_297#_c_412_n 0.00115158f $X=2.915 $Y=1.16
+ $X2=0 $Y2=0
cc_202 N_A_442_21#_c_211_n N_VPWR_M1009_d 0.00166235f $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_203 N_A_442_21#_M1000_g N_VPWR_c_442_n 0.00357877f $X=2.285 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_442_21#_M1015_g N_VPWR_c_442_n 0.00357877f $X=2.705 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_442_21#_M1010_s N_VPWR_c_437_n 0.00216833f $X=4.56 $Y=1.485 $X2=0
+ $Y2=0
cc_206 N_A_442_21#_M1000_g N_VPWR_c_437_n 0.00525237f $X=2.285 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_442_21#_M1015_g N_VPWR_c_437_n 0.00655123f $X=2.705 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_442_21#_c_202_n N_Y_c_513_n 0.0123222f $X=2.285 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_442_21#_c_202_n N_Y_c_522_n 0.00648728f $X=2.285 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_442_21#_c_203_n N_Y_c_522_n 0.0109565f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_442_21#_c_202_n N_Y_c_515_n 0.00221107f $X=2.285 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_442_21#_c_203_n N_Y_c_515_n 0.00276569f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_442_21#_c_206_n N_Y_c_515_n 0.010445f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_442_21#_c_202_n Y 0.00247781f $X=2.285 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_442_21#_M1000_g Y 0.00172567f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_442_21#_c_203_n Y 0.00208168f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_442_21#_M1015_g Y 0.00416037f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_442_21#_c_206_n Y 0.0447359f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_442_21#_c_207_n Y 0.0223265f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_442_21#_M1015_g Y 0.0041886f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_442_21#_c_211_n N_A_662_297#_M1009_s 0.00272914f $X=4.57 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_222 N_A_442_21#_c_211_n N_A_662_297#_M1019_s 0.00165831f $X=4.57 $Y=1.53
+ $X2=0 $Y2=0
cc_223 N_A_442_21#_c_211_n N_A_662_297#_c_567_n 0.0317352f $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_442_21#_c_211_n N_A_662_297#_c_568_n 0.0126919f $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_442_21#_M1010_s N_A_662_297#_c_569_n 0.00312348f $X=4.56 $Y=1.485
+ $X2=0 $Y2=0
cc_226 N_A_442_21#_c_279_p N_A_662_297#_c_569_n 0.0118865f $X=4.695 $Y=1.62
+ $X2=0 $Y2=0
cc_227 N_A_442_21#_c_211_n N_A_662_297#_c_563_n 0.00251363f $X=4.57 $Y=1.53
+ $X2=0 $Y2=0
cc_228 N_A_442_21#_c_211_n N_A_662_297#_c_564_n 0.0165158f $X=4.57 $Y=1.53 $X2=0
+ $Y2=0
cc_229 N_A_442_21#_c_204_n N_VGND_M1006_s 0.00591147f $X=3.69 $Y=0.815 $X2=0
+ $Y2=0
cc_230 N_A_442_21#_c_206_n N_VGND_M1006_s 0.00441866f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_442_21#_c_205_n N_VGND_M1017_d 0.00162089f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_232 N_A_442_21#_c_202_n N_VGND_c_598_n 0.00146339f $X=2.285 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_442_21#_c_205_n N_VGND_c_599_n 0.0122559f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_234 N_A_442_21#_c_205_n N_VGND_c_600_n 0.00830019f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_235 N_A_442_21#_c_204_n N_VGND_c_603_n 0.00198695f $X=3.69 $Y=0.815 $X2=0
+ $Y2=0
cc_236 N_A_442_21#_c_220_p N_VGND_c_603_n 0.0188551f $X=3.855 $Y=0.39 $X2=0
+ $Y2=0
cc_237 N_A_442_21#_c_205_n N_VGND_c_603_n 0.00198695f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_238 N_A_442_21#_c_205_n N_VGND_c_605_n 0.00198695f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_239 N_A_442_21#_c_226_p N_VGND_c_605_n 0.0188551f $X=4.695 $Y=0.39 $X2=0
+ $Y2=0
cc_240 N_A_442_21#_M1014_s N_VGND_c_609_n 0.00215201f $X=3.72 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_442_21#_M1012_d N_VGND_c_609_n 0.00215201f $X=4.56 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_442_21#_c_202_n N_VGND_c_609_n 0.0057435f $X=2.285 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_442_21#_c_203_n N_VGND_c_609_n 0.0108251f $X=2.705 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_442_21#_c_204_n N_VGND_c_609_n 0.00537187f $X=3.69 $Y=0.815 $X2=0
+ $Y2=0
cc_245 N_A_442_21#_c_220_p N_VGND_c_609_n 0.0122069f $X=3.855 $Y=0.39 $X2=0
+ $Y2=0
cc_246 N_A_442_21#_c_205_n N_VGND_c_609_n 0.00835832f $X=4.53 $Y=0.815 $X2=0
+ $Y2=0
cc_247 N_A_442_21#_c_226_p N_VGND_c_609_n 0.0122069f $X=4.695 $Y=0.39 $X2=0
+ $Y2=0
cc_248 N_A_442_21#_c_206_n N_VGND_c_609_n 7.36513e-19 $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_249 N_A_442_21#_c_202_n N_VGND_c_611_n 0.00423334f $X=2.285 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_442_21#_c_203_n N_VGND_c_611_n 0.00541359f $X=2.705 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_442_21#_c_203_n N_VGND_c_612_n 0.00335921f $X=2.705 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_442_21#_c_204_n N_VGND_c_612_n 0.030682f $X=3.69 $Y=0.815 $X2=0 $Y2=0
cc_253 N_A_442_21#_c_206_n N_VGND_c_612_n 0.0192004f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_254 N_A_442_21#_c_207_n N_VGND_c_612_n 0.00134655f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A1_N_c_309_n N_A2_N_c_355_n 0.023995f $X=4.065 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A1_N_M1019_g N_A2_N_M1010_g 0.023995f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_257 A1_N A2_N 0.0132033f $X=3.845 $Y=1.105 $X2=0 $Y2=0
cc_258 N_A1_N_c_311_n A2_N 2.10007e-19 $X=4.065 $Y=1.16 $X2=0 $Y2=0
cc_259 A1_N N_A2_N_c_358_n 0.00161184f $X=3.845 $Y=1.105 $X2=0 $Y2=0
cc_260 N_A1_N_c_311_n N_A2_N_c_358_n 0.023995f $X=4.065 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_N_M1009_g N_VPWR_c_441_n 0.00302074f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A1_N_M1019_g N_VPWR_c_441_n 0.00302074f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_N_M1009_g N_VPWR_c_442_n 0.00441875f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A1_N_M1019_g N_VPWR_c_443_n 0.00441875f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A1_N_M1009_g N_VPWR_c_437_n 0.00718625f $X=3.645 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A1_N_M1019_g N_VPWR_c_437_n 0.00588739f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A1_N_M1009_g N_A_662_297#_c_567_n 0.0104429f $X=3.645 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A1_N_M1019_g N_A_662_297#_c_567_n 0.0104429f $X=4.065 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A1_N_c_309_n N_VGND_c_599_n 0.00146339f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A1_N_c_308_n N_VGND_c_603_n 0.00423334f $X=3.645 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_N_c_309_n N_VGND_c_603_n 0.00423334f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_N_c_308_n N_VGND_c_609_n 0.0070399f $X=3.645 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_N_c_309_n N_VGND_c_609_n 0.0057435f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_N_c_308_n N_VGND_c_612_n 0.00335921f $X=3.645 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_N_M1010_g N_VPWR_c_443_n 0.00357877f $X=4.485 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A2_N_M1013_g N_VPWR_c_443_n 0.00357877f $X=4.905 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A2_N_M1010_g N_VPWR_c_437_n 0.00525237f $X=4.485 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A2_N_M1013_g N_VPWR_c_437_n 0.00629231f $X=4.905 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A2_N_M1010_g N_A_662_297#_c_569_n 0.0121306f $X=4.485 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A2_N_M1013_g N_A_662_297#_c_569_n 0.0121306f $X=4.905 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A2_N_M1013_g N_A_662_297#_c_563_n 7.0041e-19 $X=4.905 $Y=1.985 $X2=0
+ $Y2=0
cc_282 A2_N N_A_662_297#_c_563_n 0.0203393f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_283 N_A2_N_c_355_n N_VGND_c_599_n 0.00146448f $X=4.485 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A2_N_c_356_n N_VGND_c_600_n 0.00360182f $X=4.905 $Y=0.995 $X2=0 $Y2=0
cc_285 A2_N N_VGND_c_600_n 0.0143482f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_286 N_A2_N_c_355_n N_VGND_c_605_n 0.00423334f $X=4.485 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A2_N_c_356_n N_VGND_c_605_n 0.00541359f $X=4.905 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A2_N_c_355_n N_VGND_c_609_n 0.0057435f $X=4.485 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A2_N_c_356_n N_VGND_c_609_n 0.0105687f $X=4.905 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A_54_297#_c_399_n N_VPWR_M1004_d 0.00332635f $X=1.11 $Y=1.87 $X2=-0.19
+ $Y2=1.305
cc_291 N_A_54_297#_c_403_n N_VPWR_M1008_d 0.0032936f $X=1.95 $Y=1.87 $X2=0 $Y2=0
cc_292 N_A_54_297#_c_399_n N_VPWR_c_438_n 0.0117423f $X=1.11 $Y=1.87 $X2=0 $Y2=0
cc_293 N_A_54_297#_c_417_p N_VPWR_c_439_n 0.0142343f $X=1.235 $Y=1.96 $X2=0
+ $Y2=0
cc_294 N_A_54_297#_c_403_n N_VPWR_c_440_n 0.0117423f $X=1.95 $Y=1.87 $X2=0 $Y2=0
cc_295 N_A_54_297#_c_395_n N_VPWR_c_442_n 0.0489446f $X=2.79 $Y=2.38 $X2=0 $Y2=0
cc_296 N_A_54_297#_c_420_p N_VPWR_c_442_n 0.0143053f $X=2.2 $Y=2.38 $X2=0 $Y2=0
cc_297 N_A_54_297#_M1004_s N_VPWR_c_437_n 0.00212725f $X=0.27 $Y=1.485 $X2=0
+ $Y2=0
cc_298 N_A_54_297#_M1007_s N_VPWR_c_437_n 0.00223619f $X=1.1 $Y=1.485 $X2=0
+ $Y2=0
cc_299 N_A_54_297#_M1005_s N_VPWR_c_437_n 0.00220214f $X=1.94 $Y=1.485 $X2=0
+ $Y2=0
cc_300 N_A_54_297#_M1015_s N_VPWR_c_437_n 0.0020932f $X=2.78 $Y=1.485 $X2=0
+ $Y2=0
cc_301 N_A_54_297#_c_425_p N_VPWR_c_437_n 0.00955092f $X=0.395 $Y=1.96 $X2=0
+ $Y2=0
cc_302 N_A_54_297#_c_399_n N_VPWR_c_437_n 0.0109496f $X=1.11 $Y=1.87 $X2=0 $Y2=0
cc_303 N_A_54_297#_c_417_p N_VPWR_c_437_n 0.00955092f $X=1.235 $Y=1.96 $X2=0
+ $Y2=0
cc_304 N_A_54_297#_c_403_n N_VPWR_c_437_n 0.0109496f $X=1.95 $Y=1.87 $X2=0 $Y2=0
cc_305 N_A_54_297#_c_395_n N_VPWR_c_437_n 0.0300869f $X=2.79 $Y=2.38 $X2=0 $Y2=0
cc_306 N_A_54_297#_c_420_p N_VPWR_c_437_n 0.00962794f $X=2.2 $Y=2.38 $X2=0 $Y2=0
cc_307 N_A_54_297#_c_425_p N_VPWR_c_445_n 0.0158369f $X=0.395 $Y=1.96 $X2=0
+ $Y2=0
cc_308 N_A_54_297#_c_395_n N_Y_M1000_d 0.00312348f $X=2.79 $Y=2.38 $X2=0 $Y2=0
cc_309 N_A_54_297#_c_395_n Y 0.0118865f $X=2.79 $Y=2.38 $X2=0 $Y2=0
cc_310 N_A_54_297#_c_395_n Y 7.22078e-19 $X=2.79 $Y=2.38 $X2=0 $Y2=0
cc_311 N_A_54_297#_c_395_n N_A_662_297#_c_564_n 0.0100846f $X=2.79 $Y=2.38 $X2=0
+ $Y2=0
cc_312 N_A_54_297#_c_412_n N_A_662_297#_c_564_n 0.0280952f $X=2.915 $Y=1.96
+ $X2=0 $Y2=0
cc_313 N_VPWR_c_437_n N_Y_M1000_d 0.00216833f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_437_n N_A_662_297#_M1009_s 0.0021259f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_315 N_VPWR_c_437_n N_A_662_297#_M1019_s 0.00220079f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_437_n N_A_662_297#_M1013_d 0.00295147f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_M1009_d N_A_662_297#_c_567_n 0.00317395f $X=3.72 $Y=1.485 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_441_n N_A_662_297#_c_567_n 0.0123469f $X=3.855 $Y=2.3 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_442_n N_A_662_297#_c_567_n 0.0020229f $X=3.73 $Y=2.72 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_443_n N_A_662_297#_c_567_n 0.0020229f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_437_n N_A_662_297#_c_567_n 0.00802398f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_443_n N_A_662_297#_c_569_n 0.0330174f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_437_n N_A_662_297#_c_569_n 0.0204627f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_443_n N_A_662_297#_c_591_n 0.0143053f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_437_n N_A_662_297#_c_591_n 0.00962794f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_443_n N_A_662_297#_c_593_n 0.0159079f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_437_n N_A_662_297#_c_593_n 0.00961749f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_442_n N_A_662_297#_c_564_n 0.0158369f $X=3.73 $Y=2.72 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_437_n N_A_662_297#_c_564_n 0.00955092f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_330 N_Y_c_513_n N_VGND_M1003_s 0.00162089f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_331 N_Y_c_513_n N_VGND_c_598_n 0.0122559f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_332 N_Y_c_513_n N_VGND_c_607_n 0.00199263f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_333 N_Y_M1011_d N_VGND_c_609_n 0.00216833f $X=1.1 $Y=0.235 $X2=0 $Y2=0
cc_334 N_Y_M1001_d N_VGND_c_609_n 0.00215201f $X=2.36 $Y=0.235 $X2=0 $Y2=0
cc_335 N_Y_c_513_n N_VGND_c_609_n 0.00930722f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_336 N_Y_c_522_n N_VGND_c_609_n 0.01222f $X=2.495 $Y=0.39 $X2=0 $Y2=0
cc_337 N_Y_c_513_n N_VGND_c_611_n 0.00198695f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_338 N_Y_c_522_n N_VGND_c_611_n 0.0188977f $X=2.495 $Y=0.39 $X2=0 $Y2=0
cc_339 N_Y_c_513_n N_A_136_47#_M1016_s 0.00191752f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_340 N_Y_c_514_n N_A_136_47#_c_680_n 0.0105027f $X=1.4 $Y=0.775 $X2=0 $Y2=0
cc_341 N_Y_M1011_d N_A_136_47#_c_685_n 0.00305026f $X=1.1 $Y=0.235 $X2=0 $Y2=0
cc_342 N_Y_c_513_n N_A_136_47#_c_685_n 0.014941f $X=2.33 $Y=0.815 $X2=0 $Y2=0
cc_343 N_Y_c_514_n N_A_136_47#_c_685_n 0.0153374f $X=1.4 $Y=0.775 $X2=0 $Y2=0
cc_344 N_VGND_c_609_n N_A_136_47#_M1002_d 0.00215206f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_345 N_VGND_c_609_n N_A_136_47#_M1016_s 0.00215227f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_607_n N_A_136_47#_c_681_n 0.0151965f $X=1.99 $Y=0 $X2=0 $Y2=0
cc_347 N_VGND_c_609_n N_A_136_47#_c_681_n 0.00940324f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_597_n N_A_136_47#_c_680_n 0.0154056f $X=0.395 $Y=0.39 $X2=0
+ $Y2=0
cc_349 N_VGND_c_607_n N_A_136_47#_c_685_n 0.0504977f $X=1.99 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_609_n N_A_136_47#_c_685_n 0.0327385f $X=5.29 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__or4_1.pex.spice
* Created: Tue Sep  1 19:28:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4_1%D 3 7 9 10 17
c28 9 0 1.84467e-19 $X=0.235 $Y=0.85
r29 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r31 9 10 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.265 $Y=0.85
+ $X2=0.265 $Y2=1.16
r32 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r34 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%C 3 7 9 11 18
r37 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=1.325
r38 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r39 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r40 11 19 5.11227 $w=6.18e-07 $l=2.65e-07 $layer=LI1_cond $X=1.155 $Y=1.305
+ $X2=0.89 $Y2=1.305
r41 9 19 3.76186 $w=6.18e-07 $l=1.95e-07 $layer=LI1_cond $X=0.695 $Y=1.305
+ $X2=0.89 $Y2=1.305
r42 7 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.95 $Y=1.695
+ $X2=0.95 $Y2=1.325
r43 3 20 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.95 $Y=0.475
+ $X2=0.95 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%B 4 5 7 8 9 10 15 16
c35 15 0 1.73735e-19 $X=1.37 $Y=2.28
r36 15 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.37 $Y=2.28
+ $X2=1.37 $Y2=2.145
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=2.28 $X2=1.37 $Y2=2.28
r38 10 16 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.155 $Y=2.27
+ $X2=1.37 $Y2=2.27
r39 9 10 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=2.27
+ $X2=1.155 $Y2=2.27
r40 8 9 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=2.27
+ $X2=0.695 $Y2=2.27
r41 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.37 $Y=0.76 $X2=1.37
+ $Y2=0.475
r42 4 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.31 $Y=1.695
+ $X2=1.31 $Y2=2.145
r43 1 5 34.5933 $w=2.09e-07 $l=1.77482e-07 $layer=POLY_cond $X=1.31 $Y=0.91
+ $X2=1.37 $Y2=0.76
r44 1 4 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.31 $Y=0.91 $X2=1.31
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%A 3 7 9 12 13
r42 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.16
+ $X2=1.77 $Y2=1.325
r43 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.16
+ $X2=1.77 $Y2=0.995
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r45 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.77 $Y2=1.16
r46 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.79 $Y=1.695
+ $X2=1.79 $Y2=1.325
r47 3 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.79 $Y=0.475
+ $X2=1.79 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%A_27_297# 1 2 3 12 15 17 21 23 24 27 29 31 36
+ 38 42 43 48 49 50 53
c99 48 0 1.1436e-19 $X=2.25 $Y=1.16
c100 43 0 1.73735e-19 $X=1.595 $Y=1.58
c101 36 0 1.06604e-19 $X=2.15 $Y=1.495
r102 49 54 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.252 $Y=1.16
+ $X2=2.252 $Y2=1.325
r103 49 53 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.252 $Y=1.16
+ $X2=2.252 $Y2=0.995
r104 48 51 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.2 $Y=1.16
+ $X2=2.2 $Y2=1.325
r105 48 50 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.2 $Y=1.16
+ $X2=2.2 $Y2=0.995
r106 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r107 43 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.595 $Y=1.58
+ $X2=1.595 $Y2=1.87
r108 38 40 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=0.25 $Y=1.685
+ $X2=0.25 $Y2=1.87
r109 36 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=1.495
+ $X2=2.15 $Y2=1.325
r110 33 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=0.825
+ $X2=2.15 $Y2=0.995
r111 32 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.58
+ $X2=1.595 $Y2=1.58
r112 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=1.58
+ $X2=2.15 $Y2=1.495
r113 31 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=1.58
+ $X2=1.68 $Y2=1.58
r114 30 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.74
+ $X2=1.58 $Y2=0.74
r115 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=0.74
+ $X2=2.15 $Y2=0.825
r116 29 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.065 $Y=0.74
+ $X2=1.665 $Y2=0.74
r117 25 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.655
+ $X2=1.58 $Y2=0.74
r118 25 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.58 $Y=0.655
+ $X2=1.58 $Y2=0.47
r119 23 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=0.74
+ $X2=1.58 $Y2=0.74
r120 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.495 $Y=0.74
+ $X2=0.795 $Y2=0.74
r121 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=0.655
+ $X2=0.795 $Y2=0.74
r122 19 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.71 $Y=0.655
+ $X2=0.71 $Y2=0.47
r123 18 40 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.41 $Y=1.87
+ $X2=0.25 $Y2=1.87
r124 17 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=1.87
+ $X2=1.595 $Y2=1.87
r125 17 18 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=1.51 $Y=1.87
+ $X2=0.41 $Y2=1.87
r126 15 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.28 $Y=1.985
+ $X2=2.28 $Y2=1.325
r127 12 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.28 $Y=0.56
+ $X2=2.28 $Y2=0.995
r128 3 38 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.685
r129 2 27 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.265 $X2=1.58 $Y2=0.47
r130 1 21 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=0.71 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%VPWR 1 6 8 10 20 21 24
c26 1 0 1.06604e-19 $X=1.865 $Y=1.485
r27 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r28 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r30 18 24 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.055 $Y2=2.72
r31 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.53 $Y2=2.72
r32 17 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r33 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 12 16 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r35 10 24 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.055 $Y2=2.72
r36 10 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 8 17 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r38 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r39 4 24 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.72
r40 4 6 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2
r41 1 6 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.485 $X2=2.065 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%X 1 2 12 14 15 16
r18 14 16 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.54 $Y=1.63
+ $X2=2.54 $Y2=1.845
r19 14 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.54 $Y=1.63
+ $X2=2.54 $Y2=1.495
r20 10 12 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=2.49 $Y=0.587 $X2=2.59
+ $Y2=0.587
r21 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.59 $Y=0.76 $X2=2.59
+ $Y2=0.587
r22 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.59 $Y=0.76
+ $X2=2.59 $Y2=1.495
r23 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=1.485 $X2=2.49 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.49 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_1%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
c53 24 0 1.84467e-19 $X=0.995 $Y=0
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r55 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r56 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r57 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r58 34 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.025
+ $Y2=0
r59 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.53
+ $Y2=0
r60 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r61 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r63 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.16
+ $Y2=0
r64 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.61
+ $Y2=0
r65 29 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.025
+ $Y2=0
r66 29 32 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.61
+ $Y2=0
r67 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 25 40 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r70 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r71 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.16
+ $Y2=0
r72 24 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.69
+ $Y2=0
r73 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r74 22 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 18 46 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r76 18 20 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.4
r77 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0
r78 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0.4
r79 10 40 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r80 10 12 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.5
r81 3 20 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.265 $X2=2.05 $Y2=0.4
r82 2 16 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.265 $X2=1.16 $Y2=0.4
r83 1 12 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_684_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=3.575e+11p pd=2.4e+06u as=9.3275e+11p ps=9.37e+06u
M1001 a_115_297# C1 a_28_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.8e+11p pd=2.56e+06u as=8.65e+11p ps=7.73e+06u
M1002 a_287_297# D1 Y VPB phighvt w=1e+06u l=150000u
+  ad=2.8e+11p pd=2.56e+06u as=2.8e+11p ps=2.56e+06u
M1003 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=9.1325e+11p pd=8.01e+06u as=0p ps=0u
M1004 a_923_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1005 a_28_297# B1 a_467_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.155e+12p ps=1.031e+07u
M1006 a_467_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1007 Y D1 a_115_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_467_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_467_297# B1 a_28_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_467_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_28_297# C1 a_287_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_923_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_467_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y D1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND C1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_684_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

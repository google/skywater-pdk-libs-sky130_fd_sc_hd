* File: sky130_fd_sc_hd__a21boi_2.spice.SKY130_FD_SC_HD__A21BOI_2.pxi
* Created: Thu Aug 27 14:00:40 2020
* 
x_PM_SKY130_FD_SC_HD__A21BOI_2%B1_N N_B1_N_M1011_g N_B1_N_c_72_n N_B1_N_M1001_g
+ N_B1_N_c_73_n N_B1_N_c_74_n B1_N N_B1_N_c_76_n
+ PM_SKY130_FD_SC_HD__A21BOI_2%B1_N
x_PM_SKY130_FD_SC_HD__A21BOI_2%A_61_47# N_A_61_47#_M1001_s N_A_61_47#_M1011_d
+ N_A_61_47#_M1007_g N_A_61_47#_M1009_g N_A_61_47#_M1008_g N_A_61_47#_M1012_g
+ N_A_61_47#_c_107_n N_A_61_47#_c_108_n N_A_61_47#_c_109_n N_A_61_47#_c_110_n
+ N_A_61_47#_c_111_n N_A_61_47#_c_112_n N_A_61_47#_c_113_n
+ PM_SKY130_FD_SC_HD__A21BOI_2%A_61_47#
x_PM_SKY130_FD_SC_HD__A21BOI_2%A2 N_A2_M1002_g N_A2_M1004_g N_A2_M1013_g
+ N_A2_M1006_g N_A2_c_175_n N_A2_c_195_p N_A2_c_189_n N_A2_c_176_n N_A2_c_177_n
+ N_A2_c_178_n N_A2_c_179_n A2 N_A2_c_180_n N_A2_c_215_p
+ PM_SKY130_FD_SC_HD__A21BOI_2%A2
x_PM_SKY130_FD_SC_HD__A21BOI_2%A1 N_A1_c_256_n N_A1_M1003_g N_A1_M1000_g
+ N_A1_c_257_n N_A1_M1010_g N_A1_M1005_g A1 N_A1_c_259_n
+ PM_SKY130_FD_SC_HD__A21BOI_2%A1
x_PM_SKY130_FD_SC_HD__A21BOI_2%VPWR N_VPWR_M1011_s N_VPWR_M1002_s N_VPWR_M1005_d
+ N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n VPWR N_VPWR_c_313_n
+ N_VPWR_c_304_n PM_SKY130_FD_SC_HD__A21BOI_2%VPWR
x_PM_SKY130_FD_SC_HD__A21BOI_2%A_217_297# N_A_217_297#_M1009_d
+ N_A_217_297#_M1012_d N_A_217_297#_M1000_s N_A_217_297#_M1006_d
+ N_A_217_297#_c_368_n N_A_217_297#_c_378_n N_A_217_297#_c_369_n
+ N_A_217_297#_c_380_n N_A_217_297#_c_381_n N_A_217_297#_c_391_n
+ N_A_217_297#_c_418_n N_A_217_297#_c_394_n N_A_217_297#_c_370_n
+ N_A_217_297#_c_371_n N_A_217_297#_c_399_n
+ PM_SKY130_FD_SC_HD__A21BOI_2%A_217_297#
x_PM_SKY130_FD_SC_HD__A21BOI_2%Y N_Y_M1007_s N_Y_M1003_d N_Y_M1009_s N_Y_c_429_n
+ N_Y_c_438_n N_Y_c_446_n Y N_Y_c_461_p PM_SKY130_FD_SC_HD__A21BOI_2%Y
x_PM_SKY130_FD_SC_HD__A21BOI_2%VGND N_VGND_M1001_d N_VGND_M1008_d N_VGND_M1013_s
+ N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ N_VGND_c_475_n VGND N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ N_VGND_c_479_n VGND PM_SKY130_FD_SC_HD__A21BOI_2%VGND
cc_1 VNB N_B1_N_c_72_n 0.0194328f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.73
cc_2 VNB N_B1_N_c_73_n 0.0365526f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.805
cc_3 VNB N_B1_N_c_74_n 0.00530181f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=1.435
cc_4 VNB B1_N 0.0209655f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB N_B1_N_c_76_n 0.0337732f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=0.93
cc_6 VNB N_A_61_47#_M1007_g 0.0198506f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.88
cc_7 VNB N_A_61_47#_M1008_g 0.0177296f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.93
cc_8 VNB N_A_61_47#_c_107_n 0.0280357f $X=-0.19 $Y=-0.24 $X2=0.272 $Y2=0.93
cc_9 VNB N_A_61_47#_c_108_n 0.0250418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_61_47#_c_109_n 0.00749754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_61_47#_c_110_n 0.007816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_61_47#_c_111_n 4.45758e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_61_47#_c_112_n 0.00959726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_61_47#_c_113_n 0.00539172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_M1013_g 0.0239203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_175_n 8.46397e-19 $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.93
cc_17 VNB N_A2_c_176_n 0.00305053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_177_n 0.0192728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_178_n 0.00477698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_179_n 0.0333701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_180_n 0.0161891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_256_n 0.0157491f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.435
cc_23 VNB N_A1_c_257_n 0.0164438f $X=-0.19 $Y=-0.24 $X2=0.362 $Y2=0.805
cc_24 VNB A1 0.00456205f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_25 VNB N_A1_c_259_n 0.0309298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_304_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_429_n 0.00237487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_470_n 0.00664415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_471_n 0.0028319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_472_n 0.0145739f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=0.93
cc_31 VNB N_VGND_c_473_n 0.0303186f $X=-0.19 $Y=-0.24 $X2=0.272 $Y2=0.85
cc_32 VNB N_VGND_c_474_n 0.0294278f $X=-0.19 $Y=-0.24 $X2=0.272 $Y2=0.93
cc_33 VNB N_VGND_c_475_n 0.00461634f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_476_n 0.0198011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_477_n 0.0368771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_478_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_479_n 0.226369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_B1_N_M1011_g 0.044859f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.1
cc_39 VPB N_B1_N_c_74_n 0.0183419f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=1.435
cc_40 VPB B1_N 0.0222924f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_41 VPB N_A_61_47#_M1009_g 0.0241214f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=1.248
cc_42 VPB N_A_61_47#_M1012_g 0.0197171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_61_47#_c_107_n 0.0114994f $X=-0.19 $Y=1.305 $X2=0.272 $Y2=0.93
cc_44 VPB N_A_61_47#_c_108_n 0.00257374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_61_47#_c_111_n 0.0192563f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A2_M1002_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.1
cc_47 VPB N_A2_M1006_g 0.023393f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=1.435
cc_48 VPB N_A2_c_175_n 0.00325856f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=0.93
cc_49 VPB N_A2_c_177_n 0.00439782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A2_c_179_n 0.00546669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB A2 0.00839328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A1_M1000_g 0.0189179f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.445
cc_53 VPB N_A1_M1005_g 0.0187884f $X=-0.19 $Y=1.305 $X2=0.362 $Y2=1.248
cc_54 VPB A1 2.41965e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_55 VPB N_A1_c_259_n 0.00485795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_305_n 0.0115529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_306_n 0.0229399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_307_n 0.00407289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_308_n 4.11703e-19 $X=-0.19 $Y=1.305 $X2=0.272 $Y2=0.85
cc_60 VPB N_VPWR_c_309_n 0.0486053f $X=-0.19 $Y=1.305 $X2=0.272 $Y2=0.93
cc_61 VPB N_VPWR_c_310_n 0.00323844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_311_n 0.0147069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_312_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_313_n 0.0185595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_304_n 0.0634951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_217_297#_c_368_n 0.00487566f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_67 VPB N_A_217_297#_c_369_n 0.00283306f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=0.93
cc_68 VPB N_A_217_297#_c_370_n 0.0111305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_217_297#_c_371_n 0.0133845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_Y_c_429_n 0.00307168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_B1_N_c_72_n N_A_61_47#_M1007_g 0.0105934f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_72 N_B1_N_c_76_n N_A_61_47#_c_107_n 0.00630257f $X=0.34 $Y=0.93 $X2=0 $Y2=0
cc_73 N_B1_N_c_72_n N_A_61_47#_c_109_n 0.00598674f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_74 N_B1_N_c_73_n N_A_61_47#_c_109_n 0.00991152f $X=0.68 $Y=0.805 $X2=0 $Y2=0
cc_75 B1_N N_A_61_47#_c_109_n 0.00907806f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_76 N_B1_N_c_72_n N_A_61_47#_c_110_n 0.00593834f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_77 N_B1_N_c_73_n N_A_61_47#_c_110_n 0.0109216f $X=0.68 $Y=0.805 $X2=0 $Y2=0
cc_78 B1_N N_A_61_47#_c_110_n 0.0225548f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_79 N_B1_N_c_76_n N_A_61_47#_c_110_n 0.0041871f $X=0.34 $Y=0.93 $X2=0 $Y2=0
cc_80 N_B1_N_c_74_n N_A_61_47#_c_111_n 0.0158088f $X=0.362 $Y=1.435 $X2=0 $Y2=0
cc_81 B1_N N_A_61_47#_c_111_n 0.0400682f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_82 B1_N N_A_61_47#_c_113_n 0.0179944f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_83 N_B1_N_c_76_n N_A_61_47#_c_113_n 0.00253063f $X=0.34 $Y=0.93 $X2=0 $Y2=0
cc_84 N_B1_N_M1011_g N_VPWR_c_306_n 0.00925967f $X=0.475 $Y=2.1 $X2=0 $Y2=0
cc_85 N_B1_N_c_74_n N_VPWR_c_306_n 7.38883e-19 $X=0.362 $Y=1.435 $X2=0 $Y2=0
cc_86 B1_N N_VPWR_c_306_n 0.017703f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_87 N_B1_N_M1011_g N_VPWR_c_309_n 0.00455951f $X=0.475 $Y=2.1 $X2=0 $Y2=0
cc_88 N_B1_N_M1011_g N_VPWR_c_304_n 0.00445127f $X=0.475 $Y=2.1 $X2=0 $Y2=0
cc_89 N_B1_N_M1011_g N_A_217_297#_c_369_n 0.00257038f $X=0.475 $Y=2.1 $X2=0
+ $Y2=0
cc_90 N_B1_N_c_72_n N_VGND_c_470_n 0.00706879f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_91 N_B1_N_c_72_n N_VGND_c_474_n 0.0037867f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_92 N_B1_N_c_73_n N_VGND_c_474_n 0.00216138f $X=0.68 $Y=0.805 $X2=0 $Y2=0
cc_93 N_B1_N_c_72_n N_VGND_c_479_n 0.00713327f $X=0.68 $Y=0.73 $X2=0 $Y2=0
cc_94 N_B1_N_c_73_n N_VGND_c_479_n 0.00244058f $X=0.68 $Y=0.805 $X2=0 $Y2=0
cc_95 B1_N N_VGND_c_479_n 0.00603494f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_96 N_A_61_47#_M1012_g N_A2_M1002_g 0.0289349f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_61_47#_c_108_n N_A2_c_175_n 0.00206837f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_61_47#_M1012_g N_A2_c_189_n 0.0016751f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_61_47#_c_108_n N_A2_c_176_n 0.00148742f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_61_47#_M1008_g N_A2_c_177_n 0.0219204f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_101 N_A_61_47#_M1008_g N_A2_c_180_n 0.0218396f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_102 N_A_61_47#_M1009_g N_VPWR_c_309_n 0.0035787f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_61_47#_M1012_g N_VPWR_c_309_n 0.00357835f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_61_47#_c_111_n N_VPWR_c_309_n 0.00769913f $X=0.69 $Y=2.1 $X2=0 $Y2=0
cc_105 N_A_61_47#_M1009_g N_VPWR_c_304_n 0.00651492f $X=1.42 $Y=1.985 $X2=0
+ $Y2=0
cc_106 N_A_61_47#_M1012_g N_VPWR_c_304_n 0.00525234f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_107 N_A_61_47#_c_111_n N_VPWR_c_304_n 0.00882494f $X=0.69 $Y=2.1 $X2=0 $Y2=0
cc_108 N_A_61_47#_M1009_g N_A_217_297#_c_368_n 0.00550958f $X=1.42 $Y=1.985
+ $X2=0 $Y2=0
cc_109 N_A_61_47#_M1012_g N_A_217_297#_c_368_n 5.06027e-19 $X=1.84 $Y=1.985
+ $X2=0 $Y2=0
cc_110 N_A_61_47#_c_107_n N_A_217_297#_c_368_n 0.00527333f $X=1.345 $Y=1.16
+ $X2=0 $Y2=0
cc_111 N_A_61_47#_c_111_n N_A_217_297#_c_368_n 0.0353352f $X=0.69 $Y=2.1 $X2=0
+ $Y2=0
cc_112 N_A_61_47#_c_112_n N_A_217_297#_c_368_n 0.00886392f $X=1.16 $Y=1.16 $X2=0
+ $Y2=0
cc_113 N_A_61_47#_M1009_g N_A_217_297#_c_378_n 0.0121251f $X=1.42 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_61_47#_M1012_g N_A_217_297#_c_378_n 0.0111176f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_61_47#_M1012_g N_A_217_297#_c_380_n 0.00326762f $X=1.84 $Y=1.985
+ $X2=0 $Y2=0
cc_116 N_A_61_47#_M1009_g N_A_217_297#_c_381_n 4.65488e-19 $X=1.42 $Y=1.985
+ $X2=0 $Y2=0
cc_117 N_A_61_47#_M1012_g N_A_217_297#_c_381_n 0.00393929f $X=1.84 $Y=1.985
+ $X2=0 $Y2=0
cc_118 N_A_61_47#_M1007_g N_Y_c_429_n 0.00326511f $X=1.42 $Y=0.56 $X2=0 $Y2=0
cc_119 N_A_61_47#_M1009_g N_Y_c_429_n 0.0024934f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_61_47#_M1008_g N_Y_c_429_n 0.00316294f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_121 N_A_61_47#_M1012_g N_Y_c_429_n 0.00180214f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_61_47#_c_108_n N_Y_c_429_n 0.0199207f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_61_47#_c_111_n N_Y_c_429_n 0.0106768f $X=0.69 $Y=2.1 $X2=0 $Y2=0
cc_124 N_A_61_47#_c_112_n N_Y_c_429_n 0.0146666f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_61_47#_M1008_g N_Y_c_438_n 0.014506f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_126 N_A_61_47#_M1007_g N_VGND_c_470_n 0.0103765f $X=1.42 $Y=0.56 $X2=0 $Y2=0
cc_127 N_A_61_47#_c_107_n N_VGND_c_470_n 0.00551959f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_128 N_A_61_47#_c_110_n N_VGND_c_470_n 0.0206723f $X=0.695 $Y=1.07 $X2=0 $Y2=0
cc_129 N_A_61_47#_c_112_n N_VGND_c_470_n 0.0179109f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_61_47#_M1008_g N_VGND_c_471_n 0.00311401f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A_61_47#_c_109_n N_VGND_c_474_n 0.0188939f $X=0.595 $Y=0.445 $X2=0
+ $Y2=0
cc_132 N_A_61_47#_M1007_g N_VGND_c_476_n 0.00585385f $X=1.42 $Y=0.56 $X2=0 $Y2=0
cc_133 N_A_61_47#_M1008_g N_VGND_c_476_n 0.00422112f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_61_47#_M1001_s N_VGND_c_479_n 0.00255915f $X=0.305 $Y=0.235 $X2=0
+ $Y2=0
cc_135 N_A_61_47#_M1007_g N_VGND_c_479_n 0.0113871f $X=1.42 $Y=0.56 $X2=0 $Y2=0
cc_136 N_A_61_47#_M1008_g N_VGND_c_479_n 0.00572598f $X=1.84 $Y=0.56 $X2=0 $Y2=0
cc_137 N_A_61_47#_c_109_n N_VGND_c_479_n 0.0180144f $X=0.595 $Y=0.445 $X2=0
+ $Y2=0
cc_138 N_A2_c_180_n N_A1_c_256_n 0.0387062f $X=2.26 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_139 N_A2_M1002_g N_A1_M1000_g 0.045988f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A2_c_195_p N_A1_M1000_g 0.0108315f $X=3.385 $Y=1.585 $X2=0 $Y2=0
cc_141 N_A2_M1013_g N_A1_c_257_n 0.0393965f $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A2_M1006_g N_A1_M1005_g 0.0438039f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A2_c_195_p N_A1_M1005_g 0.0108951f $X=3.385 $Y=1.585 $X2=0 $Y2=0
cc_144 A2 N_A1_M1005_g 0.00374086f $X=3.39 $Y=1.445 $X2=0 $Y2=0
cc_145 N_A2_M1013_g A1 2.56397e-19 $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_146 N_A2_c_195_p A1 0.0392259f $X=3.385 $Y=1.585 $X2=0 $Y2=0
cc_147 N_A2_c_176_n A1 0.0197969f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_177_n A1 8.4532e-19 $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A2_c_178_n A1 0.0243499f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_179_n A1 3.16097e-19 $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_M1013_g N_A1_c_259_n 0.0171648f $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A2_c_175_n N_A1_c_259_n 0.00392425f $X=2.262 $Y=1.495 $X2=0 $Y2=0
cc_153 N_A2_c_195_p N_A1_c_259_n 0.00224497f $X=3.385 $Y=1.585 $X2=0 $Y2=0
cc_154 N_A2_c_176_n N_A1_c_259_n 8.25011e-19 $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_177_n N_A1_c_259_n 0.0387062f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_c_178_n N_A1_c_259_n 0.00101093f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_195_p N_VPWR_M1002_s 0.00602119f $X=3.385 $Y=1.585 $X2=0 $Y2=0
cc_158 N_A2_c_189_n N_VPWR_M1002_s 3.62273e-19 $X=2.425 $Y=1.585 $X2=0 $Y2=0
cc_159 N_A2_c_195_p N_VPWR_M1005_d 0.00700827f $X=3.385 $Y=1.585 $X2=0 $Y2=0
cc_160 N_A2_c_215_p N_VPWR_M1005_d 2.49555e-19 $X=3.53 $Y=1.495 $X2=0 $Y2=0
cc_161 N_A2_M1002_g N_VPWR_c_307_n 0.00268723f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A2_M1006_g N_VPWR_c_308_n 0.00785369f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_M1002_g N_VPWR_c_309_n 0.00418507f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_M1006_g N_VPWR_c_313_n 0.00351072f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A2_M1002_g N_VPWR_c_304_n 0.00572068f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A2_M1006_g N_VPWR_c_304_n 0.00510436f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A2_c_189_n N_A_217_297#_M1012_d 0.00252765f $X=2.425 $Y=1.585 $X2=0
+ $Y2=0
cc_168 N_A2_c_195_p N_A_217_297#_M1000_s 0.0033536f $X=3.385 $Y=1.585 $X2=0
+ $Y2=0
cc_169 A2 N_A_217_297#_M1006_d 3.66298e-19 $X=3.39 $Y=1.445 $X2=0 $Y2=0
cc_170 N_A2_c_215_p N_A_217_297#_M1006_d 0.00811989f $X=3.53 $Y=1.495 $X2=0
+ $Y2=0
cc_171 N_A2_M1002_g N_A_217_297#_c_378_n 0.00213389f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A2_M1002_g N_A_217_297#_c_380_n 8.93985e-19 $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A2_c_189_n N_A_217_297#_c_380_n 0.00467621f $X=2.425 $Y=1.585 $X2=0
+ $Y2=0
cc_174 N_A2_M1002_g N_A_217_297#_c_381_n 0.00409646f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A2_M1002_g N_A_217_297#_c_391_n 0.00837828f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A2_c_195_p N_A_217_297#_c_391_n 0.0182861f $X=3.385 $Y=1.585 $X2=0
+ $Y2=0
cc_177 N_A2_c_189_n N_A_217_297#_c_391_n 0.0111097f $X=2.425 $Y=1.585 $X2=0
+ $Y2=0
cc_178 N_A2_M1006_g N_A_217_297#_c_394_n 0.0115953f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_c_195_p N_A_217_297#_c_394_n 0.0202748f $X=3.385 $Y=1.585 $X2=0
+ $Y2=0
cc_180 N_A2_c_215_p N_A_217_297#_c_394_n 0.0129085f $X=3.53 $Y=1.495 $X2=0 $Y2=0
cc_181 N_A2_c_178_n N_A_217_297#_c_370_n 0.0037819f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A2_c_179_n N_A_217_297#_c_370_n 0.00212987f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A2_c_195_p N_A_217_297#_c_399_n 0.0128761f $X=3.385 $Y=1.585 $X2=0
+ $Y2=0
cc_184 N_A2_c_175_n N_Y_c_429_n 0.0107889f $X=2.262 $Y=1.495 $X2=0 $Y2=0
cc_185 N_A2_c_176_n N_Y_c_429_n 0.00712779f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_c_177_n N_Y_c_429_n 4.91324e-19 $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A2_M1013_g N_Y_c_438_n 5.07806e-19 $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A2_c_176_n N_Y_c_438_n 0.0146866f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_c_177_n N_Y_c_438_n 0.00275815f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A2_c_180_n N_Y_c_438_n 0.0119595f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_M1013_g N_Y_c_446_n 0.00107868f $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A2_c_180_n N_Y_c_446_n 0.00136667f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_180_n N_VGND_c_471_n 0.0084534f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_M1013_g N_VGND_c_473_n 0.00479037f $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A2_c_178_n N_VGND_c_473_n 0.0114864f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A2_c_179_n N_VGND_c_473_n 0.00360399f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A2_M1013_g N_VGND_c_477_n 0.00585385f $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A2_c_180_n N_VGND_c_477_n 0.00351072f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_M1013_g N_VGND_c_479_n 0.011649f $X=3.54 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A2_c_180_n N_VGND_c_479_n 0.00395482f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_M1000_g N_VPWR_c_307_n 0.00139158f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A1_M1000_g N_VPWR_c_308_n 5.31014e-19 $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A1_M1005_g N_VPWR_c_308_n 0.00643202f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A1_M1000_g N_VPWR_c_311_n 0.00433717f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A1_M1005_g N_VPWR_c_311_n 0.00351072f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A1_M1000_g N_VPWR_c_304_n 0.00586678f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A1_M1005_g N_VPWR_c_304_n 0.0040731f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A1_M1000_g N_A_217_297#_c_381_n 4.78112e-19 $X=2.68 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A1_M1000_g N_A_217_297#_c_391_n 0.0100175f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A1_M1005_g N_A_217_297#_c_394_n 0.0116015f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A1_c_256_n N_Y_c_438_n 0.00887945f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A1_c_257_n N_Y_c_438_n 0.0034662f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_213 A1 N_Y_c_438_n 0.0257864f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_214 N_A1_c_259_n N_Y_c_438_n 0.0022587f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A1_c_256_n N_Y_c_446_n 0.00614363f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A1_c_257_n N_Y_c_446_n 0.00671932f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A1_c_256_n N_VGND_c_471_n 0.00173186f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A1_c_256_n N_VGND_c_477_n 0.0041289f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A1_c_257_n N_VGND_c_477_n 0.0054895f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A1_c_256_n N_VGND_c_479_n 0.00557866f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A1_c_257_n N_VGND_c_479_n 0.00996518f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_222 N_VPWR_c_304_n N_A_217_297#_M1009_d 0.00209319f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_223 N_VPWR_c_304_n N_A_217_297#_M1012_d 0.00215201f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_304_n N_A_217_297#_M1000_s 0.00264218f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_304_n N_A_217_297#_M1006_d 0.00243803f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_306_n N_A_217_297#_c_368_n 5.73423e-19 $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_309_n N_A_217_297#_c_378_n 0.04918f $X=2.385 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_304_n N_A_217_297#_c_378_n 0.030992f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_306_n N_A_217_297#_c_369_n 0.00580963f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_309_n N_A_217_297#_c_369_n 0.0194546f $X=2.385 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_304_n N_A_217_297#_c_369_n 0.0116462f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_M1002_s N_A_217_297#_c_391_n 0.00326959f $X=2.335 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_307_n N_A_217_297#_c_391_n 0.012114f $X=2.47 $Y=2.36 $X2=0 $Y2=0
cc_234 N_VPWR_c_309_n N_A_217_297#_c_391_n 0.00211912f $X=2.385 $Y=2.72 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_311_n N_A_217_297#_c_391_n 0.00300834f $X=3.16 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_304_n N_A_217_297#_c_391_n 0.0106736f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_311_n N_A_217_297#_c_418_n 0.0116518f $X=3.16 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_304_n N_A_217_297#_c_418_n 0.00644138f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_239 N_VPWR_M1005_d N_A_217_297#_c_394_n 0.00353311f $X=3.185 $Y=1.485 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_308_n N_A_217_297#_c_394_n 0.0163189f $X=3.325 $Y=2.36 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_311_n N_A_217_297#_c_394_n 0.0027458f $X=3.16 $Y=2.72 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_313_n N_A_217_297#_c_394_n 0.00264265f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_304_n N_A_217_297#_c_394_n 0.0104634f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_313_n N_A_217_297#_c_371_n 0.0175789f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_304_n N_A_217_297#_c_371_n 0.00989761f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_304_n N_Y_M1009_s 0.00216833f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_247 N_A_217_297#_c_378_n N_Y_M1009_s 0.00312899f $X=1.885 $Y=2.375 $X2=0
+ $Y2=0
cc_248 N_A_217_297#_c_378_n N_Y_c_429_n 0.0119608f $X=1.885 $Y=2.375 $X2=0 $Y2=0
cc_249 N_Y_c_438_n N_VGND_M1008_d 0.00798906f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_250 N_Y_c_438_n N_VGND_c_471_n 0.0180367f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_251 N_Y_c_446_n N_VGND_c_471_n 0.0063569f $X=2.895 $Y=0.36 $X2=0 $Y2=0
cc_252 N_Y_c_438_n N_VGND_c_476_n 0.00327755f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_253 N_Y_c_461_p N_VGND_c_476_n 0.0124602f $X=1.63 $Y=0.42 $X2=0 $Y2=0
cc_254 N_Y_c_438_n N_VGND_c_477_n 0.00720366f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_255 N_Y_c_446_n N_VGND_c_477_n 0.0186595f $X=2.895 $Y=0.36 $X2=0 $Y2=0
cc_256 N_Y_M1007_s N_VGND_c_479_n 0.00315979f $X=1.495 $Y=0.235 $X2=0 $Y2=0
cc_257 N_Y_M1003_d N_VGND_c_479_n 0.00223231f $X=2.755 $Y=0.235 $X2=0 $Y2=0
cc_258 N_Y_c_438_n N_VGND_c_479_n 0.0189959f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_259 N_Y_c_446_n N_VGND_c_479_n 0.0121874f $X=2.895 $Y=0.36 $X2=0 $Y2=0
cc_260 N_Y_c_461_p N_VGND_c_479_n 0.00762533f $X=1.63 $Y=0.42 $X2=0 $Y2=0
cc_261 N_Y_c_438_n A_637_47# 0.00529826f $X=2.73 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_262 N_VGND_c_479_n A_637_47# 0.00239227f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_263 N_VGND_c_479_n A_479_47# 0.0119688f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o2111a_2.pxi.spice
* Created: Thu Aug 27 14:33:52 2020
* 
x_PM_SKY130_FD_SC_HD__O2111A_2%A_80_21# N_A_80_21#_M1008_s N_A_80_21#_M1010_d
+ N_A_80_21#_M1011_d N_A_80_21#_c_69_n N_A_80_21#_M1002_g N_A_80_21#_M1003_g
+ N_A_80_21#_c_70_n N_A_80_21#_M1007_g N_A_80_21#_M1012_g N_A_80_21#_c_71_n
+ N_A_80_21#_c_72_n N_A_80_21#_c_80_p N_A_80_21#_c_108_p N_A_80_21#_c_73_n
+ N_A_80_21#_c_74_n N_A_80_21#_c_94_p N_A_80_21#_c_102_p N_A_80_21#_c_116_p
+ N_A_80_21#_c_92_p PM_SKY130_FD_SC_HD__O2111A_2%A_80_21#
x_PM_SKY130_FD_SC_HD__O2111A_2%D1 N_D1_M1010_g N_D1_c_153_n N_D1_M1008_g D1 D1
+ N_D1_c_154_n PM_SKY130_FD_SC_HD__O2111A_2%D1
x_PM_SKY130_FD_SC_HD__O2111A_2%C1 N_C1_M1009_g N_C1_M1004_g C1 C1 C1 C1
+ N_C1_c_189_n PM_SKY130_FD_SC_HD__O2111A_2%C1
x_PM_SKY130_FD_SC_HD__O2111A_2%B1 N_B1_M1013_g N_B1_M1011_g B1 B1 N_B1_c_228_n
+ N_B1_c_229_n PM_SKY130_FD_SC_HD__O2111A_2%B1
x_PM_SKY130_FD_SC_HD__O2111A_2%A2 N_A2_M1001_g N_A2_M1000_g A2 A2 N_A2_c_262_n
+ N_A2_c_263_n PM_SKY130_FD_SC_HD__O2111A_2%A2
x_PM_SKY130_FD_SC_HD__O2111A_2%A1 N_A1_M1005_g N_A1_M1006_g A1 A1 A1 A1 A1
+ N_A1_c_298_n N_A1_c_299_n PM_SKY130_FD_SC_HD__O2111A_2%A1
x_PM_SKY130_FD_SC_HD__O2111A_2%VPWR N_VPWR_M1003_s N_VPWR_M1012_s N_VPWR_M1004_d
+ N_VPWR_M1006_d N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n
+ VPWR N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_327_n
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ PM_SKY130_FD_SC_HD__O2111A_2%VPWR
x_PM_SKY130_FD_SC_HD__O2111A_2%X N_X_M1002_d N_X_M1003_d X X N_X_c_395_n
+ PM_SKY130_FD_SC_HD__O2111A_2%X
x_PM_SKY130_FD_SC_HD__O2111A_2%VGND N_VGND_M1002_s N_VGND_M1007_s N_VGND_M1001_d
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n VGND
+ N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n
+ N_VGND_c_419_n PM_SKY130_FD_SC_HD__O2111A_2%VGND
x_PM_SKY130_FD_SC_HD__O2111A_2%A_566_47# N_A_566_47#_M1013_d N_A_566_47#_M1005_d
+ N_A_566_47#_c_473_n N_A_566_47#_c_485_n N_A_566_47#_c_471_n
+ N_A_566_47#_c_472_n PM_SKY130_FD_SC_HD__O2111A_2%A_566_47#
cc_1 VNB N_A_80_21#_c_69_n 0.0216086f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_70_n 0.0187937f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_A_80_21#_c_71_n 0.00459132f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_4 VNB N_A_80_21#_c_72_n 0.060617f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_5 VNB N_A_80_21#_c_73_n 0.0114657f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=0.715
cc_6 VNB N_A_80_21#_c_74_n 0.00523362f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=0.4
cc_7 VNB N_D1_c_153_n 0.019464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_D1_c_154_n 0.0314801f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_9 VNB N_C1_M1009_g 0.0168825f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=1.485
cc_10 VNB N_C1_M1004_g 3.90643e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB C1 0.00498807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_C1_c_189_n 0.0288168f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_13 VNB N_B1_M1013_g 0.0203773f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=1.485
cc_14 VNB N_B1_M1011_g 5.03674e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_228_n 0.0274126f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_16 VNB N_B1_c_229_n 0.00240549f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_17 VNB N_A2_M1001_g 0.0202587f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=1.485
cc_18 VNB N_A2_M1000_g 5.0126e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_262_n 0.0269774f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_20 VNB N_A2_c_263_n 0.00459415f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_21 VNB N_A1_M1005_g 0.0254934f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=1.485
cc_22 VNB N_A1_M1006_g 6.03208e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB A1 0.00635747f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_24 VNB N_A1_c_298_n 0.0427048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A1_c_299_n 0.021869f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=0.4
cc_26 VNB N_VPWR_c_327_n 0.193827f $X=-0.19 $Y=-0.24 $X2=3.03 $Y2=1.905
cc_27 VNB N_VGND_c_410_n 0.0105432f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_28 VNB N_VGND_c_411_n 0.00832841f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_29 VNB N_VGND_c_412_n 0.00840898f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_413_n 0.0055721f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.325
cc_31 VNB N_VGND_c_414_n 0.0184335f $X=-0.19 $Y=-0.24 $X2=1.167 $Y2=0.885
cc_32 VNB N_VGND_c_415_n 0.0550968f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.905
cc_33 VNB N_VGND_c_416_n 0.0263171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_417_n 0.254071f $X=-0.19 $Y=-0.24 $X2=2.865 $Y2=1.905
cc_35 VNB N_VGND_c_418_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=1.167 $Y2=0.8
cc_36 VNB N_VGND_c_419_n 0.00631048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_566_47#_c_471_n 0.00868775f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_38 VNB N_A_566_47#_c_472_n 0.0145675f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_39 VPB N_A_80_21#_M1003_g 0.0254232f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_40 VPB N_A_80_21#_M1012_g 0.0213167f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_41 VPB N_A_80_21#_c_71_n 0.00222257f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_42 VPB N_A_80_21#_c_72_n 0.0148772f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_43 VPB N_D1_M1010_g 0.0234078f $X=-0.19 $Y=1.305 $X2=2.83 $Y2=1.485
cc_44 VPB D1 0.00123631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_D1_c_154_n 0.00969103f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.995
cc_46 VPB N_C1_M1004_g 0.0195539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB C1 0.00248074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_B1_M1011_g 0.0218129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_B1_c_229_n 0.00127318f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_50 VPB N_A2_M1000_g 0.0226165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB A2 0.00263639f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_52 VPB N_A1_M1006_g 0.024639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB A1 0.0084504f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_54 VPB A1 0.0535117f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_55 VPB N_A1_c_299_n 4.11258e-19 $X=-0.19 $Y=1.305 $X2=1.64 $Y2=0.4
cc_56 VPB N_VPWR_c_328_n 0.0105174f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_57 VPB N_VPWR_c_329_n 0.00491148f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_58 VPB N_VPWR_c_330_n 0.00508539f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_59 VPB N_VPWR_c_331_n 0.00242814f $X=-0.19 $Y=1.305 $X2=1.167 $Y2=1.785
cc_60 VPB N_VPWR_c_332_n 0.0170865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_333_n 0.0318455f $X=-0.19 $Y=1.305 $X2=3.03 $Y2=2.34
cc_62 VPB N_VPWR_c_334_n 0.0152287f $X=-0.19 $Y=1.305 $X2=2 $Y2=1.885
cc_63 VPB N_VPWR_c_327_n 0.0519817f $X=-0.19 $Y=1.305 $X2=3.03 $Y2=1.905
cc_64 VPB N_VPWR_c_336_n 0.0184335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_337_n 0.0186467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_338_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_339_n 0.00366581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_71_n N_D1_M1010_g 0.00612424f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_80_p N_D1_M1010_g 0.0155096f $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_71_n N_D1_c_153_n 0.00287068f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_73_n N_D1_c_153_n 0.00227746f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_74_n N_D1_c_153_n 0.00516798f $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_71_n D1 0.0381098f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_72_n D1 2.86216e-19 $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_80_p D1 0.0215177f $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_73_n D1 0.0191618f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_71_n N_D1_c_154_n 0.00338293f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_72_n N_D1_c_154_n 0.0165322f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_80_p N_D1_c_154_n 7.01654e-19 $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_73_n N_D1_c_154_n 0.006842f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_92_p N_D1_c_154_n 0.00147666f $X=2 $Y=1.885 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_74_n N_C1_M1009_g 3.79543e-19 $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_94_p N_C1_M1004_g 0.0126428f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_84 N_A_80_21#_M1010_d C1 0.00195891f $X=1.86 $Y=1.485 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_73_n C1 0.012343f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_74_n C1 0.0318881f $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_94_p C1 0.0151667f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_92_p C1 0.00694246f $X=2 $Y=1.885 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_94_p N_C1_c_189_n 0.00249106f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_94_p N_B1_M1011_g 0.0159183f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_102_p N_B1_c_228_n 5.42007e-19 $X=3.03 $Y=2.025 $X2=0 $Y2=0
cc_92 N_A_80_21#_M1011_d N_B1_c_229_n 0.00429706f $X=2.83 $Y=1.485 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_94_p N_B1_c_229_n 0.0114099f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_102_p N_B1_c_229_n 0.0187931f $X=3.03 $Y=2.025 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_71_n N_VPWR_M1012_s 0.00794621f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_80_p N_VPWR_M1012_s 0.0159237f $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_108_p N_VPWR_M1012_s 0.00643789f $X=1.305 $Y=1.905 $X2=0
+ $Y2=0
cc_98 N_A_80_21#_c_94_p N_VPWR_M1004_d 0.0114464f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_99 N_A_80_21#_M1003_g N_VPWR_c_329_n 0.00440648f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_100 N_A_80_21#_c_94_p N_VPWR_c_330_n 0.0167329f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_80_p N_VPWR_c_332_n 0.00263766f $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_94_p N_VPWR_c_332_n 0.00247019f $X=2.865 $Y=1.905 $X2=0
+ $Y2=0
cc_103 N_A_80_21#_c_92_p N_VPWR_c_332_n 0.0156471f $X=2 $Y=1.885 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_94_p N_VPWR_c_333_n 0.00267952f $X=2.865 $Y=1.905 $X2=0
+ $Y2=0
cc_105 N_A_80_21#_c_116_p N_VPWR_c_333_n 0.0212535f $X=3.03 $Y=2.34 $X2=0 $Y2=0
cc_106 N_A_80_21#_M1010_d N_VPWR_c_327_n 0.00223231f $X=1.86 $Y=1.485 $X2=0
+ $Y2=0
cc_107 N_A_80_21#_M1011_d N_VPWR_c_327_n 0.00414189f $X=2.83 $Y=1.485 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_M1003_g N_VPWR_c_327_n 0.0103145f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_80_21#_M1012_g N_VPWR_c_327_n 0.011049f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_80_p N_VPWR_c_327_n 0.00623018f $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_108_p N_VPWR_c_327_n 0.00134226f $X=1.305 $Y=1.905 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_94_p N_VPWR_c_327_n 0.010802f $X=2.865 $Y=1.905 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_116_p N_VPWR_c_327_n 0.0126319f $X=3.03 $Y=2.34 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_92_p N_VPWR_c_327_n 0.0107063f $X=2 $Y=1.885 $X2=0 $Y2=0
cc_115 N_A_80_21#_M1003_g N_VPWR_c_336_n 0.00533769f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_80_21#_M1012_g N_VPWR_c_336_n 0.0054895f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_80_21#_M1012_g N_VPWR_c_337_n 0.00474014f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_80_21#_c_80_p N_VPWR_c_337_n 0.0274617f $X=1.86 $Y=1.905 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_108_p N_VPWR_c_337_n 0.022829f $X=1.305 $Y=1.905 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_69_n N_X_c_395_n 0.0135526f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_80_21#_M1003_g N_X_c_395_n 0.0206663f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_70_n N_X_c_395_n 0.0112796f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_80_21#_M1012_g N_X_c_395_n 0.0199933f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_71_n N_X_c_395_n 0.0554624f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_72_n N_X_c_395_n 0.0336136f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_74_n N_X_c_395_n 0.00505984f $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_71_n N_VGND_M1007_s 6.15036e-19 $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_73_n N_VGND_M1007_s 0.00378915f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_69_n N_VGND_c_411_n 0.00440648f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_130 N_A_80_21#_c_70_n N_VGND_c_412_n 0.00445597f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_73_n N_VGND_c_412_n 0.0193994f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_74_n N_VGND_c_412_n 0.0218711f $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_69_n N_VGND_c_414_n 0.00533769f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_70_n N_VGND_c_414_n 0.0054895f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_73_n N_VGND_c_415_n 0.0029735f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_74_n N_VGND_c_415_n 0.0205167f $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_137 N_A_80_21#_M1008_s N_VGND_c_417_n 0.00213418f $X=1.515 $Y=0.235 $X2=0
+ $Y2=0
cc_138 N_A_80_21#_c_69_n N_VGND_c_417_n 0.0103145f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_70_n N_VGND_c_417_n 0.0110515f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_73_n N_VGND_c_417_n 0.0062377f $X=1.64 $Y=0.715 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_74_n N_VGND_c_417_n 0.012325f $X=1.64 $Y=0.4 $X2=0 $Y2=0
cc_142 N_D1_c_153_n N_C1_M1009_g 0.0370577f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_143 N_D1_M1010_g N_C1_M1004_g 0.0229227f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_144 N_D1_M1010_g C1 0.0018211f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_145 N_D1_c_153_n C1 0.011208f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_146 D1 C1 0.0430216f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_147 D1 N_C1_c_189_n 4.92684e-19 $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_148 N_D1_c_154_n N_C1_c_189_n 0.0370577f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_149 D1 N_VPWR_M1012_s 0.00311713f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_150 N_D1_M1010_g N_VPWR_c_332_n 0.00433717f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_151 N_D1_M1010_g N_VPWR_c_327_n 0.00720106f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_152 N_D1_M1010_g N_VPWR_c_337_n 0.00330957f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_153 N_D1_c_153_n N_VGND_c_412_n 0.0022787f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_154 N_D1_c_153_n N_VGND_c_415_n 0.00547957f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_155 N_D1_c_153_n N_VGND_c_417_n 0.0110306f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C1_M1009_g N_B1_M1013_g 0.0254245f $X=2.215 $Y=0.56 $X2=0 $Y2=0
cc_157 C1 N_B1_M1013_g 0.00941529f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_158 N_C1_M1004_g N_B1_M1011_g 0.0335645f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_159 C1 N_B1_M1011_g 0.0022325f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_160 C1 N_B1_c_228_n 9.74588e-19 $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_161 N_C1_c_189_n N_B1_c_228_n 0.0170303f $X=2.305 $Y=1.16 $X2=0 $Y2=0
cc_162 N_C1_M1004_g N_B1_c_229_n 3.55776e-19 $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_163 C1 N_B1_c_229_n 0.028394f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_164 N_C1_c_189_n N_B1_c_229_n 8.12321e-19 $X=2.305 $Y=1.16 $X2=0 $Y2=0
cc_165 C1 N_VPWR_M1004_d 0.0019216f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_166 N_C1_M1004_g N_VPWR_c_330_n 0.00312737f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_167 N_C1_M1004_g N_VPWR_c_332_n 0.00433717f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_168 N_C1_M1004_g N_VPWR_c_327_n 0.00617618f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_169 N_C1_M1009_g N_VGND_c_415_n 0.00357668f $X=2.215 $Y=0.56 $X2=0 $Y2=0
cc_170 C1 N_VGND_c_415_n 0.02264f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_171 N_C1_M1009_g N_VGND_c_417_n 0.00543451f $X=2.215 $Y=0.56 $X2=0 $Y2=0
cc_172 C1 N_VGND_c_417_n 0.014064f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_173 C1 A_386_47# 0.00634429f $X=2.01 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_174 C1 A_458_47# 0.0091978f $X=2.01 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_175 N_B1_M1013_g N_A2_M1001_g 0.0170445f $X=2.755 $Y=0.56 $X2=0 $Y2=0
cc_176 N_B1_M1011_g N_A2_M1000_g 0.0254852f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B1_c_229_n A2 0.0135103f $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B1_c_228_n N_A2_c_262_n 0.0170867f $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B1_c_229_n N_A2_c_262_n 0.00450063f $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_c_228_n N_A2_c_263_n 5.01675e-19 $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B1_c_229_n N_A2_c_263_n 0.0179368f $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B1_M1011_g N_VPWR_c_330_n 0.0032033f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_M1011_g N_VPWR_c_333_n 0.00433717f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1011_g N_VPWR_c_327_n 0.00639348f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1013_g N_VGND_c_415_n 0.00585385f $X=2.755 $Y=0.56 $X2=0 $Y2=0
cc_186 N_B1_M1013_g N_VGND_c_417_n 0.011422f $X=2.755 $Y=0.56 $X2=0 $Y2=0
cc_187 N_B1_c_228_n N_A_566_47#_c_473_n 0.00319079f $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B1_c_229_n N_A_566_47#_c_473_n 0.0143964f $X=2.845 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_M1001_g N_A1_M1005_g 0.0229607f $X=3.295 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A2_c_263_n N_A1_M1005_g 0.00634783f $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A2_M1000_g N_A1_M1006_g 0.0308697f $X=3.295 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A2_c_262_n A1 2.41756e-19 $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A2_c_263_n A1 0.0259442f $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A2_c_263_n A1 0.00551179f $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_195 A2 N_A1_c_298_n 0.00634783f $X=3.39 $Y=2.125 $X2=0 $Y2=0
cc_196 N_A2_c_262_n N_A1_c_298_n 0.0171254f $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A2_M1000_g N_VPWR_c_331_n 0.00163679f $X=3.295 $Y=1.985 $X2=0 $Y2=0
cc_198 A2 N_VPWR_c_331_n 0.0532034f $X=3.39 $Y=2.125 $X2=0 $Y2=0
cc_199 N_A2_M1000_g N_VPWR_c_333_n 0.00585385f $X=3.295 $Y=1.985 $X2=0 $Y2=0
cc_200 A2 N_VPWR_c_333_n 0.0113688f $X=3.39 $Y=2.125 $X2=0 $Y2=0
cc_201 N_A2_M1000_g N_VPWR_c_327_n 0.0113348f $X=3.295 $Y=1.985 $X2=0 $Y2=0
cc_202 A2 N_VPWR_c_327_n 0.0105388f $X=3.39 $Y=2.125 $X2=0 $Y2=0
cc_203 A2 A_674_297# 0.0222666f $X=3.39 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_204 N_A2_M1001_g N_VGND_c_413_n 0.00326685f $X=3.295 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A2_M1001_g N_VGND_c_415_n 0.0042361f $X=3.295 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A2_M1001_g N_VGND_c_417_n 0.00614444f $X=3.295 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A2_M1001_g N_A_566_47#_c_471_n 0.0136754f $X=3.295 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A2_c_262_n N_A_566_47#_c_471_n 0.00106184f $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A2_c_263_n N_A_566_47#_c_471_n 0.0271666f $X=3.385 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A2_M1001_g N_A_566_47#_c_472_n 5.62833e-19 $X=3.295 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A1_M1006_g N_VPWR_c_331_n 0.0183966f $X=3.835 $Y=1.985 $X2=0 $Y2=0
cc_212 A1 N_VPWR_c_331_n 0.0182846f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_213 A1 N_VPWR_c_331_n 0.0664998f $X=4.31 $Y=1.445 $X2=0 $Y2=0
cc_214 N_A1_c_298_n N_VPWR_c_331_n 0.00154077f $X=4.05 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A1_M1006_g N_VPWR_c_333_n 0.00486043f $X=3.835 $Y=1.985 $X2=0 $Y2=0
cc_216 A1 N_VPWR_c_334_n 0.00855478f $X=4.31 $Y=1.445 $X2=0 $Y2=0
cc_217 N_A1_M1006_g N_VPWR_c_327_n 0.00857998f $X=3.835 $Y=1.985 $X2=0 $Y2=0
cc_218 A1 N_VPWR_c_327_n 0.00736122f $X=4.31 $Y=1.445 $X2=0 $Y2=0
cc_219 N_A1_M1005_g N_VGND_c_413_n 0.00433285f $X=3.835 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A1_M1005_g N_VGND_c_416_n 0.00414138f $X=3.835 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A1_M1005_g N_VGND_c_417_n 0.00701811f $X=3.835 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A1_M1005_g N_A_566_47#_c_471_n 0.012805f $X=3.835 $Y=0.56 $X2=0 $Y2=0
cc_223 A1 N_A_566_47#_c_471_n 0.0281659f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_224 N_A1_c_298_n N_A_566_47#_c_471_n 0.00207059f $X=4.05 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A1_M1005_g N_A_566_47#_c_472_n 0.00561561f $X=3.835 $Y=0.56 $X2=0 $Y2=0
cc_226 N_VPWR_c_327_n N_X_M1003_d 0.00223231f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_c_327_n N_X_c_395_n 0.0126068f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_336_n N_X_c_395_n 0.0196071f $X=1.035 $Y=2.5 $X2=0 $Y2=0
cc_229 N_VPWR_c_327_n A_674_297# 0.00673342f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_230 N_VPWR_c_329_n N_VGND_c_411_n 0.00713034f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_231 N_X_c_395_n N_VGND_c_414_n 0.0196071f $X=0.69 $Y=0.42 $X2=1.167 $Y2=0.885
cc_232 N_X_M1002_d N_VGND_c_417_n 0.00223231f $X=0.55 $Y=0.235 $X2=2.865
+ $Y2=1.905
cc_233 N_X_c_395_n N_VGND_c_417_n 0.0126068f $X=0.69 $Y=0.42 $X2=2.865 $Y2=1.905
cc_234 N_VGND_c_417_n A_386_47# 0.00432467f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_235 N_VGND_c_417_n A_458_47# 0.0132339f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_236 N_VGND_c_417_n N_A_566_47#_M1013_d 0.00444947f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_237 N_VGND_c_417_n N_A_566_47#_M1005_d 0.00213418f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_415_n N_A_566_47#_c_485_n 0.0210051f $X=3.385 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_417_n N_A_566_47#_c_485_n 0.012574f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_M1001_d N_A_566_47#_c_471_n 0.00708013f $X=3.37 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_VGND_c_413_n N_A_566_47#_c_471_n 0.0212136f $X=3.55 $Y=0.37 $X2=0 $Y2=0
cc_242 N_VGND_c_415_n N_A_566_47#_c_471_n 0.00292296f $X=3.385 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_416_n N_A_566_47#_c_471_n 0.00255018f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_417_n N_A_566_47#_c_471_n 0.0103582f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_245 N_VGND_c_416_n N_A_566_47#_c_472_n 0.0208048f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_246 N_VGND_c_417_n N_A_566_47#_c_472_n 0.0123922f $X=4.37 $Y=0 $X2=0 $Y2=0

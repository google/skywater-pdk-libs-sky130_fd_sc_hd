* File: sky130_fd_sc_hd__einvn_8.pex.spice
* Created: Thu Aug 27 14:20:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVN_8%TE_B 1 3 6 8 10 12 13 15 17 18 20 22 23 25
+ 27 28 30 32 33 35 37 38 40 42 43 45 47 48 51 52 53 54 55 56 57 64
c131 56 0 7.37964e-20 $X=3.465 $Y=1.395
c132 55 0 7.37964e-20 $X=3.045 $Y=1.395
c133 54 0 7.37964e-20 $X=2.625 $Y=1.395
c134 53 0 7.37964e-20 $X=2.205 $Y=1.395
c135 52 0 7.37964e-20 $X=1.785 $Y=1.395
c136 51 0 7.37964e-20 $X=1.365 $Y=1.395
c137 48 0 2.52753e-20 $X=0.945 $Y=1.25
c138 43 0 2.02538e-19 $X=3.81 $Y=1.395
c139 38 0 1.51809e-19 $X=3.39 $Y=1.395
c140 33 0 1.50694e-19 $X=2.97 $Y=1.395
c141 28 0 1.51809e-19 $X=2.55 $Y=1.395
c142 23 0 1.50694e-19 $X=2.13 $Y=1.395
c143 18 0 1.51809e-19 $X=1.71 $Y=1.395
c144 6 0 1.13048e-19 $X=0.47 $Y=1.985
r145 63 64 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.545 $Y2=1.16
r146 60 63 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r147 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r148 48 50 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.945 $Y=1.25
+ $X2=0.945 $Y2=1.395
r149 45 47 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.885 $Y=1.47
+ $X2=3.885 $Y2=2.015
r150 44 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.54 $Y=1.395
+ $X2=3.465 $Y2=1.395
r151 43 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.81 $Y=1.395
+ $X2=3.885 $Y2=1.47
r152 43 44 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.81 $Y=1.395
+ $X2=3.54 $Y2=1.395
r153 40 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.465 $Y=1.47
+ $X2=3.465 $Y2=1.395
r154 40 42 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.465 $Y=1.47
+ $X2=3.465 $Y2=2.015
r155 39 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.12 $Y=1.395
+ $X2=3.045 $Y2=1.395
r156 38 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.39 $Y=1.395
+ $X2=3.465 $Y2=1.395
r157 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.39 $Y=1.395
+ $X2=3.12 $Y2=1.395
r158 35 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.045 $Y=1.47
+ $X2=3.045 $Y2=1.395
r159 35 37 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.045 $Y=1.47
+ $X2=3.045 $Y2=2.015
r160 34 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.395
+ $X2=2.625 $Y2=1.395
r161 33 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.97 $Y=1.395
+ $X2=3.045 $Y2=1.395
r162 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.97 $Y=1.395
+ $X2=2.7 $Y2=1.395
r163 30 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.47
+ $X2=2.625 $Y2=1.395
r164 30 32 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.625 $Y=1.47
+ $X2=2.625 $Y2=2.015
r165 29 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=1.395
+ $X2=2.205 $Y2=1.395
r166 28 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.395
+ $X2=2.625 $Y2=1.395
r167 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.55 $Y=1.395
+ $X2=2.28 $Y2=1.395
r168 25 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=1.47
+ $X2=2.205 $Y2=1.395
r169 25 27 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.205 $Y=1.47
+ $X2=2.205 $Y2=2.015
r170 24 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.86 $Y=1.395
+ $X2=1.785 $Y2=1.395
r171 23 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.395
+ $X2=2.205 $Y2=1.395
r172 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.13 $Y=1.395
+ $X2=1.86 $Y2=1.395
r173 20 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.785 $Y=1.47
+ $X2=1.785 $Y2=1.395
r174 20 22 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.785 $Y=1.47
+ $X2=1.785 $Y2=2.015
r175 19 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.44 $Y=1.395
+ $X2=1.365 $Y2=1.395
r176 18 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=1.395
+ $X2=1.785 $Y2=1.395
r177 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.71 $Y=1.395
+ $X2=1.44 $Y2=1.395
r178 15 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.365 $Y=1.47
+ $X2=1.365 $Y2=1.395
r179 15 17 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.365 $Y=1.47
+ $X2=1.365 $Y2=2.015
r180 14 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.395
+ $X2=0.945 $Y2=1.395
r181 13 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.395
+ $X2=1.365 $Y2=1.395
r182 13 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.29 $Y=1.395
+ $X2=1.02 $Y2=1.395
r183 10 50 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=1.47
+ $X2=0.945 $Y2=1.395
r184 10 12 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.945 $Y=1.47
+ $X2=0.945 $Y2=2.015
r185 8 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.25
+ $X2=0.945 $Y2=1.25
r186 8 64 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.87 $Y=1.25
+ $X2=0.545 $Y2=1.25
r187 4 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r188 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r189 1 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r190 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 27 29 30 32 34 35 37 39 40 42 44 45 46 47 48 49 50 51 56 58 59 61 64 75
+ 76
c164 49 0 8.8865e-20 $X=3.51 $Y=1.035
c165 47 0 8.8865e-20 $X=2.67 $Y=1.035
c166 45 0 8.8865e-20 $X=1.83 $Y=1.035
c167 42 0 7.39636e-20 $X=4.35 $Y=0.96
c168 35 0 1.87534e-19 $X=3.855 $Y=1.035
c169 30 0 9.82445e-20 $X=3.435 $Y=1.035
c170 25 0 1.87534e-19 $X=3.015 $Y=1.035
c171 20 0 9.82445e-20 $X=2.595 $Y=1.035
c172 15 0 1.87534e-19 $X=2.175 $Y=1.035
c173 10 0 9.82445e-20 $X=1.755 $Y=1.035
r174 65 76 22.4813 $w=2.68e-07 $l=1.25e-07 $layer=POLY_cond $X=4.305 $Y=1.16
+ $X2=4.305 $Y2=1.035
r175 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=1.16 $X2=4.305 $Y2=1.16
r176 62 75 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=0.68 $Y2=1.16
r177 62 64 120.832 $w=3.28e-07 $l=3.46e-06 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=4.305 $Y2=1.16
r178 60 75 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=1.16
r179 60 61 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=1.495
r180 59 75 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.995
+ $X2=0.68 $Y2=1.16
r181 58 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=0.825
+ $X2=0.68 $Y2=0.995
r182 54 61 30.2064 $w=1.68e-07 $l=4.63e-07 $layer=LI1_cond $X=0.217 $Y=1.58
+ $X2=0.68 $Y2=1.58
r183 54 56 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=1.815
r184 51 58 30.2064 $w=1.68e-07 $l=4.63e-07 $layer=LI1_cond $X=0.217 $Y=0.74
+ $X2=0.68 $Y2=0.74
r185 51 53 4.5451 $w=2.55e-07 $l=9.5e-08 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.217 $Y2=0.56
r186 42 76 22.7584 $w=2.68e-07 $l=9.48683e-08 $layer=POLY_cond $X=4.35 $Y=0.96
+ $X2=4.305 $Y2=1.035
r187 42 44 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.35 $Y=0.96 $X2=4.35
+ $Y2=0.56
r188 41 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.005 $Y=1.035
+ $X2=3.93 $Y2=1.035
r189 40 76 16.3317 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.17 $Y=1.035
+ $X2=4.305 $Y2=1.035
r190 40 41 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.035
+ $X2=4.005 $Y2=1.035
r191 37 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.93 $Y=0.96
+ $X2=3.93 $Y2=1.035
r192 37 39 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.93 $Y=0.96 $X2=3.93
+ $Y2=0.56
r193 36 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=1.035
+ $X2=3.51 $Y2=1.035
r194 35 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.855 $Y=1.035
+ $X2=3.93 $Y2=1.035
r195 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.855 $Y=1.035
+ $X2=3.585 $Y2=1.035
r196 32 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=0.96
+ $X2=3.51 $Y2=1.035
r197 32 34 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.51 $Y=0.96 $X2=3.51
+ $Y2=0.56
r198 31 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.035
+ $X2=3.09 $Y2=1.035
r199 30 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.435 $Y=1.035
+ $X2=3.51 $Y2=1.035
r200 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.435 $Y=1.035
+ $X2=3.165 $Y2=1.035
r201 27 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.09 $Y=0.96
+ $X2=3.09 $Y2=1.035
r202 27 29 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.09 $Y=0.96 $X2=3.09
+ $Y2=0.56
r203 26 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=1.035
+ $X2=2.67 $Y2=1.035
r204 25 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=1.035
+ $X2=3.09 $Y2=1.035
r205 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.015 $Y=1.035
+ $X2=2.745 $Y2=1.035
r206 22 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=0.96
+ $X2=2.67 $Y2=1.035
r207 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.67 $Y=0.96 $X2=2.67
+ $Y2=0.56
r208 21 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.325 $Y=1.035
+ $X2=2.25 $Y2=1.035
r209 20 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.595 $Y=1.035
+ $X2=2.67 $Y2=1.035
r210 20 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.595 $Y=1.035
+ $X2=2.325 $Y2=1.035
r211 17 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=0.96
+ $X2=2.25 $Y2=1.035
r212 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.25 $Y=0.96 $X2=2.25
+ $Y2=0.56
r213 16 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.035
+ $X2=1.83 $Y2=1.035
r214 15 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.175 $Y=1.035
+ $X2=2.25 $Y2=1.035
r215 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.175 $Y=1.035
+ $X2=1.905 $Y2=1.035
r216 12 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=0.96
+ $X2=1.83 $Y2=1.035
r217 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.83 $Y=0.96 $X2=1.83
+ $Y2=0.56
r218 10 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.035
+ $X2=1.83 $Y2=1.035
r219 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.755 $Y=1.035
+ $X2=1.485 $Y2=1.035
r220 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=0.96
+ $X2=1.485 $Y2=1.035
r221 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.41 $Y=0.96 $X2=1.41
+ $Y2=0.56
r222 2 56 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.815
r223 1 53 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 45 48 50 52 55 57 58 59 60 61 62 63 85
r133 83 85 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=7.635 $Y=1.16
+ $X2=7.765 $Y2=1.16
r134 81 83 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=7.345 $Y=1.16
+ $X2=7.635 $Y2=1.16
r135 80 81 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.925 $Y=1.16
+ $X2=7.345 $Y2=1.16
r136 79 80 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.505 $Y=1.16
+ $X2=6.925 $Y2=1.16
r137 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.085 $Y=1.16
+ $X2=6.505 $Y2=1.16
r138 77 78 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.665 $Y=1.16
+ $X2=6.085 $Y2=1.16
r139 76 77 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.245 $Y=1.16
+ $X2=5.665 $Y2=1.16
r140 74 76 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.915 $Y=1.16
+ $X2=5.245 $Y2=1.16
r141 71 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.825 $Y=1.16
+ $X2=4.915 $Y2=1.16
r142 63 83 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=7.635
+ $Y=1.16 $X2=7.635 $Y2=1.16
r143 62 63 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=7.135 $Y=1.14
+ $X2=7.595 $Y2=1.14
r144 61 62 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.675 $Y=1.14
+ $X2=7.135 $Y2=1.14
r145 60 61 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.215 $Y=1.14
+ $X2=6.675 $Y2=1.14
r146 59 60 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=5.755 $Y=1.14
+ $X2=6.215 $Y2=1.14
r147 58 59 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=5.295 $Y=1.14
+ $X2=5.755 $Y2=1.14
r148 57 58 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=4.835 $Y=1.14
+ $X2=5.295 $Y2=1.14
r149 57 74 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=4.915
+ $Y=1.16 $X2=4.915 $Y2=1.16
r150 53 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=1.325
+ $X2=7.765 $Y2=1.16
r151 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.765 $Y=1.325
+ $X2=7.765 $Y2=1.985
r152 50 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=0.995
+ $X2=7.765 $Y2=1.16
r153 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.765 $Y=0.995
+ $X2=7.765 $Y2=0.56
r154 46 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.325
+ $X2=7.345 $Y2=1.16
r155 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.345 $Y=1.325
+ $X2=7.345 $Y2=1.985
r156 43 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=0.995
+ $X2=7.345 $Y2=1.16
r157 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.345 $Y=0.995
+ $X2=7.345 $Y2=0.56
r158 39 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.16
r159 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.985
r160 36 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=0.995
+ $X2=6.925 $Y2=1.16
r161 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.925 $Y=0.995
+ $X2=6.925 $Y2=0.56
r162 32 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=1.325
+ $X2=6.505 $Y2=1.16
r163 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.505 $Y=1.325
+ $X2=6.505 $Y2=1.985
r164 29 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=0.995
+ $X2=6.505 $Y2=1.16
r165 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.505 $Y=0.995
+ $X2=6.505 $Y2=0.56
r166 25 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.085 $Y=1.325
+ $X2=6.085 $Y2=1.16
r167 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.085 $Y=1.325
+ $X2=6.085 $Y2=1.985
r168 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.085 $Y=0.995
+ $X2=6.085 $Y2=1.16
r169 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.085 $Y=0.995
+ $X2=6.085 $Y2=0.56
r170 18 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.665 $Y=1.325
+ $X2=5.665 $Y2=1.16
r171 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.665 $Y=1.325
+ $X2=5.665 $Y2=1.985
r172 15 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.665 $Y=0.995
+ $X2=5.665 $Y2=1.16
r173 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.665 $Y=0.995
+ $X2=5.665 $Y2=0.56
r174 11 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.325
+ $X2=5.245 $Y2=1.16
r175 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.245 $Y=1.325
+ $X2=5.245 $Y2=1.985
r176 8 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=0.995
+ $X2=5.245 $Y2=1.16
r177 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.245 $Y=0.995
+ $X2=5.245 $Y2=0.56
r178 4 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=1.325
+ $X2=4.825 $Y2=1.16
r179 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.825 $Y=1.325
+ $X2=4.825 $Y2=1.985
r180 1 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=1.16
r181 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 47 52 71 72 75 78
r121 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 71 72 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r124 69 72 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=8.05 $Y2=2.72
r125 68 71 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=8.05 $Y2=2.72
r126 68 69 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 66 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r128 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r130 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r131 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r132 60 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r133 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=1.575 $Y2=2.72
r135 57 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 56 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 56 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 53 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r140 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.575 $Y2=2.72
r142 52 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r144 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 45 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 45 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 43 65 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.93 $Y=2.72 $X2=3.91
+ $Y2=2.72
r148 43 44 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.93 $Y=2.72
+ $X2=4.105 $Y2=2.72
r149 42 68 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.28 $Y=2.72 $X2=4.37
+ $Y2=2.72
r150 42 44 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.28 $Y=2.72
+ $X2=4.105 $Y2=2.72
r151 40 62 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.09 $Y=2.72 $X2=2.99
+ $Y2=2.72
r152 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=2.72
+ $X2=3.255 $Y2=2.72
r153 39 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.42 $Y=2.72
+ $X2=3.91 $Y2=2.72
r154 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=2.72
+ $X2=3.255 $Y2=2.72
r155 37 59 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.07 $Y2=2.72
r156 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.415 $Y2=2.72
r157 36 62 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.58 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=2.72
+ $X2=2.415 $Y2=2.72
r159 32 44 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.635
+ $X2=4.105 $Y2=2.72
r160 32 34 20.9086 $w=3.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.105 $Y=2.635
+ $X2=4.105 $Y2=2
r161 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.255 $Y=2.635
+ $X2=3.255 $Y2=2.72
r162 28 30 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.255 $Y=2.635
+ $X2=3.255 $Y2=2.02
r163 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.72
r164 24 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.02
r165 20 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.72
r166 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.02
r167 16 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r168 16 18 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.02
r169 5 34 300 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=2 $X=3.96
+ $Y=1.545 $X2=4.095 $Y2=2
r170 4 30 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.12
+ $Y=1.545 $X2=3.255 $Y2=2.02
r171 3 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.28
+ $Y=1.545 $X2=2.415 $Y2=2.02
r172 2 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.44
+ $Y=1.545 $X2=1.575 $Y2=2.02
r173 1 18 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%A_204_309# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 55 56 57 60 62 66 68 72 74 78 80 81 82 83 84 85
c123 50 0 1.87534e-19 $X=4.45 $Y=1.58
c124 44 0 3.74643e-19 $X=3.59 $Y=1.58
c125 38 0 3.74643e-19 $X=2.75 $Y=1.58
c126 33 0 1.13048e-19 $X=1.24 $Y=1.58
c127 32 0 1.8711e-19 $X=1.91 $Y=1.58
r128 76 78 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=8.042 $Y=2.295
+ $X2=8.042 $Y2=1.96
r129 75 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.38
+ $X2=7.135 $Y2=2.38
r130 74 76 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=7.89 $Y=2.38
+ $X2=8.042 $Y2=2.295
r131 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.89 $Y=2.38
+ $X2=7.22 $Y2=2.38
r132 70 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.135 $Y=2.295
+ $X2=7.135 $Y2=2.38
r133 70 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.135 $Y=2.295
+ $X2=7.135 $Y2=1.96
r134 69 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=2.38
+ $X2=6.295 $Y2=2.38
r135 68 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.05 $Y=2.38
+ $X2=7.135 $Y2=2.38
r136 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.05 $Y=2.38
+ $X2=6.38 $Y2=2.38
r137 64 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.295
+ $X2=6.295 $Y2=2.38
r138 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.295 $Y=2.295
+ $X2=6.295 $Y2=1.96
r139 63 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.54 $Y=2.38
+ $X2=5.455 $Y2=2.38
r140 62 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=2.38
+ $X2=6.295 $Y2=2.38
r141 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.21 $Y=2.38
+ $X2=5.54 $Y2=2.38
r142 58 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.455 $Y2=2.38
r143 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.455 $Y2=1.96
r144 56 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.38
+ $X2=5.455 $Y2=2.38
r145 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.37 $Y=2.38
+ $X2=4.7 $Y2=2.38
r146 53 57 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.575 $Y=2.295
+ $X2=4.7 $Y2=2.38
r147 53 55 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=4.575 $Y=2.295
+ $X2=4.575 $Y2=1.815
r148 52 55 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=4.575 $Y=1.665
+ $X2=4.575 $Y2=1.815
r149 51 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=1.58
+ $X2=3.675 $Y2=1.58
r150 50 52 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.45 $Y=1.58
+ $X2=4.575 $Y2=1.665
r151 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.45 $Y=1.58
+ $X2=3.76 $Y2=1.58
r152 46 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.665
+ $X2=3.675 $Y2=1.58
r153 46 48 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.675 $Y=1.665
+ $X2=3.675 $Y2=1.815
r154 45 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=1.58
+ $X2=2.835 $Y2=1.58
r155 44 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=1.58
+ $X2=3.675 $Y2=1.58
r156 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.59 $Y=1.58
+ $X2=2.92 $Y2=1.58
r157 40 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.835 $Y=1.665
+ $X2=2.835 $Y2=1.58
r158 40 42 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.835 $Y=1.665
+ $X2=2.835 $Y2=1.815
r159 39 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.58
+ $X2=1.995 $Y2=1.58
r160 38 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=1.58
+ $X2=2.835 $Y2=1.58
r161 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.75 $Y=1.58
+ $X2=2.08 $Y2=1.58
r162 34 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=1.665
+ $X2=1.995 $Y2=1.58
r163 34 36 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.995 $Y=1.665
+ $X2=1.995 $Y2=1.815
r164 32 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=1.58
+ $X2=1.995 $Y2=1.58
r165 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.91 $Y=1.58
+ $X2=1.24 $Y2=1.58
r166 28 33 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.127 $Y=1.665
+ $X2=1.24 $Y2=1.58
r167 28 30 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.127 $Y=1.665
+ $X2=1.127 $Y2=1.815
r168 9 78 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.84
+ $Y=1.485 $X2=7.975 $Y2=1.96
r169 8 72 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7
+ $Y=1.485 $X2=7.135 $Y2=1.96
r170 7 66 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.16
+ $Y=1.485 $X2=6.295 $Y2=1.96
r171 6 60 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.32
+ $Y=1.485 $X2=5.455 $Y2=1.96
r172 5 55 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.485 $X2=4.615 $Y2=1.815
r173 4 48 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.54
+ $Y=1.545 $X2=3.675 $Y2=1.815
r174 3 42 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=1.545 $X2=2.835 $Y2=1.815
r175 2 36 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.545 $X2=1.995 $Y2=1.815
r176 1 30 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.545 $X2=1.155 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%Z 1 2 3 4 5 6 7 8 27 29 30 33 35 37 39 41 43
+ 45 47 48 49 50 58 63 67 69
c110 49 0 7.39636e-20 $X=7.97 $Y=0.765
r111 80 82 45.4457 $w=2.03e-07 $l=8.4e-07 $layer=LI1_cond $X=6.715 $Y=0.722
+ $X2=7.555 $Y2=0.722
r112 78 80 45.4457 $w=2.03e-07 $l=8.4e-07 $layer=LI1_cond $X=5.875 $Y=0.722
+ $X2=6.715 $Y2=0.722
r113 75 78 45.4457 $w=2.03e-07 $l=8.4e-07 $layer=LI1_cond $X=5.035 $Y=0.722
+ $X2=5.875 $Y2=0.722
r114 67 69 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=8.082 $Y=0.825
+ $X2=8.082 $Y2=0.85
r115 49 67 3.27477 $w=2.25e-07 $l=1.03e-07 $layer=LI1_cond $X=8.082 $Y=0.722
+ $X2=8.082 $Y2=0.825
r116 49 82 18.6686 $w=2.63e-07 $l=4.15e-07 $layer=LI1_cond $X=7.97 $Y=0.722
+ $X2=7.555 $Y2=0.722
r117 49 50 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=8.082 $Y=0.88
+ $X2=8.082 $Y2=1.19
r118 49 69 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=8.082 $Y=0.88
+ $X2=8.082 $Y2=0.85
r119 48 63 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.555 $Y=1.87
+ $X2=7.555 $Y2=1.7
r120 47 58 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.715 $Y=1.87
+ $X2=6.715 $Y2=1.7
r121 46 50 13.5732 $w=2.23e-07 $l=2.65e-07 $layer=LI1_cond $X=8.082 $Y=1.455
+ $X2=8.082 $Y2=1.19
r122 44 63 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=7.555 $Y=1.625
+ $X2=7.555 $Y2=1.7
r123 44 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=1.625
+ $X2=7.555 $Y2=1.54
r124 42 58 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=6.715 $Y=1.625
+ $X2=6.715 $Y2=1.7
r125 42 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=1.625
+ $X2=6.715 $Y2=1.54
r126 40 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.72 $Y=1.54
+ $X2=7.555 $Y2=1.54
r127 39 46 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=7.97 $Y=1.54
+ $X2=8.082 $Y2=1.455
r128 39 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.97 $Y=1.54
+ $X2=7.72 $Y2=1.54
r129 38 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.88 $Y=1.54
+ $X2=6.715 $Y2=1.54
r130 37 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.39 $Y=1.54
+ $X2=7.555 $Y2=1.54
r131 37 38 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.39 $Y=1.54
+ $X2=6.88 $Y2=1.54
r132 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.04 $Y=1.54
+ $X2=5.875 $Y2=1.54
r133 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.55 $Y=1.54
+ $X2=6.715 $Y2=1.54
r134 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.55 $Y=1.54
+ $X2=6.04 $Y2=1.54
r135 31 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=1.625
+ $X2=5.875 $Y2=1.54
r136 31 33 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.875 $Y=1.625
+ $X2=5.875 $Y2=1.7
r137 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=1.54
+ $X2=5.875 $Y2=1.54
r138 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.71 $Y=1.54
+ $X2=5.2 $Y2=1.54
r139 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.035 $Y=1.625
+ $X2=5.2 $Y2=1.54
r140 25 27 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.035 $Y=1.625
+ $X2=5.035 $Y2=1.7
r141 8 63 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=7.42
+ $Y=1.485 $X2=7.555 $Y2=1.7
r142 7 58 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=6.58
+ $Y=1.485 $X2=6.715 $Y2=1.7
r143 6 33 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=5.74
+ $Y=1.485 $X2=5.875 $Y2=1.7
r144 5 27 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=4.9
+ $Y=1.485 $X2=5.035 $Y2=1.7
r145 4 82 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=7.42
+ $Y=0.235 $X2=7.555 $Y2=0.74
r146 3 80 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.235 $X2=6.715 $Y2=0.74
r147 2 78 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.74
+ $Y=0.235 $X2=5.875 $Y2=0.74
r148 1 75 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.9
+ $Y=0.235 $X2=5.035 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 49 54 70 71 74 77 80
r124 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r125 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r126 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r127 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r128 68 71 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=8.05
+ $Y2=0
r129 67 70 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=8.05
+ $Y2=0
r130 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r131 65 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r132 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r133 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r134 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r135 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r136 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.46
+ $Y2=0
r137 59 61 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=0
+ $X2=2.99 $Y2=0
r138 58 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r139 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r140 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r141 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r142 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r143 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.46
+ $Y2=0
r144 54 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=0
+ $X2=2.07 $Y2=0
r145 53 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r146 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r147 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r148 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r149 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r150 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r151 49 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r152 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r153 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r154 42 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r155 42 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r156 40 64 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.91
+ $Y2=0
r157 40 41 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.145
+ $Y2=0
r158 39 67 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.37
+ $Y2=0
r159 39 41 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.145
+ $Y2=0
r160 37 61 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=0
+ $X2=2.99 $Y2=0
r161 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.3
+ $Y2=0
r162 36 64 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.465 $Y=0
+ $X2=3.91 $Y2=0
r163 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.3
+ $Y2=0
r164 32 41 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=0.085
+ $X2=4.145 $Y2=0
r165 32 34 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=4.145 $Y=0.085
+ $X2=4.145 $Y2=0.36
r166 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085 $X2=3.3
+ $Y2=0
r167 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.36
r168 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r169 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.36
r170 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r171 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.36
r172 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r173 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r174 5 34 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.36
r175 4 30 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.36
r176 3 26 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.36
r177 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.36
r178 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_8%A_215_47# 1 2 3 4 5 6 7 8 9 28 31 32 33 36
+ 38 41 43 46 51 52 60 62 63 64
c98 64 0 1.50694e-19 $X=3.72 $Y=0.74
c99 63 0 1.50694e-19 $X=2.88 $Y=0.74
c100 62 0 1.50694e-19 $X=2.04 $Y=0.74
c101 46 0 5.18434e-20 $X=4.485 $Y=0.74
c102 41 0 2.99402e-19 $X=3.635 $Y=0.74
c103 36 0 2.99402e-19 $X=2.795 $Y=0.74
c104 32 0 2.52753e-20 $X=1.285 $Y=0.74
c105 31 0 2.99402e-19 $X=1.955 $Y=0.74
r106 58 60 47.7762 $w=1.93e-07 $l=8.4e-07 $layer=LI1_cond $X=7.135 $Y=0.352
+ $X2=7.975 $Y2=0.352
r107 56 58 47.7762 $w=1.93e-07 $l=8.4e-07 $layer=LI1_cond $X=6.295 $Y=0.352
+ $X2=7.135 $Y2=0.352
r108 54 56 47.7762 $w=1.93e-07 $l=8.4e-07 $layer=LI1_cond $X=5.455 $Y=0.352
+ $X2=6.295 $Y2=0.352
r109 52 54 42.9417 $w=1.93e-07 $l=7.55e-07 $layer=LI1_cond $X=4.7 $Y=0.352
+ $X2=5.455 $Y2=0.352
r110 49 51 5.09219 $w=2.13e-07 $l=9.5e-08 $layer=LI1_cond $X=4.592 $Y=0.655
+ $X2=4.592 $Y2=0.56
r111 48 52 6.83761 $w=1.95e-07 $l=1.49158e-07 $layer=LI1_cond $X=4.592 $Y=0.45
+ $X2=4.7 $Y2=0.352
r112 48 51 5.89622 $w=2.13e-07 $l=1.1e-07 $layer=LI1_cond $X=4.592 $Y=0.45
+ $X2=4.592 $Y2=0.56
r113 47 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0.74
+ $X2=3.72 $Y2=0.74
r114 46 49 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=4.485 $Y=0.74
+ $X2=4.592 $Y2=0.655
r115 46 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.485 $Y=0.74
+ $X2=3.805 $Y2=0.74
r116 43 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.655
+ $X2=3.72 $Y2=0.74
r117 43 45 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.72 $Y=0.655
+ $X2=3.72 $Y2=0.56
r118 42 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=0.74
+ $X2=2.88 $Y2=0.74
r119 41 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0.74
+ $X2=3.72 $Y2=0.74
r120 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=0.74
+ $X2=2.965 $Y2=0.74
r121 38 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.655
+ $X2=2.88 $Y2=0.74
r122 38 40 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.88 $Y=0.655
+ $X2=2.88 $Y2=0.56
r123 37 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=0.74
+ $X2=2.04 $Y2=0.74
r124 36 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.74
+ $X2=2.88 $Y2=0.74
r125 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.795 $Y=0.74
+ $X2=2.125 $Y2=0.74
r126 33 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.655
+ $X2=2.04 $Y2=0.74
r127 33 35 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.04 $Y=0.655
+ $X2=2.04 $Y2=0.56
r128 31 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=2.04 $Y2=0.74
r129 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=0.74
+ $X2=1.285 $Y2=0.74
r130 28 32 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.15 $Y=0.655
+ $X2=1.285 $Y2=0.74
r131 28 30 4.29259 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=0.655
+ $X2=1.15 $Y2=0.56
r132 9 60 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=7.84
+ $Y=0.235 $X2=7.975 $Y2=0.365
r133 8 58 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=7
+ $Y=0.235 $X2=7.135 $Y2=0.365
r134 7 56 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.235 $X2=6.295 $Y2=0.365
r135 6 54 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.235 $X2=5.455 $Y2=0.365
r136 5 51 182 $w=1.7e-07 $l=3.99061e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.59 $Y2=0.56
r137 4 45 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.56
r138 3 40 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.56
r139 2 35 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.56
r140 1 30 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.56
.ends


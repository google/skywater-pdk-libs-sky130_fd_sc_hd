* File: sky130_fd_sc_hd__o22ai_4.pex.spice
* Created: Tue Sep  1 19:23:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O22AI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 32
+ 33 35 36 39 52
c132 29 0 3.12662e-20 $X=3.275 $Y=1.53
c133 27 0 1.22518e-19 $X=3.44 $Y=1.985
c134 22 0 2.9244e-20 $X=3.44 $Y=0.995
c135 15 0 2.92312e-20 $X=1.34 $Y=0.995
r136 50 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.25 $Y=1.16 $X2=1.34
+ $Y2=1.16
r137 48 50 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=1.25 $Y2=1.16
r138 46 48 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.91 $Y=1.16 $X2=0.92
+ $Y2=1.16
r139 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.91
+ $Y=1.16 $X2=0.91 $Y2=1.16
r140 43 46 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.5 $Y=1.16
+ $X2=0.91 $Y2=1.16
r141 39 47 10.9245 $w=1.98e-07 $l=1.97e-07 $layer=LI1_cond $X=1.107 $Y=1.175
+ $X2=0.91 $Y2=1.175
r142 39 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.16 $X2=1.25 $Y2=1.16
r143 35 38 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=1.16
+ $X2=3.44 $Y2=1.245
r144 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.16 $X2=3.44 $Y2=1.16
r145 33 39 6.30458 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.282 $Y=1.445
+ $X2=1.282 $Y2=1.275
r146 32 38 7.68295 $w=2.98e-07 $l=2e-07 $layer=LI1_cond $X=3.425 $Y=1.445
+ $X2=3.425 $Y2=1.245
r147 30 33 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.415 $Y=1.53
+ $X2=1.282 $Y2=1.445
r148 29 32 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.275 $Y=1.53
+ $X2=3.425 $Y2=1.445
r149 29 30 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=3.275 $Y=1.53
+ $X2=1.415 $Y2=1.53
r150 25 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.325
+ $X2=3.44 $Y2=1.16
r151 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.44 $Y=1.325
+ $X2=3.44 $Y2=1.985
r152 22 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=1.16
r153 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=0.56
r154 18 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.16
r155 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.985
r156 15 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=0.995
+ $X2=1.34 $Y2=1.16
r157 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.34 $Y=0.995
+ $X2=1.34 $Y2=0.56
r158 11 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.16
r159 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.985
r160 8 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=0.995
+ $X2=0.92 $Y2=1.16
r161 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.92 $Y=0.995
+ $X2=0.92 $Y2=0.56
r162 4 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.325
+ $X2=0.5 $Y2=1.16
r163 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.5 $Y=1.325 $X2=0.5
+ $Y2=1.985
r164 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=0.995
+ $X2=0.5 $Y2=1.16
r165 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.5 $Y=0.995 $X2=0.5
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
c82 1 0 2.92312e-20 $X=1.76 $Y=0.995
r83 39 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.93 $Y=1.16 $X2=3.02
+ $Y2=1.16
r84 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.93
+ $Y=1.16 $X2=2.93 $Y2=1.16
r85 37 39 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.6 $Y=1.16 $X2=2.93
+ $Y2=1.16
r86 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.18 $Y=1.16 $X2=2.6
+ $Y2=1.16
r87 34 36 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.91 $Y=1.16
+ $X2=2.18 $Y2=1.16
r88 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.91
+ $Y=1.16 $X2=1.91 $Y2=1.16
r89 31 34 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.76 $Y=1.16
+ $X2=1.91 $Y2=1.16
r90 29 40 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=2.53 $Y=1.175 $X2=2.93
+ $Y2=1.175
r91 29 35 34.3818 $w=1.98e-07 $l=6.2e-07 $layer=LI1_cond $X=2.53 $Y=1.175
+ $X2=1.91 $Y2=1.175
r92 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.02 $Y=1.325
+ $X2=3.02 $Y2=1.16
r93 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.02 $Y=1.325
+ $X2=3.02 $Y2=1.985
r94 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.02 $Y=0.995
+ $X2=3.02 $Y2=1.16
r95 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.02 $Y=0.995
+ $X2=3.02 $Y2=0.56
r96 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.325
+ $X2=2.6 $Y2=1.16
r97 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.6 $Y=1.325 $X2=2.6
+ $Y2=1.985
r98 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=0.995
+ $X2=2.6 $Y2=1.16
r99 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.6 $Y=0.995 $X2=2.6
+ $Y2=0.56
r100 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=1.325
+ $X2=2.18 $Y2=1.16
r101 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.18 $Y=1.325
+ $X2=2.18 $Y2=1.985
r102 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=0.995
+ $X2=2.18 $Y2=1.16
r103 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.18 $Y=0.995
+ $X2=2.18 $Y2=0.56
r104 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.325
+ $X2=1.76 $Y2=1.16
r105 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.76 $Y=1.325
+ $X2=1.76 $Y2=1.985
r106 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=0.995
+ $X2=1.76 $Y2=1.16
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.76 $Y=0.995
+ $X2=1.76 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%B1 1 3 6 8 10 13 15 17 20 24 27 29 33 34 36
+ 44 47 53
c117 13 0 1.75548e-19 $X=4.33 $Y=1.985
c118 1 0 1.69878e-19 $X=3.91 $Y=0.995
r119 42 44 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.72 $Y=1.16 $X2=4.75
+ $Y2=1.16
r120 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.72
+ $Y=1.16 $X2=4.72 $Y2=1.16
r121 40 42 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.33 $Y=1.16
+ $X2=4.72 $Y2=1.16
r122 38 40 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.91 $Y=1.16
+ $X2=4.33 $Y2=1.16
r123 36 53 9.22546 $w=6.18e-07 $l=1.1e-07 $layer=LI1_cond $X=4.83 $Y=1.305
+ $X2=4.94 $Y2=1.305
r124 36 43 2.12207 $w=6.18e-07 $l=1.1e-07 $layer=LI1_cond $X=4.83 $Y=1.305
+ $X2=4.72 $Y2=1.305
r125 34 48 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.865 $Y=1.16
+ $X2=6.865 $Y2=1.325
r126 34 47 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.865 $Y=1.16
+ $X2=6.865 $Y2=0.995
r127 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.16 $X2=6.85 $Y2=1.16
r128 31 33 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=6.825 $Y=1.445
+ $X2=6.825 $Y2=1.16
r129 29 31 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.715 $Y=1.53
+ $X2=6.825 $Y2=1.445
r130 29 53 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=6.715 $Y=1.53
+ $X2=4.94 $Y2=1.53
r131 27 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.85 $Y=1.985
+ $X2=6.85 $Y2=1.325
r132 24 47 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.85 $Y=0.56
+ $X2=6.85 $Y2=0.995
r133 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=1.325
+ $X2=4.75 $Y2=1.16
r134 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.75 $Y=1.325
+ $X2=4.75 $Y2=1.985
r135 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.16
r136 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=0.56
r137 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.33 $Y=1.325
+ $X2=4.33 $Y2=1.16
r138 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.33 $Y=1.325
+ $X2=4.33 $Y2=1.985
r139 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=1.16
r140 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.33 $Y=0.995
+ $X2=4.33 $Y2=0.56
r141 4 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=1.325
+ $X2=3.91 $Y2=1.16
r142 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.91 $Y=1.325
+ $X2=3.91 $Y2=1.985
r143 1 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=0.995
+ $X2=3.91 $Y2=1.16
r144 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.91 $Y=0.995
+ $X2=3.91 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 41
r62 39 41 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.295 $Y=1.16
+ $X2=6.43 $Y2=1.16
r63 37 39 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=6.01 $Y=1.16
+ $X2=6.295 $Y2=1.16
r64 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.59 $Y=1.16
+ $X2=6.01 $Y2=1.16
r65 34 36 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.275 $Y=1.16
+ $X2=5.59 $Y2=1.16
r66 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.275
+ $Y=1.16 $X2=5.275 $Y2=1.16
r67 31 34 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=5.17 $Y=1.16
+ $X2=5.275 $Y2=1.16
r68 29 35 51.85 $w=1.98e-07 $l=9.35e-07 $layer=LI1_cond $X=6.21 $Y=1.175
+ $X2=5.275 $Y2=1.175
r69 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.295
+ $Y=1.16 $X2=6.295 $Y2=1.16
r70 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.16
r71 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.985
r72 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=1.16
r73 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=0.56
r74 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.01 $Y=1.325
+ $X2=6.01 $Y2=1.16
r75 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.01 $Y=1.325
+ $X2=6.01 $Y2=1.985
r76 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.01 $Y=0.995
+ $X2=6.01 $Y2=1.16
r77 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.01 $Y=0.995
+ $X2=6.01 $Y2=0.56
r78 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.59 $Y=1.325
+ $X2=5.59 $Y2=1.16
r79 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.59 $Y=1.325
+ $X2=5.59 $Y2=1.985
r80 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.59 $Y=0.995
+ $X2=5.59 $Y2=1.16
r81 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.59 $Y=0.995
+ $X2=5.59 $Y2=0.56
r82 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.17 $Y=1.325
+ $X2=5.17 $Y2=1.16
r83 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.17 $Y=1.325 $X2=5.17
+ $Y2=1.985
r84 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.16
r85 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.17 $Y=0.995 $X2=5.17
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%VPWR 1 2 3 4 5 16 18 24 28 32 34 36 39 40 42
+ 43 44 46 61 72 76
r116 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r117 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 67 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r120 64 67 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 63 66 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=6.67 $Y2=2.72
r122 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 61 75 4.22854 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=6.935 $Y=2.72
+ $X2=7.147 $Y2=2.72
r124 61 66 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.935 $Y=2.72
+ $X2=6.67 $Y2=2.72
r125 60 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r126 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r128 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 54 57 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r130 54 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 53 56 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r132 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r133 51 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.13 $Y2=2.72
r134 51 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 50 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r136 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 47 69 3.95154 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.207 $Y2=2.72
r138 47 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.69 $Y2=2.72
r139 46 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=1.13 $Y2=2.72
r140 46 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.69 $Y2=2.72
r141 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r142 44 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r143 42 59 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.37 $Y2=2.72
r144 42 43 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.545 $Y2=2.72
r145 41 63 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 41 43 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.665 $Y=2.72
+ $X2=4.545 $Y2=2.72
r147 39 56 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.565 $Y=2.72
+ $X2=3.45 $Y2=2.72
r148 39 40 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.565 $Y=2.72
+ $X2=3.675 $Y2=2.72
r149 38 59 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=4.37 $Y2=2.72
r150 38 40 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.675 $Y2=2.72
r151 34 75 3.13151 $w=2.8e-07 $l=1.15521e-07 $layer=LI1_cond $X=7.075 $Y=2.635
+ $X2=7.147 $Y2=2.72
r152 34 36 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.075 $Y=2.635
+ $X2=7.075 $Y2=2.3
r153 30 43 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=2.635
+ $X2=4.545 $Y2=2.72
r154 30 32 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=4.545 $Y=2.635
+ $X2=4.545 $Y2=2.3
r155 26 40 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=2.635
+ $X2=3.675 $Y2=2.72
r156 26 28 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=3.675 $Y=2.635
+ $X2=3.675 $Y2=2.3
r157 22 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2.72
r158 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2.3
r159 18 21 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.29 $Y=1.62
+ $X2=0.29 $Y2=2.3
r160 16 69 3.19163 $w=2.5e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.29 $Y=2.635
+ $X2=0.207 $Y2=2.72
r161 16 21 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.29 $Y=2.635
+ $X2=0.29 $Y2=2.3
r162 5 36 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.925
+ $Y=1.485 $X2=7.06 $Y2=2.3
r163 4 32 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=1.485 $X2=4.54 $Y2=2.3
r164 3 28 600 $w=1.7e-07 $l=8.98248e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.69 $Y2=2.3
r165 2 24 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.13 $Y2=2.3
r166 1 21 400 $w=1.7e-07 $l=8.89129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.29 $Y2=2.3
r167 1 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.29 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%A_115_297# 1 2 3 4 15 19 21 27 28 29 33 38
r51 38 40 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=3.25 $Y=2.3 $X2=3.25
+ $Y2=2.38
r52 33 35 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.39 $Y=2.3 $X2=2.39
+ $Y2=2.38
r53 30 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=2.38
+ $X2=2.39 $Y2=2.38
r54 29 40 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.105 $Y=2.38
+ $X2=3.25 $Y2=2.38
r55 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.105 $Y=2.38
+ $X2=2.515 $Y2=2.38
r56 27 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=2.38
+ $X2=2.39 $Y2=2.38
r57 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.265 $Y=2.38
+ $X2=1.675 $Y2=2.38
r58 24 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.55 $Y=2.295
+ $X2=1.675 $Y2=2.38
r59 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.55 $Y=2.295
+ $X2=1.55 $Y2=1.96
r60 23 26 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.55 $Y=1.955
+ $X2=1.55 $Y2=1.96
r61 22 31 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.835 $Y=1.87
+ $X2=0.71 $Y2=1.87
r62 21 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.425 $Y=1.87
+ $X2=1.55 $Y2=1.955
r63 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.425 $Y=1.87
+ $X2=0.835 $Y2=1.87
r64 17 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.955
+ $X2=0.71 $Y2=1.87
r65 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.71 $Y=1.955
+ $X2=0.71 $Y2=1.96
r66 13 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.785
+ $X2=0.71 $Y2=1.87
r67 13 15 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=1.785
+ $X2=0.71 $Y2=1.62
r68 4 38 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.485 $X2=3.23 $Y2=2.3
r69 3 33 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.255
+ $Y=1.485 $X2=2.39 $Y2=2.3
r70 2 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.485 $X2=1.55 $Y2=1.96
r71 1 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=1.485 $X2=0.71 $Y2=1.96
r72 1 15 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.485 $X2=0.71 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%Y 1 2 3 4 5 6 7 8 25 28 29 30 31 39 41 44 45
+ 52 54 57 62 67 72
c131 54 0 1.44282e-19 $X=3.745 $Y=1.87
c132 30 0 1.22518e-19 $X=4.04 $Y=1.445
r133 70 72 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.935 $Y=1.87
+ $X2=2.99 $Y2=1.87
r134 67 77 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.81 $Y=1.87 $X2=2.81
+ $Y2=1.96
r135 67 70 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.81 $Y=1.87
+ $X2=2.935 $Y2=1.87
r136 67 72 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.005 $Y=1.87
+ $X2=2.99 $Y2=1.87
r137 62 65 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=6.22 $Y=1.87 $X2=6.22
+ $Y2=1.96
r138 57 60 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.38 $Y=1.87 $X2=5.38
+ $Y2=1.96
r139 54 67 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.745 $Y=1.87
+ $X2=3.005 $Y2=1.87
r140 50 52 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.83 $Y=1.53
+ $X2=4.04 $Y2=1.53
r141 45 48 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.97 $Y=1.87 $X2=1.97
+ $Y2=1.96
r142 43 44 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.19 $Y=0.82
+ $X2=7.19 $Y2=1.785
r143 42 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.345 $Y=1.87
+ $X2=6.22 $Y2=1.87
r144 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.105 $Y=1.87
+ $X2=7.19 $Y2=1.785
r145 41 42 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.105 $Y=1.87
+ $X2=6.345 $Y2=1.87
r146 40 57 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.505 $Y=1.87
+ $X2=5.38 $Y2=1.87
r147 39 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.095 $Y=1.87
+ $X2=6.22 $Y2=1.87
r148 39 40 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.095 $Y=1.87
+ $X2=5.505 $Y2=1.87
r149 36 38 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=5.8 $Y=0.732
+ $X2=6.64 $Y2=0.732
r150 34 36 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=4.96 $Y=0.732
+ $X2=5.8 $Y2=0.732
r151 32 56 3.35006 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0.732
+ $X2=4.04 $Y2=0.732
r152 32 34 52.9195 $w=1.73e-07 $l=8.35e-07 $layer=LI1_cond $X=4.125 $Y=0.732
+ $X2=4.96 $Y2=0.732
r153 31 43 6.81835 $w=1.75e-07 $l=1.23386e-07 $layer=LI1_cond $X=7.105 $Y=0.732
+ $X2=7.19 $Y2=0.82
r154 31 38 29.4701 $w=1.73e-07 $l=4.65e-07 $layer=LI1_cond $X=7.105 $Y=0.732
+ $X2=6.64 $Y2=0.732
r155 30 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.445
+ $X2=4.04 $Y2=1.53
r156 29 56 3.4683 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=4.04 $Y=0.82 $X2=4.04
+ $Y2=0.732
r157 29 30 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.04 $Y=0.82
+ $X2=4.04 $Y2=1.445
r158 28 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.83 $Y=1.785
+ $X2=3.745 $Y2=1.87
r159 27 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=1.615
+ $X2=3.83 $Y2=1.53
r160 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.83 $Y=1.615
+ $X2=3.83 $Y2=1.785
r161 26 45 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.095 $Y=1.87
+ $X2=1.97 $Y2=1.87
r162 25 67 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.685 $Y=1.87
+ $X2=2.81 $Y2=1.87
r163 25 26 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.685 $Y=1.87
+ $X2=2.095 $Y2=1.87
r164 8 65 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.085
+ $Y=1.485 $X2=6.22 $Y2=1.96
r165 7 60 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.245
+ $Y=1.485 $X2=5.38 $Y2=1.96
r166 6 77 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.485 $X2=2.81 $Y2=1.96
r167 5 48 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.485 $X2=1.97 $Y2=1.96
r168 4 38 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.64 $Y2=0.73
r169 3 36 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.665
+ $Y=0.235 $X2=5.8 $Y2=0.73
r170 2 34 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.73
r171 1 56 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.12 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%A_797_297# 1 2 3 4 15 16 21 22 23 26 27 30
+ 35
r51 35 37 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.64 $Y=2.3 $X2=6.64
+ $Y2=2.38
r52 30 32 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.8 $Y=2.3 $X2=5.8
+ $Y2=2.38
r53 26 27 8.86878 $w=2.98e-07 $l=1.75e-07 $layer=LI1_cond $X=4.105 $Y=2.3
+ $X2=4.105 $Y2=2.125
r54 24 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.925 $Y=2.38
+ $X2=5.8 $Y2=2.38
r55 23 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.515 $Y=2.38
+ $X2=6.64 $Y2=2.38
r56 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.515 $Y=2.38
+ $X2=5.925 $Y2=2.38
r57 21 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.675 $Y=2.38
+ $X2=5.8 $Y2=2.38
r58 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.675 $Y=2.38
+ $X2=5.085 $Y2=2.38
r59 18 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.96 $Y=2.295
+ $X2=5.085 $Y2=2.38
r60 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.96 $Y=2.295
+ $X2=4.96 $Y2=1.96
r61 17 20 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.96 $Y=1.955
+ $X2=4.96 $Y2=1.96
r62 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.835 $Y=1.87
+ $X2=4.96 $Y2=1.955
r63 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.835 $Y=1.87
+ $X2=4.255 $Y2=1.87
r64 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.17 $Y=1.955
+ $X2=4.255 $Y2=1.87
r65 13 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.17 $Y=1.955
+ $X2=4.17 $Y2=2.125
r66 4 35 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.505
+ $Y=1.485 $X2=6.64 $Y2=2.3
r67 3 30 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.665
+ $Y=1.485 $X2=5.8 $Y2=2.3
r68 2 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.825
+ $Y=1.485 $X2=4.96 $Y2=1.96
r69 1 26 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.985
+ $Y=1.485 $X2=4.12 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%A_33_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 52 55 64 66 67 68
c124 68 0 2.9244e-20 $X=2.81 $Y=0.815
c125 67 0 2.92312e-20 $X=1.97 $Y=0.815
c126 66 0 2.92312e-20 $X=1.13 $Y=0.815
c127 50 0 1.69878e-19 $X=3.485 $Y=0.82
r128 62 64 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=6.22 $Y=0.365
+ $X2=7.06 $Y2=0.365
r129 60 62 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=5.38 $Y=0.365
+ $X2=6.22 $Y2=0.365
r130 58 60 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=4.54 $Y=0.365
+ $X2=5.38 $Y2=0.365
r131 56 70 4.05488 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=3.785 $Y=0.365
+ $X2=3.635 $Y2=0.365
r132 56 58 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=3.785 $Y=0.365
+ $X2=4.54 $Y2=0.365
r133 53 55 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=3.635 $Y=0.735
+ $X2=3.635 $Y2=0.73
r134 52 70 2.97358 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.635 $Y=0.475
+ $X2=3.635 $Y2=0.365
r135 52 55 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.635 $Y=0.475
+ $X2=3.635 $Y2=0.73
r136 51 68 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.975 $Y=0.82
+ $X2=2.81 $Y2=0.815
r137 50 53 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.485 $Y=0.82
+ $X2=3.635 $Y2=0.735
r138 50 51 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.485 $Y=0.82
+ $X2=2.975 $Y2=0.82
r139 46 68 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.81 $Y=0.725
+ $X2=2.81 $Y2=0.815
r140 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.81 $Y=0.725
+ $X2=2.81 $Y2=0.39
r141 45 67 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0.815
+ $X2=1.97 $Y2=0.815
r142 44 68 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0.815
+ $X2=2.81 $Y2=0.815
r143 44 45 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.645 $Y=0.815
+ $X2=2.135 $Y2=0.815
r144 40 67 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.97 $Y=0.725
+ $X2=1.97 $Y2=0.815
r145 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.97 $Y=0.725
+ $X2=1.97 $Y2=0.39
r146 39 66 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.295 $Y=0.82
+ $X2=1.13 $Y2=0.815
r147 38 67 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.805 $Y=0.82
+ $X2=1.97 $Y2=0.815
r148 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.805 $Y=0.82
+ $X2=1.295 $Y2=0.82
r149 34 66 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.13 $Y=0.725
+ $X2=1.13 $Y2=0.815
r150 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.13 $Y=0.725
+ $X2=1.13 $Y2=0.39
r151 32 66 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0.815
+ $X2=1.13 $Y2=0.815
r152 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=0.965 $Y=0.815
+ $X2=0.455 $Y2=0.815
r153 28 33 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.29 $Y=0.725
+ $X2=0.455 $Y2=0.815
r154 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.29 $Y=0.725
+ $X2=0.29 $Y2=0.39
r155 9 64 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.925
+ $Y=0.235 $X2=7.06 $Y2=0.39
r156 8 62 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.235 $X2=6.22 $Y2=0.39
r157 7 60 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.38 $Y2=0.39
r158 6 58 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.235 $X2=4.54 $Y2=0.39
r159 5 70 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.65 $Y2=0.39
r160 5 55 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.65 $Y2=0.73
r161 4 48 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.675
+ $Y=0.235 $X2=2.81 $Y2=0.39
r162 3 42 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.835
+ $Y=0.235 $X2=1.97 $Y2=0.39
r163 2 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.235 $X2=1.13 $Y2=0.39
r164 1 30 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_4%VGND 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 56 57 60
r100 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r101 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r102 54 57 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=7.13
+ $Y2=0
r103 53 56 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=7.13
+ $Y2=0
r104 53 54 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r105 51 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r106 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r107 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r108 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r109 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r110 45 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r111 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r112 42 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.71
+ $Y2=0
r113 42 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=1.15 $Y2=0
r114 40 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r115 38 50 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.145 $Y=0
+ $X2=2.99 $Y2=0
r116 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.23
+ $Y2=0
r117 37 53 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.45 $Y2=0
r118 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.23
+ $Y2=0
r119 35 47 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.07 $Y2=0
r120 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.39
+ $Y2=0
r121 34 50 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.99 $Y2=0
r122 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.39
+ $Y2=0
r123 32 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.15 $Y2=0
r124 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.55
+ $Y2=0
r125 31 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.635 $Y=0
+ $X2=2.07 $Y2=0
r126 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.55
+ $Y2=0
r127 27 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0.085
+ $X2=3.23 $Y2=0
r128 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.23 $Y=0.085
+ $X2=3.23 $Y2=0.39
r129 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0
r130 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0.39
r131 19 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r132 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.39
r133 15 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r134 15 17 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.39
r135 4 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.235 $X2=3.23 $Y2=0.39
r136 3 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.255
+ $Y=0.235 $X2=2.39 $Y2=0.39
r137 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.55 $Y2=0.39
r138 1 17 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.71 $Y2=0.39
.ends


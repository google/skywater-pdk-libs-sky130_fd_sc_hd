* File: sky130_fd_sc_hd__xnor3_2.pex.spice
* Created: Tue Sep  1 19:33:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_87_21# 1 2 7 9 12 14 16 19 21 22 23 25 26
+ 28 30 32 33 35 40 42 43
c113 19 0 1.74668e-19 $X=0.95 $Y=1.985
r114 48 49 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.93 $Y=1.16 $X2=0.95
+ $Y2=1.16
r115 47 48 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=0.53 $Y=1.16 $X2=0.93
+ $Y2=1.16
r116 45 47 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.51 $Y=1.16 $X2=0.53
+ $Y2=1.16
r117 42 43 15.2541 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=2.8 $Y=0.355
+ $X2=2.53 $Y2=0.355
r118 40 49 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.045 $Y=1.16
+ $X2=0.95 $Y2=1.16
r119 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.045
+ $Y=1.16 $X2=1.045 $Y2=1.16
r120 37 39 24.4 $w=1.9e-07 $l=3.8e-07 $layer=LI1_cond $X=1.062 $Y=0.78 $X2=1.062
+ $Y2=1.16
r121 33 35 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=1.68 $Y=2.32
+ $X2=2.725 $Y2=2.32
r122 32 43 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.565 $Y=0.34
+ $X2=2.53 $Y2=0.34
r123 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.595 $Y=2.235
+ $X2=1.68 $Y2=2.32
r124 29 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.595 $Y=2.045
+ $X2=1.595 $Y2=2.235
r125 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.48 $Y=0.425
+ $X2=1.565 $Y2=0.34
r126 27 28 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.48 $Y=0.425
+ $X2=1.48 $Y2=0.695
r127 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.51 $Y=1.96
+ $X2=1.595 $Y2=2.045
r128 25 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.51 $Y=1.96
+ $X2=1.165 $Y2=1.96
r129 24 37 1.386 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.165 $Y=0.78
+ $X2=1.062 $Y2=0.78
r130 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.395 $Y=0.78
+ $X2=1.48 $Y2=0.695
r131 23 24 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.395 $Y=0.78
+ $X2=1.165 $Y2=0.78
r132 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.08 $Y=1.875
+ $X2=1.165 $Y2=1.96
r133 21 39 10.7577 $w=1.9e-07 $l=1.73767e-07 $layer=LI1_cond $X=1.08 $Y=1.325
+ $X2=1.062 $Y2=1.16
r134 21 22 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.08 $Y=1.325
+ $X2=1.08 $Y2=1.875
r135 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.325
+ $X2=0.95 $Y2=1.16
r136 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.95 $Y=1.325
+ $X2=0.95 $Y2=1.985
r137 14 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r138 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=0.56
r139 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.325
+ $X2=0.53 $Y2=1.16
r140 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.53 $Y=1.325
+ $X2=0.53 $Y2=1.985
r141 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=1.16
r142 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=0.56
r143 2 35 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.625 $X2=2.725 $Y2=2.32
r144 1 42 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.655
+ $Y=0.245 $X2=2.8 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%C 1 3 4 6 9 11 13 15 16 17 18
c64 1 0 1.70967e-19 $X=1.465 $Y=0.995
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.16 $X2=2.375 $Y2=1.16
r66 18 22 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.53 $Y=1.2
+ $X2=2.375 $Y2=1.2
r67 16 21 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.44 $Y=1.16
+ $X2=2.375 $Y2=1.16
r68 16 17 5.03009 $w=3.3e-07 $l=1.14254e-07 $layer=POLY_cond $X=2.44 $Y=1.16
+ $X2=2.547 $Y2=1.175
r69 14 21 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=1.54 $Y=1.16
+ $X2=2.375 $Y2=1.16
r70 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=1.16
+ $X2=1.465 $Y2=1.16
r71 11 17 37.0704 $w=1.5e-07 $l=1.95806e-07 $layer=POLY_cond $X=2.58 $Y=0.995
+ $X2=2.547 $Y2=1.175
r72 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.58 $Y=0.995
+ $X2=2.58 $Y2=0.565
r73 7 17 37.0704 $w=1.5e-07 $l=1.95346e-07 $layer=POLY_cond $X=2.515 $Y=1.355
+ $X2=2.547 $Y2=1.175
r74 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.515 $Y=1.355
+ $X2=2.515 $Y2=2.045
r75 4 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.325
+ $X2=1.465 $Y2=1.16
r76 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.465 $Y=1.325
+ $X2=1.465 $Y2=1.805
r77 1 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=1.16
r78 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_308_93# 1 2 7 9 12 13 18 20 23 24 28 29 32
c75 13 0 1.74668e-19 $X=1.735 $Y=1.62
r76 29 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.16 $X2=3
+ $Y2=0.995
r77 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r78 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.895 $Y=1.16 $X2=3
+ $Y2=1.16
r79 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=1.325
+ $X2=2.895 $Y2=1.16
r80 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.895 $Y=1.325
+ $X2=2.895 $Y2=1.535
r81 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=1.62
+ $X2=1.82 $Y2=1.62
r82 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.81 $Y=1.62
+ $X2=2.895 $Y2=1.535
r83 20 21 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.81 $Y=1.62
+ $X2=1.905 $Y2=1.62
r84 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=1.535
+ $X2=1.82 $Y2=1.62
r85 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.82 $Y=1.535
+ $X2=1.82 $Y2=0.76
r86 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=1.62
+ $X2=1.82 $Y2=1.62
r87 13 15 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=1.735 $Y=1.62 $X2=1.675
+ $Y2=1.62
r88 12 32 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.02 $Y=0.565
+ $X2=3.02 $Y2=0.995
r89 7 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.325 $X2=3
+ $Y2=1.16
r90 7 9 186.373 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3 $Y=1.325 $X2=3
+ $Y2=1.905
r91 2 15 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.485 $X2=1.675 $Y2=1.62
r92 1 18 182 $w=1.7e-07 $l=4.11856e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.465 $X2=1.82 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_827_297# 1 2 9 13 15 17 19 21 22 23 27 35
+ 37 38 39 40 47 49 50 58
c169 49 0 1.83334e-19 $X=7.13 $Y=0.85
c170 27 0 1.36535e-19 $X=4.405 $Y=1.58
c171 15 0 1.24749e-19 $X=7.305 $Y=1.28
r172 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.11 $X2=7.25 $Y2=1.11
r173 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.18 $Y=0.85
+ $X2=7.18 $Y2=1.11
r174 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.85
+ $X2=7.13 $Y2=0.85
r175 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0.85
+ $X2=5.75 $Y2=0.85
r176 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0.85
+ $X2=4.37 $Y2=0.85
r177 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.895 $Y=0.85
+ $X2=5.75 $Y2=0.85
r178 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=7.13 $Y2=0.85
r179 39 40 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=5.895 $Y2=0.85
r180 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=0.85
+ $X2=4.37 $Y2=0.85
r181 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.605 $Y=0.85
+ $X2=5.75 $Y2=0.85
r182 37 38 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=5.605 $Y=0.85
+ $X2=4.515 $Y2=0.85
r183 35 47 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=5.73 $Y=0.995
+ $X2=5.73 $Y2=0.85
r184 31 35 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=5.58 $Y=1.132
+ $X2=5.73 $Y2=1.132
r185 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.58
+ $Y=1.16 $X2=5.58 $Y2=1.16
r186 28 58 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.405 $Y=1.445
+ $X2=4.405 $Y2=0.74
r187 27 28 1.42499 $w=2.4e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=1.58
+ $X2=4.405 $Y2=1.445
r188 25 27 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.27 $Y=1.58
+ $X2=4.405 $Y2=1.58
r189 22 32 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=5.84 $Y=1.16
+ $X2=5.58 $Y2=1.16
r190 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.84 $Y=1.16
+ $X2=5.915 $Y2=1.16
r191 19 55 38.945 $w=2.68e-07 $l=1.92678e-07 $layer=POLY_cond $X=7.31 $Y=0.945
+ $X2=7.25 $Y2=1.11
r192 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.31 $Y=0.945
+ $X2=7.31 $Y2=0.535
r193 15 55 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=7.305 $Y=1.28
+ $X2=7.25 $Y2=1.11
r194 15 17 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=7.305 $Y=1.28
+ $X2=7.305 $Y2=2.065
r195 11 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.325
+ $X2=5.915 $Y2=1.16
r196 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.915 $Y=1.325
+ $X2=5.915 $Y2=1.805
r197 7 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=0.995
+ $X2=5.915 $Y2=1.16
r198 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.915 $Y=0.995
+ $X2=5.915 $Y2=0.455
r199 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.27 $Y2=1.63
r200 1 58 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.44 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%B 3 7 9 10 13 18 19 20 23 27 31 34 35 37 38
+ 41
r121 37 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=1.53
+ $X2=7.13 $Y2=1.53
r122 35 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.16
+ $X2=6.77 $Y2=1.325
r123 35 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.16
+ $X2=6.77 $Y2=0.995
r124 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.16 $X2=6.77 $Y2=1.16
r125 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.77 $Y=1.445
+ $X2=6.855 $Y2=1.53
r126 32 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.77 $Y=1.445
+ $X2=6.77 $Y2=1.16
r127 28 30 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.06 $Y=1.16
+ $X2=4.23 $Y2=1.16
r128 27 42 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.79 $Y=1.965
+ $X2=6.79 $Y2=1.325
r129 25 27 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.79 $Y=2.465
+ $X2=6.79 $Y2=1.965
r130 23 41 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.71 $Y=0.565
+ $X2=6.71 $Y2=0.995
r131 19 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.715 $Y=2.54
+ $X2=6.79 $Y2=2.465
r132 19 20 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=6.715 $Y=2.54
+ $X2=5.235 $Y2=2.54
r133 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.16 $Y=2.465
+ $X2=5.235 $Y2=2.54
r134 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.16 $Y=2.465
+ $X2=5.16 $Y2=1.905
r135 15 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.16 $Y=1.235
+ $X2=5.16 $Y2=1.16
r136 15 18 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.16 $Y=1.235
+ $X2=5.16 $Y2=1.905
r137 11 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.16 $Y=1.085
+ $X2=5.16 $Y2=1.16
r138 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.16 $Y=1.085
+ $X2=5.16 $Y2=0.565
r139 10 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=1.16
+ $X2=4.23 $Y2=1.16
r140 9 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.085 $Y=1.16
+ $X2=5.16 $Y2=1.16
r141 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.085 $Y=1.16
+ $X2=4.305 $Y2=1.16
r142 5 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.23 $Y=1.085
+ $X2=4.23 $Y2=1.16
r143 5 7 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.23 $Y=1.085
+ $X2=4.23 $Y2=0.56
r144 1 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.06 $Y=1.235
+ $X2=4.06 $Y2=1.16
r145 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.06 $Y=1.235
+ $X2=4.06 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A 3 6 8 11 12 13
c44 13 0 1.83334e-19 $X=7.74 $Y=0.995
r45 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.74 $Y=1.16
+ $X2=7.74 $Y2=1.325
r46 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.74 $Y=1.16
+ $X2=7.74 $Y2=0.995
r47 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.73
+ $Y=1.16 $X2=7.73 $Y2=1.16
r48 8 12 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=7.59 $Y=1.2 $X2=7.73
+ $Y2=1.2
r49 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.81 $Y=1.985
+ $X2=7.81 $Y2=1.325
r50 3 13 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.81 $Y=0.555
+ $X2=7.81 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_933_297# 1 2 3 4 13 15 18 22 24 28 29 30
+ 31 36 37 38 41 44 45
c135 36 0 1.4656e-19 $X=8.23 $Y=1.16
c136 31 0 1.06604e-19 $X=8.17 $Y=1.495
c137 30 0 1.40536e-19 $X=8.17 $Y=1.325
r138 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0.51
+ $X2=7.59 $Y2=0.51
r139 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0.51
+ $X2=4.83 $Y2=0.51
r140 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=0.51
+ $X2=4.83 $Y2=0.51
r141 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=0.51
+ $X2=7.59 $Y2=0.51
r142 37 38 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=7.445 $Y=0.51
+ $X2=4.975 $Y2=0.51
r143 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=1.16 $X2=8.23 $Y2=1.16
r144 33 35 20.4335 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=8.2 $Y=0.82 $X2=8.2
+ $Y2=1.16
r145 32 45 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=7.62 $Y=0.735
+ $X2=7.62 $Y2=0.51
r146 30 35 10.2745 $w=2.03e-07 $l=1.79374e-07 $layer=LI1_cond $X=8.17 $Y=1.325
+ $X2=8.2 $Y2=1.16
r147 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.17 $Y=1.325
+ $X2=8.17 $Y2=1.495
r148 29 32 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.765 $Y=0.82
+ $X2=7.62 $Y2=0.735
r149 28 33 1.77774 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.085 $Y=0.82
+ $X2=8.2 $Y2=0.82
r150 28 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.085 $Y=0.82
+ $X2=7.765 $Y2=0.82
r151 24 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.085 $Y=1.6
+ $X2=8.17 $Y2=1.495
r152 24 26 25.6147 $w=2.08e-07 $l=4.85e-07 $layer=LI1_cond $X=8.085 $Y=1.6
+ $X2=7.6 $Y2=1.6
r153 20 41 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=0.595
+ $X2=4.79 $Y2=0.43
r154 20 22 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.79 $Y=0.595
+ $X2=4.79 $Y2=1.94
r155 16 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.16
r156 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.985
r157 13 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=1.16
r158 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=0.555
r159 4 26 600 $w=1.7e-07 $l=2.32164e-07 $layer=licon1_PDIFF $count=1 $X=7.38
+ $Y=1.645 $X2=7.6 $Y2=1.62
r160 3 22 600 $w=1.7e-07 $l=5.13712e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=1.485 $X2=4.79 $Y2=1.94
r161 2 45 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=7.385
+ $Y=0.235 $X2=7.6 $Y2=0.625
r162 1 41 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.245 $X2=4.95 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%VPWR 1 2 3 4 13 15 21 25 29 31 33 38 46 56
+ 57 63 66 69
c98 4 0 1.06604e-19 $X=7.885 $Y=1.485
r99 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r100 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 57 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r103 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r104 54 69 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.19 $Y=2.72
+ $X2=8.022 $Y2=2.72
r105 54 56 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.19 $Y=2.72
+ $X2=8.51 $Y2=2.72
r106 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r107 52 53 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r108 50 53 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=7.59 $Y2=2.72
r109 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r110 49 52 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=7.59 $Y2=2.72
r111 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r112 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.85 $Y2=2.72
r113 47 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.37 $Y2=2.72
r114 46 69 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.855 $Y=2.72
+ $X2=8.022 $Y2=2.72
r115 46 52 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.855 $Y=2.72
+ $X2=7.59 $Y2=2.72
r116 45 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r117 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 42 45 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 42 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 41 44 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r121 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 39 63 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.33 $Y=2.72
+ $X2=1.162 $Y2=2.72
r123 39 41 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.33 $Y=2.72
+ $X2=1.61 $Y2=2.72
r124 38 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.85 $Y2=2.72
r125 38 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 37 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r128 34 60 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.187 $Y2=2.72
r129 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 33 63 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=1.162 $Y2=2.72
r131 33 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r133 31 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r134 27 69 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.022 $Y=2.635
+ $X2=8.022 $Y2=2.72
r135 27 29 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=8.022 $Y=2.635
+ $X2=8.022 $Y2=2.36
r136 23 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.72
r137 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.32
r138 19 63 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.162 $Y=2.635
+ $X2=1.162 $Y2=2.72
r139 19 21 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.162 $Y=2.635
+ $X2=1.162 $Y2=2.3
r140 15 18 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=0.23 $Y=1.66
+ $X2=0.23 $Y2=2.34
r141 13 60 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=2.635
+ $X2=0.187 $Y2=2.72
r142 13 18 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.23 $Y=2.635
+ $X2=0.23 $Y2=2.34
r143 4 29 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.36
r144 3 25 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.725
+ $Y=2.175 $X2=3.85 $Y2=2.32
r145 2 21 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.485 $X2=1.165 $Y2=2.3
r146 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r147 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%X 1 2 9 13 14 15 16 19
r27 16 23 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.685 $Y=1.87
+ $X2=0.685 $Y2=2.3
r28 16 19 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.685 $Y=1.87
+ $X2=0.685 $Y2=1.62
r29 14 19 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=0.685 $Y=1.58
+ $X2=0.685 $Y2=1.62
r30 14 15 5.97229 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.685 $Y=1.58
+ $X2=0.685 $Y2=1.44
r31 13 15 24.2248 $w=2.43e-07 $l=5.15e-07 $layer=LI1_cond $X=0.667 $Y=0.925
+ $X2=0.667 $Y2=1.44
r32 7 13 5.81426 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.675 $Y=0.795
+ $X2=0.675 $Y2=0.925
r33 7 9 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=0.675 $Y=0.795
+ $X2=0.675 $Y2=0.56
r34 2 23 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.74 $Y2=2.3
r35 2 19 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.74 $Y2=1.62
r36 1 9 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.235 $X2=0.72 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_423_325# 1 2 3 4 13 17 22 24 25 28 29 30
+ 32 35 39 43 45 46 48
c149 29 0 1.36535e-19 $X=5.045 $Y=2.36
r150 46 47 14.9388 $w=1.96e-07 $l=2.4e-07 $layer=LI1_cond $X=5.13 $Y=0.772
+ $X2=5.37 $Y2=0.772
r151 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.68 $Y=1.12
+ $X2=3.79 $Y2=1.12
r152 37 47 1.57051 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=5.37 $Y=0.655
+ $X2=5.37 $Y2=0.772
r153 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.37 $Y=0.655
+ $X2=5.37 $Y2=0.545
r154 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=2.36
+ $X2=5.13 $Y2=2.36
r155 33 35 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=5.215 $Y=2.36
+ $X2=7.085 $Y2=2.36
r156 32 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=2.275
+ $X2=5.13 $Y2=2.36
r157 31 46 1.57051 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=5.13 $Y=0.89
+ $X2=5.13 $Y2=0.772
r158 31 32 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.13 $Y=0.89
+ $X2=5.13 $Y2=2.275
r159 29 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=2.36
+ $X2=5.13 $Y2=2.36
r160 29 30 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.045 $Y=2.36
+ $X2=4.52 $Y2=2.36
r161 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=2.275
+ $X2=4.52 $Y2=2.36
r162 27 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.435 $Y=2.065
+ $X2=4.435 $Y2=2.275
r163 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=1.98
+ $X2=3.79 $Y2=1.98
r164 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=1.98
+ $X2=4.435 $Y2=2.065
r165 25 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.35 $Y=1.98
+ $X2=3.875 $Y2=1.98
r166 24 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=1.895
+ $X2=3.79 $Y2=1.98
r167 23 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=1.205
+ $X2=3.79 $Y2=1.12
r168 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.79 $Y=1.205
+ $X2=3.79 $Y2=1.895
r169 22 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.035
+ $X2=3.68 $Y2=1.12
r170 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.68 $Y=0.455
+ $X2=3.68 $Y2=1.035
r171 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=0.37
+ $X2=3.68 $Y2=0.455
r172 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.595 $Y=0.37
+ $X2=3.3 $Y2=0.37
r173 13 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=1.98
+ $X2=3.79 $Y2=1.98
r174 13 15 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.705 $Y=1.98
+ $X2=2.305 $Y2=1.98
r175 4 35 600 $w=1.7e-07 $l=8.17634e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=1.645 $X2=7.085 $Y2=2.36
r176 3 15 600 $w=1.7e-07 $l=4.39858e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.625 $X2=2.305 $Y2=1.98
r177 2 39 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=5.235
+ $Y=0.245 $X2=5.37 $Y2=0.545
r178 1 19 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.245 $X2=3.3 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_447_49# 1 2 3 4 13 16 17 19 21 24 26 30 32
+ 33 35 36 39 42
c129 32 0 1.24749e-19 $X=6.93 $Y=0.38
r130 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.53
+ $X2=5.75 $Y2=1.53
r131 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=1.53
+ $X2=3.45 $Y2=1.53
r132 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.595 $Y=1.53
+ $X2=3.45 $Y2=1.53
r133 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.605 $Y=1.53
+ $X2=5.75 $Y2=1.53
r134 35 36 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=5.605 $Y=1.53
+ $X2=3.595 $Y2=1.53
r135 32 33 13.3743 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=6.93 $Y=0.36
+ $X2=6.685 $Y2=0.36
r136 28 30 10.6148 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=2.37 $Y=0.765
+ $X2=2.585 $Y2=0.765
r137 26 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.175 $Y=0.34
+ $X2=6.685 $Y2=0.34
r138 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.09 $Y=0.425
+ $X2=6.175 $Y2=0.34
r139 23 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.09 $Y=0.425
+ $X2=6.09 $Y2=1.445
r140 22 43 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=5.81 $Y=1.53
+ $X2=5.602 $Y2=1.53
r141 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.005 $Y=1.53
+ $X2=6.09 $Y2=1.445
r142 21 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.005 $Y=1.53
+ $X2=5.81 $Y2=1.53
r143 17 43 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.602 $Y=1.615
+ $X2=5.602 $Y2=1.53
r144 17 19 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=5.602 $Y=1.615
+ $X2=5.602 $Y2=1.62
r145 16 39 8.59825 $w=3.35e-07 $l=1.55997e-07 $layer=LI1_cond $X=3.34 $Y=1.375
+ $X2=3.342 $Y2=1.53
r146 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.34 $Y=0.795
+ $X2=3.34 $Y2=1.375
r147 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.255 $Y=0.71
+ $X2=3.34 $Y2=0.795
r148 13 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.255 $Y=0.71
+ $X2=2.585 $Y2=0.71
r149 4 19 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=5.235
+ $Y=1.485 $X2=5.57 $Y2=1.62
r150 3 39 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.485 $X2=3.315 $Y2=1.61
r151 2 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.245 $X2=6.93 $Y2=0.38
r152 1 28 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.245 $X2=2.37 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%A_1198_49# 1 2 3 4 15 18 23 26 29 31 36
c67 29 0 1.17772e-19 $X=8.17 $Y=1.99
r68 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.44 $Y=0.42
+ $X2=8.57 $Y2=0.42
r69 28 29 14.5869 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.445 $Y=1.99
+ $X2=8.17 $Y2=1.99
r70 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.57 $Y=1.875
+ $X2=8.57 $Y2=1.99
r71 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=0.585
+ $X2=8.57 $Y2=0.42
r72 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=8.57 $Y=0.585
+ $X2=8.57 $Y2=1.875
r73 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=8.507 $Y=1.99
+ $X2=8.57 $Y2=1.99
r74 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=8.507 $Y=1.99
+ $X2=8.445 $Y2=1.99
r75 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=8.507 $Y=2.105
+ $X2=8.507 $Y2=2.3
r76 20 29 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=6.58 $Y=2.02
+ $X2=8.17 $Y2=2.02
r77 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.515 $Y=2.02
+ $X2=6.58 $Y2=2.02
r78 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.43 $Y=1.935
+ $X2=6.515 $Y2=2.02
r79 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.43 $Y=1.935
+ $X2=6.43 $Y2=0.76
r80 4 28 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.445 $Y2=1.96
r81 4 23 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.445 $Y2=2.3
r82 3 20 600 $w=1.7e-07 $l=8.14709e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.485 $X2=6.58 $Y2=2.02
r83 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.42
r84 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.245 $X2=6.43 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR3_2%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34 35
+ 37 53 54 60
c108 54 0 1.70967e-19 $X=8.51 $Y=0
c109 27 0 2.87884e-20 $X=8.02 $Y=0.4
c110 4 0 1.40536e-19 $X=7.885 $Y=0.235
r111 60 61 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r112 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r113 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r114 50 51 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r115 48 51 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=7.59 $Y2=0
r116 47 50 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=7.59
+ $Y2=0
r117 47 48 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r118 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r119 45 61 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=1.15 $Y2=0
r120 44 45 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r121 42 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.1
+ $Y2=0
r122 42 44 175.171 $w=1.68e-07 $l=2.685e-06 $layer=LI1_cond $X=1.225 $Y=0
+ $X2=3.91 $Y2=0
r123 41 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r124 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r125 38 57 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r126 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.69 $Y2=0
r127 37 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.1
+ $Y2=0
r128 37 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.69 $Y2=0
r129 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r130 35 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r131 33 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.59
+ $Y2=0
r132 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=0 $X2=8.02
+ $Y2=0
r133 32 53 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=8.51 $Y2=0
r134 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.02
+ $Y2=0
r135 30 44 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=3.91
+ $Y2=0
r136 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=4.02
+ $Y2=0
r137 29 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.105 $Y=0
+ $X2=4.37 $Y2=0
r138 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.02
+ $Y2=0
r139 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0
r140 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0.4
r141 21 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r142 21 23 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.36
r143 17 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r144 17 19 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.36
r145 13 57 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.187 $Y2=0
r146 13 15 18.8762 $w=2.88e-07 $l=4.75e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.23 $Y2=0.56
r147 4 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.4
r148 3 23 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=3.865
+ $Y=0.235 $X2=4.02 $Y2=0.36
r149 2 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.36
r150 1 15 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends


* File: sky130_fd_sc_hd__o21bai_1.spice.pex
* Created: Thu Aug 27 14:36:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21BAI_1%B1_N 3 5 6 7 8 10 15 16 18 21
c42 6 0 7.39193e-20 $X=0.785 $Y=1.61
r43 16 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.45 $Y=1.16
+ $X2=0.45 $Y2=1.325
r44 16 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.45 $Y=1.16
+ $X2=0.45 $Y2=0.995
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.16 $X2=0.45 $Y2=1.16
r46 12 18 8.35926 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.22 $Y=1.345
+ $X2=0.22 $Y2=1.53
r47 11 15 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=0.22 $Y=1.17 $X2=0.45
+ $Y2=1.17
r48 11 12 2.25943 $w=2.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.22 $Y=1.17
+ $X2=0.22 $Y2=1.345
r49 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.86 $Y=1.685 $X2=0.86
+ $Y2=1.97
r50 6 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.785 $Y=1.61
+ $X2=0.86 $Y2=1.685
r51 6 7 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=0.785 $Y=1.61 $X2=0.585
+ $Y2=1.61
r52 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.51 $Y=1.535
+ $X2=0.585 $Y2=1.61
r53 5 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.51 $Y=1.535
+ $X2=0.51 $Y2=1.325
r54 3 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%A_105_352# 1 2 7 9 12 14 15 18 22 23 25 32
+ 34
r67 32 33 5.6903 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.68 $Y=0.66
+ $X2=0.805 $Y2=0.66
r68 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.16 $X2=0.93 $Y2=1.16
r69 23 25 14.6497 $w=2.93e-07 $l=3.75e-07 $layer=LI1_cond $X=0.867 $Y=1.535
+ $X2=0.867 $Y2=1.16
r70 22 34 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=0.867 $Y=1.142
+ $X2=0.867 $Y2=0.995
r71 22 25 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=0.867 $Y=1.142
+ $X2=0.867 $Y2=1.16
r72 20 33 3.40055 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=0.825
+ $X2=0.805 $Y2=0.66
r73 20 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.805 $Y=0.825
+ $X2=0.805 $Y2=0.995
r74 16 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.662 $Y=1.62
+ $X2=0.867 $Y2=1.62
r75 16 18 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=0.662 $Y=1.705
+ $X2=0.662 $Y2=1.96
r76 14 26 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=0.93 $Y2=1.16
r77 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.41 $Y2=1.16
r78 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r79 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.985
r80 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r81 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
r82 2 18 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.76 $X2=0.65 $Y2=1.96
r83 1 32 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.68 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%A2 3 7 8 11 12 13
c37 13 0 6.26376e-20 $X=1.85 $Y=0.995
r38 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=1.325
r39 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=0.995
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.16 $X2=1.85 $Y2=1.16
r41 8 12 12.6753 $w=2.08e-07 $l=2.4e-07 $layer=LI1_cond $X=1.61 $Y=1.18 $X2=1.85
+ $Y2=1.18
r42 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.87 $Y=0.56 $X2=1.87
+ $Y2=0.995
r43 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.865 $Y=1.985
+ $X2=1.865 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%A1 3 7 8 11 13
r25 11 14 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.16
+ $X2=2.37 $Y2=1.325
r26 11 13 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.16
+ $X2=2.37 $Y2=0.995
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.16 $X2=2.38 $Y2=1.16
r28 8 12 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=1.18 $X2=2.38
+ $Y2=1.18
r29 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.29 $Y=0.56 $X2=2.29
+ $Y2=0.995
r30 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.27 $Y=1.985
+ $X2=2.27 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%VPWR 1 2 9 13 15 19 21 26 32 36
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 30 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 27 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=2.72
+ $X2=1.135 $Y2=2.72
r46 27 29 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.3 $Y=2.72 $X2=2.07
+ $Y2=2.72
r47 26 35 5.14828 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.515 $Y2=2.72
r48 26 29 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.27 $Y=2.72 $X2=2.07
+ $Y2=2.72
r49 24 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 21 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=2.72
+ $X2=1.135 $Y2=2.72
r52 21 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.97 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 19 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 15 18 20.8976 $w=3.73e-07 $l=6.8e-07 $layer=LI1_cond $X=2.457 $Y=1.62
+ $X2=2.457 $Y2=2.3
r55 13 35 3.00492 $w=3.75e-07 $l=1.1025e-07 $layer=LI1_cond $X=2.457 $Y=2.635
+ $X2=2.515 $Y2=2.72
r56 13 18 10.2952 $w=3.73e-07 $l=3.35e-07 $layer=LI1_cond $X=2.457 $Y=2.635
+ $X2=2.457 $Y2=2.3
r57 9 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.135 $Y=1.96
+ $X2=1.135 $Y2=2.3
r58 7 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=2.635
+ $X2=1.135 $Y2=2.72
r59 7 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.135 $Y=2.635
+ $X2=1.135 $Y2=2.3
r60 2 18 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.485 $X2=2.48 $Y2=2.3
r61 2 15 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.485 $X2=2.48 $Y2=1.62
r62 1 12 600 $w=1.7e-07 $l=6.32139e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=1.76 $X2=1.135 $Y2=2.3
r63 1 9 600 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=1.76 $X2=1.135 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%Y 1 2 11 12 13 17 20
c47 20 0 7.39193e-20 $X=1.61 $Y=2.21
c48 13 0 6.26376e-20 $X=1.235 $Y=0.825
r49 20 25 3.19138 $w=3.23e-07 $l=9e-08 $layer=LI1_cond $X=1.632 $Y=2.21
+ $X2=1.632 $Y2=2.3
r50 17 20 20.744 $w=3.23e-07 $l=5.85e-07 $layer=LI1_cond $X=1.632 $Y=1.625
+ $X2=1.632 $Y2=2.21
r51 14 17 23.6171 $w=1.68e-07 $l=3.62e-07 $layer=LI1_cond $X=1.27 $Y=1.54
+ $X2=1.632 $Y2=1.54
r52 12 13 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=1.235 $Y=0.645
+ $X2=1.235 $Y2=0.825
r53 11 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=1.455
+ $X2=1.27 $Y2=1.54
r54 11 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.27 $Y=1.455
+ $X2=1.27 $Y2=0.825
r55 9 12 7.17647 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.2 $Y=0.545 $X2=1.2
+ $Y2=0.645
r56 2 25 400 $w=1.7e-07 $l=8.95977e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.655 $Y2=2.3
r57 2 17 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.655 $Y2=1.62
r58 1 9 182 $w=1.7e-07 $l=3.67219e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%VGND 1 2 7 9 13 15 17 24 25 31
r38 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r39 25 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r41 22 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.08
+ $Y2=0
r42 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.53
+ $Y2=0
r43 21 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r44 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 18 28 4.29305 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r46 18 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.69
+ $Y2=0
r47 17 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.08
+ $Y2=0
r48 17 20 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=1.995 $Y=0 $X2=0.69
+ $Y2=0
r49 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r50 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 11 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r52 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.39
r53 7 28 3.02899 $w=2.75e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.18 $Y2=0
r54 7 9 24.0965 $w=2.73e-07 $l=5.75e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.222 $Y2=0.66
r55 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.235 $X2=2.08 $Y2=0.39
r56 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_1%A_297_47# 1 2 10 11 12 15 18
r29 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.5 $Y=0.735
+ $X2=2.5 $Y2=0.39
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=0.82
+ $X2=2.5 $Y2=0.735
r31 11 12 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.335 $Y=0.82
+ $X2=1.74 $Y2=0.82
r32 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.655 $Y=0.735
+ $X2=1.74 $Y2=0.82
r33 8 10 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.655 $Y=0.735
+ $X2=1.655 $Y2=0.73
r34 7 18 6.0176 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.655 $Y=0.485
+ $X2=1.655 $Y2=0.39
r35 7 10 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.655 $Y=0.485
+ $X2=1.655 $Y2=0.73
r36 2 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.235 $X2=2.5 $Y2=0.39
r37 1 18 182 $w=1.7e-07 $l=2.35053e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.655 $Y2=0.39
r38 1 10 182 $w=1.7e-07 $l=5.73738e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.655 $Y2=0.73
.ends


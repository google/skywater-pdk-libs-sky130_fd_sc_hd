* NGSPICE file created from sky130_fd_sc_hd__o41ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 VGND A2 a_109_47# VNB nshort w=650000u l=150000u
+  ad=4.03e+11p pd=3.84e+06u as=7.6375e+11p ps=6.25e+06u
M1001 a_109_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_432_297# A2 a_348_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.5e+11p pd=2.7e+06u as=2.7e+11p ps=2.54e+06u
M1003 a_193_297# A4 Y VPB phighvt w=1e+06u l=150000u
+  ad=6.25e+11p pd=3.25e+06u as=2.7e+11p ps=2.54e+06u
M1004 VPWR A1 a_432_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1005 a_348_297# A3 a_193_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A4 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_109_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1009 a_109_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


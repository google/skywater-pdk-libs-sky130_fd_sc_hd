* File: sky130_fd_sc_hd__lpflow_decapkapwr_3.pxi.spice
* Created: Thu Aug 27 14:24:29 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%VGND N_VGND_M1001_s N_VGND_c_16_n
+ N_VGND_M1000_g N_VGND_c_17_n VGND N_VGND_c_18_n N_VGND_c_19_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%KAPWR N_KAPWR_M1000_s N_KAPWR_c_32_n
+ KAPWR N_KAPWR_M1001_g N_KAPWR_c_35_n N_KAPWR_c_36_n N_KAPWR_c_37_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%VPWR VPWR N_VPWR_c_52_n N_VPWR_c_51_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3%VPWR
cc_1 VNB N_VGND_c_16_n 0.0201334f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.76
cc_2 VNB N_VGND_c_17_n 0.0220173f $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=1.29
cc_3 VNB N_VGND_c_18_n 0.0862828f $X=-0.19 $Y=-0.24 $X2=1.12 $Y2=0.485
cc_4 VNB N_VGND_c_19_n 0.102847f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=0
cc_5 VNB N_KAPWR_c_32_n 0.015747f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=2.05
cc_6 VNB N_KAPWR_M1001_g 0.0972186f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0.375
cc_7 VNB N_VPWR_c_51_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=2.05
cc_8 VPB N_VGND_c_16_n 0.0842436f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.76
cc_9 VPB N_VGND_c_17_n 0.0051139f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.29
cc_10 VPB N_KAPWR_c_32_n 0.0122601f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=2.05
cc_11 VPB N_KAPWR_c_35_n 0.0679976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_12 VPB N_KAPWR_c_36_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_13 VPB N_KAPWR_c_37_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_14 VPB N_VPWR_c_52_n 0.0366162f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=2.05
cc_15 VPB N_VPWR_c_51_n 0.0418424f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=2.05
cc_16 N_VGND_c_16_n N_KAPWR_c_32_n 0.0146807f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_17 N_VGND_c_17_n N_KAPWR_c_32_n 0.0329927f $X=0.42 $Y=1.29 $X2=0 $Y2=0
cc_18 N_VGND_c_18_n N_KAPWR_c_32_n 0.0453111f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_19 N_VGND_c_16_n N_KAPWR_M1001_g 0.0377751f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_20 N_VGND_c_17_n N_KAPWR_M1001_g 0.0139364f $X=0.42 $Y=1.29 $X2=0 $Y2=0
cc_21 N_VGND_c_18_n N_KAPWR_M1001_g 0.0749649f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_22 N_VGND_c_16_n N_KAPWR_c_35_n 0.0749675f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_23 N_VGND_c_17_n N_KAPWR_c_35_n 0.0458866f $X=0.42 $Y=1.29 $X2=0 $Y2=0
cc_24 N_VGND_c_16_n N_VPWR_c_52_n 0.0140765f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_25 N_VGND_c_16_n N_VPWR_c_51_n 0.0155015f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_26 N_KAPWR_c_35_n N_VPWR_c_52_n 0.0793411f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_27 N_KAPWR_c_37_n N_VPWR_c_52_n 9.03925e-19 $X=0.215 $Y=2.21 $X2=0 $Y2=0
cc_28 N_KAPWR_M1000_s N_VPWR_c_51_n 0.00214099f $X=0.135 $Y=1.615 $X2=0 $Y2=0
cc_29 N_KAPWR_c_35_n N_VPWR_c_51_n 0.0105602f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_30 N_KAPWR_c_37_n N_VPWR_c_51_n 0.12706f $X=0.215 $Y=2.21 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o31ai_4.spice
* Created: Tue Sep  1 19:25:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o31ai_4.pex.spice"
.subckt sky130_fd_sc_hd__o31ai_4  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_31_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75007 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1008_d N_A1_M1012_g N_A_31_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A1_M1019_g N_A_31_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75006.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1019_d N_A1_M1020_g N_A_31_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75005.8 A=0.0975 P=1.6 MULT=1
MM1016 N_A_31_47#_M1020_s N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1021 N_A_31_47#_M1021_d N_A2_M1021_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1023 N_A_31_47#_M1021_d N_A2_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1029 N_A_31_47#_M1029_d N_A2_M1029_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1001 N_A_31_47#_M1029_d N_A3_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.222625 PD=0.92 PS=1.335 NRD=0 NRS=12.912 M=1 R=4.33333
+ SA=75003.5 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1002 N_A_31_47#_M1002_d N_A3_M1002_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.222625 PD=0.92 PS=1.335 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1013 N_A_31_47#_M1002_d N_A3_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75004.8 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1024 N_A_31_47#_M1024_d N_A3_M1024_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75005.3 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1003 N_A_31_47#_M1024_d N_B1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.8
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1006 N_A_31_47#_M1006_d N_B1_M1006_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1011 N_A_31_47#_M1006_d N_B1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1014 N_A_31_47#_M1014_d N_B1_M1014_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_27_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1007_d N_A1_M1022_g N_A_27_297#_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1026_d N_A1_M1026_g N_A_27_297#_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1031 N_VPWR_M1026_d N_A1_M1031_g N_A_27_297#_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1005 N_A_27_297#_M1031_s N_A2_M1005_g N_A_449_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1017 N_A_27_297#_M1017_d N_A2_M1017_g N_A_449_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1018 N_A_27_297#_M1017_d N_A2_M1018_g N_A_449_297#_M1018_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1027 N_A_27_297#_M1027_d N_A2_M1027_g N_A_449_297#_M1018_s VPB PHIGHVT L=0.15
+ W=1 AD=0.2605 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1004_d N_A3_M1004_g N_A_449_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2628 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1009 N_Y_M1009_d N_A3_M1009_g N_A_449_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1028 N_Y_M1009_d N_A3_M1028_g N_A_449_297#_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1030 N_Y_M1030_d N_A3_M1030_g N_A_449_297#_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1030_d N_B1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1010_d N_B1_M1010_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1015 N_Y_M1010_d N_B1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1025 N_Y_M1025_d N_B1_M1025_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__o31ai_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_4.pex.spice
* Created: Tue Sep  1 19:11:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%A 3 7 11 13 17 21 23 27 31 33
+ 37 41 45 47 48 49 50 51 53 54 55 56 57 58 59
r112 69 70 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r113 59 70 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=2.53 $Y=1.177
+ $X2=2.36 $Y2=1.177
r114 58 70 14.8537 $w=2.23e-07 $l=2.9e-07 $layer=LI1_cond $X=2.07 $Y=1.177
+ $X2=2.36 $Y2=1.177
r115 57 58 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=1.177
+ $X2=2.07 $Y2=1.177
r116 56 57 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.177
+ $X2=1.61 $Y2=1.177
r117 55 56 25.0976 $w=2.23e-07 $l=4.9e-07 $layer=LI1_cond $X=0.66 $Y=1.177
+ $X2=1.15 $Y2=1.177
r118 55 66 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.66
+ $Y=1.16 $X2=0.66 $Y2=1.16
r119 54 69 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.36
+ $Y2=1.16
r120 52 69 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=2.31 $Y=1.16 $X2=2.36
+ $Y2=1.16
r121 52 53 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=1.16
+ $X2=2.235 $Y2=1.16
r122 48 66 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=0.87 $Y=1.16
+ $X2=0.66 $Y2=1.16
r123 48 49 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.16
+ $X2=0.945 $Y2=1.16
r124 47 66 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=0.59 $Y=1.16 $X2=0.66
+ $Y2=1.16
r125 43 54 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.59 $Y2=1.16
r126 43 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.665 $Y2=1.985
r127 39 53 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=1.295
+ $X2=2.235 $Y2=1.16
r128 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.235 $Y=1.295
+ $X2=2.235 $Y2=1.985
r129 35 53 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=1.025
+ $X2=2.235 $Y2=1.16
r130 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.235 $Y=1.025
+ $X2=2.235 $Y2=0.445
r131 34 51 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.805 $Y2=1.16
r132 33 53 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=1.16
+ $X2=2.235 $Y2=1.16
r133 33 34 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.16 $Y=1.16
+ $X2=1.88 $Y2=1.16
r134 29 51 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.805 $Y=1.295
+ $X2=1.805 $Y2=1.16
r135 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.805 $Y=1.295
+ $X2=1.805 $Y2=1.985
r136 25 51 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.805 $Y=1.025
+ $X2=1.805 $Y2=1.16
r137 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.805 $Y=1.025
+ $X2=1.805 $Y2=0.445
r138 24 50 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.16
+ $X2=1.375 $Y2=1.16
r139 23 51 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.805 $Y2=1.16
r140 23 24 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.45 $Y2=1.16
r141 19 50 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.375 $Y=1.295
+ $X2=1.375 $Y2=1.16
r142 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.375 $Y=1.295
+ $X2=1.375 $Y2=1.985
r143 15 50 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.375 $Y=1.025
+ $X2=1.375 $Y2=1.16
r144 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.375 $Y=1.025
+ $X2=1.375 $Y2=0.445
r145 14 49 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=0.945 $Y2=1.16
r146 13 50 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.3 $Y=1.16
+ $X2=1.375 $Y2=1.16
r147 13 14 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.3 $Y=1.16
+ $X2=1.02 $Y2=1.16
r148 9 49 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.945 $Y=1.295
+ $X2=0.945 $Y2=1.16
r149 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.945 $Y=1.295
+ $X2=0.945 $Y2=1.985
r150 5 49 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.945 $Y=1.025
+ $X2=0.945 $Y2=1.16
r151 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.945 $Y=1.025
+ $X2=0.945 $Y2=0.445
r152 1 47 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.515 $Y=1.295
+ $X2=0.59 $Y2=1.16
r153 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.515 $Y=1.295
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%KAPWR 1 2 3 4 14 17 22 23 27 28
+ 32 35 42 47 52 58
r74 38 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.28 $Y=2.21
+ $X2=0.28 $Y2=2.21
r75 35 38 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.3 $Y=1.965
+ $X2=0.3 $Y2=2.21
r76 32 58 0.00150602 $w=2.49e-07 $l=3e-09 $layer=MET1_cond $X=0.252 $Y=2.21
+ $X2=0.255 $Y2=2.21
r77 31 52 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.88 $Y=2.21
+ $X2=2.88 $Y2=1.965
r78 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.92 $Y=2.21
+ $X2=2.92 $Y2=2.21
r79 26 47 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.02 $Y=2.21
+ $X2=2.02 $Y2=1.965
r80 25 28 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.04 $Y=2.21
+ $X2=2.185 $Y2=2.21
r81 25 27 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.04 $Y=2.21
+ $X2=1.895 $Y2=2.21
r82 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.04 $Y=2.21
+ $X2=2.04 $Y2=2.21
r83 23 27 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=1.285 $Y=2.24
+ $X2=1.895 $Y2=2.24
r84 21 42 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.16 $Y=2.21
+ $X2=1.16 $Y2=1.965
r85 20 23 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.14 $Y=2.21
+ $X2=1.285 $Y2=2.21
r86 20 22 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.14 $Y=2.21
+ $X2=0.995 $Y2=2.21
r87 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=2.21
+ $X2=1.14 $Y2=2.21
r88 17 30 0.0784173 $w=2.46e-07 $l=1.59295e-07 $layer=MET1_cond $X=2.775 $Y=2.24
+ $X2=2.92 $Y2=2.21
r89 17 28 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=2.775 $Y=2.24
+ $X2=2.185 $Y2=2.24
r90 14 58 0.0905443 $w=2.49e-07 $l=1.84391e-07 $layer=MET1_cond $X=0.425 $Y=2.24
+ $X2=0.255 $Y2=2.21
r91 14 22 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=0.425 $Y=2.24
+ $X2=0.995 $Y2=2.24
r92 4 52 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.485 $X2=2.88 $Y2=1.965
r93 3 47 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.88
+ $Y=1.485 $X2=2.02 $Y2=1.965
r94 2 42 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.485 $X2=1.16 $Y2=1.965
r95 1 35 300 $w=1.7e-07 $l=5.56417e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.3 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%Y 1 2 3 4 5 17 18 19 20 21 24
+ 26 30 32 36 38 42 44 48 50 52 53 54 55 56 57 58 59 65 66
r141 59 66 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=1.545
+ $X2=2.985 $Y2=1.46
r142 59 66 0.307318 $w=2.98e-07 $l=8e-09 $layer=LI1_cond $X=2.985 $Y=1.452
+ $X2=2.985 $Y2=1.46
r143 58 59 10.0647 $w=2.98e-07 $l=2.62e-07 $layer=LI1_cond $X=2.985 $Y=1.19
+ $X2=2.985 $Y2=1.452
r144 57 65 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.81
+ $X2=2.985 $Y2=0.895
r145 57 58 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=2.985 $Y=0.915
+ $X2=2.985 $Y2=1.19
r146 57 65 0.768295 $w=2.98e-07 $l=2e-08 $layer=LI1_cond $X=2.985 $Y=0.915
+ $X2=2.985 $Y2=0.895
r147 51 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=1.545
+ $X2=2.45 $Y2=1.545
r148 50 59 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.835 $Y=1.545
+ $X2=2.985 $Y2=1.545
r149 50 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.835 $Y=1.545
+ $X2=2.535 $Y2=1.545
r150 46 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=1.63
+ $X2=2.45 $Y2=1.545
r151 46 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.45 $Y=1.63 $X2=2.45
+ $Y2=1.83
r152 45 55 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.145 $Y=0.81
+ $X2=2.017 $Y2=0.81
r153 44 57 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.835 $Y=0.81
+ $X2=2.985 $Y2=0.81
r154 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.835 $Y=0.81
+ $X2=2.145 $Y2=0.81
r155 40 55 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.017 $Y=0.725
+ $X2=2.017 $Y2=0.81
r156 40 42 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=2.017 $Y=0.725
+ $X2=2.017 $Y2=0.445
r157 39 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=1.545
+ $X2=1.59 $Y2=1.545
r158 38 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=1.545
+ $X2=2.45 $Y2=1.545
r159 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.365 $Y=1.545
+ $X2=1.675 $Y2=1.545
r160 34 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=1.63
+ $X2=1.59 $Y2=1.545
r161 34 36 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.59 $Y=1.63 $X2=1.59
+ $Y2=1.83
r162 33 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.29 $Y=0.81
+ $X2=1.16 $Y2=0.81
r163 32 55 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.89 $Y=0.81
+ $X2=2.017 $Y2=0.81
r164 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.89 $Y=0.81 $X2=1.29
+ $Y2=0.81
r165 28 53 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.725
+ $X2=1.16 $Y2=0.81
r166 28 30 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.16 $Y=0.725
+ $X2=1.16 $Y2=0.445
r167 27 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=1.545
+ $X2=0.73 $Y2=1.545
r168 26 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.545
+ $X2=1.59 $Y2=1.545
r169 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.505 $Y=1.545
+ $X2=0.815 $Y2=1.545
r170 22 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.63
+ $X2=0.73 $Y2=1.545
r171 22 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.73 $Y=1.63 $X2=0.73
+ $Y2=1.83
r172 20 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=1.545
+ $X2=0.73 $Y2=1.545
r173 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.645 $Y=1.545
+ $X2=0.275 $Y2=1.545
r174 18 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.03 $Y=0.81
+ $X2=1.16 $Y2=0.81
r175 18 19 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.03 $Y=0.81
+ $X2=0.275 $Y2=0.81
r176 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.19 $Y=1.46
+ $X2=0.275 $Y2=1.545
r177 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.19 $Y=0.895
+ $X2=0.275 $Y2=0.81
r178 16 17 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.19 $Y=0.895
+ $X2=0.19 $Y2=1.46
r179 5 48 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=2.31
+ $Y=1.485 $X2=2.45 $Y2=1.83
r180 4 36 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=1.485 $X2=1.59 $Y2=1.83
r181 3 24 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.73 $Y2=1.83
r182 2 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.02 $Y2=0.445
r183 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.16 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%VGND 1 2 3 12 16 20 22 24 29 34
+ 41 42 45 48 51
r45 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r47 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r49 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r50 39 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.465
+ $Y2=0
r51 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.99
+ $Y2=0
r52 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r53 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r54 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r55 35 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=1.59
+ $Y2=0
r56 35 37 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=2.07
+ $Y2=0
r57 34 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.465
+ $Y2=0
r58 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.07
+ $Y2=0
r59 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r60 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r61 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 30 45 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.712
+ $Y2=0
r63 30 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.15
+ $Y2=0
r64 29 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.59
+ $Y2=0
r65 29 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.15
+ $Y2=0
r66 24 45 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.712
+ $Y2=0
r67 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.23
+ $Y2=0
r68 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 18 51 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.085
+ $X2=2.465 $Y2=0
r71 18 20 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0.085
+ $X2=2.465 $Y2=0.39
r72 14 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r73 14 16 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.39
r74 10 45 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0
r75 10 12 11.9151 $w=2.93e-07 $l=3.05e-07 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0.39
r76 3 20 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.235 $X2=2.45 $Y2=0.39
r77 2 16 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.59 $Y2=0.39
r78 1 12 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=0.54
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%VPWR 1 8 9
r42 8 9 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 4 8 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=2.99
+ $Y2=2.72
r44 1 9 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 1 4 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


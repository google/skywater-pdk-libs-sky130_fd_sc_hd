* File: sky130_fd_sc_hd__buf_16.pxi.spice
* Created: Tue Sep  1 18:59:00 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_16%A N_A_M1018_g N_A_M1007_g N_A_M1022_g N_A_M1011_g
+ N_A_M1025_g N_A_M1012_g N_A_M1028_g N_A_M1026_g N_A_M1035_g N_A_M1030_g
+ N_A_M1039_g N_A_M1037_g A A N_A_c_209_n N_A_c_210_n
+ PM_SKY130_FD_SC_HD__BUF_16%A
x_PM_SKY130_FD_SC_HD__BUF_16%A_109_47# N_A_109_47#_M1018_s N_A_109_47#_M1025_s
+ N_A_109_47#_M1035_s N_A_109_47#_M1007_d N_A_109_47#_M1012_d
+ N_A_109_47#_M1030_d N_A_109_47#_M1000_g N_A_109_47#_M1001_g
+ N_A_109_47#_M1005_g N_A_109_47#_M1002_g N_A_109_47#_M1006_g
+ N_A_109_47#_M1003_g N_A_109_47#_M1008_g N_A_109_47#_M1004_g
+ N_A_109_47#_M1010_g N_A_109_47#_M1009_g N_A_109_47#_M1013_g
+ N_A_109_47#_M1014_g N_A_109_47#_M1015_g N_A_109_47#_M1017_g
+ N_A_109_47#_M1016_g N_A_109_47#_M1019_g N_A_109_47#_M1023_g
+ N_A_109_47#_M1020_g N_A_109_47#_M1029_g N_A_109_47#_M1021_g
+ N_A_109_47#_M1031_g N_A_109_47#_M1024_g N_A_109_47#_M1032_g
+ N_A_109_47#_M1027_g N_A_109_47#_M1036_g N_A_109_47#_M1033_g
+ N_A_109_47#_M1040_g N_A_109_47#_M1034_g N_A_109_47#_M1041_g
+ N_A_109_47#_M1038_g N_A_109_47#_M1043_g N_A_109_47#_M1042_g
+ N_A_109_47#_c_388_n N_A_109_47#_c_391_n N_A_109_47#_c_354_n
+ N_A_109_47#_c_355_n N_A_109_47#_c_380_n N_A_109_47#_c_381_n
+ N_A_109_47#_c_410_n N_A_109_47#_c_414_n N_A_109_47#_c_356_n
+ N_A_109_47#_c_382_n N_A_109_47#_c_426_n N_A_109_47#_c_429_n
+ N_A_109_47#_c_357_n N_A_109_47#_c_358_n N_A_109_47#_c_359_n
+ N_A_109_47#_c_360_n N_A_109_47#_c_384_n N_A_109_47#_c_361_n
+ N_A_109_47#_c_385_n N_A_109_47#_c_362_n N_A_109_47#_c_363_n
+ PM_SKY130_FD_SC_HD__BUF_16%A_109_47#
x_PM_SKY130_FD_SC_HD__BUF_16%VPWR N_VPWR_M1007_s N_VPWR_M1011_s N_VPWR_M1026_s
+ N_VPWR_M1037_s N_VPWR_M1002_s N_VPWR_M1004_s N_VPWR_M1014_s N_VPWR_M1019_s
+ N_VPWR_M1021_s N_VPWR_M1027_s N_VPWR_M1034_s N_VPWR_M1042_s N_VPWR_c_786_n
+ N_VPWR_c_787_n N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_791_n
+ N_VPWR_c_792_n N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n N_VPWR_c_796_n
+ N_VPWR_c_797_n N_VPWR_c_798_n N_VPWR_c_799_n N_VPWR_c_800_n N_VPWR_c_801_n
+ N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_805_n N_VPWR_c_806_n
+ N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n
+ N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n
+ N_VPWR_c_817_n N_VPWR_c_818_n VPWR N_VPWR_c_819_n N_VPWR_c_785_n
+ N_VPWR_c_821_n N_VPWR_c_822_n PM_SKY130_FD_SC_HD__BUF_16%VPWR
x_PM_SKY130_FD_SC_HD__BUF_16%X N_X_M1000_s N_X_M1006_s N_X_M1010_s N_X_M1015_s
+ N_X_M1023_s N_X_M1031_s N_X_M1036_s N_X_M1041_s N_X_M1001_d N_X_M1003_d
+ N_X_M1009_d N_X_M1017_d N_X_M1020_d N_X_M1024_d N_X_M1033_d N_X_M1038_d
+ N_X_c_988_n N_X_c_986_n N_X_c_987_n N_X_c_949_n N_X_c_950_n N_X_c_967_n
+ N_X_c_968_n N_X_c_1016_n N_X_c_1018_n N_X_c_1022_n N_X_c_951_n N_X_c_969_n
+ N_X_c_1034_n N_X_c_1036_n N_X_c_1040_n N_X_c_952_n N_X_c_970_n N_X_c_1052_n
+ N_X_c_1056_n N_X_c_953_n N_X_c_971_n N_X_c_1068_n N_X_c_1072_n N_X_c_954_n
+ N_X_c_972_n N_X_c_1084_n N_X_c_1088_n N_X_c_955_n N_X_c_973_n N_X_c_1100_n
+ N_X_c_1104_n N_X_c_956_n N_X_c_974_n N_X_c_1116_n N_X_c_1119_n N_X_c_957_n
+ N_X_c_975_n N_X_c_958_n N_X_c_976_n N_X_c_959_n N_X_c_977_n N_X_c_960_n
+ N_X_c_978_n N_X_c_961_n N_X_c_979_n N_X_c_962_n N_X_c_980_n N_X_c_963_n
+ N_X_c_981_n N_X_c_964_n N_X_c_982_n N_X_c_965_n X X N_X_c_985_n
+ PM_SKY130_FD_SC_HD__BUF_16%X
x_PM_SKY130_FD_SC_HD__BUF_16%VGND N_VGND_M1018_d N_VGND_M1022_d N_VGND_M1028_d
+ N_VGND_M1039_d N_VGND_M1005_d N_VGND_M1008_d N_VGND_M1013_d N_VGND_M1016_d
+ N_VGND_M1029_d N_VGND_M1032_d N_VGND_M1040_d N_VGND_M1043_d N_VGND_c_1297_n
+ N_VGND_c_1298_n N_VGND_c_1299_n N_VGND_c_1300_n N_VGND_c_1301_n
+ N_VGND_c_1302_n N_VGND_c_1303_n N_VGND_c_1304_n N_VGND_c_1305_n
+ N_VGND_c_1306_n N_VGND_c_1307_n N_VGND_c_1308_n N_VGND_c_1309_n
+ N_VGND_c_1310_n N_VGND_c_1311_n N_VGND_c_1312_n N_VGND_c_1313_n
+ N_VGND_c_1314_n N_VGND_c_1315_n N_VGND_c_1316_n N_VGND_c_1317_n
+ N_VGND_c_1318_n N_VGND_c_1319_n N_VGND_c_1320_n N_VGND_c_1321_n
+ N_VGND_c_1322_n N_VGND_c_1323_n N_VGND_c_1324_n N_VGND_c_1325_n
+ N_VGND_c_1326_n N_VGND_c_1327_n N_VGND_c_1328_n N_VGND_c_1329_n VGND
+ N_VGND_c_1330_n N_VGND_c_1331_n N_VGND_c_1332_n N_VGND_c_1333_n
+ PM_SKY130_FD_SC_HD__BUF_16%VGND
cc_1 VNB N_A_M1018_g 0.0237664f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1007_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_A_M1022_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_A_M1011_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB N_A_M1025_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_6 VNB N_A_M1012_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_7 VNB N_A_M1028_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_A_M1026_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB N_A_M1035_g 0.0172827f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=0.56
cc_10 VNB N_A_M1030_g 4.49807e-19 $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_11 VNB N_A_M1039_g 0.017512f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.56
cc_12 VNB N_A_M1037_g 4.62853e-19 $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.985
cc_13 VNB N_A_c_209_n 0.0220589f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=1.16
cc_14 VNB N_A_c_210_n 0.100238f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.16
cc_15 VNB N_A_109_47#_M1000_g 0.0176384f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.295
cc_16 VNB N_A_109_47#_M1001_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.025
cc_17 VNB N_A_109_47#_M1005_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.295
cc_18 VNB N_A_109_47#_M1002_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.025
cc_19 VNB N_A_109_47#_M1006_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.295
cc_20 VNB N_A_109_47#_M1003_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.025
cc_21 VNB N_A_109_47#_M1008_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.295
cc_22 VNB N_A_109_47#_M1004_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_23 VNB N_A_109_47#_M1010_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_24 VNB N_A_109_47#_M1009_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_25 VNB N_A_109_47#_M1013_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.16
cc_26 VNB N_A_109_47#_M1014_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.16
cc_27 VNB N_A_109_47#_M1015_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.175
cc_28 VNB N_A_109_47#_M1017_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=1.175
cc_29 VNB N_A_109_47#_M1016_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_109_47#_M1019_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_109_47#_M1023_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_109_47#_M1020_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_109_47#_M1029_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_109_47#_M1021_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_109_47#_M1031_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_109_47#_M1024_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_109_47#_M1032_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_109_47#_M1027_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_109_47#_M1036_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_109_47#_M1033_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_109_47#_M1040_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_109_47#_M1034_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_109_47#_M1041_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_109_47#_M1038_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_109_47#_M1043_g 0.0211164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_109_47#_M1042_g 5.14212e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_109_47#_c_354_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_109_47#_c_355_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_109_47#_c_356_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_109_47#_c_357_n 0.00356912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_109_47#_c_358_n 5.27693e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_109_47#_c_359_n 0.00639236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_109_47#_c_360_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_109_47#_c_361_n 0.00344553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_109_47#_c_362_n 0.00154098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_109_47#_c_363_n 0.259182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_785_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_X_c_949_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_59 VNB N_X_c_950_n 0.00223017f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_60 VNB N_X_c_951_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.175
cc_61 VNB N_X_c_952_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_X_c_953_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_X_c_954_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_X_c_955_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_X_c_956_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_X_c_957_n 0.00429963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_X_c_958_n 0.00223011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_X_c_959_n 0.00223011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_X_c_960_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_X_c_961_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_X_c_962_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_X_c_963_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_X_c_964_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_X_c_965_n 0.0333467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB X 0.0244967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1297_n 0.0110515f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.295
cc_77 VNB N_VGND_c_1298_n 0.00661728f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_78 VNB N_VGND_c_1299_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.56
cc_79 VNB N_VGND_c_1300_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.985
cc_80 VNB N_VGND_c_1301_n 0.00358349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1302_n 0.00357798f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_82 VNB N_VGND_c_1303_n 0.00357798f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_83 VNB N_VGND_c_1304_n 0.0168382f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.16
cc_84 VNB N_VGND_c_1305_n 0.00358349f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.16
cc_85 VNB N_VGND_c_1306_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.175
cc_86 VNB N_VGND_c_1307_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=1.175
cc_87 VNB N_VGND_c_1308_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1309_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1310_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1311_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1312_n 0.0174747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1313_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1314_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1315_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1316_n 0.0168651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1317_n 0.00323787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1318_n 0.0173761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1319_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1320_n 0.0168382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1321_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1322_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1323_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1324_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1325_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1326_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1327_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1328_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1329_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1330_n 0.0164504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1331_n 0.471029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1332_n 0.00323972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1333_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VPB N_A_M1007_g 0.0264483f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_114 VPB N_A_M1011_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_115 VPB N_A_M1012_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_116 VPB N_A_M1026_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_117 VPB N_A_M1030_g 0.0191652f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_118 VPB N_A_M1037_g 0.0194265f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.985
cc_119 VPB N_A_109_47#_M1001_g 0.0196632f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_120 VPB N_A_109_47#_M1002_g 0.0191654f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.025
cc_121 VPB N_A_109_47#_M1003_g 0.0191843f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.025
cc_122 VPB N_A_109_47#_M1004_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_123 VPB N_A_109_47#_M1009_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_124 VPB N_A_109_47#_M1014_g 0.0191843f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.16
cc_125 VPB N_A_109_47#_M1017_g 0.0191843f $X=-0.19 $Y=1.305 $X2=2.3 $Y2=1.175
cc_126 VPB N_A_109_47#_M1019_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_109_47#_M1020_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_109_47#_M1021_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_109_47#_M1024_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_109_47#_M1027_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_109_47#_M1033_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_109_47#_M1034_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_109_47#_M1038_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_109_47#_M1042_g 0.0234647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_109_47#_c_380_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_109_47#_c_381_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_109_47#_c_382_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_109_47#_c_358_n 0.00304142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_109_47#_c_384_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_109_47#_c_385_n 0.00359185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_786_n 0.0110239f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.295
cc_142 VPB N_VPWR_c_787_n 0.00753744f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_143 VPB N_VPWR_c_788_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.295
cc_144 VPB N_VPWR_c_789_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_145 VPB N_VPWR_c_790_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_146 VPB N_VPWR_c_791_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_147 VPB N_VPWR_c_792_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.16
cc_148 VPB N_VPWR_c_793_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.3 $Y2=1.16
cc_149 VPB N_VPWR_c_794_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.175
cc_150 VPB N_VPWR_c_795_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.075 $Y2=1.175
cc_151 VPB N_VPWR_c_796_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_797_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_798_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_799_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_800_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_801_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_802_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_803_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_804_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_805_n 0.0178722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_806_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_807_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_808_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_809_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_810_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_811_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_812_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_813_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_814_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_815_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_816_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_817_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_818_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_819_n 0.0170604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_785_n 0.0532876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_821_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_822_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_X_c_967_n 0.00218965f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_179 VPB N_X_c_968_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_180 VPB N_X_c_969_n 0.00218965f $X=-0.19 $Y=1.305 $X2=2.075 $Y2=1.175
cc_181 VPB N_X_c_970_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_X_c_971_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_X_c_972_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_X_c_973_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_X_c_974_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_X_c_975_n 0.0049359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_X_c_976_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_X_c_977_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_X_c_978_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_X_c_979_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_X_c_980_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_X_c_981_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_X_c_982_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB X 0.00883532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB X 0.014331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_X_c_985_n 0.0433978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 N_A_M1039_g N_A_109_47#_M1000_g 0.0214679f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_M1037_g N_A_109_47#_M1001_g 0.0214679f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_M1018_g N_A_109_47#_c_388_n 0.00545788f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_M1022_g N_A_109_47#_c_388_n 0.00636826f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_M1025_g N_A_109_47#_c_388_n 5.23702e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_M1007_g N_A_109_47#_c_391_n 0.0095746f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_M1011_g N_A_109_47#_c_391_n 0.0106215f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_M1012_g N_A_109_47#_c_391_n 7.66249e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_M1022_g N_A_109_47#_c_354_n 0.00850187f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_M1025_g N_A_109_47#_c_354_n 0.00850187f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_c_209_n N_A_109_47#_c_354_n 0.0359512f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_c_210_n N_A_109_47#_c_354_n 0.00205431f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_M1018_g N_A_109_47#_c_355_n 0.00251756f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_210 N_A_M1022_g N_A_109_47#_c_355_n 0.00110541f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A_c_209_n N_A_109_47#_c_355_n 0.0265235f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_c_210_n N_A_109_47#_c_355_n 0.00213376f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_M1011_g N_A_109_47#_c_380_n 0.0107189f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_M1012_g N_A_109_47#_c_380_n 0.0107189f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_c_209_n N_A_109_47#_c_380_n 0.0359514f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_c_210_n N_A_109_47#_c_380_n 0.00198252f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_M1007_g N_A_109_47#_c_381_n 0.00276634f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_M1011_g N_A_109_47#_c_381_n 0.00135419f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_c_209_n N_A_109_47#_c_381_n 0.026643f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_c_210_n N_A_109_47#_c_381_n 0.00206439f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_M1022_g N_A_109_47#_c_410_n 5.23702e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_M1025_g N_A_109_47#_c_410_n 0.00636826f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A_M1028_g N_A_109_47#_c_410_n 0.00636826f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_M1035_g N_A_109_47#_c_410_n 5.23702e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A_M1011_g N_A_109_47#_c_414_n 7.66249e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_M1012_g N_A_109_47#_c_414_n 0.0106215f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_M1026_g N_A_109_47#_c_414_n 0.0106215f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_M1030_g N_A_109_47#_c_414_n 7.66249e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_M1028_g N_A_109_47#_c_356_n 0.00850187f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_M1035_g N_A_109_47#_c_356_n 0.00850187f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_c_209_n N_A_109_47#_c_356_n 0.0568321f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_c_210_n N_A_109_47#_c_356_n 0.00205431f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_M1026_g N_A_109_47#_c_382_n 0.0107189f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_M1030_g N_A_109_47#_c_382_n 0.0107189f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_c_209_n N_A_109_47#_c_382_n 0.0568326f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_c_210_n N_A_109_47#_c_382_n 0.00198252f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_M1028_g N_A_109_47#_c_426_n 5.24491e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A_M1035_g N_A_109_47#_c_426_n 0.00647394f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_239 N_A_M1039_g N_A_109_47#_c_426_n 0.00647394f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_240 N_A_M1026_g N_A_109_47#_c_429_n 7.67038e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A_M1030_g N_A_109_47#_c_429_n 0.0107272f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A_M1037_g N_A_109_47#_c_429_n 0.0107272f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_M1039_g N_A_109_47#_c_357_n 0.00417409f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A_c_210_n N_A_109_47#_c_358_n 0.00412038f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_M1025_g N_A_109_47#_c_360_n 0.00110541f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A_M1028_g N_A_109_47#_c_360_n 0.00110541f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A_c_209_n N_A_109_47#_c_360_n 0.0265235f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_c_210_n N_A_109_47#_c_360_n 0.00213376f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A_M1012_g N_A_109_47#_c_384_n 0.00135419f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_M1026_g N_A_109_47#_c_384_n 0.00135419f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A_c_209_n N_A_109_47#_c_384_n 0.026643f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_c_210_n N_A_109_47#_c_384_n 0.00206439f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_M1035_g N_A_109_47#_c_361_n 0.00123754f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_M1039_g N_A_109_47#_c_361_n 0.0110598f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A_c_210_n N_A_109_47#_c_361_n 0.00205431f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_M1030_g N_A_109_47#_c_385_n 0.00139111f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A_M1037_g N_A_109_47#_c_385_n 0.0134729f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_c_210_n N_A_109_47#_c_385_n 0.00198252f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_c_209_n N_A_109_47#_c_362_n 0.015316f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A_c_210_n N_A_109_47#_c_362_n 0.00217042f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_c_210_n N_A_109_47#_c_363_n 0.0214679f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_M1007_g N_VPWR_c_787_n 0.0040429f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_c_209_n N_VPWR_c_787_n 0.0143482f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_M1011_g N_VPWR_c_788_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_M1012_g N_VPWR_c_788_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_M1026_g N_VPWR_c_789_n 0.00146448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A_M1030_g N_VPWR_c_789_n 0.00146448f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A_M1037_g N_VPWR_c_790_n 0.00146448f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_M1007_g N_VPWR_c_801_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_M1011_g N_VPWR_c_801_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_M1012_g N_VPWR_c_803_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_M1026_g N_VPWR_c_803_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_M1030_g N_VPWR_c_805_n 0.00541359f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_M1037_g N_VPWR_c_805_n 0.00541359f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A_M1007_g N_VPWR_c_785_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_M1011_g N_VPWR_c_785_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_M1012_g N_VPWR_c_785_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A_M1026_g N_VPWR_c_785_n 0.00950154f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A_M1030_g N_VPWR_c_785_n 0.00950154f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A_M1037_g N_VPWR_c_785_n 0.00952874f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_M1039_g N_X_c_986_n 4.74777e-19 $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_M1037_g N_X_c_987_n 7.66249e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A_M1018_g N_VGND_c_1298_n 0.00360182f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_c_209_n N_VGND_c_1298_n 0.0143482f $X=2.3 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_M1022_g N_VGND_c_1299_n 0.00146448f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_M1025_g N_VGND_c_1299_n 0.00146448f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_M1028_g N_VGND_c_1300_n 0.00146448f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_M1035_g N_VGND_c_1300_n 0.00146448f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_M1039_g N_VGND_c_1301_n 0.00146448f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_M1018_g N_VGND_c_1312_n 0.00541562f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_M1022_g N_VGND_c_1312_n 0.00424619f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A_M1025_g N_VGND_c_1314_n 0.00424619f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_M1028_g N_VGND_c_1314_n 0.00424619f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A_M1035_g N_VGND_c_1316_n 0.00423644f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_295 N_A_M1039_g N_VGND_c_1316_n 0.00423644f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_296 N_A_M1018_g N_VGND_c_1331_n 0.0104559f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A_M1022_g N_VGND_c_1331_n 0.00573624f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A_M1025_g N_VGND_c_1331_n 0.00573624f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A_M1028_g N_VGND_c_1331_n 0.00573624f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_300 N_A_M1035_g N_VGND_c_1331_n 0.00575105f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A_M1039_g N_VGND_c_1331_n 0.00577825f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_302 N_A_109_47#_c_380_n N_VPWR_M1011_s 0.00185611f $X=1.355 $Y=1.53 $X2=0
+ $Y2=0
cc_303 N_A_109_47#_c_382_n N_VPWR_M1026_s 0.00185611f $X=2.195 $Y=1.53 $X2=0
+ $Y2=0
cc_304 N_A_109_47#_c_385_n N_VPWR_M1037_s 0.00207031f $X=2.777 $Y=1.53 $X2=0
+ $Y2=0
cc_305 N_A_109_47#_c_381_n N_VPWR_c_787_n 0.00863458f $X=0.845 $Y=1.53 $X2=0
+ $Y2=0
cc_306 N_A_109_47#_c_380_n N_VPWR_c_788_n 0.0104788f $X=1.355 $Y=1.53 $X2=0
+ $Y2=0
cc_307 N_A_109_47#_c_382_n N_VPWR_c_789_n 0.0104788f $X=2.195 $Y=1.53 $X2=0
+ $Y2=0
cc_308 N_A_109_47#_M1001_g N_VPWR_c_790_n 0.00146448f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_109_47#_c_385_n N_VPWR_c_790_n 0.0104788f $X=2.777 $Y=1.53 $X2=0
+ $Y2=0
cc_310 N_A_109_47#_M1002_g N_VPWR_c_791_n 0.00146448f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_109_47#_M1003_g N_VPWR_c_791_n 0.00146448f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_109_47#_M1004_g N_VPWR_c_792_n 0.00146448f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_109_47#_M1009_g N_VPWR_c_792_n 0.00146448f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_109_47#_M1009_g N_VPWR_c_793_n 0.00541359f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_109_47#_M1014_g N_VPWR_c_793_n 0.00541359f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_109_47#_M1014_g N_VPWR_c_794_n 0.00146448f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_317 N_A_109_47#_M1017_g N_VPWR_c_794_n 0.00146448f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_109_47#_M1019_g N_VPWR_c_795_n 0.00146448f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_319 N_A_109_47#_M1020_g N_VPWR_c_795_n 0.00146448f $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_320 N_A_109_47#_M1021_g N_VPWR_c_796_n 0.00146448f $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_321 N_A_109_47#_M1024_g N_VPWR_c_796_n 0.00146448f $X=7.19 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A_109_47#_M1027_g N_VPWR_c_797_n 0.00146448f $X=7.61 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_109_47#_M1033_g N_VPWR_c_797_n 0.00146448f $X=8.03 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_109_47#_M1034_g N_VPWR_c_798_n 0.00146448f $X=8.45 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_109_47#_M1038_g N_VPWR_c_798_n 0.00146448f $X=8.87 $Y=1.985 $X2=0
+ $Y2=0
cc_326 N_A_109_47#_M1038_g N_VPWR_c_799_n 0.00541359f $X=8.87 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A_109_47#_M1042_g N_VPWR_c_799_n 0.00541359f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_328 N_A_109_47#_M1042_g N_VPWR_c_800_n 0.00316354f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A_109_47#_c_391_n N_VPWR_c_801_n 0.0189039f $X=0.68 $Y=1.63 $X2=0 $Y2=0
cc_330 N_A_109_47#_c_414_n N_VPWR_c_803_n 0.0189039f $X=1.52 $Y=1.63 $X2=0 $Y2=0
cc_331 N_A_109_47#_c_429_n N_VPWR_c_805_n 0.0189039f $X=2.36 $Y=1.63 $X2=0 $Y2=0
cc_332 N_A_109_47#_M1001_g N_VPWR_c_807_n 0.00541359f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_333 N_A_109_47#_M1002_g N_VPWR_c_807_n 0.00541359f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_A_109_47#_M1003_g N_VPWR_c_809_n 0.00541359f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_109_47#_M1004_g N_VPWR_c_809_n 0.00541359f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_109_47#_M1017_g N_VPWR_c_811_n 0.00541359f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A_109_47#_M1019_g N_VPWR_c_811_n 0.00541359f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_109_47#_M1020_g N_VPWR_c_813_n 0.00541359f $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_109_47#_M1021_g N_VPWR_c_813_n 0.00541359f $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_109_47#_M1024_g N_VPWR_c_815_n 0.00541359f $X=7.19 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_109_47#_M1027_g N_VPWR_c_815_n 0.00541359f $X=7.61 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_109_47#_M1033_g N_VPWR_c_817_n 0.00541359f $X=8.03 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_109_47#_M1034_g N_VPWR_c_817_n 0.00541359f $X=8.45 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_109_47#_M1007_d N_VPWR_c_785_n 0.00215201f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_345 N_A_109_47#_M1012_d N_VPWR_c_785_n 0.00215201f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_346 N_A_109_47#_M1030_d N_VPWR_c_785_n 0.00215201f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_347 N_A_109_47#_M1001_g N_VPWR_c_785_n 0.00952874f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_A_109_47#_M1002_g N_VPWR_c_785_n 0.00950154f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_109_47#_M1003_g N_VPWR_c_785_n 0.00950154f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A_109_47#_M1004_g N_VPWR_c_785_n 0.00950154f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A_109_47#_M1009_g N_VPWR_c_785_n 0.00950154f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_109_47#_M1014_g N_VPWR_c_785_n 0.00950154f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A_109_47#_M1017_g N_VPWR_c_785_n 0.00950154f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_109_47#_M1019_g N_VPWR_c_785_n 0.00950154f $X=5.93 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_109_47#_M1020_g N_VPWR_c_785_n 0.00950154f $X=6.35 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A_109_47#_M1021_g N_VPWR_c_785_n 0.00950154f $X=6.77 $Y=1.985 $X2=0
+ $Y2=0
cc_357 N_A_109_47#_M1024_g N_VPWR_c_785_n 0.00950154f $X=7.19 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A_109_47#_M1027_g N_VPWR_c_785_n 0.00950154f $X=7.61 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A_109_47#_M1033_g N_VPWR_c_785_n 0.00950154f $X=8.03 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_109_47#_M1034_g N_VPWR_c_785_n 0.00950154f $X=8.45 $Y=1.985 $X2=0
+ $Y2=0
cc_361 N_A_109_47#_M1038_g N_VPWR_c_785_n 0.00950154f $X=8.87 $Y=1.985 $X2=0
+ $Y2=0
cc_362 N_A_109_47#_M1042_g N_VPWR_c_785_n 0.0108276f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_363 N_A_109_47#_c_391_n N_VPWR_c_785_n 0.0122217f $X=0.68 $Y=1.63 $X2=0 $Y2=0
cc_364 N_A_109_47#_c_414_n N_VPWR_c_785_n 0.0122217f $X=1.52 $Y=1.63 $X2=0 $Y2=0
cc_365 N_A_109_47#_c_429_n N_VPWR_c_785_n 0.0122217f $X=2.36 $Y=1.63 $X2=0 $Y2=0
cc_366 N_A_109_47#_M1000_g N_X_c_988_n 0.00202914f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A_109_47#_M1005_g N_X_c_988_n 0.00198339f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_109_47#_M1000_g N_X_c_986_n 0.00439074f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_369 N_A_109_47#_M1005_g N_X_c_986_n 0.00439074f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_109_47#_M1006_g N_X_c_986_n 4.74777e-19 $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_109_47#_c_426_n N_X_c_986_n 0.00518536f $X=2.36 $Y=0.4 $X2=0 $Y2=0
cc_372 N_A_109_47#_M1001_g N_X_c_987_n 0.0106215f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_373 N_A_109_47#_M1002_g N_X_c_987_n 0.0106215f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A_109_47#_M1003_g N_X_c_987_n 7.66249e-19 $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A_109_47#_c_429_n N_X_c_987_n 0.00671496f $X=2.36 $Y=1.63 $X2=0 $Y2=0
cc_376 N_A_109_47#_M1005_g N_X_c_949_n 0.00850187f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A_109_47#_M1006_g N_X_c_949_n 0.00850187f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_378 N_A_109_47#_c_359_n N_X_c_949_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_109_47#_c_363_n N_X_c_949_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_380 N_A_109_47#_M1000_g N_X_c_950_n 0.00241717f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_381 N_A_109_47#_M1005_g N_X_c_950_n 0.0011083f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_382 N_A_109_47#_c_359_n N_X_c_950_n 0.0265361f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_109_47#_c_361_n N_X_c_950_n 0.00795337f $X=2.777 $Y=0.82 $X2=0 $Y2=0
cc_384 N_A_109_47#_c_363_n N_X_c_950_n 0.00213429f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A_109_47#_M1002_g N_X_c_967_n 0.0107189f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_386 N_A_109_47#_M1003_g N_X_c_967_n 0.0107189f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_387 N_A_109_47#_c_359_n N_X_c_967_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_388 N_A_109_47#_c_363_n N_X_c_967_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_109_47#_M1001_g N_X_c_968_n 0.00265135f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_390 N_A_109_47#_M1002_g N_X_c_968_n 0.00134262f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A_109_47#_c_359_n N_X_c_968_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_392 N_A_109_47#_c_385_n N_X_c_968_n 0.0088897f $X=2.777 $Y=1.53 $X2=0 $Y2=0
cc_393 N_A_109_47#_c_363_n N_X_c_968_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_394 N_A_109_47#_M1006_g N_X_c_1016_n 0.00198339f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_395 N_A_109_47#_M1008_g N_X_c_1016_n 0.00198339f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_396 N_A_109_47#_M1005_g N_X_c_1018_n 4.74777e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_397 N_A_109_47#_M1006_g N_X_c_1018_n 0.00439074f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_398 N_A_109_47#_M1008_g N_X_c_1018_n 0.00439074f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_399 N_A_109_47#_M1010_g N_X_c_1018_n 4.74777e-19 $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_400 N_A_109_47#_M1002_g N_X_c_1022_n 7.66249e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A_109_47#_M1003_g N_X_c_1022_n 0.0106215f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A_109_47#_M1004_g N_X_c_1022_n 0.0106215f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_403 N_A_109_47#_M1009_g N_X_c_1022_n 7.66249e-19 $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_404 N_A_109_47#_M1008_g N_X_c_951_n 0.00850187f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_405 N_A_109_47#_M1010_g N_X_c_951_n 0.00850187f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_406 N_A_109_47#_c_359_n N_X_c_951_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_407 N_A_109_47#_c_363_n N_X_c_951_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_408 N_A_109_47#_M1004_g N_X_c_969_n 0.0107189f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_409 N_A_109_47#_M1009_g N_X_c_969_n 0.0107189f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_410 N_A_109_47#_c_359_n N_X_c_969_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_411 N_A_109_47#_c_363_n N_X_c_969_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_412 N_A_109_47#_M1010_g N_X_c_1034_n 0.00198339f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A_109_47#_M1013_g N_X_c_1034_n 0.00198339f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_414 N_A_109_47#_M1008_g N_X_c_1036_n 4.74777e-19 $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_415 N_A_109_47#_M1010_g N_X_c_1036_n 0.00439074f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_416 N_A_109_47#_M1013_g N_X_c_1036_n 0.00439074f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_417 N_A_109_47#_M1015_g N_X_c_1036_n 4.74777e-19 $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_418 N_A_109_47#_M1004_g N_X_c_1040_n 7.66249e-19 $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_419 N_A_109_47#_M1009_g N_X_c_1040_n 0.0106215f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_420 N_A_109_47#_M1014_g N_X_c_1040_n 0.0106215f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_421 N_A_109_47#_M1017_g N_X_c_1040_n 7.66249e-19 $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_422 N_A_109_47#_M1013_g N_X_c_952_n 0.00850187f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A_109_47#_M1015_g N_X_c_952_n 0.00850187f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_424 N_A_109_47#_c_359_n N_X_c_952_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_425 N_A_109_47#_c_363_n N_X_c_952_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_426 N_A_109_47#_M1014_g N_X_c_970_n 0.0107189f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_427 N_A_109_47#_M1017_g N_X_c_970_n 0.0107189f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_428 N_A_109_47#_c_359_n N_X_c_970_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_429 N_A_109_47#_c_363_n N_X_c_970_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_430 N_A_109_47#_M1013_g N_X_c_1052_n 5.23702e-19 $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_431 N_A_109_47#_M1015_g N_X_c_1052_n 0.00636826f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_432 N_A_109_47#_M1016_g N_X_c_1052_n 0.00636826f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_433 N_A_109_47#_M1023_g N_X_c_1052_n 5.23702e-19 $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_434 N_A_109_47#_M1014_g N_X_c_1056_n 7.66249e-19 $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_435 N_A_109_47#_M1017_g N_X_c_1056_n 0.0106215f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_436 N_A_109_47#_M1019_g N_X_c_1056_n 0.0106215f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_437 N_A_109_47#_M1020_g N_X_c_1056_n 7.66249e-19 $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_438 N_A_109_47#_M1016_g N_X_c_953_n 0.00850187f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A_109_47#_M1023_g N_X_c_953_n 0.00850187f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A_109_47#_c_359_n N_X_c_953_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_441 N_A_109_47#_c_363_n N_X_c_953_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_442 N_A_109_47#_M1019_g N_X_c_971_n 0.0107189f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_443 N_A_109_47#_M1020_g N_X_c_971_n 0.0107189f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_444 N_A_109_47#_c_359_n N_X_c_971_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_445 N_A_109_47#_c_363_n N_X_c_971_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_109_47#_M1016_g N_X_c_1068_n 5.23702e-19 $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_447 N_A_109_47#_M1023_g N_X_c_1068_n 0.00636826f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_448 N_A_109_47#_M1029_g N_X_c_1068_n 0.00636826f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_449 N_A_109_47#_M1031_g N_X_c_1068_n 5.23702e-19 $X=7.19 $Y=0.56 $X2=0 $Y2=0
cc_450 N_A_109_47#_M1019_g N_X_c_1072_n 7.66249e-19 $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_451 N_A_109_47#_M1020_g N_X_c_1072_n 0.0106215f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_452 N_A_109_47#_M1021_g N_X_c_1072_n 0.0106215f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_453 N_A_109_47#_M1024_g N_X_c_1072_n 7.66249e-19 $X=7.19 $Y=1.985 $X2=0 $Y2=0
cc_454 N_A_109_47#_M1029_g N_X_c_954_n 0.00850187f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_455 N_A_109_47#_M1031_g N_X_c_954_n 0.00850187f $X=7.19 $Y=0.56 $X2=0 $Y2=0
cc_456 N_A_109_47#_c_359_n N_X_c_954_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_109_47#_c_363_n N_X_c_954_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_458 N_A_109_47#_M1021_g N_X_c_972_n 0.0107189f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_459 N_A_109_47#_M1024_g N_X_c_972_n 0.0107189f $X=7.19 $Y=1.985 $X2=0 $Y2=0
cc_460 N_A_109_47#_c_359_n N_X_c_972_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_461 N_A_109_47#_c_363_n N_X_c_972_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_109_47#_M1029_g N_X_c_1084_n 5.23702e-19 $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_463 N_A_109_47#_M1031_g N_X_c_1084_n 0.00636826f $X=7.19 $Y=0.56 $X2=0 $Y2=0
cc_464 N_A_109_47#_M1032_g N_X_c_1084_n 0.00636826f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_465 N_A_109_47#_M1036_g N_X_c_1084_n 5.23702e-19 $X=8.03 $Y=0.56 $X2=0 $Y2=0
cc_466 N_A_109_47#_M1021_g N_X_c_1088_n 7.66249e-19 $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_467 N_A_109_47#_M1024_g N_X_c_1088_n 0.0106215f $X=7.19 $Y=1.985 $X2=0 $Y2=0
cc_468 N_A_109_47#_M1027_g N_X_c_1088_n 0.0106215f $X=7.61 $Y=1.985 $X2=0 $Y2=0
cc_469 N_A_109_47#_M1033_g N_X_c_1088_n 7.66249e-19 $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_470 N_A_109_47#_M1032_g N_X_c_955_n 0.00850187f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_471 N_A_109_47#_M1036_g N_X_c_955_n 0.00850187f $X=8.03 $Y=0.56 $X2=0 $Y2=0
cc_472 N_A_109_47#_c_359_n N_X_c_955_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_473 N_A_109_47#_c_363_n N_X_c_955_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_474 N_A_109_47#_M1027_g N_X_c_973_n 0.0107189f $X=7.61 $Y=1.985 $X2=0 $Y2=0
cc_475 N_A_109_47#_M1033_g N_X_c_973_n 0.0107189f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_476 N_A_109_47#_c_359_n N_X_c_973_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_477 N_A_109_47#_c_363_n N_X_c_973_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_478 N_A_109_47#_M1032_g N_X_c_1100_n 5.23702e-19 $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_479 N_A_109_47#_M1036_g N_X_c_1100_n 0.00636826f $X=8.03 $Y=0.56 $X2=0 $Y2=0
cc_480 N_A_109_47#_M1040_g N_X_c_1100_n 0.00636826f $X=8.45 $Y=0.56 $X2=0 $Y2=0
cc_481 N_A_109_47#_M1041_g N_X_c_1100_n 5.23702e-19 $X=8.87 $Y=0.56 $X2=0 $Y2=0
cc_482 N_A_109_47#_M1027_g N_X_c_1104_n 7.66249e-19 $X=7.61 $Y=1.985 $X2=0 $Y2=0
cc_483 N_A_109_47#_M1033_g N_X_c_1104_n 0.0106215f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_484 N_A_109_47#_M1034_g N_X_c_1104_n 0.0106215f $X=8.45 $Y=1.985 $X2=0 $Y2=0
cc_485 N_A_109_47#_M1038_g N_X_c_1104_n 7.66249e-19 $X=8.87 $Y=1.985 $X2=0 $Y2=0
cc_486 N_A_109_47#_M1040_g N_X_c_956_n 0.00850187f $X=8.45 $Y=0.56 $X2=0 $Y2=0
cc_487 N_A_109_47#_M1041_g N_X_c_956_n 0.00850187f $X=8.87 $Y=0.56 $X2=0 $Y2=0
cc_488 N_A_109_47#_c_359_n N_X_c_956_n 0.0359512f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_489 N_A_109_47#_c_363_n N_X_c_956_n 0.00205431f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_490 N_A_109_47#_M1034_g N_X_c_974_n 0.0107189f $X=8.45 $Y=1.985 $X2=0 $Y2=0
cc_491 N_A_109_47#_M1038_g N_X_c_974_n 0.0107189f $X=8.87 $Y=1.985 $X2=0 $Y2=0
cc_492 N_A_109_47#_c_359_n N_X_c_974_n 0.0359514f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_493 N_A_109_47#_c_363_n N_X_c_974_n 0.00198252f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_494 N_A_109_47#_M1040_g N_X_c_1116_n 5.23702e-19 $X=8.45 $Y=0.56 $X2=0 $Y2=0
cc_495 N_A_109_47#_M1041_g N_X_c_1116_n 0.00636826f $X=8.87 $Y=0.56 $X2=0 $Y2=0
cc_496 N_A_109_47#_M1043_g N_X_c_1116_n 0.0068957f $X=9.29 $Y=0.56 $X2=0 $Y2=0
cc_497 N_A_109_47#_M1034_g N_X_c_1119_n 7.66249e-19 $X=8.45 $Y=1.985 $X2=0 $Y2=0
cc_498 N_A_109_47#_M1038_g N_X_c_1119_n 0.0106215f $X=8.87 $Y=1.985 $X2=0 $Y2=0
cc_499 N_A_109_47#_M1042_g N_X_c_1119_n 0.011433f $X=9.29 $Y=1.985 $X2=0 $Y2=0
cc_500 N_A_109_47#_M1043_g N_X_c_957_n 0.0105322f $X=9.29 $Y=0.56 $X2=0 $Y2=0
cc_501 N_A_109_47#_c_359_n N_X_c_957_n 0.0116336f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_502 N_A_109_47#_M1042_g N_X_c_975_n 0.0127492f $X=9.29 $Y=1.985 $X2=0 $Y2=0
cc_503 N_A_109_47#_c_359_n N_X_c_975_n 0.0116336f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_504 N_A_109_47#_M1006_g N_X_c_958_n 0.00111988f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_505 N_A_109_47#_M1008_g N_X_c_958_n 0.00111988f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_506 N_A_109_47#_c_359_n N_X_c_958_n 0.0265319f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_507 N_A_109_47#_c_363_n N_X_c_958_n 0.00213429f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_508 N_A_109_47#_M1003_g N_X_c_976_n 0.00135419f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_509 N_A_109_47#_M1004_g N_X_c_976_n 0.00135419f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_510 N_A_109_47#_c_359_n N_X_c_976_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_511 N_A_109_47#_c_363_n N_X_c_976_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_512 N_A_109_47#_M1010_g N_X_c_959_n 0.00111988f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_513 N_A_109_47#_M1013_g N_X_c_959_n 0.00111988f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_514 N_A_109_47#_c_359_n N_X_c_959_n 0.0265319f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_515 N_A_109_47#_c_363_n N_X_c_959_n 0.00213429f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_516 N_A_109_47#_M1009_g N_X_c_977_n 0.00135419f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_517 N_A_109_47#_M1014_g N_X_c_977_n 0.00135419f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_518 N_A_109_47#_c_359_n N_X_c_977_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_519 N_A_109_47#_c_363_n N_X_c_977_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_520 N_A_109_47#_M1015_g N_X_c_960_n 0.00110541f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_521 N_A_109_47#_M1016_g N_X_c_960_n 0.00110541f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_522 N_A_109_47#_c_359_n N_X_c_960_n 0.0265235f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_523 N_A_109_47#_c_363_n N_X_c_960_n 0.00213376f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_524 N_A_109_47#_M1017_g N_X_c_978_n 0.00135419f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_525 N_A_109_47#_M1019_g N_X_c_978_n 0.00135419f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_526 N_A_109_47#_c_359_n N_X_c_978_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_527 N_A_109_47#_c_363_n N_X_c_978_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_528 N_A_109_47#_M1023_g N_X_c_961_n 0.00110541f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_529 N_A_109_47#_M1029_g N_X_c_961_n 0.00110541f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_530 N_A_109_47#_c_359_n N_X_c_961_n 0.0265235f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_531 N_A_109_47#_c_363_n N_X_c_961_n 0.00213376f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_532 N_A_109_47#_M1020_g N_X_c_979_n 0.00135419f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_533 N_A_109_47#_M1021_g N_X_c_979_n 0.00135419f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_534 N_A_109_47#_c_359_n N_X_c_979_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_535 N_A_109_47#_c_363_n N_X_c_979_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_536 N_A_109_47#_M1031_g N_X_c_962_n 0.00110541f $X=7.19 $Y=0.56 $X2=0 $Y2=0
cc_537 N_A_109_47#_M1032_g N_X_c_962_n 0.00110541f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_538 N_A_109_47#_c_359_n N_X_c_962_n 0.0265235f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_539 N_A_109_47#_c_363_n N_X_c_962_n 0.00213376f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_540 N_A_109_47#_M1024_g N_X_c_980_n 0.00135419f $X=7.19 $Y=1.985 $X2=0 $Y2=0
cc_541 N_A_109_47#_M1027_g N_X_c_980_n 0.00135419f $X=7.61 $Y=1.985 $X2=0 $Y2=0
cc_542 N_A_109_47#_c_359_n N_X_c_980_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_543 N_A_109_47#_c_363_n N_X_c_980_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_544 N_A_109_47#_M1036_g N_X_c_963_n 0.00110541f $X=8.03 $Y=0.56 $X2=0 $Y2=0
cc_545 N_A_109_47#_M1040_g N_X_c_963_n 0.00110541f $X=8.45 $Y=0.56 $X2=0 $Y2=0
cc_546 N_A_109_47#_c_359_n N_X_c_963_n 0.0265235f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_547 N_A_109_47#_c_363_n N_X_c_963_n 0.00213376f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_548 N_A_109_47#_M1033_g N_X_c_981_n 0.00135419f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_549 N_A_109_47#_M1034_g N_X_c_981_n 0.00135419f $X=8.45 $Y=1.985 $X2=0 $Y2=0
cc_550 N_A_109_47#_c_359_n N_X_c_981_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_551 N_A_109_47#_c_363_n N_X_c_981_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_552 N_A_109_47#_M1041_g N_X_c_964_n 0.00110541f $X=8.87 $Y=0.56 $X2=0 $Y2=0
cc_553 N_A_109_47#_M1043_g N_X_c_964_n 0.00110541f $X=9.29 $Y=0.56 $X2=0 $Y2=0
cc_554 N_A_109_47#_c_359_n N_X_c_964_n 0.0265235f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_555 N_A_109_47#_c_363_n N_X_c_964_n 0.00213376f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_556 N_A_109_47#_M1038_g N_X_c_982_n 0.00135419f $X=8.87 $Y=1.985 $X2=0 $Y2=0
cc_557 N_A_109_47#_M1042_g N_X_c_982_n 0.00135419f $X=9.29 $Y=1.985 $X2=0 $Y2=0
cc_558 N_A_109_47#_c_359_n N_X_c_982_n 0.026643f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_559 N_A_109_47#_c_363_n N_X_c_982_n 0.00206439f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_560 N_A_109_47#_M1043_g N_X_c_965_n 0.00292435f $X=9.29 $Y=0.56 $X2=0 $Y2=0
cc_561 N_A_109_47#_M1043_g X 0.00597224f $X=9.29 $Y=0.56 $X2=0 $Y2=0
cc_562 N_A_109_47#_c_359_n X 0.0136932f $X=9.22 $Y=1.16 $X2=0 $Y2=0
cc_563 N_A_109_47#_c_363_n X 0.00703263f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_564 N_A_109_47#_M1042_g N_X_c_985_n 0.00432902f $X=9.29 $Y=1.985 $X2=0 $Y2=0
cc_565 N_A_109_47#_c_354_n N_VGND_M1022_d 0.00162006f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_566 N_A_109_47#_c_356_n N_VGND_M1028_d 0.00162006f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_567 N_A_109_47#_c_361_n N_VGND_M1039_d 0.00186748f $X=2.777 $Y=0.82 $X2=0
+ $Y2=0
cc_568 N_A_109_47#_c_355_n N_VGND_c_1298_n 0.00787895f $X=0.845 $Y=0.82 $X2=0
+ $Y2=0
cc_569 N_A_109_47#_c_354_n N_VGND_c_1299_n 0.0122414f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_570 N_A_109_47#_c_356_n N_VGND_c_1300_n 0.0122414f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_571 N_A_109_47#_M1000_g N_VGND_c_1301_n 0.00146448f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_572 N_A_109_47#_c_361_n N_VGND_c_1301_n 0.0122414f $X=2.777 $Y=0.82 $X2=0
+ $Y2=0
cc_573 N_A_109_47#_M1005_g N_VGND_c_1302_n 0.00146448f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_574 N_A_109_47#_M1006_g N_VGND_c_1302_n 0.00146448f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_575 N_A_109_47#_M1008_g N_VGND_c_1303_n 0.00146448f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_576 N_A_109_47#_M1010_g N_VGND_c_1303_n 0.00146448f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_577 N_A_109_47#_M1010_g N_VGND_c_1304_n 0.00423108f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_578 N_A_109_47#_M1013_g N_VGND_c_1304_n 0.00423108f $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_579 N_A_109_47#_M1013_g N_VGND_c_1305_n 0.00146448f $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_580 N_A_109_47#_M1015_g N_VGND_c_1305_n 0.00146448f $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_581 N_A_109_47#_M1016_g N_VGND_c_1306_n 0.00146448f $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_582 N_A_109_47#_M1023_g N_VGND_c_1306_n 0.00146448f $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_583 N_A_109_47#_M1029_g N_VGND_c_1307_n 0.00146448f $X=6.77 $Y=0.56 $X2=0
+ $Y2=0
cc_584 N_A_109_47#_M1031_g N_VGND_c_1307_n 0.00146448f $X=7.19 $Y=0.56 $X2=0
+ $Y2=0
cc_585 N_A_109_47#_M1032_g N_VGND_c_1308_n 0.00146448f $X=7.61 $Y=0.56 $X2=0
+ $Y2=0
cc_586 N_A_109_47#_M1036_g N_VGND_c_1308_n 0.00146448f $X=8.03 $Y=0.56 $X2=0
+ $Y2=0
cc_587 N_A_109_47#_M1040_g N_VGND_c_1309_n 0.00146448f $X=8.45 $Y=0.56 $X2=0
+ $Y2=0
cc_588 N_A_109_47#_M1041_g N_VGND_c_1309_n 0.00146448f $X=8.87 $Y=0.56 $X2=0
+ $Y2=0
cc_589 N_A_109_47#_M1041_g N_VGND_c_1310_n 0.00424619f $X=8.87 $Y=0.56 $X2=0
+ $Y2=0
cc_590 N_A_109_47#_M1043_g N_VGND_c_1310_n 0.00424619f $X=9.29 $Y=0.56 $X2=0
+ $Y2=0
cc_591 N_A_109_47#_M1043_g N_VGND_c_1311_n 0.00316354f $X=9.29 $Y=0.56 $X2=0
+ $Y2=0
cc_592 N_A_109_47#_c_388_n N_VGND_c_1312_n 0.0182681f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_593 N_A_109_47#_c_354_n N_VGND_c_1312_n 0.00193763f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_594 N_A_109_47#_c_354_n N_VGND_c_1314_n 0.00193763f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_595 N_A_109_47#_c_410_n N_VGND_c_1314_n 0.0182681f $X=1.52 $Y=0.4 $X2=0 $Y2=0
cc_596 N_A_109_47#_c_356_n N_VGND_c_1314_n 0.00193763f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_597 N_A_109_47#_c_356_n N_VGND_c_1316_n 0.00390702f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_598 N_A_109_47#_c_426_n N_VGND_c_1316_n 0.0179571f $X=2.36 $Y=0.4 $X2=0 $Y2=0
cc_599 N_A_109_47#_M1000_g N_VGND_c_1318_n 0.00539841f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_600 N_A_109_47#_M1005_g N_VGND_c_1318_n 0.00423108f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_601 N_A_109_47#_M1006_g N_VGND_c_1320_n 0.00423108f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_602 N_A_109_47#_M1008_g N_VGND_c_1320_n 0.00423108f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_603 N_A_109_47#_M1015_g N_VGND_c_1322_n 0.00424619f $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_604 N_A_109_47#_M1016_g N_VGND_c_1322_n 0.00424619f $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_605 N_A_109_47#_M1023_g N_VGND_c_1324_n 0.00424619f $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_606 N_A_109_47#_M1029_g N_VGND_c_1324_n 0.00424619f $X=6.77 $Y=0.56 $X2=0
+ $Y2=0
cc_607 N_A_109_47#_M1031_g N_VGND_c_1326_n 0.00424619f $X=7.19 $Y=0.56 $X2=0
+ $Y2=0
cc_608 N_A_109_47#_M1032_g N_VGND_c_1326_n 0.00424619f $X=7.61 $Y=0.56 $X2=0
+ $Y2=0
cc_609 N_A_109_47#_M1036_g N_VGND_c_1328_n 0.00424619f $X=8.03 $Y=0.56 $X2=0
+ $Y2=0
cc_610 N_A_109_47#_M1040_g N_VGND_c_1328_n 0.00424619f $X=8.45 $Y=0.56 $X2=0
+ $Y2=0
cc_611 N_A_109_47#_M1018_s N_VGND_c_1331_n 0.00215347f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_612 N_A_109_47#_M1025_s N_VGND_c_1331_n 0.00215347f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_613 N_A_109_47#_M1035_s N_VGND_c_1331_n 0.00215347f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_614 N_A_109_47#_M1000_g N_VGND_c_1331_n 0.00949176f $X=2.99 $Y=0.56 $X2=0
+ $Y2=0
cc_615 N_A_109_47#_M1005_g N_VGND_c_1331_n 0.00574532f $X=3.41 $Y=0.56 $X2=0
+ $Y2=0
cc_616 N_A_109_47#_M1006_g N_VGND_c_1331_n 0.00574532f $X=3.83 $Y=0.56 $X2=0
+ $Y2=0
cc_617 N_A_109_47#_M1008_g N_VGND_c_1331_n 0.00574532f $X=4.25 $Y=0.56 $X2=0
+ $Y2=0
cc_618 N_A_109_47#_M1010_g N_VGND_c_1331_n 0.00574532f $X=4.67 $Y=0.56 $X2=0
+ $Y2=0
cc_619 N_A_109_47#_M1013_g N_VGND_c_1331_n 0.00574532f $X=5.09 $Y=0.56 $X2=0
+ $Y2=0
cc_620 N_A_109_47#_M1015_g N_VGND_c_1331_n 0.00573624f $X=5.51 $Y=0.56 $X2=0
+ $Y2=0
cc_621 N_A_109_47#_M1016_g N_VGND_c_1331_n 0.00573624f $X=5.93 $Y=0.56 $X2=0
+ $Y2=0
cc_622 N_A_109_47#_M1023_g N_VGND_c_1331_n 0.00573624f $X=6.35 $Y=0.56 $X2=0
+ $Y2=0
cc_623 N_A_109_47#_M1029_g N_VGND_c_1331_n 0.00573624f $X=6.77 $Y=0.56 $X2=0
+ $Y2=0
cc_624 N_A_109_47#_M1031_g N_VGND_c_1331_n 0.00573624f $X=7.19 $Y=0.56 $X2=0
+ $Y2=0
cc_625 N_A_109_47#_M1032_g N_VGND_c_1331_n 0.00573624f $X=7.61 $Y=0.56 $X2=0
+ $Y2=0
cc_626 N_A_109_47#_M1036_g N_VGND_c_1331_n 0.00573624f $X=8.03 $Y=0.56 $X2=0
+ $Y2=0
cc_627 N_A_109_47#_M1040_g N_VGND_c_1331_n 0.00573624f $X=8.45 $Y=0.56 $X2=0
+ $Y2=0
cc_628 N_A_109_47#_M1041_g N_VGND_c_1331_n 0.00573624f $X=8.87 $Y=0.56 $X2=0
+ $Y2=0
cc_629 N_A_109_47#_M1043_g N_VGND_c_1331_n 0.00706231f $X=9.29 $Y=0.56 $X2=0
+ $Y2=0
cc_630 N_A_109_47#_c_388_n N_VGND_c_1331_n 0.0121741f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_631 N_A_109_47#_c_354_n N_VGND_c_1331_n 0.00825759f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_632 N_A_109_47#_c_410_n N_VGND_c_1331_n 0.0121741f $X=1.52 $Y=0.4 $X2=0 $Y2=0
cc_633 N_A_109_47#_c_356_n N_VGND_c_1331_n 0.012122f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_634 N_A_109_47#_c_426_n N_VGND_c_1331_n 0.0120759f $X=2.36 $Y=0.4 $X2=0 $Y2=0
cc_635 N_A_109_47#_c_361_n N_VGND_c_1331_n 6.28727e-19 $X=2.777 $Y=0.82 $X2=0
+ $Y2=0
cc_636 N_VPWR_c_785_n N_X_M1001_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_637 N_VPWR_c_785_n N_X_M1003_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_638 N_VPWR_c_785_n N_X_M1009_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_639 N_VPWR_c_785_n N_X_M1017_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_640 N_VPWR_c_785_n N_X_M1020_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_641 N_VPWR_c_785_n N_X_M1024_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_642 N_VPWR_c_785_n N_X_M1033_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_643 N_VPWR_c_785_n N_X_M1038_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_644 N_VPWR_c_807_n N_X_c_987_n 0.0189039f $X=3.535 $Y=2.72 $X2=0 $Y2=0
cc_645 N_VPWR_c_785_n N_X_c_987_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_646 N_VPWR_M1002_s N_X_c_967_n 0.00185611f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_647 N_VPWR_c_791_n N_X_c_967_n 0.0104788f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_648 N_VPWR_c_809_n N_X_c_1022_n 0.0189039f $X=4.375 $Y=2.72 $X2=0 $Y2=0
cc_649 N_VPWR_c_785_n N_X_c_1022_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_650 N_VPWR_M1004_s N_X_c_969_n 0.00185611f $X=4.325 $Y=1.485 $X2=0 $Y2=0
cc_651 N_VPWR_c_792_n N_X_c_969_n 0.0104788f $X=4.46 $Y=2 $X2=0 $Y2=0
cc_652 N_VPWR_c_793_n N_X_c_1040_n 0.0189039f $X=5.215 $Y=2.72 $X2=0 $Y2=0
cc_653 N_VPWR_c_785_n N_X_c_1040_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_654 N_VPWR_M1014_s N_X_c_970_n 0.00185611f $X=5.165 $Y=1.485 $X2=0 $Y2=0
cc_655 N_VPWR_c_794_n N_X_c_970_n 0.0104788f $X=5.3 $Y=2 $X2=0 $Y2=0
cc_656 N_VPWR_c_811_n N_X_c_1056_n 0.0189039f $X=6.055 $Y=2.72 $X2=0 $Y2=0
cc_657 N_VPWR_c_785_n N_X_c_1056_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_658 N_VPWR_M1019_s N_X_c_971_n 0.00185611f $X=6.005 $Y=1.485 $X2=0 $Y2=0
cc_659 N_VPWR_c_795_n N_X_c_971_n 0.0104788f $X=6.14 $Y=2 $X2=0 $Y2=0
cc_660 N_VPWR_c_813_n N_X_c_1072_n 0.0189039f $X=6.895 $Y=2.72 $X2=0 $Y2=0
cc_661 N_VPWR_c_785_n N_X_c_1072_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_662 N_VPWR_M1021_s N_X_c_972_n 0.00185611f $X=6.845 $Y=1.485 $X2=0 $Y2=0
cc_663 N_VPWR_c_796_n N_X_c_972_n 0.0104788f $X=6.98 $Y=2 $X2=0 $Y2=0
cc_664 N_VPWR_c_815_n N_X_c_1088_n 0.0189039f $X=7.735 $Y=2.72 $X2=0 $Y2=0
cc_665 N_VPWR_c_785_n N_X_c_1088_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_666 N_VPWR_M1027_s N_X_c_973_n 0.00185611f $X=7.685 $Y=1.485 $X2=0 $Y2=0
cc_667 N_VPWR_c_797_n N_X_c_973_n 0.0104788f $X=7.82 $Y=2 $X2=0 $Y2=0
cc_668 N_VPWR_c_817_n N_X_c_1104_n 0.0189039f $X=8.575 $Y=2.72 $X2=0 $Y2=0
cc_669 N_VPWR_c_785_n N_X_c_1104_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_670 N_VPWR_M1034_s N_X_c_974_n 0.00185611f $X=8.525 $Y=1.485 $X2=0 $Y2=0
cc_671 N_VPWR_c_798_n N_X_c_974_n 0.0104788f $X=8.66 $Y=2 $X2=0 $Y2=0
cc_672 N_VPWR_c_799_n N_X_c_1119_n 0.0189039f $X=9.415 $Y=2.72 $X2=0 $Y2=0
cc_673 N_VPWR_c_785_n N_X_c_1119_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_674 N_VPWR_M1042_s N_X_c_975_n 0.00406309f $X=9.365 $Y=1.485 $X2=0 $Y2=0
cc_675 N_VPWR_c_800_n N_X_c_975_n 0.0108818f $X=9.5 $Y=2 $X2=0 $Y2=0
cc_676 N_VPWR_c_800_n N_X_c_985_n 0.0396024f $X=9.5 $Y=2 $X2=0 $Y2=0
cc_677 N_VPWR_c_819_n N_X_c_985_n 0.0117463f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_678 N_VPWR_c_785_n N_X_c_985_n 0.00998997f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_679 N_X_c_949_n N_VGND_M1005_d 0.00162006f $X=3.875 $Y=0.82 $X2=0 $Y2=0
cc_680 N_X_c_951_n N_VGND_M1008_d 0.00162006f $X=4.715 $Y=0.82 $X2=0 $Y2=0
cc_681 N_X_c_952_n N_VGND_M1013_d 0.00162006f $X=5.555 $Y=0.82 $X2=0 $Y2=0
cc_682 N_X_c_953_n N_VGND_M1016_d 0.00162006f $X=6.395 $Y=0.82 $X2=0 $Y2=0
cc_683 N_X_c_954_n N_VGND_M1029_d 0.00162006f $X=7.235 $Y=0.82 $X2=0 $Y2=0
cc_684 N_X_c_955_n N_VGND_M1032_d 0.00162006f $X=8.075 $Y=0.82 $X2=0 $Y2=0
cc_685 N_X_c_956_n N_VGND_M1040_d 0.00162006f $X=8.915 $Y=0.82 $X2=0 $Y2=0
cc_686 N_X_c_957_n N_VGND_M1043_d 0.0031176f $X=9.655 $Y=0.82 $X2=0 $Y2=0
cc_687 N_X_c_949_n N_VGND_c_1302_n 0.0122414f $X=3.875 $Y=0.82 $X2=0 $Y2=0
cc_688 N_X_c_951_n N_VGND_c_1303_n 0.0122414f $X=4.715 $Y=0.82 $X2=0 $Y2=0
cc_689 N_X_c_951_n N_VGND_c_1304_n 0.00193763f $X=4.715 $Y=0.82 $X2=0 $Y2=0
cc_690 N_X_c_1034_n N_VGND_c_1304_n 0.0187595f $X=4.88 $Y=0.425 $X2=0 $Y2=0
cc_691 N_X_c_952_n N_VGND_c_1304_n 0.00193763f $X=5.555 $Y=0.82 $X2=0 $Y2=0
cc_692 N_X_c_952_n N_VGND_c_1305_n 0.0122414f $X=5.555 $Y=0.82 $X2=0 $Y2=0
cc_693 N_X_c_953_n N_VGND_c_1306_n 0.0122414f $X=6.395 $Y=0.82 $X2=0 $Y2=0
cc_694 N_X_c_954_n N_VGND_c_1307_n 0.0122414f $X=7.235 $Y=0.82 $X2=0 $Y2=0
cc_695 N_X_c_955_n N_VGND_c_1308_n 0.0122414f $X=8.075 $Y=0.82 $X2=0 $Y2=0
cc_696 N_X_c_956_n N_VGND_c_1309_n 0.0122414f $X=8.915 $Y=0.82 $X2=0 $Y2=0
cc_697 N_X_c_956_n N_VGND_c_1310_n 0.00193763f $X=8.915 $Y=0.82 $X2=0 $Y2=0
cc_698 N_X_c_1116_n N_VGND_c_1310_n 0.0182681f $X=9.08 $Y=0.4 $X2=0 $Y2=0
cc_699 N_X_c_957_n N_VGND_c_1310_n 0.00193763f $X=9.655 $Y=0.82 $X2=0 $Y2=0
cc_700 N_X_c_957_n N_VGND_c_1311_n 0.0127122f $X=9.655 $Y=0.82 $X2=0 $Y2=0
cc_701 N_X_c_965_n N_VGND_c_1311_n 0.0150442f $X=9.845 $Y=0.82 $X2=0 $Y2=0
cc_702 N_X_c_988_n N_VGND_c_1318_n 0.0188753f $X=3.2 $Y=0.425 $X2=0 $Y2=0
cc_703 N_X_c_949_n N_VGND_c_1318_n 0.00193763f $X=3.875 $Y=0.82 $X2=0 $Y2=0
cc_704 N_X_c_949_n N_VGND_c_1320_n 0.00193763f $X=3.875 $Y=0.82 $X2=0 $Y2=0
cc_705 N_X_c_1016_n N_VGND_c_1320_n 0.0187595f $X=4.04 $Y=0.425 $X2=0 $Y2=0
cc_706 N_X_c_951_n N_VGND_c_1320_n 0.00193763f $X=4.715 $Y=0.82 $X2=0 $Y2=0
cc_707 N_X_c_952_n N_VGND_c_1322_n 0.00193763f $X=5.555 $Y=0.82 $X2=0 $Y2=0
cc_708 N_X_c_1052_n N_VGND_c_1322_n 0.0182681f $X=5.72 $Y=0.4 $X2=0 $Y2=0
cc_709 N_X_c_953_n N_VGND_c_1322_n 0.00193763f $X=6.395 $Y=0.82 $X2=0 $Y2=0
cc_710 N_X_c_953_n N_VGND_c_1324_n 0.00193763f $X=6.395 $Y=0.82 $X2=0 $Y2=0
cc_711 N_X_c_1068_n N_VGND_c_1324_n 0.0182681f $X=6.56 $Y=0.4 $X2=0 $Y2=0
cc_712 N_X_c_954_n N_VGND_c_1324_n 0.00193763f $X=7.235 $Y=0.82 $X2=0 $Y2=0
cc_713 N_X_c_954_n N_VGND_c_1326_n 0.00193763f $X=7.235 $Y=0.82 $X2=0 $Y2=0
cc_714 N_X_c_1084_n N_VGND_c_1326_n 0.0182681f $X=7.4 $Y=0.4 $X2=0 $Y2=0
cc_715 N_X_c_955_n N_VGND_c_1326_n 0.00193763f $X=8.075 $Y=0.82 $X2=0 $Y2=0
cc_716 N_X_c_955_n N_VGND_c_1328_n 0.00193763f $X=8.075 $Y=0.82 $X2=0 $Y2=0
cc_717 N_X_c_1100_n N_VGND_c_1328_n 0.0182681f $X=8.24 $Y=0.4 $X2=0 $Y2=0
cc_718 N_X_c_956_n N_VGND_c_1328_n 0.00193763f $X=8.915 $Y=0.82 $X2=0 $Y2=0
cc_719 N_X_c_957_n N_VGND_c_1330_n 0.0010013f $X=9.655 $Y=0.82 $X2=0 $Y2=0
cc_720 N_X_c_965_n N_VGND_c_1330_n 0.0132595f $X=9.845 $Y=0.82 $X2=0 $Y2=0
cc_721 N_X_M1000_s N_VGND_c_1331_n 0.00215228f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_722 N_X_M1006_s N_VGND_c_1331_n 0.00215254f $X=3.905 $Y=0.235 $X2=0 $Y2=0
cc_723 N_X_M1010_s N_VGND_c_1331_n 0.00215254f $X=4.745 $Y=0.235 $X2=0 $Y2=0
cc_724 N_X_M1015_s N_VGND_c_1331_n 0.00215347f $X=5.585 $Y=0.235 $X2=0 $Y2=0
cc_725 N_X_M1023_s N_VGND_c_1331_n 0.00215347f $X=6.425 $Y=0.235 $X2=0 $Y2=0
cc_726 N_X_M1031_s N_VGND_c_1331_n 0.00215347f $X=7.265 $Y=0.235 $X2=0 $Y2=0
cc_727 N_X_M1036_s N_VGND_c_1331_n 0.00215347f $X=8.105 $Y=0.235 $X2=0 $Y2=0
cc_728 N_X_M1041_s N_VGND_c_1331_n 0.00215347f $X=8.945 $Y=0.235 $X2=0 $Y2=0
cc_729 N_X_c_988_n N_VGND_c_1331_n 0.0122666f $X=3.2 $Y=0.425 $X2=0 $Y2=0
cc_730 N_X_c_949_n N_VGND_c_1331_n 0.00825759f $X=3.875 $Y=0.82 $X2=0 $Y2=0
cc_731 N_X_c_1016_n N_VGND_c_1331_n 0.0122584f $X=4.04 $Y=0.425 $X2=0 $Y2=0
cc_732 N_X_c_951_n N_VGND_c_1331_n 0.00825759f $X=4.715 $Y=0.82 $X2=0 $Y2=0
cc_733 N_X_c_1034_n N_VGND_c_1331_n 0.0122584f $X=4.88 $Y=0.425 $X2=0 $Y2=0
cc_734 N_X_c_952_n N_VGND_c_1331_n 0.00825759f $X=5.555 $Y=0.82 $X2=0 $Y2=0
cc_735 N_X_c_1052_n N_VGND_c_1331_n 0.0121741f $X=5.72 $Y=0.4 $X2=0 $Y2=0
cc_736 N_X_c_953_n N_VGND_c_1331_n 0.00825759f $X=6.395 $Y=0.82 $X2=0 $Y2=0
cc_737 N_X_c_1068_n N_VGND_c_1331_n 0.0121741f $X=6.56 $Y=0.4 $X2=0 $Y2=0
cc_738 N_X_c_954_n N_VGND_c_1331_n 0.00825759f $X=7.235 $Y=0.82 $X2=0 $Y2=0
cc_739 N_X_c_1084_n N_VGND_c_1331_n 0.0121741f $X=7.4 $Y=0.4 $X2=0 $Y2=0
cc_740 N_X_c_955_n N_VGND_c_1331_n 0.00825759f $X=8.075 $Y=0.82 $X2=0 $Y2=0
cc_741 N_X_c_1100_n N_VGND_c_1331_n 0.0121741f $X=8.24 $Y=0.4 $X2=0 $Y2=0
cc_742 N_X_c_956_n N_VGND_c_1331_n 0.00825759f $X=8.915 $Y=0.82 $X2=0 $Y2=0
cc_743 N_X_c_1116_n N_VGND_c_1331_n 0.0121741f $X=9.08 $Y=0.4 $X2=0 $Y2=0
cc_744 N_X_c_957_n N_VGND_c_1331_n 0.00631085f $X=9.655 $Y=0.82 $X2=0 $Y2=0
cc_745 N_X_c_965_n N_VGND_c_1331_n 0.012834f $X=9.845 $Y=0.82 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dfrtp_2.spice.pex
* Created: Thu Aug 27 14:14:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFRTP_2%CLK 1 2 3 5 6 8 11 13 14
c40 6 0 9.23148e-20 $X=0.47 $Y=1.74
c41 1 0 2.71124e-20 $X=0.305 $Y=1.325
r42 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r43 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r47 3 18 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r50 1 18 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_27_47# 1 2 9 13 17 20 21 22 25 27 29 33 37
+ 41 42 43 46 49 50 51 52 55 61 68 71 72 77
c236 77 0 4.56546e-20 $X=6.07 $Y=1.11
c237 61 0 1.76704e-20 $X=6.11 $Y=1.19
c238 51 0 1.58851e-19 $X=5.965 $Y=1.19
c239 29 0 4.11863e-20 $X=5.845 $Y=2.275
c240 22 0 1.90473e-19 $X=2.72 $Y=1.32
r241 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.11 $X2=6.07 $Y2=1.11
r242 71 74 47.4498 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=1.095
r243 71 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=0.765
r244 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.93 $X2=2.585 $Y2=0.93
r245 65 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r246 61 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.19
+ $X2=6.11 $Y2=1.19
r247 59 72 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.56 $Y=1.19
+ $X2=2.56 $Y2=0.93
r248 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r249 55 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r250 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.19
+ $X2=0.695 $Y2=1.19
r251 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.19
+ $X2=2.53 $Y2=1.19
r252 51 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=6.11 $Y2=1.19
r253 51 52 4.07177 $w=1.4e-07 $l=3.29e-06 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=2.675 $Y2=1.19
r254 50 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.19
+ $X2=0.695 $Y2=1.19
r255 49 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r256 49 50 1.91213 $w=1.4e-07 $l=1.545e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.84 $Y2=1.19
r257 48 55 30.3143 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.19
r258 47 55 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.19
r259 44 46 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r260 43 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.795
r261 43 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r262 41 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r263 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r264 35 42 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.345 $Y2=0.72
r265 35 37 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.51
r266 31 76 38.5991 $w=2.92e-07 $l=1.76125e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=5.987 $Y2=1.11
r267 31 33 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=6.01 $Y2=0.415
r268 27 76 58.4073 $w=2.92e-07 $l=3.48848e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.987 $Y2=1.11
r269 27 29 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.845 $Y2=2.275
r270 23 25 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.18 $Y=1.395
+ $X2=3.18 $Y2=2.275
r271 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=3.18 $Y2=1.395
r272 21 22 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=2.72 $Y2=1.32
r273 20 22 26.9401 $w=1.5e-07 $l=1.09243e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.72 $Y2=1.32
r274 20 74 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.642 $Y2=1.095
r275 17 73 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.64 $Y=0.415
+ $X2=2.64 $Y2=0.765
r276 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r277 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r278 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r279 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r280 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r281 1 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%D 3 7 9 10 15 19
c53 10 0 1.85993e-19 $X=2.09 $Y=1.3
c54 7 0 1.77283e-19 $X=2.225 $Y=2.275
r55 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.465 $X2=1.79 $Y2=1.465
r56 15 19 1.96287 $w=4.04e-07 $l=6.5e-08 $layer=LI1_cond $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.465
r57 9 18 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.09 $Y=1.465 $X2=1.79
+ $Y2=1.465
r58 9 10 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.465
+ $X2=2.09 $Y2=1.3
r59 5 10 37.0704 $w=1.5e-07 $l=3.91727e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.09 $Y2=1.3
r60 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.225 $Y2=2.275
r61 1 10 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=1.3 $X2=2.09
+ $Y2=1.3
r62 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.165 $Y=1.3
+ $X2=2.165 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_193_47# 1 2 9 13 15 17 20 23 26 27 29 30
+ 34 35 37 38 39 40 47 49 53 65 66 70
c212 66 0 3.94709e-20 $X=6.265 $Y=1.74
c213 47 0 1.77283e-19 $X=2.99 $Y=1.87
c214 39 0 1.36782e-20 $X=5.965 $Y=1.87
c215 38 0 9.23148e-20 $X=1.245 $Y=1.87
c216 37 0 1.20979e-19 $X=2.845 $Y=1.87
c217 35 0 1.61046e-19 $X=3.095 $Y=0.9
c218 29 0 1.76704e-20 $X=5.97 $Y=1.58
c219 26 0 1.28114e-19 $X=5.59 $Y=0.87
r220 65 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.74
+ $X2=6.265 $Y2=1.905
r221 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.265
+ $Y=1.74 $X2=6.265 $Y2=1.74
r222 53 56 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.695 $Y=1.74
+ $X2=2.695 $Y2=1.875
r223 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.74 $X2=2.695 $Y2=1.74
r224 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.87
+ $X2=6.11 $Y2=1.87
r225 47 54 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=1.77
+ $X2=2.695 $Y2=1.77
r226 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.87
+ $X2=2.99 $Y2=1.87
r227 43 70 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.1 $Y=1.87
+ $X2=1.1 $Y2=0.51
r228 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.87 $X2=1.1
+ $Y2=1.87
r229 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.87
+ $X2=2.99 $Y2=1.87
r230 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=6.11 $Y2=1.87
r231 39 40 3.50247 $w=1.4e-07 $l=2.83e-06 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=3.135 $Y2=1.87
r232 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.87
+ $X2=1.1 $Y2=1.87
r233 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=2.99 $Y2=1.87
r234 37 38 1.98019 $w=1.4e-07 $l=1.6e-06 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=1.245 $Y2=1.87
r235 35 58 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.095 $Y=0.9
+ $X2=3.095 $Y2=0.765
r236 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=0.9 $X2=3.095 $Y2=0.9
r237 31 34 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.875
+ $X2=3.095 $Y2=0.875
r238 29 66 5.43733 $w=3.59e-07 $l=2.995e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=6.2 $Y2=1.74
r239 29 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.675 $Y2=1.58
r240 27 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.59 $Y=0.87
+ $X2=5.465 $Y2=0.87
r241 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=0.87 $X2=5.59 $Y2=0.87
r242 24 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.675 $Y2=1.58
r243 24 26 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.57 $Y2=0.87
r244 23 47 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.99 $Y=1.575
+ $X2=2.99 $Y2=1.77
r245 22 31 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=0.875
r246 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=1.575
r247 20 68 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.275 $Y=2.275
+ $X2=6.275 $Y2=1.905
r248 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.87
r249 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.415
r250 13 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.12 $Y=0.415
+ $X2=3.12 $Y2=0.765
r251 9 56 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.685 $Y=2.275
+ $X2=2.685 $Y2=1.875
r252 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r253 1 70 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_761_289# 1 2 9 13 15 18 21 23 25 26 27 30
+ 33 36 37
c109 36 0 1.00332e-19 $X=5.145 $Y=0.835
c110 23 0 4.11863e-20 $X=5.19 $Y=1.525
r111 33 35 3.58511 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.36
+ $X2=5.19 $Y2=0.445
r112 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.58 $Y=2.005
+ $X2=5.58 $Y2=2.3
r113 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.58 $Y2=2.005
r114 26 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.275 $Y2=1.92
r115 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.19 $Y=1.835
+ $X2=5.275 $Y2=1.92
r116 24 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.61
r117 24 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.835
r118 23 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=1.61
r119 23 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=0.835
r120 21 36 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.835
r121 21 35 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.445
r122 18 40 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.775
r123 18 39 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.445
r124 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.61 $X2=3.94 $Y2=1.61
r125 15 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=5.19 $Y2=1.61
r126 15 17 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=3.94 $Y2=1.61
r127 13 39 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.95 $Y=0.445
+ $X2=3.95 $Y2=1.445
r128 9 40 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.88 $Y=2.275 $X2=3.88
+ $Y2=1.775
r129 2 30 600 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.645 $X2=5.58 $Y2=2.3
r130 1 33 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.2 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%RESET_B 3 6 10 14 16 17 20 23 25 26 27 29 37
+ 39 42 57
c154 37 0 1.00332e-19 $X=4.37 $Y=0.93
c155 29 0 4.83118e-21 $X=7.19 $Y=1.165
c156 23 0 6.10372e-20 $X=4.25 $Y=0.85
c157 14 0 1.03533e-19 $X=7.235 $Y=2.275
c158 10 0 4.70414e-20 $X=7.235 $Y=0.445
r159 49 57 3.2703 $w=2.4e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=1.035
+ $X2=7.525 $Y2=1.22
r160 42 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=1.285
r161 42 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=0.955
r162 37 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=1.095
r163 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=0.765
r164 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.12 $X2=7.27 $Y2=1.12
r165 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.19 $Y=1.165
+ $X2=7.19 $Y2=1.165
r166 27 34 0.181159 $w=2.07e-07 $l=3e-07 $layer=MET1_cond $X=7.19 $Y=0.85
+ $X2=7.49 $Y2=0.85
r167 27 29 0.0979621 $w=2.9e-07 $l=2e-07 $layer=MET1_cond $X=7.19 $Y=0.965
+ $X2=7.19 $Y2=1.165
r168 25 27 0.10072 $w=2.07e-07 $l=1.45e-07 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=7.19 $Y2=0.85
r169 25 26 3.2797 $w=1.4e-07 $l=2.65e-06 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=4.395 $Y2=0.85
r170 23 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=0.93 $X2=4.37 $Y2=0.93
r171 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.25 $Y=0.85
+ $X2=4.25 $Y2=0.85
r172 20 26 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.395 $Y2=0.85
r173 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.25 $Y2=0.85
r174 17 57 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.49 $Y=1.22
+ $X2=7.525 $Y2=1.22
r175 17 30 9.34413 $w=3.68e-07 $l=3e-07 $layer=LI1_cond $X=7.49 $Y=1.22 $X2=7.19
+ $Y2=1.22
r176 16 49 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=0.85
+ $X2=7.525 $Y2=1.035
r177 16 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.49 $Y=0.85
+ $X2=7.49 $Y2=0.85
r178 14 45 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=7.235 $Y=2.275
+ $X2=7.235 $Y2=1.285
r179 10 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.235 $Y=0.445
+ $X2=7.235 $Y2=0.955
r180 6 40 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.365 $Y=2.275
+ $X2=4.365 $Y2=1.095
r181 3 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.31 $Y=0.445
+ $X2=4.31 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_543_47# 1 2 9 11 13 15 16 20 25 27 28 29
+ 34 35
c126 35 0 6.10372e-20 $X=4.85 $Y=1.17
c127 29 0 1.61046e-19 $X=3.6 $Y=1.27
c128 11 0 1.36782e-20 $X=5.275 $Y=1.495
c129 9 0 1.28114e-19 $X=4.97 $Y=0.555
r130 34 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.85 $Y=1.17 $X2=4.85
+ $Y2=1.27
r131 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.17 $X2=4.85 $Y2=1.17
r132 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.33 $Y=1.27
+ $X2=3.515 $Y2=1.27
r133 29 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.27
+ $X2=3.515 $Y2=1.27
r134 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=4.85 $Y2=1.27
r135 28 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=3.6 $Y2=1.27
r136 27 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=1.27
r137 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.515 $Y=0.475
+ $X2=3.515 $Y2=1.185
r138 24 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=1.27
r139 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=2.135
r140 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=3.515 $Y2=0.475
r141 20 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=2.91 $Y2=0.39
r142 16 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=3.33 $Y2=2.135
r143 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=2.9 $Y2=2.3
r144 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.35 $Y=1.57
+ $X2=5.35 $Y2=2.065
r145 12 35 61.4314 $w=2.55e-07 $l=3.99061e-07 $layer=POLY_cond $X=5.045 $Y=1.495
+ $X2=4.88 $Y2=1.17
r146 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.35 $Y2=1.57
r147 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.045 $Y2=1.495
r148 7 35 39.2931 $w=2.55e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.88 $Y2=1.17
r149 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.97 $Y2=0.555
r150 2 18 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.065 $X2=2.9 $Y2=2.33
r151 1 22 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.91 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_1283_21# 1 2 9 13 15 17 20 22 24 27 31 35
+ 36 37 40 42 43 44 45 47 50 55 59 61 66
c161 66 0 3.00828e-19 $X=9.15 $Y=1.16
c162 61 0 6.15427e-20 $X=6.695 $Y=0.98
c163 59 0 1.99375e-19 $X=7.815 $Y=0.82
c164 55 0 1.94811e-19 $X=7.15 $Y=0.78
c165 13 0 2.35828e-20 $X=6.695 $Y=2.275
r166 65 66 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.73 $Y=1.16
+ $X2=9.15 $Y2=1.16
r167 51 65 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=8.645 $Y=1.16
+ $X2=8.73 $Y2=1.16
r168 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.645
+ $Y=1.16 $X2=8.645 $Y2=1.16
r169 48 59 0.295496 $w=3.3e-07 $l=4.86133e-07 $layer=LI1_cond $X=8.16 $Y=1.16
+ $X2=7.815 $Y2=0.82
r170 48 50 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=8.16 $Y=1.16
+ $X2=8.645 $Y2=1.16
r171 46 59 6.56857 $w=2.45e-07 $l=6.2155e-07 $layer=LI1_cond $X=8.075 $Y=1.325
+ $X2=7.815 $Y2=0.82
r172 46 47 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.075 $Y=1.325
+ $X2=8.075 $Y2=1.915
r173 45 59 6.56857 $w=2.45e-07 $l=1.6e-07 $layer=LI1_cond $X=7.975 $Y=0.82
+ $X2=7.815 $Y2=0.82
r174 44 58 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=0.465
+ $X2=7.975 $Y2=0.38
r175 44 45 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=7.975 $Y=0.465
+ $X2=7.975 $Y2=0.82
r176 42 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.99 $Y=2
+ $X2=8.075 $Y2=1.915
r177 42 43 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.99 $Y=2 $X2=7.53
+ $Y2=2
r178 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.53 $Y2=2
r179 38 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.445 $Y2=2.21
r180 36 58 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.975 $Y2=0.38
r181 36 37 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.235 $Y2=0.38
r182 35 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=0.695
+ $X2=7.15 $Y2=0.78
r183 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.235 $Y2=0.38
r184 34 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.15 $Y2=0.695
r185 32 61 17.8171 $w=2.57e-07 $l=9.5e-08 $layer=POLY_cond $X=6.79 $Y=0.98
+ $X2=6.695 $Y2=0.98
r186 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=0.98 $X2=6.79 $Y2=0.98
r187 29 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0.78
+ $X2=7.15 $Y2=0.78
r188 29 31 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=6.815 $Y=0.865
+ $X2=6.815 $Y2=0.98
r189 25 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.15 $Y=1.325
+ $X2=9.15 $Y2=1.16
r190 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.15 $Y=1.325
+ $X2=9.15 $Y2=1.985
r191 22 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.15 $Y=0.995
+ $X2=9.15 $Y2=1.16
r192 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.15 $Y=0.995
+ $X2=9.15 $Y2=0.56
r193 18 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=1.325
+ $X2=8.73 $Y2=1.16
r194 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.73 $Y=1.325
+ $X2=8.73 $Y2=1.985
r195 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=0.995
+ $X2=8.73 $Y2=1.16
r196 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.73 $Y=0.995
+ $X2=8.73 $Y2=0.56
r197 11 61 15.359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=0.98
r198 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=2.275
r199 7 61 38.4475 $w=2.57e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.695 $Y2=0.98
r200 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.49 $Y2=0.445
r201 2 40 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=2.065 $X2=7.445 $Y2=2.21
r202 1 58 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=7.765
+ $Y=0.235 $X2=7.9 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_1108_47# 1 2 9 13 15 19 24 25 26 29 30
c103 25 0 2.04429e-20 $X=6.685 $Y=1.745
c104 24 0 1.60161e-19 $X=6.45 $Y=1.315
c105 19 0 1.03533e-19 $X=6.6 $Y=2.295
c106 15 0 4.70414e-20 $X=6.365 $Y=0.395
c107 13 0 1.79199e-19 $X=7.69 $Y=0.445
r108 30 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.66
+ $X2=7.655 $Y2=1.495
r109 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.655
+ $Y=1.66 $X2=7.655 $Y2=1.66
r110 27 32 3.26844 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.77 $Y=1.66 $X2=6.6
+ $Y2=1.66
r111 27 29 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.77 $Y=1.66
+ $X2=7.655 $Y2=1.66
r112 25 32 5.45986 $w=2.62e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.6 $Y2=1.66
r113 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.685 $Y2=2.125
r114 24 32 17.5667 $w=2.62e-07 $l=4.13249e-07 $layer=LI1_cond $X=6.45 $Y=1.315
+ $X2=6.6 $Y2=1.66
r115 23 24 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.45 $Y=0.535
+ $X2=6.45 $Y2=1.315
r116 19 26 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.685 $Y2=2.125
r117 19 21 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.065 $Y2=2.295
r118 15 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=6.45 $Y2=0.535
r119 15 17 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=5.75 $Y2=0.395
r120 13 34 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=7.69 $Y=0.445
+ $X2=7.69 $Y2=1.495
r121 7 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=1.66
r122 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=2.275
r123 2 21 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=2.065 $X2=6.065 $Y2=2.335
r124 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.54
+ $Y=0.235 $X2=5.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 53
+ 55 60 61 63 64 66 67 68 70 75 84 95 99 105 108 111 114 118
r155 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r156 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r157 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r158 108 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r160 103 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r161 103 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r162 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r163 100 114 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.685 $Y=2.72
+ $X2=8.532 $Y2=2.72
r164 100 102 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.685 $Y=2.72
+ $X2=8.97 $Y2=2.72
r165 99 117 3.98688 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=9.275 $Y=2.72
+ $X2=9.467 $Y2=2.72
r166 99 102 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.275 $Y=2.72
+ $X2=8.97 $Y2=2.72
r167 98 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r168 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r169 95 114 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.38 $Y=2.72
+ $X2=8.532 $Y2=2.72
r170 95 97 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.38 $Y=2.72
+ $X2=8.05 $Y2=2.72
r171 94 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r172 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r173 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r174 91 112 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.29 $Y2=2.72
r175 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r176 88 111 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.14 $Y2=2.72
r177 88 90 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=6.67 $Y2=2.72
r178 87 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r179 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r180 84 111 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.14 $Y2=2.72
r181 84 86 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.83 $Y2=2.72
r182 83 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r183 83 109 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.07 $Y2=2.72
r184 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r185 80 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=1.975 $Y2=2.72
r186 80 82 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=3.91 $Y2=2.72
r187 79 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r188 79 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r189 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r190 76 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r191 76 78 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r192 75 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.975 $Y2=2.72
r193 75 78 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r194 70 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r195 70 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r196 68 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r197 68 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r198 66 93 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.59 $Y2=2.72
r199 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.875 $Y2=2.72
r200 65 97 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=8.05 $Y2=2.72
r201 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=7.875 $Y2=2.72
r202 63 90 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=6.67 $Y2=2.72
r203 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=7.065 $Y2=2.72
r204 62 93 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.19 $Y=2.72 $X2=7.59
+ $Y2=2.72
r205 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.065 $Y2=2.72
r206 60 82 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.99 $Y=2.72 $X2=3.91
+ $Y2=2.72
r207 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=2.72
+ $X2=4.155 $Y2=2.72
r208 59 86 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.83 $Y2=2.72
r209 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.155 $Y2=2.72
r210 55 58 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=9.4 $Y=1.66 $X2=9.4
+ $Y2=2.34
r211 53 117 3.15628 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=9.4 $Y=2.635
+ $X2=9.467 $Y2=2.72
r212 53 58 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.4 $Y=2.635
+ $X2=9.4 $Y2=2.34
r213 49 114 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.532 $Y=2.635
+ $X2=8.532 $Y2=2.72
r214 49 51 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=8.532 $Y=2.635
+ $X2=8.532 $Y2=2
r215 45 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.72
r216 45 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.34
r217 41 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.72
r218 41 43 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.34
r219 37 111 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.72
r220 37 39 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.34
r221 33 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.72
r222 33 35 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.29
r223 29 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.72
r224 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.34
r225 25 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r226 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r227 8 58 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.225
+ $Y=1.485 $X2=9.36 $Y2=2.34
r228 8 55 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.225
+ $Y=1.485 $X2=9.36 $Y2=1.66
r229 7 51 300 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=1.845 $X2=8.52 $Y2=2
r230 6 47 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=2.065 $X2=7.875 $Y2=2.34
r231 5 43 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=2.065 $X2=7.025 $Y2=2.34
r232 4 39 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.645 $X2=5.14 $Y2=2.34
r233 3 35 600 $w=1.7e-07 $l=3.09233e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=2.065 $X2=4.155 $Y2=2.29
r234 2 31 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=2.065 $X2=2.015 $Y2=2.34
r235 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_448_47# 1 2 8 9 11
c34 8 0 6.94938e-20 $X=2.13 $Y=1.835
r35 9 11 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.215 $Y=0.39
+ $X2=2.375 $Y2=0.39
r36 8 14 22.5629 $w=2.72e-07 $l=5.35635e-07 $layer=LI1_cond $X=2.13 $Y=1.835
+ $X2=2.282 $Y2=2.3
r37 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.215 $Y2=0.39
r38 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.13 $Y2=1.835
r39 2 14 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.065 $X2=2.435 $Y2=2.3
r40 1 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.375 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%A_651_413# 1 2 9 11 12 15
c36 12 0 1.58851e-19 $X=3.755 $Y=1.95
r37 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.035
+ $X2=4.575 $Y2=2.21
r38 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=4.575 $Y2=2.035
r39 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=3.755 $Y2=1.95
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.755 $Y2=1.95
r41 7 9 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.67 $Y2=2.21
r42 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=2.065 $X2=4.575 $Y2=2.21
r43 1 9 600 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=2.065 $X2=3.67 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%Q 1 2 9 10 11 12 13 38
c16 11 0 1.60027e-19 $X=8.88 $Y=1.445
c17 9 0 1.408e-19 $X=8.98 $Y=0.795
r18 25 38 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=8.98 $Y=1.57 $X2=8.98
+ $Y2=1.53
r19 12 13 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=8.98 $Y=1.82
+ $X2=8.98 $Y2=2.21
r20 11 38 1.06025 $w=2.48e-07 $l=2.3e-08 $layer=LI1_cond $X=8.98 $Y=1.507
+ $X2=8.98 $Y2=1.53
r21 11 12 10.5103 $w=2.48e-07 $l=2.28e-07 $layer=LI1_cond $X=8.98 $Y=1.592
+ $X2=8.98 $Y2=1.82
r22 11 25 1.01415 $w=2.48e-07 $l=2.2e-08 $layer=LI1_cond $X=8.98 $Y=1.592
+ $X2=8.98 $Y2=1.57
r23 10 24 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=8.98 $Y=0.51
+ $X2=8.98 $Y2=0.63
r24 9 11 22.3451 $w=3.53e-07 $l=6.5e-07 $layer=LI1_cond $X=9.002 $Y=0.795
+ $X2=9.002 $Y2=1.445
r25 7 24 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=8.98 $Y=0.67 $X2=8.98
+ $Y2=0.63
r26 7 9 6.16968 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.98 $Y=0.67 $X2=8.98
+ $Y2=0.795
r27 2 12 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=8.805
+ $Y=1.485 $X2=8.94 $Y2=1.82
r28 1 24 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=8.805
+ $Y=0.235 $X2=8.94 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_2%VGND 1 2 3 4 5 6 21 23 27 31 35 39 41 43 46
+ 47 49 50 51 53 71 78 84 87 90 94
c142 94 0 2.26487e-19 $X=9.43 $Y=0
r143 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r144 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r145 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r146 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r147 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r148 82 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.43
+ $Y2=0
r149 82 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=8.51
+ $Y2=0
r150 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r151 79 90 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.685 $Y=0
+ $X2=8.532 $Y2=0
r152 79 81 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.685 $Y=0
+ $X2=8.97 $Y2=0
r153 78 93 3.98688 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=9.275 $Y=0
+ $X2=9.467 $Y2=0
r154 78 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.275 $Y=0
+ $X2=8.97 $Y2=0
r155 77 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.51
+ $Y2=0
r156 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r157 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r158 73 76 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r159 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r160 71 90 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.38 $Y=0 $X2=8.532
+ $Y2=0
r161 71 76 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.38 $Y=0 $X2=8.05
+ $Y2=0
r162 70 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r163 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r164 67 70 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.67 $Y2=0
r165 66 69 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.67
+ $Y2=0
r166 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r167 64 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r168 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r169 61 64 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r170 61 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r171 60 63 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r172 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r173 58 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r174 58 60 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.07 $Y2=0
r175 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r176 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r177 51 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r178 51 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r179 49 69 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.67
+ $Y2=0
r180 49 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.8
+ $Y2=0
r181 48 73 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.895 $Y=0
+ $X2=7.13 $Y2=0
r182 48 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.8
+ $Y2=0
r183 46 63 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r184 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r185 45 66 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.83
+ $Y2=0
r186 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r187 41 93 3.15628 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=9.4 $Y=0.085
+ $X2=9.467 $Y2=0
r188 41 43 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=9.4 $Y=0.085
+ $X2=9.4 $Y2=0.55
r189 37 90 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.532 $Y=0.085
+ $X2=8.532 $Y2=0
r190 37 39 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=8.532 $Y=0.085
+ $X2=8.532 $Y2=0.38
r191 33 50 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0
r192 33 35 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0.36
r193 29 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r194 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.38
r195 25 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r196 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.36
r197 24 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r198 23 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r199 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=0.845
+ $Y2=0
r200 19 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r201 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r202 6 43 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=9.225
+ $Y=0.235 $X2=9.36 $Y2=0.55
r203 5 39 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.235 $X2=8.52 $Y2=0.38
r204 4 35 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.81 $Y2=0.36
r205 3 31 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.64 $Y2=0.38
r206 2 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.71 $Y2=0.36
r207 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_615_93# C a_515_93# VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.58e+06u as=1.47e+11p ps=1.54e+06u
M1001 a_515_93# a_223_47# a_429_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1002 VPWR a_223_47# a_343_93# VPB phighvt w=420000u l=150000u
+  ad=7.304e+11p pd=7.28e+06u as=2.73e+11p ps=2.98e+06u
M1003 VPWR D a_343_93# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_343_93# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_343_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.654e+11p pd=1.82e+06u as=3.706e+11p ps=3.62e+06u
M1006 VPWR A_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.68e+11p ps=1.64e+06u
M1007 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.68e+11p ps=1.64e+06u
M1008 a_343_93# a_27_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_223_47# B_N VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1010 VGND D a_615_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_429_93# a_27_47# a_343_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1012 a_223_47# B_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1013 X a_343_93# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__nand3b_2.spice
* Created: Thu Aug 27 14:29:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand3b_2.pex.spice"
.subckt sky130_fd_sc_hd__nand3b_2  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0940093 AS=0.1092 PD=0.820374 PS=1.36 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1013_d N_C_M1005_g N_A_218_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.145491 AS=0.08775 PD=1.26963 PS=0.92 NRD=10.152 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_C_M1008_g N_A_218_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_218_47#_M1000_d N_B_M1000_g N_A_408_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 N_A_218_47#_M1000_d N_B_M1002_g N_A_408_47#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 N_A_408_47#_M1002_s N_A_27_47#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_408_47#_M1009_d N_A_27_47#_M1009_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.103965 AS=0.1092 PD=0.825211 PS=1.36 NRD=29.3136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1004_d N_C_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.247535
+ AS=0.135 PD=1.96479 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75000.4
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_C_M1011_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.9 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1001 N_VPWR_M1011_d N_B_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.3 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.7 SB=75000.2
+ A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_47#_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A_27_47#_M1012_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_41 VNB 0 9.80354e-20 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__nand3b_2.pxi.spice"
*
.ends
*
*

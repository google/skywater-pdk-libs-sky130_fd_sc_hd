* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_109_47# VNB nshort w=650000u l=150000u
+  ad=3.055e+11p pd=2.24e+06u as=1.495e+11p ps=1.76e+06u
M1001 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=9.7e+11p pd=7.94e+06u as=2.7e+11p ps=2.54e+06u
M1002 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.3e+11p pd=5.06e+06u as=0p ps=0u
M1003 a_309_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.43e+11p pd=1.74e+06u as=0p ps=0u
M1004 a_383_47# A2 a_309_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=0p ps=0u
M1005 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_109_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.38e+11p ps=3.64e+06u
M1009 VGND A3 a_383_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__o21ba_2.spice
* Created: Thu Aug 27 14:36:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21ba_2.spice.pex"
.subckt sky130_fd_sc_hd__o21ba_2  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_B1_N_M1010_g N_A_27_93#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1010_d N_A_174_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.08775 PD=1.18458 PS=0.92 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_174_21#_M1011_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_478_47#_M1003_d N_A_27_93#_M1003_g N_A_174_21#_M1003_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.105625 AS=0.169 PD=0.975 PS=1.82 NRD=9.228 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_478_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.105625 PD=0.92 PS=0.975 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_478_47#_M1008_d N_A1_M1008_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_B1_N_M1006_g N_A_27_93#_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=70.4866 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1006_d N_A_174_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.205282 AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_174_21#_M1009_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.395 AS=0.135 PD=1.79 PS=1.27 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1004 N_A_174_21#_M1004_d N_A_27_93#_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1 AD=0.165 AS=0.395 PD=1.33 PS=1.79 NRD=10.8153 NRS=6.8753 M=1 R=6.66667
+ SA=75001.7 SB=75001 A=0.15 P=2.3 MULT=1
MM1000 A_574_297# N_A2_M1000_g N_A_174_21#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.165 PD=1.21 PS=1.33 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75002.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_574_297# VPB PHIGHVT L=0.15 W=1 AD=0.28
+ AS=0.105 PD=2.56 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.6 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_73 VPB 0 7.75504e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__o21ba_2.spice.SKY130_FD_SC_HD__O21BA_2.pxi"
*
.ends
*
*

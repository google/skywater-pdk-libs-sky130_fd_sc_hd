* File: sky130_fd_sc_hd__edfxtp_1.spice.pex
* Created: Thu Aug 27 14:19:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%CLK 1 2 3 5 6 8 11 13
c40 1 0 2.71124e-20 $X=0.31 $Y=1.325
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r42 9 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.47 $Y2=1.665
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r44 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r45 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r46 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r47 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r48 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r49 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_27_47# 1 2 9 13 17 21 25 27 31 35 39 40
+ 41 44 46 48 51 54 56 57 58 59 60 67 69 74 82 85 89
c251 89 0 1.92554e-19 $X=7.875 $Y=1.41
c252 51 0 1.74912e-19 $X=4.98 $Y=0.87
c253 48 0 1.43548e-19 $X=5.15 $Y=0.845
c254 44 0 1.8506e-19 $X=0.73 $Y=1.795
c255 41 0 5.65522e-20 $X=0.615 $Y=1.88
r256 88 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.875 $Y=1.41
+ $X2=7.875 $Y2=1.575
r257 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.875
+ $Y=1.41 $X2=7.875 $Y2=1.41
r258 85 88 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.875 $Y=1.32
+ $X2=7.875 $Y2=1.41
r259 79 82 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.31 $Y=1.74
+ $X2=5.405 $Y2=1.74
r260 70 89 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=7.885 $Y=1.87
+ $X2=7.885 $Y2=1.41
r261 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.885 $Y=1.87
+ $X2=7.885 $Y2=1.87
r262 67 96 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=5.295 $Y=1.83
+ $X2=5.235 $Y2=1.83
r263 67 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.405
+ $Y=1.74 $X2=5.405 $Y2=1.74
r264 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.295 $Y=1.87
+ $X2=5.295 $Y2=1.87
r265 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=1.87
r266 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.44 $Y=1.87
+ $X2=5.295 $Y2=1.87
r267 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.74 $Y=1.87
+ $X2=7.885 $Y2=1.87
r268 59 60 2.84653 $w=1.4e-07 $l=2.3e-06 $layer=MET1_cond $X=7.74 $Y=1.87
+ $X2=5.44 $Y2=1.87
r269 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=1.87
+ $X2=0.72 $Y2=1.87
r270 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.15 $Y=1.87
+ $X2=5.295 $Y2=1.87
r271 57 58 5.30321 $w=1.4e-07 $l=4.285e-06 $layer=MET1_cond $X=5.15 $Y=1.87
+ $X2=0.865 $Y2=1.87
r272 54 96 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.235 $Y=1.655
+ $X2=5.235 $Y2=1.83
r273 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.235 $Y=0.955
+ $X2=5.235 $Y2=1.655
r274 51 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.98 $Y=0.87
+ $X2=4.98 $Y2=0.735
r275 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=0.87 $X2=4.98 $Y2=0.87
r276 48 53 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.15 $Y=0.845
+ $X2=5.235 $Y2=0.955
r277 48 50 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=5.15 $Y=0.845
+ $X2=4.98 $Y2=0.845
r278 47 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r279 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r280 44 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r281 44 46 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r282 43 46 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.73 $Y=0.805
+ $X2=0.73 $Y2=1.235
r283 42 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r284 41 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r285 41 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.345 $Y2=1.88
r286 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.73 $Y2=0.805
r287 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r288 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r289 33 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r290 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=8.51 $Y=1.245
+ $X2=8.51 $Y2=0.415
r291 28 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.01 $Y=1.32
+ $X2=7.875 $Y2=1.32
r292 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.435 $Y=1.32
+ $X2=8.51 $Y2=1.245
r293 27 28 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=8.435 $Y=1.32
+ $X2=8.01 $Y2=1.32
r294 25 90 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=7.88 $Y=2.275
+ $X2=7.88 $Y2=1.575
r295 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.905
+ $X2=5.31 $Y2=1.74
r296 19 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.31 $Y=1.905
+ $X2=5.31 $Y2=2.275
r297 17 77 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.99 $Y=0.415
+ $X2=4.99 $Y2=0.735
r298 11 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r299 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r300 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r301 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r302 2 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r303 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%D 3 7 9 12 13 16
c51 7 0 5.26342e-20 $X=1.83 $Y=2.165
r52 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.78
+ $Y=1.145 $X2=1.78 $Y2=1.145
r53 11 16 70.9845 $w=3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.765 $Y=1.5
+ $X2=1.765 $Y2=1.145
r54 11 12 43.217 $w=3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.765 $Y=1.5 $X2=1.765
+ $Y2=1.65
r55 9 16 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.765 $Y=1.13 $X2=1.765
+ $Y2=1.145
r56 9 10 43.217 $w=3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.765 $Y=1.13 $X2=1.765
+ $Y2=0.98
r57 7 12 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.83 $Y=2.165
+ $X2=1.83 $Y2=1.65
r58 3 10 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_423_343# 1 2 7 9 12 16 20 23 26 27 36
c88 27 0 1.67735e-19 $X=3.55 $Y=1.01
c89 23 0 5.26342e-20 $X=2.932 $Y=1.355
c90 20 0 1.1082e-19 $X=2.92 $Y=0.51
r91 30 33 10.7351 $w=3.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.58 $Y=1.537
+ $X2=2.92 $Y2=1.537
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.52 $X2=2.58 $Y2=1.52
r93 27 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.01
+ $X2=3.55 $Y2=0.845
r94 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.01 $X2=3.55 $Y2=1.01
r95 24 36 0.565906 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=3.085 $Y=1.01
+ $X2=2.932 $Y2=1.01
r96 24 26 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.085 $Y=1.01
+ $X2=3.55 $Y2=1.01
r97 23 33 0.378885 $w=3.63e-07 $l=1.2e-08 $layer=LI1_cond $X=2.932 $Y=1.537
+ $X2=2.92 $Y2=1.537
r98 22 36 6.17543 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=2.932 $Y=1.175
+ $X2=2.932 $Y2=1.01
r99 22 23 6.8013 $w=3.03e-07 $l=1.8e-07 $layer=LI1_cond $X=2.932 $Y=1.175
+ $X2=2.932 $Y2=1.355
r100 18 36 6.17543 $w=2.65e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.892 $Y=0.845
+ $X2=2.932 $Y2=1.01
r101 18 20 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=2.892 $Y=0.845
+ $X2=2.892 $Y2=0.51
r102 14 33 1.32393 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=2.92 $Y=1.72
+ $X2=2.92 $Y2=1.537
r103 14 16 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.92 $Y=1.72
+ $X2=2.92 $Y2=1.99
r104 12 40 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.57 $Y=0.445
+ $X2=3.57 $Y2=0.845
r105 7 31 69.3653 $w=2.71e-07 $l=4.76833e-07 $layer=POLY_cond $X=2.19 $Y=1.77
+ $X2=2.58 $Y2=1.577
r106 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.19 $Y=1.77
+ $X2=2.19 $Y2=2.165
r107 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=1.845 $X2=2.92 $Y2=1.99
r108 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.92 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%DE 3 5 6 9 12 15 17 21 23 24 25
c85 6 0 1.1082e-19 $X=2.455 $Y=0.925
r86 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.01 $X2=2.29 $Y2=1.01
r87 27 29 13.5393 $w=3.56e-07 $l=1e-07 $layer=POLY_cond $X=2.19 $Y=0.992
+ $X2=2.29 $Y2=0.992
r88 25 30 5.12336 $w=3.81e-07 $l=1.6e-07 $layer=LI1_cond $X=2.337 $Y=0.85
+ $X2=2.337 $Y2=1.01
r89 19 21 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.57 $Y=1.61
+ $X2=3.57 $Y2=2.165
r90 18 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.205 $Y=1.535
+ $X2=3.13 $Y2=1.535
r91 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.495 $Y=1.535
+ $X2=3.57 $Y2=1.61
r92 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.495 $Y=1.535
+ $X2=3.205 $Y2=1.535
r93 13 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.61
+ $X2=3.13 $Y2=1.535
r94 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.13 $Y=1.61
+ $X2=3.13 $Y2=2.165
r95 12 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.46
+ $X2=3.13 $Y2=1.535
r96 11 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1 $X2=3.13
+ $Y2=0.925
r97 11 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.13 $Y=1 $X2=3.13
+ $Y2=1.46
r98 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=0.85 $X2=3.13
+ $Y2=0.925
r99 7 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.13 $Y=0.85 $X2=3.13
+ $Y2=0.445
r100 6 29 38.8573 $w=3.56e-07 $l=1.95653e-07 $layer=POLY_cond $X=2.455 $Y=0.925
+ $X2=2.29 $Y2=0.992
r101 5 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=0.925
+ $X2=3.13 $Y2=0.925
r102 5 6 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.055 $Y=0.925 $X2=2.455
+ $Y2=0.925
r103 1 27 23.0368 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.19 $Y=0.81
+ $X2=2.19 $Y2=0.992
r104 1 3 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.19 $Y=0.81 $X2=2.19
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_791_264# 1 2 9 13 17 21 23 26 30 34 40 41
+ 44 46 47 48 51 54 55
c167 21 0 2.06462e-20 $X=8.985 $Y=0.445
r168 60 62 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=8.87 $Y=1.74
+ $X2=8.985 $Y2=1.74
r169 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.785 $Y=0.85
+ $X2=9.785 $Y2=0.85
r170 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.89 $Y=0.85
+ $X2=3.89 $Y2=0.85
r171 48 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.035 $Y=0.85
+ $X2=3.89 $Y2=0.85
r172 47 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.64 $Y=0.85
+ $X2=9.785 $Y2=0.85
r173 47 48 6.93687 $w=1.4e-07 $l=5.605e-06 $layer=MET1_cond $X=9.64 $Y=0.85
+ $X2=4.035 $Y2=0.85
r174 46 55 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=9.785 $Y=0.825
+ $X2=9.785 $Y2=0.85
r175 43 55 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=9.785 $Y=1.53
+ $X2=9.785 $Y2=0.85
r176 43 44 6.82437 $w=2.65e-07 $l=2.21346e-07 $layer=LI1_cond $X=9.785 $Y=1.53
+ $X2=9.71 $Y2=1.717
r177 41 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.485
+ $X2=4.09 $Y2=1.65
r178 41 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.485
+ $X2=4.09 $Y2=1.32
r179 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.485 $X2=4.09 $Y2=1.485
r180 37 51 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.89 $Y=1.32
+ $X2=3.89 $Y2=0.85
r181 36 40 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.89 $Y=1.485 $X2=4.09
+ $Y2=1.485
r182 36 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=1.485
+ $X2=3.89 $Y2=1.32
r183 32 46 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.715 $Y=0.66
+ $X2=9.715 $Y2=0.825
r184 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.715 $Y=0.66
+ $X2=9.715 $Y2=0.385
r185 28 44 6.82437 $w=2.65e-07 $l=1.88e-07 $layer=LI1_cond $X=9.71 $Y=1.905
+ $X2=9.71 $Y2=1.717
r186 28 30 2.88111 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=9.71 $Y=1.905
+ $X2=9.71 $Y2=1.99
r187 26 62 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=9.065 $Y=1.74
+ $X2=8.985 $Y2=1.74
r188 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.065
+ $Y=1.74 $X2=9.065 $Y2=1.74
r189 23 44 0.127723 $w=3.75e-07 $l=1.7e-07 $layer=LI1_cond $X=9.54 $Y=1.717
+ $X2=9.71 $Y2=1.717
r190 23 25 14.5976 $w=3.73e-07 $l=4.75e-07 $layer=LI1_cond $X=9.54 $Y=1.717
+ $X2=9.065 $Y2=1.717
r191 19 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.985 $Y=1.575
+ $X2=8.985 $Y2=1.74
r192 19 21 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=8.985 $Y=1.575
+ $X2=8.985 $Y2=0.445
r193 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.87 $Y=1.905
+ $X2=8.87 $Y2=1.74
r194 15 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.87 $Y=1.905
+ $X2=8.87 $Y2=2.275
r195 13 59 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.08 $Y=2.165
+ $X2=4.08 $Y2=1.65
r196 9 58 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.08 $Y=0.445
+ $X2=4.08 $Y2=1.32
r197 2 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.58
+ $Y=1.845 $X2=9.705 $Y2=1.99
r198 1 34 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=9.59
+ $Y=0.235 $X2=9.715 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_193_47# 1 2 9 11 15 17 19 22 26 27 30 31
+ 32 33 42 43 45 49 58 62
c196 43 0 2.06462e-20 $X=8.305 $Y=1.53
c197 33 0 1.37287e-19 $X=5.03 $Y=1.53
c198 32 0 3.76247e-20 $X=8.16 $Y=1.53
c199 22 0 1.92554e-19 $X=8.3 $Y=2.275
c200 11 0 1.43548e-19 $X=5.355 $Y=1.29
r201 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.385
+ $Y=1.74 $X2=8.385 $Y2=1.74
r202 55 58 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=8.3 $Y=1.74
+ $X2=8.385 $Y2=1.74
r203 48 50 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.88 $Y=1.35
+ $X2=4.88 $Y2=1.485
r204 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.88
+ $Y=1.35 $X2=4.88 $Y2=1.35
r205 45 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.88 $Y=1.29 $X2=4.88
+ $Y2=1.35
r206 43 59 7.56291 $w=3.18e-07 $l=2.1e-07 $layer=LI1_cond $X=8.31 $Y=1.53
+ $X2=8.31 $Y2=1.74
r207 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.305 $Y=1.53
+ $X2=8.305 $Y2=1.53
r208 40 49 10.7912 $w=1.83e-07 $l=1.8e-07 $layer=LI1_cond $X=4.887 $Y=1.53
+ $X2=4.887 $Y2=1.35
r209 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.885 $Y=1.53
+ $X2=4.885 $Y2=1.53
r210 36 66 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.1 $Y=1.53 $X2=1.1
+ $Y2=1.96
r211 36 62 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.1 $Y=1.53
+ $X2=1.1 $Y2=0.51
r212 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.53 $X2=1.1
+ $Y2=1.53
r213 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.03 $Y=1.53
+ $X2=4.885 $Y2=1.53
r214 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.16 $Y=1.53
+ $X2=8.305 $Y2=1.53
r215 32 33 3.87375 $w=1.4e-07 $l=3.13e-06 $layer=MET1_cond $X=8.16 $Y=1.53
+ $X2=5.03 $Y2=1.53
r216 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.53
+ $X2=1.1 $Y2=1.53
r217 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.74 $Y=1.53
+ $X2=4.885 $Y2=1.53
r218 30 31 4.32549 $w=1.4e-07 $l=3.495e-06 $layer=MET1_cond $X=4.74 $Y=1.53
+ $X2=1.245 $Y2=1.53
r219 29 43 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=8.31 $Y=1.035
+ $X2=8.31 $Y2=1.53
r220 27 51 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.09 $Y=0.87
+ $X2=7.98 $Y2=0.87
r221 26 29 5.41706 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.237 $Y=0.87
+ $X2=8.237 $Y2=1.035
r222 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=0.87 $X2=8.09 $Y2=0.87
r223 20 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.3 $Y=1.875
+ $X2=8.3 $Y2=1.74
r224 20 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.3 $Y=1.875 $X2=8.3
+ $Y2=2.275
r225 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.98 $Y=0.705
+ $X2=7.98 $Y2=0.87
r226 17 19 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.98 $Y=0.705
+ $X2=7.98 $Y2=0.415
r227 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.43 $Y=1.215
+ $X2=5.43 $Y2=0.415
r228 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.045 $Y=1.29
+ $X2=4.88 $Y2=1.29
r229 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.355 $Y=1.29
+ $X2=5.43 $Y2=1.215
r230 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=5.355 $Y=1.29
+ $X2=5.045 $Y2=1.29
r231 9 50 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.855 $Y=2.275
+ $X2=4.855 $Y2=1.485
r232 2 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r233 1 62 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_1150_159# 1 2 9 13 17 21 25 27 28 32 36
+ 40 41 47 55
c118 40 0 6.28645e-20 $X=7.36 $Y=1.21
r119 49 50 5.12431 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=6.732 $Y=1.21
+ $X2=6.732 $Y2=1.375
r120 45 55 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=5.955 $Y=0.93
+ $X2=5.96 $Y2=0.93
r121 45 52 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=5.955 $Y=0.93
+ $X2=5.825 $Y2=0.93
r122 44 47 4.13427 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.955 $Y=0.93
+ $X2=6.07 $Y2=0.93
r123 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.955
+ $Y=0.93 $X2=5.955 $Y2=0.93
r124 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.36
+ $Y=1.21 $X2=7.36 $Y2=1.21
r125 38 49 1.93884 $w=3.3e-07 $l=2.03e-07 $layer=LI1_cond $X=6.935 $Y=1.21
+ $X2=6.732 $Y2=1.21
r126 38 40 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=6.935 $Y=1.21
+ $X2=7.36 $Y2=1.21
r127 36 50 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.695 $Y=1.88
+ $X2=6.695 $Y2=1.375
r128 30 32 10.6708 $w=4.03e-07 $l=3.75e-07 $layer=LI1_cond $X=6.732 $Y=0.765
+ $X2=6.732 $Y2=0.39
r129 28 49 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=6.732 $Y=0.915
+ $X2=6.732 $Y2=1.21
r130 28 30 4.26831 $w=4.03e-07 $l=1.5e-07 $layer=LI1_cond $X=6.732 $Y=0.915
+ $X2=6.732 $Y2=0.765
r131 28 47 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.53 $Y=0.915
+ $X2=6.07 $Y2=0.915
r132 26 41 6.10776 $w=2.75e-07 $l=2.8e-08 $layer=POLY_cond $X=7.362 $Y=1.238
+ $X2=7.362 $Y2=1.21
r133 26 27 42.1909 $w=2.75e-07 $l=1.37e-07 $layer=POLY_cond $X=7.362 $Y=1.238
+ $X2=7.362 $Y2=1.375
r134 25 41 35.9921 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.362 $Y=1.045
+ $X2=7.362 $Y2=1.21
r135 24 25 45.0266 $w=2.75e-07 $l=1.5e-07 $layer=POLY_cond $X=7.397 $Y=0.895
+ $X2=7.397 $Y2=1.045
r136 21 24 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.495 $Y=0.445
+ $X2=7.495 $Y2=0.895
r137 17 27 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=7.425 $Y=2.275
+ $X2=7.425 $Y2=1.375
r138 11 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.96 $Y=0.795
+ $X2=5.96 $Y2=0.93
r139 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.96 $Y=0.795
+ $X2=5.96 $Y2=0.445
r140 7 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.825 $Y=1.065
+ $X2=5.825 $Y2=0.93
r141 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.825 $Y=1.065
+ $X2=5.825 $Y2=2.275
r142 2 36 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.56
+ $Y=1.735 $X2=6.695 $Y2=1.88
r143 1 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.63
+ $Y=0.235 $X2=6.765 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_986_413# 1 2 8 11 15 16 17 18 19 20 24 29
+ 31 33
c106 29 0 1.40584e-19 $X=5.595 $Y=1.315
c107 17 0 6.28645e-20 $X=6.52 $Y=1.1
r108 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.275
+ $Y=1.41 $X2=6.275 $Y2=1.41
r109 33 35 20.25 $w=2.44e-07 $l=4.05e-07 $layer=LI1_cond $X=5.87 $Y=1.41
+ $X2=6.275 $Y2=1.41
r110 30 33 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.87 $Y=1.575
+ $X2=5.87 $Y2=1.41
r111 30 31 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.87 $Y=1.575
+ $X2=5.87 $Y2=2.175
r112 29 33 13.75 $w=2.44e-07 $l=2.75e-07 $layer=LI1_cond $X=5.595 $Y=1.41
+ $X2=5.87 $Y2=1.41
r113 28 29 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.595 $Y=0.565
+ $X2=5.595 $Y2=1.315
r114 24 28 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.51 $Y=0.41
+ $X2=5.595 $Y2=0.565
r115 24 26 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=5.51 $Y=0.41
+ $X2=5.2 $Y2=0.41
r116 20 31 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.785 $Y=2.275
+ $X2=5.87 $Y2=2.175
r117 20 22 39.0955 $w=1.98e-07 $l=7.05e-07 $layer=LI1_cond $X=5.785 $Y=2.275
+ $X2=5.08 $Y2=2.275
r118 18 36 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.41 $Y=1.41
+ $X2=6.275 $Y2=1.41
r119 18 19 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.41 $Y=1.41
+ $X2=6.485 $Y2=1.41
r120 16 17 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.52 $Y=0.95
+ $X2=6.52 $Y2=1.1
r121 15 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.555 $Y=0.555
+ $X2=6.555 $Y2=0.95
r122 9 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.485 $Y=1.545
+ $X2=6.485 $Y2=1.41
r123 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.485 $Y=1.545
+ $X2=6.485 $Y2=2.11
r124 8 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.485 $Y=1.275
+ $X2=6.485 $Y2=1.41
r125 8 17 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.485 $Y=1.275
+ $X2=6.485 $Y2=1.1
r126 2 22 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=2.065 $X2=5.08 $Y2=2.275
r127 1 26 182 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_NDIFF $count=1 $X=5.065
+ $Y=0.235 $X2=5.2 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_1591_413# 1 2 9 13 15 17 19 22 24 25 26
+ 27 31 36 38 41 44
c110 44 0 1.78258e-19 $X=8.725 $Y=1.16
r111 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.425
+ $Y=1.16 $X2=9.425 $Y2=1.16
r112 39 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=1.16
+ $X2=8.725 $Y2=1.16
r113 39 41 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=8.81 $Y=1.16
+ $X2=9.425 $Y2=1.16
r114 37 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=1.325
+ $X2=8.725 $Y2=1.16
r115 37 38 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.725 $Y=1.325
+ $X2=8.725 $Y2=2.165
r116 36 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=0.995
+ $X2=8.725 $Y2=1.16
r117 35 36 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.725 $Y=0.535
+ $X2=8.725 $Y2=0.995
r118 31 35 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=8.64 $Y=0.432
+ $X2=8.725 $Y2=0.535
r119 31 33 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=8.64 $Y=0.432
+ $X2=8.205 $Y2=0.432
r120 27 38 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.64 $Y=2.26
+ $X2=8.725 $Y2=2.165
r121 27 29 32.1053 $w=1.88e-07 $l=5.5e-07 $layer=LI1_cond $X=8.64 $Y=2.26
+ $X2=8.09 $Y2=2.26
r122 24 42 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=9.85 $Y=1.16
+ $X2=9.425 $Y2=1.16
r123 24 25 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.85 $Y=1.16
+ $X2=9.925 $Y2=1.16
r124 20 26 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.41 $Y=1.325
+ $X2=10.41 $Y2=1.16
r125 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.41 $Y=1.325
+ $X2=10.41 $Y2=1.985
r126 17 26 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.41 $Y=0.995
+ $X2=10.41 $Y2=1.16
r127 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.41 $Y=0.995
+ $X2=10.41 $Y2=0.56
r128 16 25 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10 $Y=1.16
+ $X2=9.925 $Y2=1.16
r129 15 26 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.335 $Y=1.16
+ $X2=10.41 $Y2=1.16
r130 15 16 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=10.335 $Y=1.16
+ $X2=10 $Y2=1.16
r131 11 25 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.925 $Y=1.325
+ $X2=9.925 $Y2=1.16
r132 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.925 $Y=1.325
+ $X2=9.925 $Y2=2.165
r133 7 25 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.925 $Y=0.995
+ $X2=9.925 $Y2=1.16
r134 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=9.925 $Y=0.995
+ $X2=9.925 $Y2=0.445
r135 2 29 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=7.955
+ $Y=2.065 $X2=8.09 $Y2=2.26
r136 1 33 182 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_NDIFF $count=1 $X=8.055
+ $Y=0.235 $X2=8.205 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 38 42 46 50
+ 55 56 58 59 61 62 63 65 77 81 97 98 101 104 107 110
c156 98 0 1.8506e-19 $X=10.81 $Y=2.72
c157 32 0 1.67735e-19 $X=3.35 $Y=1.99
c158 1 0 5.65522e-20 $X=0.545 $Y=1.815
r159 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r160 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r161 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r162 104 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r163 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r164 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r165 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r166 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r167 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r168 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r169 89 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.97 $Y2=2.72
r170 89 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r171 88 91 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=8.97 $Y2=2.72
r172 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r173 86 110 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.36 $Y=2.72
+ $X2=7.215 $Y2=2.72
r174 86 88 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.36 $Y=2.72
+ $X2=7.59 $Y2=2.72
r175 85 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r176 85 105 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.45 $Y2=2.72
r177 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r178 82 104 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.46 $Y=2.72
+ $X2=3.362 $Y2=2.72
r179 82 84 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=3.46 $Y=2.72
+ $X2=5.75 $Y2=2.72
r180 81 107 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.125 $Y=2.72
+ $X2=6.242 $Y2=2.72
r181 81 84 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.125 $Y=2.72
+ $X2=5.75 $Y2=2.72
r182 80 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r183 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r184 77 104 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.362 $Y2=2.72
r185 77 79 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=2.99 $Y2=2.72
r186 76 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r187 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r188 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r189 73 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r190 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r191 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r192 70 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r193 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r194 65 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r195 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r196 63 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r197 63 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r198 61 94 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=10.05 $Y=2.72
+ $X2=9.89 $Y2=2.72
r199 61 62 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=10.05 $Y=2.72
+ $X2=10.172 $Y2=2.72
r200 60 97 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=10.295 $Y=2.72
+ $X2=10.81 $Y2=2.72
r201 60 62 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=10.295 $Y=2.72
+ $X2=10.172 $Y2=2.72
r202 58 91 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.98 $Y=2.72
+ $X2=8.97 $Y2=2.72
r203 58 59 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.98 $Y=2.72
+ $X2=9.11 $Y2=2.72
r204 57 94 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.24 $Y=2.72
+ $X2=9.89 $Y2=2.72
r205 57 59 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.24 $Y=2.72
+ $X2=9.11 $Y2=2.72
r206 55 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r207 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.4 $Y2=2.72
r208 54 79 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.99 $Y2=2.72
r209 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.4 $Y2=2.72
r210 50 53 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=10.172 $Y=1.63
+ $X2=10.172 $Y2=1.97
r211 48 62 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.172 $Y=2.635
+ $X2=10.172 $Y2=2.72
r212 48 53 31.2806 $w=2.43e-07 $l=6.65e-07 $layer=LI1_cond $X=10.172 $Y=2.635
+ $X2=10.172 $Y2=1.97
r213 44 59 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.11 $Y=2.635
+ $X2=9.11 $Y2=2.72
r214 44 46 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=9.11 $Y=2.635
+ $X2=9.11 $Y2=2.3
r215 40 110 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=2.635
+ $X2=7.215 $Y2=2.72
r216 40 42 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.215 $Y=2.635
+ $X2=7.215 $Y2=2.275
r217 39 107 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.242 $Y2=2.72
r218 38 110 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.07 $Y=2.72
+ $X2=7.215 $Y2=2.72
r219 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.07 $Y=2.72
+ $X2=6.36 $Y2=2.72
r220 34 107 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.242 $Y=2.635
+ $X2=6.242 $Y2=2.72
r221 34 36 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=6.242 $Y=2.635
+ $X2=6.242 $Y2=2
r222 30 104 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.362 $Y=2.635
+ $X2=3.362 $Y2=2.72
r223 30 32 36.6853 $w=1.93e-07 $l=6.45e-07 $layer=LI1_cond $X=3.362 $Y=2.635
+ $X2=3.362 $Y2=1.99
r224 26 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.635 $X2=2.4
+ $Y2=2.72
r225 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2
r226 22 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r227 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r228 7 53 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=10
+ $Y=1.845 $X2=10.2 $Y2=1.97
r229 7 50 600 $w=1.7e-07 $l=2.98706e-07 $layer=licon1_PDIFF $count=1 $X=10
+ $Y=1.845 $X2=10.2 $Y2=1.63
r230 6 46 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=2.065 $X2=9.085 $Y2=2.3
r231 5 42 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=7.09
+ $Y=2.065 $X2=7.215 $Y2=2.275
r232 4 36 300 $w=1.7e-07 $l=3.76098e-07 $layer=licon1_PDIFF $count=2 $X=5.9
+ $Y=2.065 $X2=6.245 $Y2=2
r233 3 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=1.845 $X2=3.35 $Y2=1.99
r234 2 28 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.845 $X2=2.4 $Y2=2
r235 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%A_299_47# 1 2 3 4 20 21 24 25 29 36 38 40
+ 43 48
c120 38 0 1.82232e-19 $X=4.27 $Y=0.51
r121 38 40 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.27 $Y=0.51
+ $X2=4.125 $Y2=0.51
r122 38 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.27 $Y=0.51
+ $X2=4.27 $Y2=0.51
r123 36 40 2.17465 $w=1.85e-07 $l=2.54e-06 $layer=MET1_cond $X=1.585 $Y=0.487
+ $X2=4.125 $Y2=0.487
r124 34 48 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.44 $Y=0.385
+ $X2=1.62 $Y2=0.385
r125 33 36 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.44 $Y=0.51
+ $X2=1.585 $Y2=0.51
r126 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.44 $Y=0.51
+ $X2=1.44 $Y2=0.51
r127 28 43 22.8354 $w=2.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.28 $Y=0.98
+ $X2=4.28 $Y2=0.445
r128 28 29 8.82932 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.33 $Y=0.98
+ $X2=4.33 $Y2=1.15
r129 25 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.43 $Y=1.82
+ $X2=4.43 $Y2=1.15
r130 24 25 9.05087 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=4.32 $Y=2 $X2=4.32
+ $Y2=1.82
r131 20 21 7.04283 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=1.57 $Y=1.99 $X2=1.57
+ $Y2=1.89
r132 13 34 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.44 $Y=0.515
+ $X2=1.44 $Y2=0.385
r133 13 21 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=1.44 $Y=0.515
+ $X2=1.44 $Y2=1.89
r134 4 24 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=4.155
+ $Y=1.845 $X2=4.29 $Y2=2
r135 3 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r136 2 43 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.235 $X2=4.29 $Y2=0.445
r137 1 48 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%Q 1 2 7 10
r17 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.63 $Y=1.63
+ $X2=10.63 $Y2=2.31
r18 7 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=10.63 $Y=1.19
+ $X2=10.63 $Y2=1.63
r19 7 10 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=10.63 $Y=1.19
+ $X2=10.63 $Y2=0.395
r20 2 17 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.485
+ $Y=1.485 $X2=10.63 $Y2=2.31
r21 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.485
+ $Y=1.485 $X2=10.63 $Y2=1.63
r22 1 10 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=10.485
+ $Y=0.235 $X2=10.63 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__EDFXTP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 48 53
+ 54 56 57 59 60 62 63 64 66 78 82 101 102 105 108 111
c170 102 0 2.71124e-20 $X=10.81 $Y=0
c171 82 0 1.82232e-19 $X=5.945 $Y=0
r172 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r173 108 109 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r174 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r175 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r176 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r177 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r178 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r179 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r180 93 96 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.97 $Y2=0
r181 92 95 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.59 $Y=0 $X2=8.97
+ $Y2=0
r182 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r183 90 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r184 90 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.21 $Y2=0
r185 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r186 87 111 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.142 $Y2=0
r187 87 89 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=7.13
+ $Y2=0
r188 86 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r189 86 109 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=3.45 $Y2=0
r190 85 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r191 83 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=3.35 $Y2=0
r192 83 85 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=5.75 $Y2=0
r193 82 111 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=6.142 $Y2=0
r194 82 85 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=5.75 $Y2=0
r195 81 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.45 $Y2=0
r196 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r197 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.35 $Y2=0
r198 78 80 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=2.99 $Y2=0
r199 77 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r200 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r201 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r202 74 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r203 73 76 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r204 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r205 71 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r206 71 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r207 66 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r208 66 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r209 64 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r210 64 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r211 62 98 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=10.05 $Y=0 $X2=9.89
+ $Y2=0
r212 62 63 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=10.05 $Y=0
+ $X2=10.172 $Y2=0
r213 61 101 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=10.295 $Y=0
+ $X2=10.81 $Y2=0
r214 61 63 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=10.295 $Y=0
+ $X2=10.172 $Y2=0
r215 59 95 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=9.05 $Y=0 $X2=8.97
+ $Y2=0
r216 59 60 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=9.05 $Y=0 $X2=9.207
+ $Y2=0
r217 58 98 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.365 $Y=0
+ $X2=9.89 $Y2=0
r218 58 60 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=9.365 $Y=0
+ $X2=9.207 $Y2=0
r219 56 89 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.165 $Y=0 $X2=7.13
+ $Y2=0
r220 56 57 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=7.302 $Y2=0
r221 55 92 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.59
+ $Y2=0
r222 55 57 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.302
+ $Y2=0
r223 53 76 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0
+ $X2=2.07 $Y2=0
r224 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.4
+ $Y2=0
r225 52 80 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=0
+ $X2=2.99 $Y2=0
r226 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.4
+ $Y2=0
r227 48 50 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=10.172 $Y=0.395
+ $X2=10.172 $Y2=0.735
r228 46 63 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.172 $Y=0.085
+ $X2=10.172 $Y2=0
r229 46 48 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=10.172 $Y=0.085
+ $X2=10.172 $Y2=0.395
r230 42 60 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=9.207 $Y=0.085
+ $X2=9.207 $Y2=0
r231 42 44 13.3537 $w=3.13e-07 $l=3.65e-07 $layer=LI1_cond $X=9.207 $Y=0.085
+ $X2=9.207 $Y2=0.45
r232 38 57 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.302 $Y=0.085
+ $X2=7.302 $Y2=0
r233 38 40 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=7.302 $Y=0.085
+ $X2=7.302 $Y2=0.45
r234 34 111 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.142 $Y=0.085
+ $X2=6.142 $Y2=0
r235 34 36 9.77388 $w=3.93e-07 $l=3.35e-07 $layer=LI1_cond $X=6.142 $Y=0.085
+ $X2=6.142 $Y2=0.42
r236 30 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r237 30 32 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.445
r238 26 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=0.085 $X2=2.4
+ $Y2=0
r239 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.4 $Y=0.085
+ $X2=2.4 $Y2=0.38
r240 22 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r241 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r242 7 50 182 $w=1.7e-07 $l=5.91608e-07 $layer=licon1_NDIFF $count=1 $X=10
+ $Y=0.235 $X2=10.2 $Y2=0.735
r243 7 48 182 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_NDIFF $count=1 $X=10
+ $Y=0.235 $X2=10.2 $Y2=0.395
r244 6 44 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=9.06
+ $Y=0.235 $X2=9.195 $Y2=0.45
r245 5 40 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.235 $X2=7.285 $Y2=0.45
r246 4 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.035
+ $Y=0.235 $X2=6.175 $Y2=0.42
r247 3 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.35 $Y2=0.445
r248 2 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.38
r249 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


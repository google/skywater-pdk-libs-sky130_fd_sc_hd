* File: sky130_fd_sc_hd__o311a_2.spice
* Created: Thu Aug 27 14:39:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o311a_2.pex.spice"
.subckt sky130_fd_sc_hd__o311a_2  VNB VPB A1 A2 A3 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_91_21#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.208 AS=0.08775 PD=1.94 PS=0.92 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_91_21#_M1011_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.203125 AS=0.08775 PD=1.275 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1013 N_A_360_47#_M1013_d N_A1_M1013_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.203125 PD=1 PS=1.275 NRD=5.532 NRS=1.836 M=1 R=4.33333
+ SA=75001.4 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g N_A_360_47#_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1365 AS=0.11375 PD=1.07 PS=1 NRD=12.912 NRS=7.38 M=1 R=4.33333 SA=75001.9
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_A_360_47#_M1005_d N_A3_M1005_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.1365 PD=1.015 PS=1.07 NRD=8.304 NRS=12.912 M=1 R=4.33333
+ SA=75002.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 A_677_47# N_B1_M1006_g N_A_360_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.118625 PD=0.86 PS=1.015 NRD=9.228 NRS=7.38 M=1 R=4.33333
+ SA=75003 SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1008 N_A_91_21#_M1008_d N_C1_M1008_g A_677_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.06825 PD=1.82 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75003.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_91_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.32 AS=0.135 PD=2.64 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.3 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_91_21#_M1007_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3125 AS=0.135 PD=1.625 PS=1.27 NRD=25.5903 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1000 A_360_297# N_A1_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1 AD=0.175
+ AS=0.3125 PD=1.35 PS=1.625 NRD=23.6203 NRS=42.3353 M=1 R=6.66667 SA=75001.4
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1004 A_460_297# N_A2_M1004_g A_360_297# VPB PHIGHVT L=0.15 W=1 AD=0.21
+ AS=0.175 PD=1.42 PS=1.35 NRD=30.5153 NRS=23.6203 M=1 R=6.66667 SA=75001.9
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1001 N_A_91_21#_M1001_d N_A3_M1001_g A_460_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.21 PD=1.275 PS=1.42 NRD=0 NRS=30.5153 M=1 R=6.66667 SA=75002.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_B1_M1010_g N_A_91_21#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.1375 PD=1.3 PS=1.275 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_91_21#_M1003_d N_C1_M1003_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.15 PD=2.52 PS=1.3 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75003.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__o311a_2.pxi.spice"
*
.ends
*
*

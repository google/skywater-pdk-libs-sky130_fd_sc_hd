* File: sky130_fd_sc_hd__dlxbn_1.spice.pex
* Created: Thu Aug 27 14:17:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLXBN_1%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39414e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.21 $Y=1.19
+ $X2=0.21 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%A_27_47# 1 2 9 13 15 17 21 25 29 30 31 35 43
+ 46 48 51 52 55 58 59 63 67 72
c157 72 0 1.70289e-19 $X=3.12 $Y=1.415
c158 35 0 1.57777e-19 $X=2.95 $Y=0.87
c159 13 0 2.69707e-20 $X=0.89 $Y=2.135
c160 9 0 2.69707e-20 $X=0.89 $Y=0.445
r161 67 69 16.1264 $w=2.69e-07 $l=9e-08 $layer=POLY_cond $X=3.205 $Y=1.745
+ $X2=3.295 $Y2=1.745
r162 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.745 $X2=3.205 $Y2=1.745
r163 59 68 7.28751 $w=3.38e-07 $l=2.15e-07 $layer=LI1_cond $X=3.12 $Y=1.53
+ $X2=3.12 $Y2=1.745
r164 59 72 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.53
+ $X2=3.12 $Y2=1.415
r165 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.04 $Y=1.53
+ $X2=3.04 $Y2=1.53
r166 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r167 52 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r168 51 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.895 $Y=1.53
+ $X2=3.04 $Y2=1.53
r169 51 52 2.54331 $w=1.4e-07 $l=2.055e-06 $layer=MET1_cond $X=2.895 $Y=1.53
+ $X2=0.84 $Y2=1.53
r170 50 55 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r171 49 55 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r172 47 63 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r173 46 49 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r174 46 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r175 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r176 40 72 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.035 $Y=1.035
+ $X2=3.035 $Y2=1.415
r177 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=0.91 $X2=2.75 $Y2=0.91
r178 35 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.95 $Y=0.87
+ $X2=3.035 $Y2=1.035
r179 35 37 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.95 $Y=0.87 $X2=2.75
+ $Y2=0.87
r180 33 48 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r181 32 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r182 31 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r183 31 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r184 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r185 29 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r186 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r187 23 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r188 19 69 16.4183 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.295 $Y=1.88
+ $X2=3.295 $Y2=1.745
r189 19 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.295 $Y=1.88
+ $X2=3.295 $Y2=2.275
r190 15 38 40.7934 $w=3.34e-07 $l=1.8735e-07 $layer=POLY_cond $X=2.725 $Y=0.73
+ $X2=2.74 $Y2=0.91
r191 15 17 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.725 $Y=0.73
+ $X2=2.725 $Y2=0.415
r192 11 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r193 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r194 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r195 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r196 2 43 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r197 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%D 1 3 5 8 10 11 12 16
c49 11 0 1.27156e-19 $X=1.822 $Y=1.715
c50 1 0 1.29183e-19 $X=1.79 $Y=1.205
r51 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.04 $X2=1.61 $Y2=1.04
r52 12 16 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.615 $Y=1.19
+ $X2=1.615 $Y2=1.04
r53 10 11 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=1.822 $Y=1.565
+ $X2=1.822 $Y2=1.715
r54 8 11 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.855 $Y=2.165
+ $X2=1.855 $Y2=1.715
r55 3 15 60.1993 $w=3.23e-07 $l=3.73497e-07 $layer=POLY_cond $X=1.83 $Y=0.73
+ $X2=1.69 $Y2=1.04
r56 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.73 $X2=1.83
+ $Y2=0.445
r57 1 15 38.5615 $w=3.23e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.79 $Y=1.205
+ $X2=1.69 $Y2=1.04
r58 1 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.79 $Y=1.205
+ $X2=1.79 $Y2=1.565
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%A_299_47# 1 2 9 11 13 17 19 21 22 23 24 26
c91 23 0 1.52561e-19 $X=2.08 $Y=1.235
c92 11 0 1.57777e-19 $X=2.275 $Y=1.235
r93 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.215
+ $Y=1.07 $X2=2.215 $Y2=1.07
r94 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r95 23 32 9.08131 $w=2.76e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.08 $Y=1.235
+ $X2=2.18 $Y2=1.07
r96 23 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.08 $Y=1.235
+ $X2=2.08 $Y2=1.495
r97 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.995 $Y=1.58
+ $X2=2.08 $Y2=1.495
r98 21 22 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.995 $Y=1.58
+ $X2=1.81 $Y2=1.58
r99 20 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r100 19 32 16.3551 $w=2.76e-07 $l=4.53156e-07 $layer=LI1_cond $X=1.995 $Y=0.7
+ $X2=2.18 $Y2=1.07
r101 19 20 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.995 $Y=0.7
+ $X2=1.705 $Y2=0.7
r102 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.81 $Y2=1.58
r103 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.99
r104 11 33 38.9235 $w=2.69e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.275 $Y=1.235
+ $X2=2.215 $Y2=1.07
r105 11 13 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.275 $Y=1.235
+ $X2=2.275 $Y2=2.165
r106 7 33 38.9235 $w=2.69e-07 $l=1.81659e-07 $layer=POLY_cond $X=2.25 $Y=0.905
+ $X2=2.215 $Y2=1.07
r107 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.25 $Y=0.905
+ $X2=2.25 $Y2=0.445
r108 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.52
+ $Y=1.845 $X2=1.645 $Y2=1.99
r109 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%A_193_47# 1 2 9 11 13 15 18 20 22 23 26 29
+ 34 35
c105 35 0 1.52561e-19 $X=2.755 $Y=1.42
c106 20 0 1.27156e-19 $X=1.127 $Y=1.797
r107 33 35 10.791 $w=2.68e-07 $l=6e-08 $layer=POLY_cond $X=2.695 $Y=1.42
+ $X2=2.755 $Y2=1.42
r108 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.52 $X2=2.695 $Y2=1.52
r109 30 34 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.637 $Y=1.87
+ $X2=2.637 $Y2=1.52
r110 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.58 $Y=1.87
+ $X2=2.58 $Y2=1.87
r111 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r112 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r113 22 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.435 $Y=1.87
+ $X2=2.58 $Y2=1.87
r114 22 23 1.4047 $w=1.4e-07 $l=1.135e-06 $layer=MET1_cond $X=2.435 $Y=1.87
+ $X2=1.3 $Y2=1.87
r115 20 26 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r116 20 21 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r117 18 21 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r118 15 35 82.7313 $w=2.68e-07 $l=5.69473e-07 $layer=POLY_cond $X=3.215 $Y=1.175
+ $X2=2.755 $Y2=1.42
r119 14 15 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.215 $Y=0.785
+ $X2=3.215 $Y2=1.175
r120 11 14 28.5207 $w=1.69e-07 $l=1.16189e-07 $layer=POLY_cond $X=3.18 $Y=0.685
+ $X2=3.215 $Y2=0.785
r121 11 13 86.76 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.18 $Y=0.685
+ $X2=3.18 $Y2=0.415
r122 7 35 16.3317 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.755 $Y=1.685
+ $X2=2.755 $Y2=1.42
r123 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.755 $Y=1.685
+ $X2=2.755 $Y2=2.275
r124 2 26 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r125 1 18 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%A_716_21# 1 2 9 13 15 17 20 22 24 26 28 31
+ 33 34 35 38 42 44 45 47 50 51 56 57
c112 51 0 1.10692e-19 $X=5.055 $Y=1.16
c113 34 0 1.94082e-19 $X=5.952 $Y=1.77
c114 24 0 7.57733e-20 $X=5.95 $Y=1.325
r115 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.16 $X2=5.055 $Y2=1.16
r116 48 57 0.63164 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=4.58 $Y=1.16
+ $X2=4.487 $Y2=1.16
r117 48 50 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=4.58 $Y=1.16
+ $X2=5.055 $Y2=1.16
r118 47 56 7.19657 $w=2.17e-07 $l=1.87e-07 $layer=LI1_cond $X=4.487 $Y=1.535
+ $X2=4.3 $Y2=1.535
r119 46 57 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=4.487 $Y=1.325
+ $X2=4.487 $Y2=1.16
r120 46 47 12.5897 $w=1.83e-07 $l=2.1e-07 $layer=LI1_cond $X=4.487 $Y=1.325
+ $X2=4.487 $Y2=1.535
r121 45 57 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=4.487 $Y=0.995
+ $X2=4.487 $Y2=1.16
r122 44 54 14.9708 $w=2.16e-07 $l=2.82524e-07 $layer=LI1_cond $X=4.487 $Y=0.84
+ $X2=4.44 $Y2=0.58
r123 44 45 9.29238 $w=1.83e-07 $l=1.55e-07 $layer=LI1_cond $X=4.487 $Y=0.84
+ $X2=4.487 $Y2=0.995
r124 40 56 7.19657 $w=2.17e-07 $l=3.87492e-07 $layer=LI1_cond $X=4.425 $Y=1.865
+ $X2=4.3 $Y2=1.535
r125 40 42 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=4.425 $Y=1.865
+ $X2=4.425 $Y2=2.27
r126 38 58 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.885 $Y=1.7
+ $X2=3.655 $Y2=1.7
r127 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.885
+ $Y=1.7 $X2=3.885 $Y2=1.7
r128 35 56 0.105856 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=1.7 $X2=4.3
+ $Y2=1.535
r129 35 37 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.3 $Y=1.7
+ $X2=3.885 $Y2=1.7
r130 33 34 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=5.952 $Y=1.62
+ $X2=5.952 $Y2=1.77
r131 31 34 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.955 $Y=2.165
+ $X2=5.955 $Y2=1.77
r132 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.955 $Y=0.73
+ $X2=5.955 $Y2=0.445
r133 24 33 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.62
r134 23 51 5.03009 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.005 $Y2=1.16
r135 22 24 52.6689 $w=1.51e-07 $l=1.65997e-07 $layer=POLY_cond $X=5.952 $Y=1.16
+ $X2=5.95 $Y2=1.325
r136 22 26 137.258 $w=1.51e-07 $l=4.31497e-07 $layer=POLY_cond $X=5.952 $Y=1.16
+ $X2=5.955 $Y2=0.73
r137 22 23 137.266 $w=3.3e-07 $l=7.85e-07 $layer=POLY_cond $X=5.875 $Y=1.16
+ $X2=5.09 $Y2=1.16
r138 18 51 37.0704 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=5.015 $Y=1.325
+ $X2=5.005 $Y2=1.16
r139 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.015 $Y=1.325
+ $X2=5.015 $Y2=1.985
r140 15 51 37.0704 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=5.015 $Y=0.995
+ $X2=5.005 $Y2=1.16
r141 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.015 $Y=0.995
+ $X2=5.015 $Y2=0.56
r142 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.865
+ $X2=3.655 $Y2=1.7
r143 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.655 $Y=1.865
+ $X2=3.655 $Y2=2.275
r144 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.535
+ $X2=3.655 $Y2=1.7
r145 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.655 $Y=1.535
+ $X2=3.655 $Y2=0.445
r146 2 56 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.26
+ $Y=1.485 $X2=4.385 $Y2=1.755
r147 2 42 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.26
+ $Y=1.485 $X2=4.385 $Y2=2.27
r148 1 54 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.235 $X2=4.385 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%A_560_47# 1 2 7 9 12 14 15 16 20 25 27 30 33
c87 33 0 1.56164e-19 $X=3.355 $Y=0.995
c88 30 0 1.10692e-19 $X=4.14 $Y=1.16
c89 15 0 1.26672e-19 $X=4.595 $Y=1.16
r90 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.16 $X2=4.14 $Y2=1.16
r91 28 33 0.89609 $w=3.3e-07 $l=3.47851e-07 $layer=LI1_cond $X=3.63 $Y=1.16
+ $X2=3.355 $Y2=0.995
r92 28 30 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.63 $Y=1.16
+ $X2=4.14 $Y2=1.16
r93 27 34 2.65936 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.545 $Y=2.015
+ $X2=3.545 $Y2=2.145
r94 26 33 8.61065 $w=1.7e-07 $l=4.14246e-07 $layer=LI1_cond $X=3.545 $Y=1.325
+ $X2=3.355 $Y2=0.995
r95 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.545 $Y=1.325
+ $X2=3.545 $Y2=2.015
r96 25 33 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0.995
+ $X2=3.355 $Y2=0.995
r97 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.44 $Y=0.535
+ $X2=3.44 $Y2=0.995
r98 20 34 10.5376 $w=2.36e-07 $l=2.06277e-07 $layer=LI1_cond $X=3.36 $Y=2.19
+ $X2=3.545 $Y2=2.145
r99 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.36 $Y=2.19
+ $X2=3.085 $Y2=2.19
r100 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.355 $Y=0.45
+ $X2=3.44 $Y2=0.535
r101 16 18 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.355 $Y=0.45
+ $X2=2.955 $Y2=0.45
r102 14 31 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=4.52 $Y=1.16
+ $X2=4.14 $Y2=1.16
r103 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.52 $Y=1.16
+ $X2=4.595 $Y2=1.16
r104 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=1.325
+ $X2=4.595 $Y2=1.16
r105 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.595 $Y=1.325
+ $X2=4.595 $Y2=1.985
r106 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=0.995
+ $X2=4.595 $Y2=1.16
r107 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.595 $Y=0.995
+ $X2=4.595 $Y2=0.56
r108 2 22 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=2.065 $X2=3.085 $Y2=2.19
r109 1 18 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.955 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%A_1124_47# 1 2 9 12 16 20 24 25 27 29
c45 24 0 1.94082e-19 $X=6.37 $Y=1.16
r46 25 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=1.16
+ $X2=6.37 $Y2=1.325
r47 25 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=1.16
+ $X2=6.37 $Y2=0.995
r48 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.37
+ $Y=1.16 $X2=6.37 $Y2=1.16
r49 22 27 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.91 $Y=1.16
+ $X2=5.785 $Y2=1.16
r50 22 24 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.91 $Y=1.16
+ $X2=6.37 $Y2=1.16
r51 18 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=1.325
+ $X2=5.785 $Y2=1.16
r52 18 20 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=5.785 $Y=1.325
+ $X2=5.785 $Y2=2.165
r53 14 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0.995
+ $X2=5.785 $Y2=1.16
r54 14 16 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=5.785 $Y=0.995
+ $X2=5.785 $Y2=0.51
r55 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.985
+ $X2=6.43 $Y2=1.325
r56 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.56 $X2=6.43
+ $Y2=0.995
r57 2 20 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=1.845 $X2=5.745 $Y2=2.165
r58 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=5.62
+ $Y=0.235 $X2=5.745 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 39 41 46
+ 58 62 69 70 73 76 79 82
r106 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r107 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r110 70 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r112 67 82 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.237 $Y2=2.72
r113 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.67 $Y2=2.72
r114 66 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 66 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r116 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r117 63 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.97 $Y=2.72
+ $X2=4.845 $Y2=2.72
r118 63 65 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.97 $Y=2.72
+ $X2=5.75 $Y2=2.72
r119 62 82 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=6.237 $Y2=2.72
r120 62 65 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=5.75 $Y2=2.72
r121 61 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r122 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r123 58 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.845 $Y2=2.72
r124 58 60 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 57 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r126 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r127 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 54 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r129 53 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r130 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r131 51 76 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.137 $Y2=2.72
r132 51 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.53 $Y2=2.72
r133 50 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 50 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r136 47 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r137 47 49 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r138 46 76 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=2.137 $Y2=2.72
r139 46 49 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 41 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r141 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r142 39 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r143 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r144 37 56 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.45 $Y2=2.72
r145 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.865 $Y2=2.72
r146 36 60 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.95 $Y=2.72
+ $X2=4.37 $Y2=2.72
r147 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=2.72
+ $X2=3.865 $Y2=2.72
r148 32 82 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.237 $Y=2.635
+ $X2=6.237 $Y2=2.72
r149 32 34 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=6.237 $Y=2.635
+ $X2=6.237 $Y2=2
r150 28 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.845 $Y=2.635
+ $X2=4.845 $Y2=2.72
r151 28 30 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=4.845 $Y=2.635
+ $X2=4.845 $Y2=1.995
r152 24 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=2.635
+ $X2=3.865 $Y2=2.72
r153 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.865 $Y=2.635
+ $X2=3.865 $Y2=2.34
r154 20 76 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=2.635
+ $X2=2.137 $Y2=2.72
r155 20 22 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.137 $Y=2.635
+ $X2=2.137 $Y2=2
r156 16 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r157 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r158 5 34 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=6.03
+ $Y=1.845 $X2=6.22 $Y2=2
r159 4 30 300 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=2 $X=4.67
+ $Y=1.485 $X2=4.805 $Y2=1.995
r160 3 26 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=2.065 $X2=3.865 $Y2=2.34
r161 2 22 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.845 $X2=2.065 $Y2=2
r162 1 18 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%Q 1 2 9 10 11 18 27 30
c25 30 0 1.26672e-19 $X=5.31 $Y=1.67
c26 27 0 6.43759e-20 $X=5.395 $Y=0.58
r27 16 18 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=5.31 $Y=1.84 $X2=5.31
+ $Y2=1.87
r28 10 16 0.949071 $w=3.38e-07 $l=2.8e-08 $layer=LI1_cond $X=5.31 $Y=1.812
+ $X2=5.31 $Y2=1.84
r29 10 30 7.69232 $w=3.38e-07 $l=1.42e-07 $layer=LI1_cond $X=5.31 $Y=1.812
+ $X2=5.31 $Y2=1.67
r30 10 11 10.6093 $w=3.38e-07 $l=3.13e-07 $layer=LI1_cond $X=5.31 $Y=1.897
+ $X2=5.31 $Y2=2.21
r31 10 18 0.915175 $w=3.38e-07 $l=2.7e-08 $layer=LI1_cond $X=5.31 $Y=1.897
+ $X2=5.31 $Y2=1.87
r32 9 27 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.225 $Y=0.58
+ $X2=5.395 $Y2=0.58
r33 7 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=0.745
+ $X2=5.395 $Y2=0.58
r34 7 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.395 $Y=0.745
+ $X2=5.395 $Y2=1.67
r35 2 10 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.09
+ $Y=1.485 $X2=5.225 $Y2=1.835
r36 1 9 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.235 $X2=5.225 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%Q_N 1 2 10 11 12 13 14 15
r14 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=6.685 $Y=1.82
+ $X2=6.685 $Y2=2.21
r15 11 14 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=6.685 $Y=1.635
+ $X2=6.685 $Y2=1.82
r16 11 12 6.61899 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=6.685 $Y=1.635
+ $X2=6.685 $Y2=1.505
r17 10 12 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=6.72 $Y=0.825
+ $X2=6.72 $Y2=1.505
r18 9 13 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=6.685 $Y=0.695
+ $X2=6.685 $Y2=0.51
r19 9 10 6.61899 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=6.685 $Y=0.695
+ $X2=6.685 $Y2=0.825
r20 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=6.505
+ $Y=1.485 $X2=6.64 $Y2=1.82
r21 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.64 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLXBN_1%VGND 1 2 3 4 5 18 22 26 30 34 36 38 43 48 56
+ 61 68 69 72 75 78 81 84
c103 69 0 2.71124e-20 $X=6.67 $Y=0
c104 61 0 1.13975e-20 $X=6.09 $Y=0
c105 43 0 1.29183e-19 $X=1.875 $Y=0
r106 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r107 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r108 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r110 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r111 69 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r112 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r113 66 84 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.237 $Y2=0
r114 66 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.67 $Y2=0
r115 65 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r116 65 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=4.83
+ $Y2=0
r117 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r118 62 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=0 $X2=4.805
+ $Y2=0
r119 62 64 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.97 $Y=0 $X2=5.75
+ $Y2=0
r120 61 84 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=6.237
+ $Y2=0
r121 61 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=5.75
+ $Y2=0
r122 60 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r123 60 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r124 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r125 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0 $X2=3.93
+ $Y2=0
r126 57 59 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=4.37 $Y2=0
r127 56 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.805
+ $Y2=0
r128 56 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.37
+ $Y2=0
r129 55 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r130 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r131 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r132 52 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r133 51 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r134 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r135 49 75 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.23 $Y=0 $X2=2.052
+ $Y2=0
r136 49 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.23 $Y=0 $X2=2.53
+ $Y2=0
r137 48 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.93
+ $Y2=0
r138 48 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.765 $Y=0
+ $X2=3.45 $Y2=0
r139 47 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r140 47 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r141 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r142 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r143 44 46 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r144 43 75 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.052 $Y2=0
r145 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r146 38 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r147 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r148 36 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r149 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r150 32 84 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.237 $Y=0.085
+ $X2=6.237 $Y2=0
r151 32 34 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=6.237 $Y=0.085
+ $X2=6.237 $Y2=0.38
r152 28 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.805 $Y=0.085
+ $X2=4.805 $Y2=0
r153 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.805 $Y=0.085
+ $X2=4.805 $Y2=0.38
r154 24 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=0.085
+ $X2=3.93 $Y2=0
r155 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.93 $Y=0.085
+ $X2=3.93 $Y2=0.445
r156 20 75 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.052 $Y=0.085
+ $X2=2.052 $Y2=0
r157 20 22 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=2.052 $Y=0.085
+ $X2=2.052 $Y2=0.36
r158 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r159 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r160 5 34 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=6.03
+ $Y=0.235 $X2=6.22 $Y2=0.38
r161 4 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.235 $X2=4.805 $Y2=0.38
r162 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.865 $Y2=0.445
r163 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r164 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o41a_2.spice.pex
* Created: Thu Aug 27 14:41:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O41A_2%A_79_21# 1 2 7 9 12 14 16 19 21 25 28 31 34
+ 37 40 42 46 48
c74 28 0 1.30817e-19 $X=1.13 $Y=1.16
r75 40 46 17.9412 $w=4.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.92 $Y=2.34
+ $X2=1.92 $Y2=1.665
r76 37 42 6.01496 $w=2.07e-07 $l=1.42741e-07 $layer=LI1_cond $X=1.515 $Y=1.075
+ $X2=1.477 $Y2=1.2
r77 37 48 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.515 $Y=1.075
+ $X2=1.515 $Y2=0.85
r78 32 48 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=1.607 $Y=0.673
+ $X2=1.607 $Y2=0.85
r79 32 34 9.51171 $w=3.53e-07 $l=2.93e-07 $layer=LI1_cond $X=1.607 $Y=0.673
+ $X2=1.607 $Y2=0.38
r80 31 46 24.9872 $w=1.68e-07 $l=3.83e-07 $layer=LI1_cond $X=1.477 $Y=1.58
+ $X2=1.86 $Y2=1.58
r81 30 42 6.01496 $w=2.07e-07 $l=1.25e-07 $layer=LI1_cond $X=1.477 $Y=1.325
+ $X2=1.477 $Y2=1.2
r82 30 31 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=1.477 $Y=1.325
+ $X2=1.477 $Y2=1.495
r83 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.16 $X2=1.13 $Y2=1.16
r84 25 42 0.681005 $w=2.5e-07 $l=1.22e-07 $layer=LI1_cond $X=1.355 $Y=1.2
+ $X2=1.477 $Y2=1.2
r85 25 27 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=1.355 $Y=1.2
+ $X2=1.13 $Y2=1.2
r86 22 24 65.5021 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r87 21 28 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=1.13 $Y2=1.16
r88 21 24 16.0178 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=0.89 $Y2=1.16
r89 17 24 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.89 $Y=1.345
+ $X2=0.89 $Y2=1.16
r90 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.89 $Y=1.345
+ $X2=0.89 $Y2=1.985
r91 14 24 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.89 $Y=0.975
+ $X2=0.89 $Y2=1.16
r92 14 16 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.89 $Y=0.975
+ $X2=0.89 $Y2=0.56
r93 10 22 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.47 $Y=1.345
+ $X2=0.47 $Y2=1.16
r94 10 12 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.47 $Y=1.345
+ $X2=0.47 $Y2=1.985
r95 7 22 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.47 $Y=0.975
+ $X2=0.47 $Y2=1.16
r96 7 9 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.47 $Y=0.975
+ $X2=0.47 $Y2=0.56
r97 2 46 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.485 $X2=1.86 $Y2=1.66
r98 2 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.485 $X2=1.86 $Y2=2.34
r99 1 34 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%B1 3 7 9 15
c36 9 0 1.30817e-19 $X=2.07 $Y=1.19
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=1.16 $X2=1.94 $Y2=1.16
r38 13 15 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=1.89 $Y=1.16 $X2=1.94
+ $Y2=1.16
r39 11 13 53.3217 $w=2.7e-07 $l=2.4e-07 $layer=POLY_cond $X=1.65 $Y=1.16
+ $X2=1.89 $Y2=1.16
r40 9 16 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.07 $Y=1.2 $X2=1.94
+ $Y2=1.2
r41 5 13 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.89 $Y=1.025
+ $X2=1.89 $Y2=1.16
r42 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.89 $Y=1.025
+ $X2=1.89 $Y2=0.56
r43 1 11 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.65 $Y=1.295
+ $X2=1.65 $Y2=1.16
r44 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.65 $Y=1.295 $X2=1.65
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%A4 3 6 8 9 13 15
r34 13 16 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.477 $Y=1.16
+ $X2=2.477 $Y2=1.325
r35 13 15 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.477 $Y=1.16
+ $X2=2.477 $Y2=0.995
r36 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.49 $Y=1.16 $X2=2.49
+ $Y2=1.53
r37 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.16 $X2=2.49 $Y2=1.16
r38 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.405 $Y=1.985
+ $X2=2.405 $Y2=1.325
r39 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.405 $Y=0.56
+ $X2=2.405 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%A3 3 6 8 9 10 11 17 19
c34 8 0 1.19851e-19 $X=2.99 $Y=1.19
r35 17 20 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=1.16
+ $X2=2.98 $Y2=1.325
r36 17 19 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=1.16
+ $X2=2.98 $Y2=0.995
r37 10 11 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.99 $Y=1.87
+ $X2=2.99 $Y2=2.21
r38 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.99 $Y=1.53 $X2=2.99
+ $Y2=1.87
r39 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.99 $Y=1.16 $X2=2.99
+ $Y2=1.53
r40 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.16 $X2=2.99 $Y2=1.16
r41 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.91 $Y=1.985
+ $X2=2.91 $Y2=1.325
r42 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.91 $Y=0.56 $X2=2.91
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%A2 3 6 8 9 10 11 17 19
c31 6 0 1.19851e-19 $X=3.41 $Y=1.985
r32 17 20 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.48 $Y2=1.325
r33 17 19 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.48 $Y2=0.995
r34 10 11 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.49 $Y=1.87
+ $X2=3.49 $Y2=2.21
r35 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.49 $Y=1.53 $X2=3.49
+ $Y2=1.87
r36 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.49 $Y=1.16 $X2=3.49
+ $Y2=1.53
r37 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.16 $X2=3.49 $Y2=1.16
r38 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.985
+ $X2=3.41 $Y2=1.325
r39 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.56 $X2=3.41
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%A1 3 6 8 11 13
r24 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.16
+ $X2=3.98 $Y2=1.325
r25 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.16
+ $X2=3.98 $Y2=0.995
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.99
+ $Y=1.16 $X2=3.99 $Y2=1.16
r27 8 12 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.37 $Y=1.2 $X2=3.99
+ $Y2=1.2
r28 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.91 $Y=1.985
+ $X2=3.91 $Y2=1.325
r29 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.91 $Y=0.56 $X2=3.91
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%VPWR 1 2 3 10 12 18 21 22 24 29 31 33 38 50
+ 54
r57 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r58 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 45 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r60 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 42 45 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 42 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 41 44 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 39 50 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.525 $Y=2.72
+ $X2=1.27 $Y2=2.72
r66 39 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=2.72
+ $X2=1.61 $Y2=2.72
r67 38 53 4.56733 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=4.332 $Y2=2.72
r68 38 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 37 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 34 47 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r72 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 33 50 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.27 $Y2=2.72
r74 33 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 31 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 29 30 9.57885 $w=5.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.27 $Y=2 $X2=1.27
+ $Y2=1.835
r78 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.23 $Y=1.66
+ $X2=4.23 $Y2=2.34
r79 22 53 3.19884 $w=3.3e-07 $l=1.38109e-07 $layer=LI1_cond $X=4.23 $Y=2.635
+ $X2=4.332 $Y2=2.72
r80 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.23 $Y=2.635
+ $X2=4.23 $Y2=2.34
r81 21 50 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2.72
r82 20 29 2.11073 $w=5.08e-07 $l=9e-08 $layer=LI1_cond $X=1.27 $Y=2.09 $X2=1.27
+ $Y2=2
r83 20 21 12.7816 $w=5.08e-07 $l=5.45e-07 $layer=LI1_cond $X=1.27 $Y=2.09
+ $X2=1.27 $Y2=2.635
r84 18 30 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.1 $Y=1.66 $X2=1.1
+ $Y2=1.835
r85 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r86 10 47 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r87 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r88 3 27 400 $w=1.7e-07 $l=9.69794e-07 $layer=licon1_PDIFF $count=1 $X=3.985
+ $Y=1.485 $X2=4.23 $Y2=2.34
r89 3 24 400 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_PDIFF $count=1 $X=3.985
+ $Y=1.485 $X2=4.23 $Y2=1.66
r90 2 29 150 $w=1.7e-07 $l=7.14038e-07 $layer=licon1_PDIFF $count=4 $X=0.965
+ $Y=1.485 $X2=1.44 $Y2=2
r91 2 18 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.66
r92 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r93 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%X 1 2 7 8 9 10 11 12 23 45 48
r22 48 49 1.57638 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.68 $Y=1.53
+ $X2=0.68 $Y2=1.495
r23 45 46 1.40177 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.68 $Y=0.85 $X2=0.68
+ $Y2=0.88
r24 12 41 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=2.21
+ $X2=0.68 $Y2=2.34
r25 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=2.21
r26 11 35 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=1.66
r27 10 35 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.68 $Y=1.555
+ $X2=0.68 $Y2=1.66
r28 10 48 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.68 $Y=1.555
+ $X2=0.68 $Y2=1.53
r29 10 49 1.04768 $w=2.73e-07 $l=2.5e-08 $layer=LI1_cond $X=0.652 $Y=1.47
+ $X2=0.652 $Y2=1.495
r30 9 10 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=0.652 $Y=1.19
+ $X2=0.652 $Y2=1.47
r31 8 45 0.97783 $w=3.28e-07 $l=2.8e-08 $layer=LI1_cond $X=0.68 $Y=0.822
+ $X2=0.68 $Y2=0.85
r32 8 21 3.73671 $w=3.28e-07 $l=1.07e-07 $layer=LI1_cond $X=0.68 $Y=0.822
+ $X2=0.68 $Y2=0.715
r33 8 9 11.8597 $w=2.73e-07 $l=2.83e-07 $layer=LI1_cond $X=0.652 $Y=0.907
+ $X2=0.652 $Y2=1.19
r34 8 46 1.13149 $w=2.73e-07 $l=2.7e-08 $layer=LI1_cond $X=0.652 $Y=0.907
+ $X2=0.652 $Y2=0.88
r35 7 21 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.68 $Y=0.51
+ $X2=0.68 $Y2=0.715
r36 7 23 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=0.51 $X2=0.68
+ $Y2=0.38
r37 2 41 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r38 2 35 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r39 1 23 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 39 49
+ 50 56 59
r65 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r66 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r68 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r69 47 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r70 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r71 44 59 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.617
+ $Y2=0
r72 44 46 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=3.45
+ $Y2=0
r73 43 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r74 43 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r75 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r76 40 56 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.137
+ $Y2=0
r77 40 42 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.61
+ $Y2=0
r78 39 59 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.485 $Y=0 $X2=2.617
+ $Y2=0
r79 39 42 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.485 $Y=0 $X2=1.61
+ $Y2=0
r80 38 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r81 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r82 35 53 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r83 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r84 34 56 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.137
+ $Y2=0
r85 34 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.69
+ $Y2=0
r86 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r87 32 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r88 30 46 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.45
+ $Y2=0
r89 30 31 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.64
+ $Y2=0
r90 29 49 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.775 $Y=0 $X2=4.37
+ $Y2=0
r91 29 31 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.775 $Y=0 $X2=3.64
+ $Y2=0
r92 25 31 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r93 25 27 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.38
r94 21 59 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.617 $Y=0.085
+ $X2=2.617 $Y2=0
r95 21 23 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=2.617 $Y=0.085
+ $X2=2.617 $Y2=0.38
r96 17 56 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0
r97 17 19 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0.38
r98 13 53 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r99 13 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.38
r100 4 27 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.64 $Y2=0.38
r101 3 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.615 $Y2=0.38
r102 2 19 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r103 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_2%A_393_47# 1 2 3 12 14 15 18 20 24 26
r46 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.23 $Y=0.715
+ $X2=4.23 $Y2=0.38
r47 21 26 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=0.81
+ $X2=3.12 $Y2=0.81
r48 20 22 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.065 $Y=0.81
+ $X2=4.23 $Y2=0.715
r49 20 21 45.5311 $w=1.88e-07 $l=7.8e-07 $layer=LI1_cond $X=4.065 $Y=0.81
+ $X2=3.285 $Y2=0.81
r50 16 26 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.12 $Y=0.715
+ $X2=3.12 $Y2=0.81
r51 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=0.715
+ $X2=3.12 $Y2=0.38
r52 14 26 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0.81
+ $X2=3.12 $Y2=0.81
r53 14 15 37.3589 $w=1.88e-07 $l=6.4e-07 $layer=LI1_cond $X=2.955 $Y=0.81
+ $X2=2.315 $Y2=0.81
r54 10 15 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.15 $Y=0.715
+ $X2=2.315 $Y2=0.81
r55 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.15 $Y=0.715
+ $X2=2.15 $Y2=0.38
r56 3 24 91 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=2 $X=3.985
+ $Y=0.235 $X2=4.23 $Y2=0.38
r57 2 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.985
+ $Y=0.235 $X2=3.12 $Y2=0.38
r58 1 12 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.235 $X2=2.15 $Y2=0.38
.ends


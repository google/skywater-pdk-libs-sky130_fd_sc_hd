* File: sky130_fd_sc_hd__a21o_1.spice.pex
* Created: Thu Aug 27 14:00:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21O_1%A_81_21# 1 2 7 9 12 17 18 19 20 21 23 25
r55 25 27 3.34516 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.635
+ $X2=1.62 $Y2=0.55
r56 21 23 3.62806 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=1.725
+ $X2=1.18 $Y2=1.81
r57 19 25 7.23722 $w=2e-07 $l=1.98809e-07 $layer=LI1_cond $X=1.465 $Y=0.735
+ $X2=1.62 $Y2=0.635
r58 19 20 34.9364 $w=1.98e-07 $l=6.3e-07 $layer=LI1_cond $X=1.465 $Y=0.735
+ $X2=0.835 $Y2=0.735
r59 18 32 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.695 $Y=1.16
+ $X2=0.48 $Y2=1.16
r60 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.16 $X2=0.695 $Y2=1.16
r61 15 21 25.668 $w=2.18e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=1.615
+ $X2=1.18 $Y2=1.615
r62 15 17 13.7101 $w=2.88e-07 $l=3.45e-07 $layer=LI1_cond $X=0.69 $Y=1.505
+ $X2=0.69 $Y2=1.16
r63 14 20 7.11991 $w=2e-07 $l=1.88481e-07 $layer=LI1_cond $X=0.69 $Y=0.835
+ $X2=0.835 $Y2=0.735
r64 14 17 12.9153 $w=2.88e-07 $l=3.25e-07 $layer=LI1_cond $X=0.69 $Y=0.835
+ $X2=0.69 $Y2=1.16
r65 10 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r66 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.985
r67 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r68 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995 $X2=0.48
+ $Y2=0.56
r69 2 23 300 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.485 $X2=1.21 $Y2=1.81
r70 1 27 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.63 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%B1 1 3 6 8 14
c32 14 0 8.83951e-20 $X=1.42 $Y=1.16
r33 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.205 $Y=1.16
+ $X2=1.42 $Y2=1.16
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.205
+ $Y=1.16 $X2=1.205 $Y2=1.16
r35 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.325
+ $X2=1.42 $Y2=1.16
r36 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.42 $Y=1.325 $X2=1.42
+ $Y2=1.985
r37 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=0.995
+ $X2=1.42 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.42 $Y=0.995 $X2=1.42
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%A1 1 3 6 8 9 10 15
c38 8 0 8.83951e-20 $X=2.07 $Y=0.51
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.16 $X2=1.845 $Y2=1.16
r40 10 16 8.36451 $w=3.08e-07 $l=2.25e-07 $layer=LI1_cond $X=2.07 $Y=1.17
+ $X2=1.845 $Y2=1.17
r41 10 17 2.48709 $w=2.3e-07 $l=1.55e-07 $layer=LI1_cond $X=2.07 $Y=1.17
+ $X2=2.07 $Y2=1.015
r42 9 17 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0.85
+ $X2=2.07 $Y2=1.015
r43 8 9 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.07 $Y=0.51 $X2=2.07
+ $Y2=0.85
r44 4 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.16
r45 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.985
r46 1 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=0.995
+ $X2=1.845 $Y2=1.16
r47 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.845 $Y=0.995
+ $X2=1.845 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%A2 1 3 6 8 13
r26 10 13 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.275 $Y=1.16
+ $X2=2.485 $Y2=1.16
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.16 $X2=2.485 $Y2=1.16
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.325
+ $X2=2.275 $Y2=1.16
r29 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.275 $Y=1.325
+ $X2=2.275 $Y2=1.985
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%X 1 2 7 8 9 10 11 12
r10 11 12 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=2.21
r11 11 30 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.77
r12 10 30 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=0.225 $Y=1.53
+ $X2=0.225 $Y2=1.77
r13 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=1.19
+ $X2=0.225 $Y2=1.53
r14 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=0.85
+ $X2=0.225 $Y2=1.19
r15 7 8 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.225 $Y=0.51
+ $X2=0.225 $Y2=0.85
r16 2 30 300 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.77
r17 1 7 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r40 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.06 $Y2=2.72
r45 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 23 33 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.695 $Y2=2.72
r50 23 25 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.06 $Y2=2.72
r52 22 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 17 33 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.695 $Y2=2.72
r54 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=2.635
+ $X2=2.06 $Y2=2.72
r58 11 13 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.06 $Y=2.635
+ $X2=2.06 $Y2=2.02
r59 7 33 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r60 7 9 21.5236 $w=3.38e-07 $l=6.35e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2
r61 2 13 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.485 $X2=2.06 $Y2=2.02
r62 1 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.69 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%A_299_297# 1 2 9 11 12 15
r20 13 15 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.745
+ $X2=2.525 $Y2=1.83
r21 11 13 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=2.395 $Y=1.625
+ $X2=2.525 $Y2=1.745
r22 11 12 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=2.395 $Y=1.625
+ $X2=1.725 $Y2=1.625
r23 7 12 6.82051 $w=2.4e-07 $l=1.67929e-07 $layer=LI1_cond $X=1.61 $Y=1.745
+ $X2=1.725 $Y2=1.625
r24 7 9 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.745 $X2=1.61
+ $Y2=1.83
r25 2 15 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=2.35
+ $Y=1.485 $X2=2.49 $Y2=1.83
r26 1 9 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.63 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_1%VGND 1 2 9 11 13 15 21 29 32
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r40 27 29 9.10347 $w=5.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.15 $Y=0.185
+ $X2=1.285 $Y2=0.185
r41 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r42 25 27 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=1.12 $Y=0.185
+ $X2=1.15 $Y2=0.185
r43 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r44 21 25 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=0.69 $Y=0.185
+ $X2=1.12 $Y2=0.185
r45 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r46 19 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r47 19 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r48 18 29 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.285
+ $Y2=0
r49 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r50 15 31 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.562
+ $Y2=0
r51 15 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.07
+ $Y2=0
r52 13 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r53 9 31 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.562 $Y2=0
r54 9 11 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0.53
r55 2 11 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.49 $Y2=0.53
r56 1 25 91 $w=1.7e-07 $l=6.2438e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=1.12 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__lpflow_inputiso1n_1.spice
* Created: Thu Aug 27 14:25:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_inputiso1n_1.spice.pex"
.subckt sky130_fd_sc_hd__lpflow_inputiso1n_1  VNB VPB SLEEP_B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* SLEEP_B	SLEEP_B
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_SLEEP_B_M1003_g N_A_27_53#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1575 AS=0.1092 PD=1.17 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 N_A_219_297#_M1002_d N_A_27_53#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1575 PD=0.69 PS=1.17 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_219_297#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_219_297#_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.123773 PD=1.84 PS=1.2028 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_53#_M1007_d N_SLEEP_B_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1176 AS=0.1092 PD=1.4 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_301_297# N_A_27_53#_M1005_g N_A_219_297#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_301_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.0441 PD=0.792676 PS=0.63 NRD=72.1217 NRS=23.443 M=1 R=2.8
+ SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_219_297#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.208803 PD=2.54 PS=1.88732 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__lpflow_inputiso1n_1.spice.SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__o31ai_1.spice.SKY130_FD_SC_HD__O31AI_1.pxi
* Created: Thu Aug 27 14:40:18 2020
* 
x_PM_SKY130_FD_SC_HD__O31AI_1%A1 N_A1_c_47_n N_A1_M1007_g N_A1_M1004_g A1
+ N_A1_c_49_n PM_SKY130_FD_SC_HD__O31AI_1%A1
x_PM_SKY130_FD_SC_HD__O31AI_1%A2 N_A2_c_71_n N_A2_M1002_g N_A2_M1001_g A2 A2 A2
+ A2 N_A2_c_72_n N_A2_c_73_n PM_SKY130_FD_SC_HD__O31AI_1%A2
x_PM_SKY130_FD_SC_HD__O31AI_1%A3 N_A3_M1003_g N_A3_M1000_g A3 N_A3_c_110_n
+ N_A3_c_111_n N_A3_c_115_n PM_SKY130_FD_SC_HD__O31AI_1%A3
x_PM_SKY130_FD_SC_HD__O31AI_1%B1 N_B1_M1005_g N_B1_M1006_g N_B1_c_144_n
+ N_B1_c_145_n B1 N_B1_c_147_n PM_SKY130_FD_SC_HD__O31AI_1%B1
x_PM_SKY130_FD_SC_HD__O31AI_1%VPWR N_VPWR_M1004_s N_VPWR_M1006_d N_VPWR_c_173_n
+ N_VPWR_c_174_n N_VPWR_c_175_n N_VPWR_c_176_n VPWR N_VPWR_c_177_n
+ N_VPWR_c_172_n PM_SKY130_FD_SC_HD__O31AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O31AI_1%Y N_Y_M1005_d N_Y_M1000_d Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_HD__O31AI_1%Y
x_PM_SKY130_FD_SC_HD__O31AI_1%VGND N_VGND_M1007_s N_VGND_M1002_d N_VGND_c_232_n
+ N_VGND_c_233_n N_VGND_c_234_n VGND N_VGND_c_235_n N_VGND_c_236_n
+ N_VGND_c_237_n N_VGND_c_238_n PM_SKY130_FD_SC_HD__O31AI_1%VGND
x_PM_SKY130_FD_SC_HD__O31AI_1%A_109_47# N_A_109_47#_M1007_d N_A_109_47#_M1003_d
+ N_A_109_47#_c_269_n N_A_109_47#_c_267_n N_A_109_47#_c_268_n
+ N_A_109_47#_c_278_n PM_SKY130_FD_SC_HD__O31AI_1%A_109_47#
cc_1 VNB N_A1_c_47_n 0.0215757f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A1 0.00931883f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A1_c_49_n 0.0401281f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A2_c_71_n 0.0162239f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_A2_c_72_n 0.0190122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A2_c_73_n 0.00438076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB A3 0.00388336f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_8 VNB N_A3_c_110_n 0.0277597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A3_c_111_n 0.0186412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_144_n 0.0204279f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_B1_c_145_n 0.0218583f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_12 VNB B1 0.0147977f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_13 VNB N_B1_c_147_n 0.0293418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_172_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB Y 0.0294353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB Y 0.00785375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_232_n 0.0110498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_233_n 0.00602085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_234_n 0.00415222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_235_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_236_n 0.0415265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_237_n 0.164378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_238_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_109_47#_c_267_n 0.00890875f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_25 VNB N_A_109_47#_c_268_n 0.00437869f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_26 VPB N_A1_M1004_g 0.0252861f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_27 VPB A1 0.00355152f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_28 VPB N_A1_c_49_n 0.00995901f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_29 VPB N_A2_M1001_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_30 VPB N_A2_c_72_n 0.00440081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A2_c_73_n 0.00320885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A3_M1000_g 0.0221902f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB A3 8.28589e-19 $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_34 VPB N_A3_c_110_n 0.00990406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A3_c_115_n 0.00276082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_B1_M1006_g 0.029338f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_B1_c_144_n 0.00624757f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_38 VPB B1 0.00392453f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_39 VPB N_B1_c_147_n 0.011053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_173_n 0.0104466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_174_n 0.0418125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_175_n 0.0115225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_176_n 0.0450372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_177_n 0.050688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_172_n 0.0429195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB Y 0.00295379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 N_A1_c_47_n N_A2_c_71_n 0.0124239f $X=0.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_48 N_A1_M1004_g N_A2_M1001_g 0.0556174f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_49 A1 N_A2_c_72_n 2.02389e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A1_c_49_n N_A2_c_72_n 0.021722f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_51 A1 N_A2_c_73_n 0.0203479f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_52 N_A1_c_49_n N_A2_c_73_n 0.013826f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A1_M1004_g N_VPWR_c_174_n 0.0185404f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_54 A1 N_VPWR_c_174_n 0.0257559f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A1_c_49_n N_VPWR_c_174_n 0.00208296f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A1_M1004_g N_VPWR_c_177_n 0.00407992f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A1_M1004_g N_VPWR_c_172_n 0.0070745f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A1_c_47_n N_VGND_c_233_n 0.00360182f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_59 A1 N_VGND_c_233_n 0.0139721f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_60 N_A1_c_49_n N_VGND_c_233_n 0.00431028f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A1_c_47_n N_VGND_c_235_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A1_c_47_n N_VGND_c_237_n 0.0104829f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A1_c_47_n N_A_109_47#_c_269_n 0.00550646f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A1_c_47_n N_A_109_47#_c_268_n 0.00359092f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A2_M1001_g N_A3_M1000_g 0.0564456f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A2_c_72_n A3 8.11543e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A2_c_73_n A3 0.021802f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A2_c_72_n N_A3_c_110_n 0.0221546f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A2_c_73_n N_A3_c_110_n 0.0120353f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A2_c_71_n N_A3_c_111_n 0.0254185f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A2_c_73_n N_A3_c_115_n 0.0461381f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A2_M1001_g N_VPWR_c_174_n 0.00193777f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A2_c_73_n N_VPWR_c_174_n 0.0773983f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A2_M1001_g N_VPWR_c_177_n 0.00357668f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A2_c_73_n N_VPWR_c_177_n 0.0268592f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A2_M1001_g N_VPWR_c_172_n 0.00532039f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A2_c_73_n N_VPWR_c_172_n 0.0163747f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A2_c_73_n A_109_297# 0.0105526f $X=0.89 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_79 N_A2_c_73_n A_193_297# 0.012549f $X=0.89 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_80 N_A2_c_71_n N_VGND_c_234_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A2_c_71_n N_VGND_c_235_n 0.00424416f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A2_c_71_n N_VGND_c_237_n 0.00579048f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A2_c_71_n N_A_109_47#_c_269_n 0.00645631f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A2_c_71_n N_A_109_47#_c_267_n 0.00845282f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A2_c_72_n N_A_109_47#_c_267_n 0.001478f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A2_c_73_n N_A_109_47#_c_267_n 0.0163508f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A2_c_71_n N_A_109_47#_c_268_n 0.00109929f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A2_c_72_n N_A_109_47#_c_268_n 0.00153445f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A2_c_73_n N_A_109_47#_c_268_n 0.0213077f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A2_c_71_n N_A_109_47#_c_278_n 5.1881e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_91 A3 N_B1_c_144_n 9.4839e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A3_c_110_n N_B1_c_144_n 0.0103284f $X=1.46 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A3_c_111_n N_B1_c_145_n 0.00828535f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A3_M1000_g N_VPWR_c_177_n 0.00585385f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A3_c_115_n N_VPWR_c_177_n 0.0120564f $X=1.58 $Y=1.2 $X2=0 $Y2=0
cc_96 N_A3_M1000_g N_VPWR_c_172_n 0.0122169f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A3_c_115_n N_VPWR_c_172_n 0.00888736f $X=1.58 $Y=1.2 $X2=0 $Y2=0
cc_98 N_A3_c_115_n N_Y_M1000_d 0.0355153f $X=1.58 $Y=1.2 $X2=0 $Y2=0
cc_99 N_A3_M1000_g Y 0.00313406f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_100 A3 Y 0.0160006f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A3_c_110_n Y 0.00236864f $X=1.46 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A3_c_111_n Y 0.00143362f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A3_c_115_n Y 0.0630645f $X=1.58 $Y=1.2 $X2=0 $Y2=0
cc_104 N_A3_c_111_n N_VGND_c_234_n 0.00268723f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A3_c_111_n N_VGND_c_236_n 0.0043257f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A3_c_111_n N_VGND_c_237_n 0.00650358f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A3_c_111_n N_A_109_47#_c_269_n 5.28455e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_108 A3 N_A_109_47#_c_267_n 0.0376087f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_109 N_A3_c_110_n N_A_109_47#_c_267_n 0.00614237f $X=1.46 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A3_c_111_n N_A_109_47#_c_267_n 0.0100204f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A3_c_111_n N_A_109_47#_c_278_n 0.00594327f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B1_M1006_g N_VPWR_c_176_n 0.00492552f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_113 B1 N_VPWR_c_176_n 0.0265665f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_114 N_B1_c_147_n N_VPWR_c_176_n 0.00242497f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B1_M1006_g N_VPWR_c_177_n 0.00585385f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_M1006_g N_VPWR_c_172_n 0.0127575f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B1_c_144_n Y 0.00699713f $X=2.157 $Y=1.16 $X2=0 $Y2=0
cc_118 N_B1_c_145_n Y 0.01546f $X=2.157 $Y=0.995 $X2=0 $Y2=0
cc_119 B1 Y 0.0283093f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B1_c_147_n Y 0.00250861f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B1_M1006_g Y 0.0122042f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_c_144_n Y 0.0161495f $X=2.157 $Y=1.16 $X2=0 $Y2=0
cc_123 N_B1_c_145_n Y 0.00610087f $X=2.157 $Y=0.995 $X2=0 $Y2=0
cc_124 B1 Y 0.024062f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_125 N_B1_c_145_n N_VGND_c_236_n 0.00358923f $X=2.157 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_c_145_n N_VGND_c_237_n 0.00701436f $X=2.157 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_c_145_n N_A_109_47#_c_267_n 7.7232e-19 $X=2.157 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_c_145_n N_A_109_47#_c_278_n 0.00203805f $X=2.157 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_VPWR_c_172_n A_109_297# 0.00445931f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_130 N_VPWR_c_172_n A_193_297# 0.00845161f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_131 N_VPWR_c_172_n N_Y_M1000_d 0.0179667f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_132 N_VPWR_c_177_n Y 0.0133757f $X=2.33 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_172_n Y 0.008203f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_134 Y N_VGND_c_236_n 0.0451839f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_135 N_Y_M1005_d N_VGND_c_237_n 0.00275131f $X=2.145 $Y=0.235 $X2=0 $Y2=0
cc_136 Y N_VGND_c_237_n 0.0271339f $X=2.45 $Y=0.425 $X2=0 $Y2=0
cc_137 Y N_A_109_47#_c_267_n 0.00335198f $X=2.075 $Y=0.85 $X2=0 $Y2=0
cc_138 N_VGND_c_237_n N_A_109_47#_M1007_d 0.00215201f $X=2.53 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_139 N_VGND_c_237_n N_A_109_47#_M1003_d 0.0134646f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_140 N_VGND_c_235_n N_A_109_47#_c_269_n 0.0188551f $X=1.015 $Y=0 $X2=0 $Y2=0
cc_141 N_VGND_c_237_n N_A_109_47#_c_269_n 0.0122069f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_142 N_VGND_M1002_d N_A_109_47#_c_267_n 0.00162006f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_VGND_c_234_n N_A_109_47#_c_267_n 0.0122414f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_144 N_VGND_c_235_n N_A_109_47#_c_267_n 0.00193763f $X=1.015 $Y=0 $X2=0 $Y2=0
cc_145 N_VGND_c_236_n N_A_109_47#_c_267_n 0.00213422f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_146 N_VGND_c_237_n N_A_109_47#_c_267_n 0.00857624f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_147 N_VGND_c_233_n N_A_109_47#_c_268_n 0.00787895f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_148 N_VGND_c_236_n N_A_109_47#_c_278_n 0.020954f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_149 N_VGND_c_237_n N_A_109_47#_c_278_n 0.0124805f $X=2.53 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__mux4_4.spice.pex
* Created: Thu Aug 27 14:28:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX4_4%S0 3 7 9 11 13 17 21 23 24 27 29 30 33 34 35
+ 36 43 45 46 52 58
c201 46 0 7.62213e-20 $X=6.215 $Y=1.53
c202 43 0 9.63205e-21 $X=1.155 $Y=1.53
c203 35 0 7.52734e-20 $X=6.07 $Y=1.53
c204 17 0 1.33206e-19 $X=1.915 $Y=0.415
r205 61 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.385 $Y=1.41
+ $X2=6.385 $Y2=1.575
r206 58 61 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.385 $Y=1.32
+ $X2=6.385 $Y2=1.41
r207 54 56 24.3813 $w=2.57e-07 $l=1.3e-07 $layer=POLY_cond $X=1.31 $Y=1.32
+ $X2=1.31 $Y2=1.45
r208 49 52 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r209 46 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.385
+ $Y=1.41 $X2=6.385 $Y2=1.41
r210 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=1.53
+ $X2=6.215 $Y2=1.53
r211 43 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.45 $X2=1.31 $Y2=1.45
r212 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.53
+ $X2=1.155 $Y2=1.53
r213 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.53
+ $X2=1.155 $Y2=1.53
r214 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.07 $Y=1.53
+ $X2=6.215 $Y2=1.53
r215 35 36 5.90345 $w=1.4e-07 $l=4.77e-06 $layer=MET1_cond $X=6.07 $Y=1.53
+ $X2=1.3 $Y2=1.53
r216 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.38 $Y=1.53
+ $X2=0.235 $Y2=1.53
r217 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.01 $Y=1.53
+ $X2=1.155 $Y2=1.53
r218 33 34 0.779701 $w=1.4e-07 $l=6.3e-07 $layer=MET1_cond $X=1.01 $Y=1.53
+ $X2=0.38 $Y2=1.53
r219 30 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.53
+ $X2=0.235 $Y2=1.53
r220 29 30 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.16
+ $X2=0.24 $Y2=1.53
r221 29 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r222 27 63 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.325 $Y=2.275
+ $X2=6.325 $Y2=1.575
r223 23 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.25 $Y=1.32
+ $X2=6.385 $Y2=1.32
r224 23 24 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.25 $Y=1.32
+ $X2=5.86 $Y2=1.32
r225 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.785 $Y=1.245
+ $X2=5.86 $Y2=1.32
r226 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.785 $Y=1.245
+ $X2=5.785 $Y2=0.415
r227 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.915 $Y=1.245
+ $X2=1.915 $Y2=0.415
r228 14 54 15.359 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.445 $Y=1.32
+ $X2=1.31 $Y2=1.32
r229 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.84 $Y=1.32
+ $X2=1.915 $Y2=1.245
r230 13 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.84 $Y=1.32
+ $X2=1.445 $Y2=1.32
r231 9 56 39.2307 $w=2.57e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.37 $Y=1.615
+ $X2=1.31 $Y2=1.45
r232 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.37 $Y=1.615
+ $X2=1.37 $Y2=2.275
r233 5 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r234 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=2.165
r235 1 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r236 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A2 3 6 8 9 14 16
c57 9 0 1.60284e-19 $X=1.155 $Y=0.85
r58 15 25 7.22896 $w=3.28e-07 $l=2.07e-07 $layer=LI1_cond $X=0.925 $Y=0.93
+ $X2=1.132 $Y2=0.93
r59 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=0.93
+ $X2=0.925 $Y2=1.095
r60 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=0.93
+ $X2=0.925 $Y2=0.765
r61 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=0.93 $X2=0.925 $Y2=0.93
r62 9 25 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=1.155 $Y=0.93
+ $X2=1.132 $Y2=0.93
r63 9 25 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.132 $Y=0.765
+ $X2=1.132 $Y2=0.93
r64 8 9 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.132 $Y=0.51
+ $X2=1.132 $Y2=0.765
r65 6 17 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.89 $Y=2.165
+ $X2=0.89 $Y2=1.095
r66 3 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A_27_47# 1 2 7 9 12 16 18 20 23 27 30 31 32
+ 37 43 45 51 54 55 61 69 70 74 75 80 85
c241 69 0 9.63205e-21 $X=1.82 $Y=1.74
c242 51 0 3.21039e-20 $X=6.205 $Y=0.87
r243 74 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.875 $Y=1.74
+ $X2=5.875 $Y2=1.875
r244 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.875
+ $Y=1.74 $X2=5.875 $Y2=1.74
r245 70 85 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.74
+ $X2=1.735 $Y2=1.575
r246 69 72 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.82 $Y=1.74
+ $X2=1.82 $Y2=1.875
r247 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.74 $X2=1.82 $Y2=1.74
r248 61 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.755 $Y=1.87
+ $X2=5.755 $Y2=1.87
r249 58 70 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.735 $Y=1.87
+ $X2=1.735 $Y2=1.74
r250 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=1.87
+ $X2=1.615 $Y2=1.87
r251 55 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=1.87
+ $X2=1.615 $Y2=1.87
r252 54 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.61 $Y=1.87
+ $X2=5.755 $Y2=1.87
r253 54 55 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=5.61 $Y=1.87
+ $X2=1.76 $Y2=1.87
r254 52 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=6.205 $Y=0.87
+ $X2=6.335 $Y2=0.87
r255 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.205
+ $Y=0.87 $X2=6.205 $Y2=0.87
r256 48 75 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5.815 $Y=1.035
+ $X2=5.815 $Y2=1.74
r257 47 51 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.815 $Y=0.87
+ $X2=6.205 $Y2=0.87
r258 47 48 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0.87
+ $X2=5.815 $Y2=1.035
r259 43 64 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.495 $Y=0.87
+ $X2=1.365 $Y2=0.87
r260 42 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.495 $Y=0.87
+ $X2=1.65 $Y2=0.87
r261 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=0.87 $X2=1.495 $Y2=0.87
r262 39 40 19.9479 $w=2.11e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.935
+ $X2=0.585 $Y2=1.935
r263 33 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=1.035
+ $X2=1.65 $Y2=0.87
r264 33 85 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.65 $Y=1.035
+ $X2=1.65 $Y2=1.575
r265 32 40 5.41085 $w=2.11e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.67 $Y=1.87
+ $X2=0.585 $Y2=1.935
r266 31 58 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.565 $Y=1.87
+ $X2=1.735 $Y2=1.87
r267 31 32 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.565 $Y=1.87
+ $X2=0.67 $Y2=1.87
r268 30 40 2.00497 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.585 $Y=1.785
+ $X2=0.585 $Y2=1.935
r269 29 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=0.805
+ $X2=0.585 $Y2=0.72
r270 29 30 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.585 $Y=0.805
+ $X2=0.585 $Y2=1.785
r271 25 39 0.745451 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=2.085
+ $X2=0.24 $Y2=1.935
r272 25 27 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.085
+ $X2=0.24 $Y2=2.21
r273 21 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=0.72
+ $X2=0.585 $Y2=0.72
r274 21 23 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.635
+ $X2=0.24 $Y2=0.51
r275 18 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=0.705
+ $X2=6.335 $Y2=0.87
r276 18 20 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.335 $Y=0.705
+ $X2=6.335 $Y2=0.415
r277 16 77 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.905 $Y=2.275
+ $X2=5.905 $Y2=1.875
r278 12 72 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.79 $Y=2.275
+ $X2=1.79 $Y2=1.875
r279 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.705
+ $X2=1.365 $Y2=0.87
r280 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.365 $Y=0.705
+ $X2=1.365 $Y2=0.415
r281 2 27 600 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.21
r282 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A3 3 5 6 8 11 13 14 18 20
c59 20 0 1.3041e-19 $X=2.41 $Y=0.765
c60 18 0 1.47056e-19 $X=2.41 $Y=0.93
c61 13 0 4.84598e-20 $X=2.535 $Y=0.85
r62 19 30 4.96365 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.432 $Y=0.93
+ $X2=2.432 $Y2=1.015
r63 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=0.93
+ $X2=2.41 $Y2=1.095
r64 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=0.93
+ $X2=2.41 $Y2=0.765
r65 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=0.93 $X2=2.41 $Y2=0.93
r66 14 30 9.46785 $w=2.03e-07 $l=1.75e-07 $layer=LI1_cond $X=2.517 $Y=1.19
+ $X2=2.517 $Y2=1.015
r67 13 19 2.45854 $w=3.73e-07 $l=8e-08 $layer=LI1_cond $X=2.432 $Y=0.85
+ $X2=2.432 $Y2=0.93
r68 9 11 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=2.395 $Y=1.575
+ $X2=2.51 $Y2=1.575
r69 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.51 $Y=1.65 $X2=2.51
+ $Y2=1.575
r70 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.51 $Y=1.65 $X2=2.51
+ $Y2=2.045
r71 5 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.395 $Y=1.5 $X2=2.395
+ $Y2=1.575
r72 5 21 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.395 $Y=1.5
+ $X2=2.395 $Y2=1.095
r73 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.395 $Y=0.445
+ $X2=2.395 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%S1 1 4 5 7 8 9 10 12 14 17 19 20
c86 19 0 1.3041e-19 $X=2.995 $Y=0.85
c87 5 0 4.84598e-20 $X=2.935 $Y=0.73
c88 1 0 3.58022e-19 $X=2.93 $Y=1.095
r89 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.89
+ $Y=0.93 $X2=2.89 $Y2=0.93
r90 23 25 23.1731 $w=2.6e-07 $l=1.25e-07 $layer=POLY_cond $X=2.89 $Y=0.805
+ $X2=2.89 $Y2=0.93
r91 20 26 10.3322 $w=2.88e-07 $l=2.6e-07 $layer=LI1_cond $X=2.935 $Y=1.19
+ $X2=2.935 $Y2=0.93
r92 19 26 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=2.935 $Y=0.85
+ $X2=2.935 $Y2=0.93
r93 15 17 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.29 $Y=2.465
+ $X2=4.29 $Y2=1.85
r94 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.885 $Y=0.73
+ $X2=3.885 $Y2=0.445
r95 11 23 15.628 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.025 $Y=0.805
+ $X2=2.89 $Y2=0.805
r96 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.81 $Y=0.805
+ $X2=3.885 $Y2=0.73
r97 10 11 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.81 $Y=0.805
+ $X2=3.025 $Y2=0.805
r98 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.215 $Y=2.54
+ $X2=4.29 $Y2=2.465
r99 8 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=4.215 $Y=2.54
+ $X2=3.005 $Y2=2.54
r100 5 23 22.4589 $w=2.6e-07 $l=9.48683e-08 $layer=POLY_cond $X=2.935 $Y=0.73
+ $X2=2.89 $Y2=0.805
r101 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.935 $Y=0.73
+ $X2=2.935 $Y2=0.445
r102 2 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.93 $Y=2.465
+ $X2=3.005 $Y2=2.54
r103 2 4 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.93 $Y=2.465
+ $X2=2.93 $Y2=2.045
r104 1 25 39.1435 $w=2.6e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.93 $Y=1.095
+ $X2=2.89 $Y2=0.93
r105 1 4 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.93 $Y=1.095
+ $X2=2.93 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A_601_345# 1 2 9 11 15 17 18 20 22 29
c69 22 0 2.63684e-19 $X=3.4 $Y=1.225
r70 27 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.155 $Y=0.38
+ $X2=3.335 $Y2=0.38
r71 22 25 31.9878 $w=2.46e-07 $l=7.25034e-07 $layer=LI1_cond $X=3.4 $Y=1.225
+ $X2=3.23 $Y2=1.87
r72 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.225 $X2=3.4 $Y2=1.225
r73 20 22 9.35836 $w=2.46e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.335 $Y=1.06
+ $X2=3.4 $Y2=1.225
r74 19 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.465
+ $X2=3.335 $Y2=0.38
r75 19 20 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.335 $Y=0.465
+ $X2=3.335 $Y2=1.06
r76 17 23 87.7586 $w=2.7e-07 $l=3.95e-07 $layer=POLY_cond $X=3.795 $Y=1.225
+ $X2=3.4 $Y2=1.225
r77 17 18 15.2969 $w=2.1e-07 $l=7.5e-08 $layer=POLY_cond $X=3.795 $Y=1.225
+ $X2=3.87 $Y2=1.225
r78 13 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.31 $Y=1.09
+ $X2=4.31 $Y2=0.445
r79 12 18 15.2969 $w=2.1e-07 $l=1.00623e-07 $layer=POLY_cond $X=3.945 $Y=1.165
+ $X2=3.87 $Y2=1.225
r80 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.235 $Y=1.165
+ $X2=4.31 $Y2=1.09
r81 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.235 $Y=1.165
+ $X2=3.945 $Y2=1.165
r82 7 18 10.1846 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.87 $Y=1.36
+ $X2=3.87 $Y2=1.225
r83 7 9 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.87 $Y=1.36 $X2=3.87
+ $Y2=1.85
r84 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.725 $X2=3.14 $Y2=1.87
r85 1 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.235 $X2=3.155 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A1 3 7 9 10 16
r40 16 17 3.00312 $w=3.21e-07 $l=2e-08 $layer=POLY_cond $X=5.23 $Y=1.23 $X2=5.25
+ $Y2=1.23
r41 14 16 29.2804 $w=3.21e-07 $l=1.95e-07 $layer=POLY_cond $X=5.035 $Y=1.23
+ $X2=5.23 $Y2=1.23
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.035
+ $Y=1.23 $X2=5.035 $Y2=1.23
r43 10 15 1.24588 $w=3.68e-07 $l=4e-08 $layer=LI1_cond $X=4.935 $Y=1.19
+ $X2=4.935 $Y2=1.23
r44 9 10 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.935 $Y=0.85 $X2=4.935
+ $Y2=1.19
r45 5 17 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.25 $Y=1.065
+ $X2=5.25 $Y2=1.23
r46 5 7 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.25 $Y=1.065 $X2=5.25
+ $Y2=0.445
r47 1 16 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.23 $Y=1.395
+ $X2=5.23 $Y2=1.23
r48 1 3 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.23 $Y=1.395 $X2=5.23
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A0 3 7 9 12 13 14
c49 12 0 3.21168e-19 $X=6.865 $Y=1.16
c50 9 0 4.70922e-20 $X=6.695 $Y=0.995
r51 13 14 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=6.695 $Y=0.51
+ $X2=6.695 $Y2=0.85
r52 12 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.865 $Y=1.16
+ $X2=6.865 $Y2=1.325
r53 12 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.865 $Y=1.16
+ $X2=6.865 $Y2=0.995
r54 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.865
+ $Y=1.16 $X2=6.865 $Y2=1.16
r55 9 14 5.39046 $w=3.08e-07 $l=1.45e-07 $layer=LI1_cond $X=6.695 $Y=0.995
+ $X2=6.695 $Y2=0.85
r56 9 11 6.10881 $w=3.34e-07 $l=1.88348e-07 $layer=LI1_cond $X=6.695 $Y=0.995
+ $X2=6.745 $Y2=1.16
r57 7 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.83 $Y=2.165
+ $X2=6.83 $Y2=1.325
r58 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.81 $Y=0.445
+ $X2=6.81 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A_789_316# 1 2 7 9 12 14 16 19 21 22 23 25 28
+ 30 32 35 38 42 47 48 49 51 52 56 59 60 63 66 77
c186 51 0 1.33968e-19 $X=7.205 $Y=1.495
c187 49 0 1.93706e-19 $X=6.85 $Y=1.58
c188 42 0 1.35566e-19 $X=4.1 $Y=0.51
r189 67 77 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.675 $Y=2.21
+ $X2=6.765 $Y2=2.21
r190 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.675 $Y=2.21
+ $X2=6.675 $Y2=2.21
r191 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.375 $Y=2.21
+ $X2=4.375 $Y2=2.21
r192 60 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.52 $Y=2.21
+ $X2=4.375 $Y2=2.21
r193 59 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.53 $Y=2.21
+ $X2=6.675 $Y2=2.21
r194 59 60 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=6.53 $Y=2.21
+ $X2=4.52 $Y2=2.21
r195 57 72 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=7.345 $Y=1.16
+ $X2=7.735 $Y2=1.16
r196 57 69 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=7.345 $Y=1.16
+ $X2=7.315 $Y2=1.16
r197 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.345
+ $Y=1.16 $X2=7.345 $Y2=1.16
r198 53 56 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.205 $Y=1.16
+ $X2=7.345 $Y2=1.16
r199 52 63 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=2.21
+ $X2=4.375 $Y2=2.21
r200 50 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.205 $Y=1.325
+ $X2=7.205 $Y2=1.16
r201 50 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.205 $Y=1.325
+ $X2=7.205 $Y2=1.495
r202 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.12 $Y=1.58
+ $X2=7.205 $Y2=1.495
r203 48 49 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.12 $Y=1.58
+ $X2=6.85 $Y2=1.58
r204 47 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.765 $Y=2.125
+ $X2=6.765 $Y2=2.21
r205 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.765 $Y=1.665
+ $X2=6.85 $Y2=1.58
r206 46 47 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.765 $Y=1.665
+ $X2=6.765 $Y2=2.125
r207 42 45 70.9234 $w=1.88e-07 $l=1.215e-06 $layer=LI1_cond $X=4.09 $Y=0.51
+ $X2=4.09 $Y2=1.725
r208 40 52 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.09 $Y=2.125
+ $X2=4.185 $Y2=2.21
r209 40 45 23.3493 $w=1.88e-07 $l=4e-07 $layer=LI1_cond $X=4.09 $Y=2.125
+ $X2=4.09 $Y2=1.725
r210 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.235 $Y=1.16
+ $X2=8.655 $Y2=1.16
r211 33 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=1.325
+ $X2=8.655 $Y2=1.16
r212 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.655 $Y=1.325
+ $X2=8.655 $Y2=1.985
r213 30 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=0.995
+ $X2=8.655 $Y2=1.16
r214 30 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.655 $Y=0.995
+ $X2=8.655 $Y2=0.56
r215 26 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=1.325
+ $X2=8.235 $Y2=1.16
r216 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.235 $Y=1.325
+ $X2=8.235 $Y2=1.985
r217 23 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=0.995
+ $X2=8.235 $Y2=1.16
r218 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.235 $Y=0.995
+ $X2=8.235 $Y2=0.56
r219 22 72 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.81 $Y=1.16
+ $X2=7.735 $Y2=1.16
r220 21 37 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.16 $Y=1.16
+ $X2=8.235 $Y2=1.16
r221 21 22 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=8.16 $Y=1.16
+ $X2=7.81 $Y2=1.16
r222 17 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.735 $Y=1.325
+ $X2=7.735 $Y2=1.16
r223 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.735 $Y=1.325
+ $X2=7.735 $Y2=1.985
r224 14 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.735 $Y=0.995
+ $X2=7.735 $Y2=1.16
r225 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.735 $Y=0.995
+ $X2=7.735 $Y2=0.56
r226 10 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.315 $Y=1.325
+ $X2=7.315 $Y2=1.16
r227 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.315 $Y=1.325
+ $X2=7.315 $Y2=1.985
r228 7 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.315 $Y=0.995
+ $X2=7.315 $Y2=1.16
r229 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.315 $Y=0.995
+ $X2=7.315 $Y2=0.56
r230 2 45 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.58 $X2=4.08 $Y2=1.725
r231 1 42 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.235 $X2=4.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 43 48 49
+ 51 52 53 55 67 78 82 88 91 94 98
c146 4 0 1.33968e-19 $X=6.905 $Y=1.845
r147 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r148 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r149 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r150 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 86 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r152 86 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r153 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r154 83 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=2.72
+ $X2=8.065 $Y2=2.72
r155 83 85 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.19 $Y=2.72
+ $X2=8.51 $Y2=2.72
r156 82 97 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=9.027 $Y2=2.72
r157 82 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=8.51 $Y2=2.72
r158 81 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r159 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r160 78 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.94 $Y=2.72
+ $X2=8.065 $Y2=2.72
r161 78 80 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.94 $Y=2.72
+ $X2=7.59 $Y2=2.72
r162 77 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r163 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r164 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.67 $Y2=2.72
r165 74 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r166 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=6.67 $Y2=2.72
r167 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r168 71 91 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=4.932 $Y2=2.72
r169 71 73 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=5.29 $Y2=2.72
r170 70 92 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r171 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r172 67 91 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.76 $Y=2.72
+ $X2=4.932 $Y2=2.72
r173 67 69 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=4.76 $Y=2.72
+ $X2=2.99 $Y2=2.72
r174 66 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r175 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r176 63 66 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 63 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r178 62 65 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r179 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r180 60 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r181 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r182 55 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r183 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r184 53 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r185 53 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r186 51 76 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.02 $Y=2.72
+ $X2=6.67 $Y2=2.72
r187 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.02 $Y=2.72
+ $X2=7.105 $Y2=2.72
r188 50 80 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.19 $Y=2.72 $X2=7.59
+ $Y2=2.72
r189 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.105 $Y2=2.72
r190 48 65 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.6 $Y=2.72 $X2=2.53
+ $Y2=2.72
r191 48 49 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.6 $Y=2.72
+ $X2=2.715 $Y2=2.72
r192 47 69 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.83 $Y=2.72
+ $X2=2.99 $Y2=2.72
r193 47 49 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.83 $Y=2.72
+ $X2=2.715 $Y2=2.72
r194 43 46 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.98 $Y=1.66
+ $X2=8.98 $Y2=2.34
r195 41 97 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=8.98 $Y=2.635
+ $X2=9.027 $Y2=2.72
r196 41 46 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=2.635
+ $X2=8.98 $Y2=2.34
r197 37 40 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.065 $Y=1.66
+ $X2=8.065 $Y2=2.34
r198 35 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=2.635
+ $X2=8.065 $Y2=2.72
r199 35 40 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.065 $Y=2.635
+ $X2=8.065 $Y2=2.34
r200 31 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.105 $Y=2.635
+ $X2=7.105 $Y2=2.72
r201 31 33 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.105 $Y=2.635
+ $X2=7.105 $Y2=2
r202 27 91 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.932 $Y=2.635
+ $X2=4.932 $Y2=2.72
r203 27 29 15.5329 $w=3.43e-07 $l=4.65e-07 $layer=LI1_cond $X=4.932 $Y=2.635
+ $X2=4.932 $Y2=2.17
r204 23 49 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=2.635
+ $X2=2.715 $Y2=2.72
r205 23 25 20.7941 $w=2.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.715 $Y=2.635
+ $X2=2.715 $Y2=2.22
r206 19 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r207 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r208 6 46 400 $w=1.7e-07 $l=9.54241e-07 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.485 $X2=8.94 $Y2=2.34
r209 6 43 400 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.485 $X2=8.94 $Y2=1.66
r210 5 40 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=1.485 $X2=8.025 $Y2=2.34
r211 5 37 400 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=1.485 $X2=8.025 $Y2=1.66
r212 4 33 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=6.905
+ $Y=1.845 $X2=7.105 $Y2=2
r213 3 29 600 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.845 $X2=5.02 $Y2=2.17
r214 2 25 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.725 $X2=2.72 $Y2=2.22
r215 1 21 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A_288_47# 1 2 3 4 13 17 22 24 25 26 28 33 35
+ 37 40 41 47
c132 47 0 2.0604e-19 $X=3.455 $Y=2.21
c133 22 0 2.70784e-20 $X=1.99 $Y=1.235
c134 13 0 7.52734e-20 $X=2.075 $Y=2.21
r135 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.455 $Y=2.21
+ $X2=3.455 $Y2=2.21
r136 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.075 $Y=2.21
+ $X2=2.075 $Y2=2.21
r137 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.22 $Y=2.21
+ $X2=2.075 $Y2=2.21
r138 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.31 $Y=2.21
+ $X2=3.455 $Y2=2.21
r139 40 41 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=3.31 $Y=2.21
+ $X2=2.22 $Y2=2.21
r140 37 39 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=3.707 $Y=0.51
+ $X2=3.707 $Y2=0.675
r141 35 39 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=3.74 $Y=1.81
+ $X2=3.74 $Y2=0.675
r142 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.99 $Y=1.32
+ $X2=2.16 $Y2=1.32
r143 26 48 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.7 $Y=2.21
+ $X2=3.455 $Y2=2.21
r144 26 28 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.7 $Y=2.125
+ $X2=3.7 $Y2=1.975
r145 25 35 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.7 $Y=1.935
+ $X2=3.7 $Y2=1.81
r146 25 28 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.7 $Y=1.935 $X2=3.7
+ $Y2=1.975
r147 24 44 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.125
+ $X2=2.16 $Y2=2.21
r148 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.405
+ $X2=2.16 $Y2=1.32
r149 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.16 $Y=1.405
+ $X2=2.16 $Y2=2.125
r150 22 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=1.235
+ $X2=1.99 $Y2=1.32
r151 21 22 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.99 $Y=0.535
+ $X2=1.99 $Y2=1.235
r152 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.905 $Y=0.45
+ $X2=1.99 $Y2=0.535
r153 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.905 $Y=0.45
+ $X2=1.64 $Y2=0.45
r154 13 44 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=2.21
+ $X2=2.16 $Y2=2.21
r155 13 15 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.075 $Y=2.21
+ $X2=1.58 $Y2=2.21
r156 4 28 600 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=1.58 $X2=3.66 $Y2=1.975
r157 3 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=2.065 $X2=1.58 $Y2=2.21
r158 2 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.235 $X2=3.675 $Y2=0.51
r159 1 19 182 $w=1.7e-07 $l=2.98706e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.64 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%A_873_316# 1 2 3 4 14 15 18 20 21 23 25 27 30
+ 35
r87 30 32 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=4.502 $Y=0.42
+ $X2=4.502 $Y2=0.585
r88 25 27 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.5 $Y=2.24
+ $X2=6.115 $Y2=2.24
r89 21 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.5 $Y=0.38 $X2=6.06
+ $Y2=0.38
r90 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=2.155
+ $X2=5.5 $Y2=2.24
r91 19 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=1.735
+ $X2=5.415 $Y2=1.65
r92 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.415 $Y=1.735
+ $X2=5.415 $Y2=2.155
r93 18 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=1.565
+ $X2=5.415 $Y2=1.65
r94 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=0.465
+ $X2=5.5 $Y2=0.38
r95 17 18 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=5.415 $Y=0.465
+ $X2=5.415 $Y2=1.565
r96 16 34 3.40825 $w=1.7e-07 $l=1.28938e-07 $layer=LI1_cond $X=4.59 $Y=1.65
+ $X2=4.495 $Y2=1.73
r97 15 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=1.65
+ $X2=5.415 $Y2=1.65
r98 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.33 $Y=1.65
+ $X2=4.59 $Y2=1.65
r99 14 34 3.40825 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=4.485 $Y=1.565
+ $X2=4.495 $Y2=1.73
r100 14 32 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.485 $Y=1.565
+ $X2=4.485 $Y2=0.585
r101 4 27 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.98
+ $Y=2.065 $X2=6.115 $Y2=2.24
r102 3 34 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=4.365
+ $Y=1.58 $X2=4.5 $Y2=1.73
r103 2 23 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=5.86
+ $Y=0.235 $X2=6.06 $Y2=0.38
r104 1 30 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.52 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%X 1 2 3 4 15 18 21 24 25 29 31 32 33 34 35 36
+ 37 38
c58 31 0 2.84211e-20 $X=7.615 $Y=1.495
c59 18 0 3.78084e-20 $X=7.685 $Y=1.065
r60 37 38 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=8.522 $Y=1.87
+ $X2=8.522 $Y2=2.21
r61 37 56 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=8.522 $Y=1.87
+ $X2=8.522 $Y2=1.66
r62 36 56 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=8.522 $Y=1.53
+ $X2=8.522 $Y2=1.66
r63 36 52 7.97845 $w=3.23e-07 $l=2.25e-07 $layer=LI1_cond $X=8.522 $Y=1.53
+ $X2=8.522 $Y2=1.305
r64 35 45 3.98661 $w=3.25e-07 $l=1.2e-07 $layer=LI1_cond $X=8.522 $Y=1.185
+ $X2=8.522 $Y2=1.065
r65 35 52 3.98661 $w=3.25e-07 $l=1.2e-07 $layer=LI1_cond $X=8.522 $Y=1.185
+ $X2=8.522 $Y2=1.305
r66 34 45 7.62385 $w=3.23e-07 $l=2.15e-07 $layer=LI1_cond $X=8.522 $Y=0.85
+ $X2=8.522 $Y2=1.065
r67 33 34 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=8.522 $Y=0.51
+ $X2=8.522 $Y2=0.85
r68 27 29 4.16027 $w=4.58e-07 $l=1.6e-07 $layer=LI1_cond $X=7.525 $Y=0.495
+ $X2=7.685 $Y2=0.495
r69 24 25 3.10188 $w=4.08e-07 $l=8.5e-08 $layer=LI1_cond $X=7.565 $Y=1.92
+ $X2=7.565 $Y2=1.835
r70 22 32 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=1.185
+ $X2=7.685 $Y2=1.185
r71 21 35 2.45386 $w=2.4e-07 $l=1.62e-07 $layer=LI1_cond $X=8.36 $Y=1.185
+ $X2=8.522 $Y2=1.185
r72 21 22 28.3309 $w=2.38e-07 $l=5.9e-07 $layer=LI1_cond $X=8.36 $Y=1.185
+ $X2=7.77 $Y2=1.185
r73 19 32 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.685 $Y=1.305
+ $X2=7.685 $Y2=1.185
r74 19 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.685 $Y=1.305
+ $X2=7.685 $Y2=1.495
r75 18 32 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.685 $Y=1.065
+ $X2=7.685 $Y2=1.185
r76 17 29 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.685 $Y=0.725
+ $X2=7.685 $Y2=0.495
r77 17 18 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.685 $Y=0.725
+ $X2=7.685 $Y2=1.065
r78 15 31 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=7.615 $Y=1.65
+ $X2=7.615 $Y2=1.495
r79 15 25 6.87748 $w=3.08e-07 $l=1.85e-07 $layer=LI1_cond $X=7.615 $Y=1.65
+ $X2=7.615 $Y2=1.835
r80 4 56 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=1.485 $X2=8.445 $Y2=1.66
r81 3 24 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=7.39
+ $Y=1.485 $X2=7.525 $Y2=1.92
r82 2 33 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.235 $X2=8.445 $Y2=0.56
r83 1 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=7.39
+ $Y=0.235 $X2=7.525 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 43 45
+ 50 55 60 68 73 79 82 85 88 91 95
c147 95 0 1.64811e-19 $X=8.97 $Y=0
c148 50 0 1.47056e-19 $X=2.455 $Y=0
r149 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r150 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r151 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r152 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r153 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r154 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r155 77 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.97
+ $Y2=0
r156 77 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.05
+ $Y2=0
r157 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r158 74 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.065
+ $Y2=0
r159 74 76 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.51
+ $Y2=0
r160 73 94 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=8.855 $Y=0
+ $X2=9.027 $Y2=0
r161 73 76 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.855 $Y=0 $X2=8.51
+ $Y2=0
r162 72 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r163 72 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r164 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r165 69 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.27 $Y=0 $X2=7.145
+ $Y2=0
r166 69 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.27 $Y=0 $X2=7.59
+ $Y2=0
r167 68 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.94 $Y=0 $X2=8.065
+ $Y2=0
r168 68 71 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.94 $Y=0 $X2=7.59
+ $Y2=0
r169 67 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r170 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r171 64 67 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r172 64 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r173 63 66 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=6.67
+ $Y2=0
r174 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r175 61 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=0 $X2=4.965
+ $Y2=0
r176 61 63 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.13 $Y=0 $X2=5.29
+ $Y2=0
r177 60 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.02 $Y=0 $X2=7.145
+ $Y2=0
r178 60 66 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.02 $Y=0 $X2=6.67
+ $Y2=0
r179 59 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.83 $Y2=0
r180 59 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r181 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r182 56 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=2.62
+ $Y2=0
r183 56 58 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.785 $Y=0
+ $X2=2.99 $Y2=0
r184 55 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.965
+ $Y2=0
r185 55 58 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=4.8 $Y=0 $X2=2.99
+ $Y2=0
r186 54 83 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.53 $Y2=0
r187 54 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r188 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r189 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r190 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r191 50 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.62
+ $Y2=0
r192 50 53 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=2.455 $Y=0
+ $X2=1.15 $Y2=0
r193 45 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r194 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r195 43 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r196 43 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r197 39 94 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=9.027 $Y2=0
r198 39 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0.38
r199 35 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=0.085
+ $X2=8.065 $Y2=0
r200 35 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.065 $Y=0.085
+ $X2=8.065 $Y2=0.38
r201 31 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=0.085
+ $X2=7.145 $Y2=0
r202 31 33 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=7.145 $Y=0.085
+ $X2=7.145 $Y2=0.51
r203 27 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=0.085
+ $X2=4.965 $Y2=0
r204 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.965 $Y=0.085
+ $X2=4.965 $Y2=0.38
r205 23 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0
r206 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0.38
r207 19 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r208 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r209 6 41 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.235 $X2=8.94 $Y2=0.38
r210 5 37 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=7.81
+ $Y=0.235 $X2=8.025 $Y2=0.38
r211 4 33 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=6.885
+ $Y=0.235 $X2=7.105 $Y2=0.51
r212 3 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.235 $X2=5.04 $Y2=0.38
r213 2 25 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.66 $Y2=0.38
r214 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__maj3_1.pxi.spice
* Created: Tue Sep  1 19:13:59 2020
* 
x_PM_SKY130_FD_SC_HD__MAJ3_1%A N_A_M1005_g N_A_M1006_g N_A_M1007_g N_A_M1003_g A
+ A A A N_A_c_70_n N_A_c_71_n PM_SKY130_FD_SC_HD__MAJ3_1%A
x_PM_SKY130_FD_SC_HD__MAJ3_1%B N_B_M1008_g N_B_M1004_g N_B_M1001_g N_B_M1011_g B
+ B N_B_c_115_n N_B_c_116_n PM_SKY130_FD_SC_HD__MAJ3_1%B
x_PM_SKY130_FD_SC_HD__MAJ3_1%C N_C_M1013_g N_C_M1010_g N_C_c_167_n N_C_c_168_n
+ N_C_M1002_g N_C_M1012_g C C N_C_c_165_n PM_SKY130_FD_SC_HD__MAJ3_1%C
x_PM_SKY130_FD_SC_HD__MAJ3_1%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1008_d
+ N_A_27_47#_M1010_s N_A_27_47#_M1004_d N_A_27_47#_M1009_g N_A_27_47#_M1000_g
+ N_A_27_47#_c_314_p N_A_27_47#_c_224_n N_A_27_47#_c_241_n N_A_27_47#_c_242_n
+ N_A_27_47#_c_225_n N_A_27_47#_c_235_n N_A_27_47#_c_236_n N_A_27_47#_c_237_n
+ N_A_27_47#_c_226_n N_A_27_47#_c_227_n N_A_27_47#_c_228_n N_A_27_47#_c_265_n
+ N_A_27_47#_c_229_n N_A_27_47#_c_230_n N_A_27_47#_c_231_n
+ PM_SKY130_FD_SC_HD__MAJ3_1%A_27_47#
x_PM_SKY130_FD_SC_HD__MAJ3_1%VPWR N_VPWR_M1006_d N_VPWR_M1012_d N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n VPWR N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_334_n N_VPWR_c_342_n VPWR
+ PM_SKY130_FD_SC_HD__MAJ3_1%VPWR
x_PM_SKY130_FD_SC_HD__MAJ3_1%X N_X_M1009_d N_X_M1000_d N_X_c_383_n X X X X X
+ N_X_c_381_n X X PM_SKY130_FD_SC_HD__MAJ3_1%X
x_PM_SKY130_FD_SC_HD__MAJ3_1%VGND N_VGND_M1005_d N_VGND_M1002_d N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n VGND N_VGND_c_414_n
+ N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n VGND
+ PM_SKY130_FD_SC_HD__MAJ3_1%VGND
cc_1 VNB N_A_M1005_g 0.0249701f $X=-0.19 $Y=-0.24 $X2=0.83 $Y2=0.445
cc_2 VNB N_A_M1007_g 0.024996f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=0.445
cc_3 VNB N_A_c_70_n 0.00331023f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=1.16
cc_4 VNB N_A_c_71_n 0.0292864f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.16
cc_5 VNB N_B_M1008_g 0.0251904f $X=-0.19 $Y=-0.24 $X2=0.83 $Y2=0.445
cc_6 VNB N_B_M1001_g 0.0241487f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=0.445
cc_7 VNB N_B_c_115_n 0.0036505f $X=-0.19 $Y=-0.24 $X2=0.83 $Y2=1.16
cc_8 VNB N_B_c_116_n 0.027614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_M1013_g 0.0477881f $X=-0.19 $Y=-0.24 $X2=0.83 $Y2=0.445
cc_10 VNB N_C_M1002_g 0.0304296f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=0.445
cc_11 VNB C 0.00821185f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_12 VNB N_C_c_165_n 0.0301464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_224_n 0.0242776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_225_n 0.00316856f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_226_n 0.00743298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_227_n 0.021153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_228_n 0.00543147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_229_n 0.00281267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_230_n 0.0297614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_231_n 0.0216819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_334_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.53
cc_22 VNB X 0.00666696f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.325
cc_23 VNB N_X_c_381_n 0.0160045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB X 0.0235973f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.53
cc_25 VNB N_VGND_c_410_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=0.995
cc_26 VNB N_VGND_c_411_n 0.00567158f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.325
cc_27 VNB N_VGND_c_412_n 0.0351383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_413_n 0.0064108f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_29 VNB N_VGND_c_414_n 0.0244556f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=2.125
cc_30 VNB N_VGND_c_415_n 0.0244211f $X=-0.19 $Y=-0.24 $X2=1.25 $Y2=1.16
cc_31 VNB N_VGND_c_416_n 0.201216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_417_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.87
cc_33 VPB N_A_M1006_g 0.0242965f $X=-0.19 $Y=1.305 $X2=0.83 $Y2=1.915
cc_34 VPB N_A_M1003_g 0.0268222f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.915
cc_35 VPB A 0.00872573f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_36 VPB N_A_c_70_n 5.31834e-19 $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.16
cc_37 VPB N_A_c_71_n 0.00427902f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.16
cc_38 VPB N_B_M1004_g 0.0246619f $X=-0.19 $Y=1.305 $X2=0.83 $Y2=1.915
cc_39 VPB N_B_M1011_g 0.0252101f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.915
cc_40 VPB N_B_c_115_n 0.00862027f $X=-0.19 $Y=1.305 $X2=0.83 $Y2=1.16
cc_41 VPB N_B_c_116_n 0.00417904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_C_M1013_g 0.0490381f $X=-0.19 $Y=1.305 $X2=0.83 $Y2=0.445
cc_43 VPB N_C_c_167_n 0.138382f $X=-0.19 $Y=1.305 $X2=0.83 $Y2=1.915
cc_44 VPB N_C_c_168_n 0.0129123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_C_M1012_g 0.0471165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB C 0.00282153f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_47 VPB N_C_c_165_n 0.00929012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_M1000_g 0.0250016f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_49 VPB N_A_27_47#_c_224_n 0.0233219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_225_n 0.00165755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_235_n 3.55719e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_236_n 0.00837238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_237_n 0.00204768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_230_n 0.00837392f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_335_n 0.0105088f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=0.995
cc_56 VPB N_VPWR_c_336_n 0.00976536f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=1.325
cc_57 VPB N_VPWR_c_337_n 0.039244f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_58 VPB N_VPWR_c_338_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.785
cc_59 VPB N_VPWR_c_339_n 0.0286522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_340_n 0.024262f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_61 VPB N_VPWR_c_334_n 0.0515307f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.53
cc_62 VPB N_VPWR_c_342_n 0.00330333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_X_c_383_n 0.0123181f $X=-0.19 $Y=1.305 $X2=1.25 $Y2=0.995
cc_64 VPB X 0.0194623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB X 0.00938312f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.53
cc_66 VPB X 0.00644835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 N_A_M1007_g N_B_M1008_g 0.0442567f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_B_M1004_g 0.0442567f $X=1.25 $Y=1.915 $X2=0 $Y2=0
cc_69 N_A_c_70_n N_B_c_115_n 0.0151361f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_c_71_n N_B_c_115_n 0.00978496f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_70_n N_B_c_116_n 2.95512e-19 $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_71_n N_B_c_116_n 0.0442567f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1005_g N_C_M1013_g 0.12866f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_74 A N_C_M1013_g 0.0160523f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_75 N_A_c_70_n N_C_M1013_g 0.00246976f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_C_c_167_n 0.0101565f $X=0.83 $Y=1.915 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_C_c_167_n 0.0102879f $X=1.25 $Y=1.915 $X2=0 $Y2=0
cc_78 A N_C_c_167_n 0.00315449f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_79 A N_A_27_47#_c_224_n 0.0511096f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_80 N_A_c_70_n N_A_27_47#_c_224_n 0.023622f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_A_27_47#_c_241_n 0.00141465f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_A_27_47#_c_242_n 7.174e-19 $X=1.25 $Y=1.915 $X2=0 $Y2=0
cc_83 N_A_M1005_g N_A_27_47#_c_227_n 0.0110822f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_M1007_g N_A_27_47#_c_227_n 0.0156634f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_c_70_n N_A_27_47#_c_227_n 0.0387448f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_c_71_n N_A_27_47#_c_227_n 0.00201785f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_87 A A_109_341# 0.00374721f $X=0.61 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_88 N_A_M1006_g N_VPWR_c_335_n 0.00102427f $X=0.83 $Y=1.915 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VPWR_c_335_n 0.01208f $X=1.25 $Y=1.915 $X2=0 $Y2=0
cc_90 A N_VPWR_c_335_n 0.0385015f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_91 N_A_c_70_n N_VPWR_c_335_n 0.00704809f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_c_71_n N_VPWR_c_335_n 0.00182924f $X=1.25 $Y=1.16 $X2=0 $Y2=0
cc_93 A N_VPWR_c_339_n 0.0116727f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_VPWR_c_334_n 7.83281e-19 $X=0.83 $Y=1.915 $X2=0 $Y2=0
cc_95 N_A_M1003_g N_VPWR_c_334_n 7.52198e-19 $X=1.25 $Y=1.915 $X2=0 $Y2=0
cc_96 A N_VPWR_c_334_n 0.00578509f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_97 N_A_M1005_g N_VGND_c_410_n 0.00946659f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_M1007_g N_VGND_c_410_n 0.00934722f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_M1007_g N_VGND_c_412_n 0.00341689f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_M1005_g N_VGND_c_414_n 0.00341689f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_M1005_g N_VGND_c_416_n 0.00389164f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_M1007_g N_VGND_c_416_n 0.00389164f $X=1.25 $Y=0.445 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_C_c_167_n 0.0102915f $X=1.61 $Y=1.915 $X2=0 $Y2=0
cc_104 N_B_M1011_g N_C_c_167_n 0.00979168f $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_105 N_B_M1001_g N_C_M1002_g 0.0434688f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_106 N_B_M1011_g N_C_M1012_g 0.0434688f $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_107 N_B_M1001_g C 4.57524e-19 $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B_c_116_n N_C_c_165_n 0.0434688f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B_M1008_g N_A_27_47#_c_241_n 0.00676611f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_110 N_B_M1001_g N_A_27_47#_c_241_n 0.00717733f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_111 N_B_M1004_g N_A_27_47#_c_242_n 0.00514254f $X=1.61 $Y=1.915 $X2=0 $Y2=0
cc_112 N_B_M1011_g N_A_27_47#_c_242_n 0.0129294f $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_113 N_B_c_115_n N_A_27_47#_c_242_n 0.0163922f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B_c_116_n N_A_27_47#_c_242_n 3.48906e-19 $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B_M1008_g N_A_27_47#_c_225_n 8.43412e-19 $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_116 N_B_M1001_g N_A_27_47#_c_225_n 0.00394364f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_117 N_B_M1011_g N_A_27_47#_c_225_n 0.00267261f $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_118 N_B_c_115_n N_A_27_47#_c_225_n 0.0369492f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B_c_116_n N_A_27_47#_c_225_n 0.00719527f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_M1004_g N_A_27_47#_c_235_n 5.39025e-19 $X=1.61 $Y=1.915 $X2=0 $Y2=0
cc_121 N_B_M1011_g N_A_27_47#_c_235_n 0.0033736f $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_122 N_B_M1008_g N_A_27_47#_c_227_n 0.00780314f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B_c_115_n N_A_27_47#_c_227_n 0.0316492f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_124 N_B_M1008_g N_A_27_47#_c_228_n 0.00339145f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_125 N_B_M1001_g N_A_27_47#_c_228_n 0.0141438f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_126 N_B_c_116_n N_A_27_47#_c_228_n 6.38322e-19 $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B_M1004_g N_A_27_47#_c_265_n 3.3453e-19 $X=1.61 $Y=1.915 $X2=0 $Y2=0
cc_128 N_B_M1011_g N_A_27_47#_c_265_n 0.00379481f $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_129 N_B_c_115_n N_A_27_47#_c_265_n 0.0102261f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_M1004_g N_VPWR_c_335_n 0.00213046f $X=1.61 $Y=1.915 $X2=0 $Y2=0
cc_131 N_B_M1004_g N_VPWR_c_334_n 9.32477e-19 $X=1.61 $Y=1.915 $X2=0 $Y2=0
cc_132 N_B_M1011_g N_VPWR_c_334_n 9.32477e-19 $X=2.03 $Y=1.915 $X2=0 $Y2=0
cc_133 N_B_M1008_g N_VGND_c_410_n 0.00185594f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_134 N_B_M1008_g N_VGND_c_412_n 0.00414405f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_135 N_B_M1001_g N_VGND_c_412_n 0.00412653f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_136 N_B_M1008_g N_VGND_c_416_n 0.00564955f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_137 N_B_M1001_g N_VGND_c_416_n 0.00563363f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_138 N_C_M1012_g N_A_27_47#_M1000_g 0.0205353f $X=2.39 $Y=1.915 $X2=0 $Y2=0
cc_139 N_C_M1013_g N_A_27_47#_c_224_n 0.0254711f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_140 N_C_M1002_g N_A_27_47#_c_241_n 0.00148577f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_141 N_C_c_167_n N_A_27_47#_c_242_n 0.00680145f $X=2.315 $Y=2.54 $X2=0 $Y2=0
cc_142 N_C_M1012_g N_A_27_47#_c_242_n 0.00305168f $X=2.39 $Y=1.915 $X2=0 $Y2=0
cc_143 N_C_M1002_g N_A_27_47#_c_225_n 0.00699791f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_144 C N_A_27_47#_c_225_n 0.0376219f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_145 N_C_M1012_g N_A_27_47#_c_235_n 0.00333437f $X=2.39 $Y=1.915 $X2=0 $Y2=0
cc_146 N_C_M1012_g N_A_27_47#_c_236_n 0.0187991f $X=2.39 $Y=1.915 $X2=0 $Y2=0
cc_147 C N_A_27_47#_c_236_n 0.0262136f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_148 N_C_c_165_n N_A_27_47#_c_236_n 0.00193861f $X=2.575 $Y=1.16 $X2=0 $Y2=0
cc_149 N_C_M1012_g N_A_27_47#_c_237_n 0.00277534f $X=2.39 $Y=1.915 $X2=0 $Y2=0
cc_150 N_C_M1013_g N_A_27_47#_c_226_n 0.00327202f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_151 N_C_M1013_g N_A_27_47#_c_227_n 0.0139477f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_152 N_C_M1002_g N_A_27_47#_c_228_n 0.00412704f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_153 C N_A_27_47#_c_228_n 0.00498519f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_154 C N_A_27_47#_c_229_n 0.02712f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_155 N_C_c_165_n N_A_27_47#_c_229_n 0.00100653f $X=2.575 $Y=1.16 $X2=0 $Y2=0
cc_156 C N_A_27_47#_c_230_n 0.00101797f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_157 N_C_c_165_n N_A_27_47#_c_230_n 0.0214498f $X=2.575 $Y=1.16 $X2=0 $Y2=0
cc_158 N_C_M1002_g N_A_27_47#_c_231_n 0.0167376f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_159 C N_A_27_47#_c_231_n 0.00316041f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_160 N_C_M1013_g N_VPWR_c_335_n 4.47339e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_161 N_C_c_167_n N_VPWR_c_335_n 0.0212715f $X=2.315 $Y=2.54 $X2=0 $Y2=0
cc_162 N_C_M1012_g N_VPWR_c_336_n 0.0178089f $X=2.39 $Y=1.915 $X2=0 $Y2=0
cc_163 N_C_c_167_n N_VPWR_c_337_n 0.0390544f $X=2.315 $Y=2.54 $X2=0 $Y2=0
cc_164 N_C_c_168_n N_VPWR_c_339_n 0.018084f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_165 N_C_c_167_n N_VPWR_c_334_n 0.0640247f $X=2.315 $Y=2.54 $X2=0 $Y2=0
cc_166 N_C_c_168_n N_VPWR_c_334_n 0.0110038f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_167 C X 0.00226641f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_168 C X 0.00398774f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_169 N_C_M1013_g N_VGND_c_410_n 0.00186677f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_170 N_C_M1002_g N_VGND_c_411_n 0.00700322f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_171 C N_VGND_c_411_n 0.0111716f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_172 N_C_c_165_n N_VGND_c_411_n 9.07191e-19 $X=2.575 $Y=1.16 $X2=0 $Y2=0
cc_173 N_C_M1002_g N_VGND_c_412_n 0.00585385f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_174 N_C_M1013_g N_VGND_c_414_n 0.00428022f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_175 N_C_M1013_g N_VGND_c_416_n 0.00678186f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_176 N_C_M1002_g N_VGND_c_416_n 0.00973615f $X=2.39 $Y=0.445 $X2=0 $Y2=0
cc_177 C N_VGND_c_416_n 0.00606394f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_236_n N_VPWR_M1012_d 0.0170332f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_242_n N_VPWR_c_335_n 0.00921613f $X=2.075 $Y=1.947 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_M1000_g N_VPWR_c_336_n 0.0105018f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_242_n N_VPWR_c_336_n 0.0126928f $X=2.075 $Y=1.947 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_236_n N_VPWR_c_336_n 0.0255687f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_242_n N_VPWR_c_337_n 0.00900861f $X=2.075 $Y=1.947 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_224_n N_VPWR_c_339_n 0.00487678f $X=0.26 $Y=1.915 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_M1000_g N_VPWR_c_340_n 0.00585385f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_M1000_g N_VPWR_c_334_n 0.0125071f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_224_n N_VPWR_c_334_n 0.0079931f $X=0.26 $Y=1.915 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_242_n N_VPWR_c_334_n 0.0146039f $X=2.075 $Y=1.947 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_242_n A_421_341# 0.00417044f $X=2.075 $Y=1.947 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_27_47#_c_235_n A_421_341# 0.0012025f $X=2.16 $Y=1.815 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_27_47#_M1000_g N_X_c_383_n 0.00761163f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_230_n X 8.46963e-19 $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_231_n N_X_c_381_n 0.0191414f $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_27_47#_M1000_g X 0.00238576f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_237_n X 0.006117f $X=3.01 $Y=1.495 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_229_n X 0.0249708f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_230_n X 0.00819657f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_231_n X 0.00279048f $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1000_g X 0.0187679f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_236_n X 0.0139683f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_230_n X 4.22311e-19 $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_314_p N_VGND_c_410_n 0.00817147f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_241_n N_VGND_c_410_n 0.00784134f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_227_n N_VGND_c_410_n 0.020154f $X=1.655 $Y=0.732 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_241_n N_VGND_c_411_n 0.00655764f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_231_n N_VGND_c_411_n 0.00568126f $X=3.115 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_241_n N_VGND_c_412_n 0.0183123f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_227_n N_VGND_c_412_n 0.0074151f $X=1.655 $Y=0.732 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_228_n N_VGND_c_412_n 0.0039792f $X=2.16 $Y=0.732 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_314_p N_VGND_c_414_n 0.0161917f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_227_n N_VGND_c_414_n 0.00788392f $X=1.655 $Y=0.732 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_231_n N_VGND_c_415_n 0.00585385f $X=3.115 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_M1013_s N_VGND_c_416_n 0.00208516f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1008_d N_VGND_c_416_n 0.00216807f $X=1.685 $Y=0.235 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_314_p N_VGND_c_416_n 0.00993603f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_241_n N_VGND_c_416_n 0.01217f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_227_n N_VGND_c_416_n 0.0248377f $X=1.655 $Y=0.732 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_228_n N_VGND_c_416_n 0.00681187f $X=2.16 $Y=0.732 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_231_n N_VGND_c_416_n 0.0125071f $X=3.115 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_228_n A_421_47# 0.00163974f $X=2.16 $Y=0.732 $X2=-0.19
+ $Y2=-0.24
cc_221 N_VPWR_c_334_n N_X_M1000_d 0.0056004f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_336_n N_X_c_383_n 0.013822f $X=2.72 $Y=1.93 $X2=0 $Y2=0
cc_223 N_VPWR_c_340_n N_X_c_383_n 0.0238006f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_334_n N_X_c_383_n 0.0130102f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_336_n X 0.0139407f $X=2.72 $Y=1.93 $X2=0 $Y2=0
cc_226 N_X_c_381_n N_VGND_c_411_n 0.00965721f $X=3.42 $Y=0.38 $X2=0 $Y2=0
cc_227 N_X_c_381_n N_VGND_c_415_n 0.0237331f $X=3.42 $Y=0.38 $X2=0 $Y2=0
cc_228 N_X_M1009_d N_VGND_c_416_n 0.0056004f $X=3.18 $Y=0.235 $X2=0 $Y2=0
cc_229 N_X_c_381_n N_VGND_c_416_n 0.0129969f $X=3.42 $Y=0.38 $X2=0 $Y2=0
cc_230 A_109_47# N_VGND_c_416_n 0.00251327f $X=0.545 $Y=0.235 $X2=3.45 $Y2=0
cc_231 N_VGND_c_416_n A_265_47# 0.00251327f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_232 N_VGND_c_416_n A_421_47# 0.00462548f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__or3b_2.pxi.spice
* Created: Tue Sep  1 19:28:08 2020
* 
x_PM_SKY130_FD_SC_HD__OR3B_2%C_N N_C_N_M1009_g N_C_N_M1010_g C_N C_N
+ N_C_N_c_72_n PM_SKY130_FD_SC_HD__OR3B_2%C_N
x_PM_SKY130_FD_SC_HD__OR3B_2%A_176_21# N_A_176_21#_M1005_d N_A_176_21#_M1006_d
+ N_A_176_21#_M1008_d N_A_176_21#_c_98_n N_A_176_21#_M1002_g N_A_176_21#_M1007_g
+ N_A_176_21#_c_99_n N_A_176_21#_M1004_g N_A_176_21#_M1011_g N_A_176_21#_c_100_n
+ N_A_176_21#_c_101_n N_A_176_21#_c_102_n N_A_176_21#_c_188_p
+ N_A_176_21#_c_103_n N_A_176_21#_c_104_n N_A_176_21#_c_105_n
+ N_A_176_21#_c_106_n N_A_176_21#_c_107_n N_A_176_21#_c_112_n
+ N_A_176_21#_c_108_n PM_SKY130_FD_SC_HD__OR3B_2%A_176_21#
x_PM_SKY130_FD_SC_HD__OR3B_2%A N_A_M1005_g N_A_M1001_g A A N_A_c_202_n
+ N_A_c_203_n PM_SKY130_FD_SC_HD__OR3B_2%A
x_PM_SKY130_FD_SC_HD__OR3B_2%B N_B_M1003_g N_B_M1000_g B B N_B_c_249_n
+ PM_SKY130_FD_SC_HD__OR3B_2%B
x_PM_SKY130_FD_SC_HD__OR3B_2%A_27_47# N_A_27_47#_M1009_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1006_g N_A_27_47#_M1008_g N_A_27_47#_c_277_n N_A_27_47#_c_278_n
+ N_A_27_47#_c_279_n N_A_27_47#_c_297_n N_A_27_47#_c_280_n N_A_27_47#_c_285_n
+ N_A_27_47#_c_286_n N_A_27_47#_c_287_n N_A_27_47#_c_311_n N_A_27_47#_c_312_n
+ N_A_27_47#_c_288_n N_A_27_47#_c_281_n N_A_27_47#_c_282_n
+ PM_SKY130_FD_SC_HD__OR3B_2%A_27_47#
x_PM_SKY130_FD_SC_HD__OR3B_2%VPWR N_VPWR_M1010_d N_VPWR_M1011_d N_VPWR_c_377_n
+ N_VPWR_c_378_n VPWR N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n
+ N_VPWR_c_376_n N_VPWR_c_383_n N_VPWR_c_384_n PM_SKY130_FD_SC_HD__OR3B_2%VPWR
x_PM_SKY130_FD_SC_HD__OR3B_2%X N_X_M1002_s N_X_M1007_s N_X_c_423_n N_X_c_433_n X
+ PM_SKY130_FD_SC_HD__OR3B_2%X
x_PM_SKY130_FD_SC_HD__OR3B_2%VGND N_VGND_M1009_d N_VGND_M1004_d N_VGND_M1003_d
+ N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n
+ N_VGND_c_462_n N_VGND_c_463_n VGND N_VGND_c_464_n N_VGND_c_465_n
+ N_VGND_c_466_n N_VGND_c_467_n PM_SKY130_FD_SC_HD__OR3B_2%VGND
cc_1 VNB N_C_N_M1009_g 0.0359264f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB C_N 0.00882738f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_72_n 0.0383384f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_176_21#_c_98_n 0.0163075f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_176_21#_c_99_n 0.0166084f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_6 VNB N_A_176_21#_c_100_n 3.67994e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_176_21#_c_101_n 0.00617416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_176_21#_c_102_n 0.00455355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_176_21#_c_103_n 0.00650435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_176_21#_c_104_n 0.0116331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_176_21#_c_105_n 0.0228353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_176_21#_c_106_n 0.00292732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_176_21#_c_107_n 0.0125721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_176_21#_c_108_n 0.0361096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_M1005_g 0.0265668f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_16 VNB N_A_c_202_n 0.0193541f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_17 VNB N_A_c_203_n 0.00397264f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_18 VNB N_B_M1003_g 0.0389657f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_19 VNB N_A_27_47#_M1006_g 0.0309843f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A_27_47#_c_277_n 0.0182008f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_21 VNB N_A_27_47#_c_278_n 0.00373709f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_22 VNB N_A_27_47#_c_279_n 0.00930805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_280_n 0.00665521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_281_n 0.00311094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_282_n 0.0221007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_376_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_423_n 6.68115e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_457_n 0.00467885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_458_n 0.00418552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_459_n 0.00107531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_460_n 0.0178916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_461_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_462_n 0.0203929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_463_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_464_n 0.0161844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_465_n 0.0159724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_466_n 0.186066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_467_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_C_N_M1010_g 0.0489853f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.01
cc_40 VPB C_N 0.0160532f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_41 VPB N_C_N_c_72_n 0.0100411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_42 VPB N_A_176_21#_M1007_g 0.0202141f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_43 VPB N_A_176_21#_M1011_g 0.0209504f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.53
cc_44 VPB N_A_176_21#_c_105_n 0.00921272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_176_21#_c_112_n 0.0206507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_176_21#_c_108_n 0.00569201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_M1001_g 0.0189131f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.01
cc_48 VPB N_A_c_202_n 0.00442471f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_A_c_203_n 0.00175482f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_50 VPB N_B_M1003_g 0.0258583f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_51 VPB B 0.0350186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_B_c_249_n 0.0385933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_M1008_g 0.0217657f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_54 VPB N_A_27_47#_c_280_n 0.00552992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_285_n 0.00503197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_286_n 0.0013109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_287_n 0.0187262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_288_n 9.06945e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_281_n 3.5559e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_282_n 0.00573807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_377_n 0.00980336f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_62 VPB N_VPWR_c_378_n 0.00773614f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_63 VPB N_VPWR_c_379_n 0.0172683f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_64 VPB N_VPWR_c_380_n 0.0121472f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.53
cc_65 VPB N_VPWR_c_381_n 0.0394927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_376_n 0.0602099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_383_n 0.00565096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_384_n 0.00510392f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_X_c_423_n 0.00152849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 N_C_N_M1009_g N_A_176_21#_c_98_n 0.0203819f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_71 N_C_N_M1010_g N_A_176_21#_M1007_g 0.0203819f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_72 N_C_N_c_72_n N_A_176_21#_c_108_n 0.0203819f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_73 N_C_N_M1009_g N_A_27_47#_c_277_n 0.00233406f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_74 N_C_N_M1009_g N_A_27_47#_c_278_n 0.0170801f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_75 C_N N_A_27_47#_c_278_n 0.0060742f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_C_N_c_72_n N_A_27_47#_c_278_n 0.0012291f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_77 C_N N_A_27_47#_c_279_n 0.0227094f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 N_C_N_c_72_n N_A_27_47#_c_279_n 0.00599978f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C_N_M1010_g N_A_27_47#_c_297_n 0.0151922f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_80 C_N N_A_27_47#_c_297_n 0.00445498f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_81 N_C_N_M1009_g N_A_27_47#_c_280_n 0.0130087f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_82 C_N N_A_27_47#_c_280_n 0.042517f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 C_N N_A_27_47#_c_287_n 0.0223722f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_84 N_C_N_c_72_n N_A_27_47#_c_287_n 8.87396e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_85 N_C_N_M1010_g N_VPWR_c_377_n 0.00394846f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_86 N_C_N_M1010_g N_VPWR_c_379_n 0.00378081f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_87 N_C_N_M1010_g N_VPWR_c_376_n 0.00502381f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_88 N_C_N_M1009_g N_X_c_423_n 8.17584e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_89 N_C_N_M1009_g N_VGND_c_457_n 0.00278284f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_90 N_C_N_M1009_g N_VGND_c_460_n 0.00439206f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_91 N_C_N_M1009_g N_VGND_c_466_n 0.00712566f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_176_21#_c_99_n N_A_M1005_g 0.0183242f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_176_21#_c_100_n N_A_M1005_g 3.49988e-19 $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_176_21#_c_101_n N_A_M1005_g 0.0122183f $X=1.99 $Y=0.82 $X2=0 $Y2=0
cc_95 N_A_176_21#_c_102_n N_A_M1005_g 7.00739e-19 $X=1.595 $Y=0.82 $X2=0 $Y2=0
cc_96 N_A_176_21#_c_106_n N_A_M1005_g 0.00164017f $X=2.075 $Y=0.78 $X2=0 $Y2=0
cc_97 N_A_176_21#_M1011_g N_A_M1001_g 0.0239964f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_176_21#_c_100_n N_A_c_202_n 7.76354e-19 $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_176_21#_c_101_n N_A_c_202_n 0.00270709f $X=1.99 $Y=0.82 $X2=0 $Y2=0
cc_100 N_A_176_21#_c_106_n N_A_c_202_n 2.55256e-19 $X=2.075 $Y=0.78 $X2=0 $Y2=0
cc_101 N_A_176_21#_c_108_n N_A_c_202_n 0.01929f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_176_21#_M1011_g N_A_c_203_n 0.00284284f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_176_21#_c_100_n N_A_c_203_n 0.0147766f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_176_21#_c_101_n N_A_c_203_n 0.0226185f $X=1.99 $Y=0.82 $X2=0 $Y2=0
cc_105 N_A_176_21#_c_103_n N_A_c_203_n 0.00417568f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_176_21#_c_106_n N_A_c_203_n 0.0154664f $X=2.075 $Y=0.78 $X2=0 $Y2=0
cc_107 N_A_176_21#_c_108_n N_A_c_203_n 0.00188403f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_176_21#_c_103_n N_B_M1003_g 0.0151583f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_176_21#_c_106_n N_B_M1003_g 0.00253635f $X=2.075 $Y=0.78 $X2=0 $Y2=0
cc_110 N_A_176_21#_c_112_n B 0.0214764f $X=3.05 $Y=1.71 $X2=0 $Y2=0
cc_111 N_A_176_21#_c_103_n N_A_27_47#_M1006_g 0.0128071f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_112 N_A_176_21#_c_105_n N_A_27_47#_M1006_g 0.00569309f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_113 N_A_176_21#_c_105_n N_A_27_47#_M1008_g 0.00334083f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_114 N_A_176_21#_c_112_n N_A_27_47#_M1008_g 9.05821e-19 $X=3.05 $Y=1.71 $X2=0
+ $Y2=0
cc_115 N_A_176_21#_c_98_n N_A_27_47#_c_278_n 0.00131401f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_116 N_A_176_21#_c_98_n N_A_27_47#_c_280_n 0.00846484f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_117 N_A_176_21#_c_112_n N_A_27_47#_c_285_n 0.00663023f $X=3.05 $Y=1.71 $X2=0
+ $Y2=0
cc_118 N_A_176_21#_c_105_n N_A_27_47#_c_286_n 0.00783501f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_119 N_A_176_21#_M1007_g N_A_27_47#_c_311_n 0.00162764f $X=0.955 $Y=1.985
+ $X2=0 $Y2=0
cc_120 N_A_176_21#_M1007_g N_A_27_47#_c_312_n 0.0135693f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_176_21#_M1011_g N_A_27_47#_c_312_n 0.0133355f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_176_21#_c_100_n N_A_27_47#_c_312_n 0.00327749f $X=1.36 $Y=1.16 $X2=0
+ $Y2=0
cc_123 N_A_176_21#_M1011_g N_A_27_47#_c_288_n 0.00257575f $X=1.375 $Y=1.985
+ $X2=0 $Y2=0
cc_124 N_A_176_21#_c_103_n N_A_27_47#_c_281_n 0.0223157f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_125 N_A_176_21#_c_105_n N_A_27_47#_c_281_n 0.0240581f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_126 N_A_176_21#_c_103_n N_A_27_47#_c_282_n 0.00305475f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_127 N_A_176_21#_c_105_n N_A_27_47#_c_282_n 0.00753642f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_128 N_A_176_21#_c_107_n N_A_27_47#_c_282_n 2.9537e-19 $X=2.982 $Y=0.715 $X2=0
+ $Y2=0
cc_129 N_A_176_21#_c_112_n N_A_27_47#_c_282_n 2.2867e-19 $X=3.05 $Y=1.71 $X2=0
+ $Y2=0
cc_130 N_A_176_21#_M1007_g N_VPWR_c_377_n 0.010086f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_176_21#_M1011_g N_VPWR_c_377_n 0.00124016f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_176_21#_M1007_g N_VPWR_c_378_n 0.0012252f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_176_21#_M1011_g N_VPWR_c_378_n 0.0097367f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_176_21#_M1007_g N_VPWR_c_380_n 0.00344532f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_176_21#_M1011_g N_VPWR_c_380_n 0.00358919f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_176_21#_M1007_g N_VPWR_c_376_n 0.00407565f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_176_21#_M1011_g N_VPWR_c_376_n 0.00422197f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_176_21#_c_98_n N_X_c_423_n 0.00958406f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_176_21#_M1007_g N_X_c_423_n 0.00362416f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_176_21#_c_99_n N_X_c_423_n 0.00358135f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_176_21#_M1011_g N_X_c_423_n 0.00153756f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_176_21#_c_100_n N_X_c_423_n 0.0268466f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_176_21#_c_102_n N_X_c_423_n 0.0098479f $X=1.595 $Y=0.82 $X2=0 $Y2=0
cc_144 N_A_176_21#_c_108_n N_X_c_423_n 0.0116158f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_176_21#_M1007_g N_X_c_433_n 0.00460053f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_176_21#_M1011_g N_X_c_433_n 0.00426043f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_176_21#_c_100_n N_X_c_433_n 0.00322481f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_176_21#_c_108_n N_X_c_433_n 0.00344981f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_176_21#_c_98_n X 0.0062773f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_176_21#_c_108_n X 0.00285198f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_176_21#_c_101_n N_VGND_M1004_d 0.00145046f $X=1.99 $Y=0.82 $X2=0
+ $Y2=0
cc_152 N_A_176_21#_c_102_n N_VGND_M1004_d 0.00102401f $X=1.595 $Y=0.82 $X2=0
+ $Y2=0
cc_153 N_A_176_21#_c_103_n N_VGND_M1003_d 0.00160115f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_176_21#_c_98_n N_VGND_c_457_n 0.00514031f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_A_176_21#_c_99_n N_VGND_c_458_n 0.00466764f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_156 N_A_176_21#_c_101_n N_VGND_c_458_n 0.00734233f $X=1.99 $Y=0.82 $X2=0
+ $Y2=0
cc_157 N_A_176_21#_c_102_n N_VGND_c_458_n 0.00590088f $X=1.595 $Y=0.82 $X2=0
+ $Y2=0
cc_158 N_A_176_21#_c_103_n N_VGND_c_459_n 0.0160613f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_176_21#_c_98_n N_VGND_c_462_n 0.00442618f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_176_21#_c_99_n N_VGND_c_462_n 0.00560999f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A_176_21#_c_102_n N_VGND_c_462_n 9.64229e-19 $X=1.595 $Y=0.82 $X2=0
+ $Y2=0
cc_162 N_A_176_21#_c_101_n N_VGND_c_464_n 0.00417479f $X=1.99 $Y=0.82 $X2=0
+ $Y2=0
cc_163 N_A_176_21#_c_188_p N_VGND_c_464_n 0.00854817f $X=2.075 $Y=0.47 $X2=0
+ $Y2=0
cc_164 N_A_176_21#_c_103_n N_VGND_c_464_n 0.00232396f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_165 N_A_176_21#_c_103_n N_VGND_c_465_n 0.00232396f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_176_21#_c_104_n N_VGND_c_465_n 0.0132221f $X=2.915 $Y=0.47 $X2=0
+ $Y2=0
cc_167 N_A_176_21#_c_107_n N_VGND_c_465_n 0.00108171f $X=2.982 $Y=0.715 $X2=0
+ $Y2=0
cc_168 N_A_176_21#_c_98_n N_VGND_c_466_n 0.00743728f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_176_21#_c_99_n N_VGND_c_466_n 0.00647293f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_176_21#_c_101_n N_VGND_c_466_n 0.00750204f $X=1.99 $Y=0.82 $X2=0
+ $Y2=0
cc_171 N_A_176_21#_c_102_n N_VGND_c_466_n 0.00745835f $X=1.595 $Y=0.82 $X2=0
+ $Y2=0
cc_172 N_A_176_21#_c_188_p N_VGND_c_466_n 0.00628404f $X=2.075 $Y=0.47 $X2=0
+ $Y2=0
cc_173 N_A_176_21#_c_103_n N_VGND_c_466_n 0.00970544f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_176_21#_c_104_n N_VGND_c_466_n 0.00945913f $X=2.915 $Y=0.47 $X2=0
+ $Y2=0
cc_175 N_A_176_21#_c_107_n N_VGND_c_466_n 0.00153781f $X=2.982 $Y=0.715 $X2=0
+ $Y2=0
cc_176 N_A_M1005_g N_B_M1003_g 0.0221593f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_177 N_A_M1001_g N_B_M1003_g 0.0338134f $X=1.865 $Y=1.695 $X2=0 $Y2=0
cc_178 N_A_c_202_n N_B_M1003_g 0.0213853f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_203_n N_B_M1003_g 0.0124924f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_203_n N_A_27_47#_M1008_g 2.50323e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_M1001_g N_A_27_47#_c_285_n 0.011183f $X=1.865 $Y=1.695 $X2=0 $Y2=0
cc_182 N_A_c_202_n N_A_27_47#_c_285_n 3.01349e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_c_203_n N_A_27_47#_c_286_n 0.0162706f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_M1001_g N_A_27_47#_c_288_n 0.0025456f $X=1.865 $Y=1.695 $X2=0 $Y2=0
cc_185 N_A_c_203_n N_A_27_47#_c_288_n 0.0280576f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_203_n N_A_27_47#_c_281_n 0.0148056f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_c_203_n N_A_27_47#_c_282_n 2.25713e-19 $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_203_n N_VPWR_M1011_d 0.00201923f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_M1001_g N_VPWR_c_381_n 0.00317443f $X=1.865 $Y=1.695 $X2=0 $Y2=0
cc_190 N_A_M1001_g N_VPWR_c_376_n 0.00403572f $X=1.865 $Y=1.695 $X2=0 $Y2=0
cc_191 N_A_c_203_n N_X_c_423_n 0.00581448f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_M1001_g N_X_c_433_n 5.16539e-19 $X=1.865 $Y=1.695 $X2=0 $Y2=0
cc_193 N_A_c_203_n N_X_c_433_n 0.00542099f $X=1.865 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_c_203_n A_388_297# 0.00168094f $X=1.865 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_195 N_A_M1005_g N_VGND_c_458_n 0.00279433f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_196 N_A_M1005_g N_VGND_c_459_n 5.73165e-19 $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_197 N_A_M1005_g N_VGND_c_464_n 0.00413798f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_198 N_A_M1005_g N_VGND_c_466_n 0.00598057f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_199 N_B_M1003_g N_A_27_47#_M1006_g 0.0247458f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_200 N_B_M1003_g N_A_27_47#_M1008_g 0.0316547f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_201 B N_A_27_47#_M1008_g 0.00649556f $X=2.91 $Y=2.125 $X2=0 $Y2=0
cc_202 N_B_M1003_g N_A_27_47#_c_285_n 0.0142699f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_203 B N_A_27_47#_c_285_n 0.0543392f $X=2.91 $Y=2.125 $X2=0 $Y2=0
cc_204 N_B_c_249_n N_A_27_47#_c_285_n 0.00120401f $X=2.285 $Y=2.28 $X2=0 $Y2=0
cc_205 N_B_M1003_g N_A_27_47#_c_286_n 0.00568321f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_206 N_B_M1003_g N_A_27_47#_c_288_n 2.62061e-19 $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_207 N_B_M1003_g N_A_27_47#_c_281_n 0.00354236f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_208 N_B_M1003_g N_A_27_47#_c_282_n 0.019405f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_209 B N_VPWR_c_378_n 0.0130812f $X=2.91 $Y=2.125 $X2=0 $Y2=0
cc_210 N_B_c_249_n N_VPWR_c_378_n 0.00158436f $X=2.285 $Y=2.28 $X2=0 $Y2=0
cc_211 B N_VPWR_c_381_n 0.0477704f $X=2.91 $Y=2.125 $X2=0 $Y2=0
cc_212 N_B_c_249_n N_VPWR_c_381_n 0.00749157f $X=2.285 $Y=2.28 $X2=0 $Y2=0
cc_213 B N_VPWR_c_376_n 0.0420525f $X=2.91 $Y=2.125 $X2=0 $Y2=0
cc_214 N_B_c_249_n N_VPWR_c_376_n 0.0106165f $X=2.285 $Y=2.28 $X2=0 $Y2=0
cc_215 N_B_M1003_g N_VGND_c_459_n 0.00712901f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_216 N_B_M1003_g N_VGND_c_464_n 0.00322006f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_217 N_B_M1003_g N_VGND_c_466_n 0.00390029f $X=2.285 $Y=0.475 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_280_n N_VPWR_M1010_d 0.00417632f $X=0.68 $Y=1.81 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_27_47#_c_311_n N_VPWR_M1010_d 0.0024773f $X=0.68 $Y=1.925 $X2=-0.19
+ $Y2=-0.24
cc_220 N_A_27_47#_c_312_n N_VPWR_M1010_d 0.00276232f $X=1.55 $Y=1.912 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_27_47#_c_312_n N_VPWR_M1011_d 0.00203539f $X=1.55 $Y=1.912 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_288_n N_VPWR_M1011_d 0.0089384f $X=1.72 $Y=1.912 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_311_n N_VPWR_c_377_n 0.0138837f $X=0.68 $Y=1.925 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_312_n N_VPWR_c_377_n 0.0065098f $X=1.55 $Y=1.912 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_285_n N_VPWR_c_378_n 0.00196088f $X=2.49 $Y=1.87 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_312_n N_VPWR_c_378_n 0.0185039f $X=1.55 $Y=1.912 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_297_n N_VPWR_c_379_n 0.00272266f $X=0.595 $Y=1.925 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_287_n N_VPWR_c_379_n 0.00662803f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_312_n N_VPWR_c_380_n 0.00707194f $X=1.55 $Y=1.912 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_297_n N_VPWR_c_376_n 0.00572244f $X=0.595 $Y=1.925 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_285_n N_VPWR_c_376_n 0.00710536f $X=2.49 $Y=1.87 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_287_n N_VPWR_c_376_n 0.00838075f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_311_n N_VPWR_c_376_n 7.87123e-19 $X=0.68 $Y=1.925 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_312_n N_VPWR_c_376_n 0.0147317f $X=1.55 $Y=1.912 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_312_n N_X_M1007_s 0.00442755f $X=1.55 $Y=1.912 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_277_n N_X_c_423_n 0.00299513f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_278_n N_X_c_423_n 0.0134531f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_280_n N_X_c_423_n 0.0420777f $X=0.68 $Y=1.81 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_280_n N_X_c_433_n 0.0152771f $X=0.68 $Y=1.81 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_312_n N_X_c_433_n 0.0199837f $X=1.55 $Y=1.912 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_285_n A_388_297# 0.00162642f $X=2.49 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_242 N_A_27_47#_c_285_n A_472_297# 0.0027472f $X=2.49 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_27_47#_c_286_n A_472_297# 0.00318603f $X=2.575 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_c_278_n N_VGND_M1009_d 0.00309755f $X=0.595 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_245 N_A_27_47#_c_278_n N_VGND_c_457_n 0.0143363f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_246 N_A_27_47#_M1006_g N_VGND_c_459_n 0.00953333f $X=2.705 $Y=0.475 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_277_n N_VGND_c_460_n 0.014595f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_278_n N_VGND_c_460_n 0.00343878f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1006_g N_VGND_c_465_n 0.00322006f $X=2.705 $Y=0.475 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1009_s N_VGND_c_466_n 0.00236396f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1006_g N_VGND_c_466_n 0.00468173f $X=2.705 $Y=0.475 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_277_n N_VGND_c_466_n 0.00973659f $X=0.26 $Y=0.455 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_278_n N_VGND_c_466_n 0.00645338f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_376_n N_X_M1007_s 0.00333025f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_255 X N_VGND_c_457_n 0.0222902f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_256 X N_VGND_c_462_n 0.0187386f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_257 N_X_M1002_s N_VGND_c_466_n 0.00223333f $X=1.03 $Y=0.235 $X2=0 $Y2=0
cc_258 X N_VGND_c_466_n 0.0126517f $X=1.07 $Y=0.425 $X2=0 $Y2=0

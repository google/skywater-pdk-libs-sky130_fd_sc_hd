* File: sky130_fd_sc_hd__a2111o_1.spice
* Created: Thu Aug 27 13:58:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111o_1.pex.spice"
.subckt sky130_fd_sc_hd__a2111o_1  VNB VPB D1 C1 B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_85_193#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.274625 AS=0.2145 PD=1.495 PS=1.96 NRD=8.304 NRS=4.608 M=1 R=4.33333
+ SA=75000.3 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1011 N_A_85_193#_M1011_d N_D1_M1011_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.274625 PD=0.96 PS=1.495 NRD=0 NRS=32.304 M=1 R=4.33333
+ SA=75001.2 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_C1_M1004_g N_A_85_193#_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.10075 PD=1.01 PS=0.96 NRD=7.38 NRS=5.532 M=1 R=4.33333
+ SA=75001.7 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_85_193#_M1009_d N_B1_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.117 PD=1.22 PS=1.01 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75002.2
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1007 A_660_47# N_A1_M1007_g N_A_85_193#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.082875 AS=0.18525 PD=0.905 PS=1.22 NRD=13.38 NRS=53.532 M=1 R=4.33333
+ SA=75002.9 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g A_660_47# VNB NSHORT L=0.15 W=0.65 AD=0.1885
+ AS=0.082875 PD=1.88 PS=0.905 NRD=0 NRS=13.38 M=1 R=4.33333 SA=75003.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_85_193#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.29 PD=2.53 PS=2.58 NRD=0 NRS=0.9653 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 A_334_297# N_D1_M1006_g N_A_85_193#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.125 AS=0.385 PD=1.25 PS=2.77 NRD=13.7703 NRS=23.6203 M=1 R=6.66667
+ SA=75000.3 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1002 A_414_297# N_C1_M1002_g A_334_297# VPB PHIGHVT L=0.15 W=1 AD=0.18
+ AS=0.125 PD=1.36 PS=1.25 NRD=24.6053 NRS=13.7703 M=1 R=6.66667 SA=75000.7
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_A_516_297#_M1003_d N_B1_M1003_g A_414_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.18 PD=1.56 PS=1.36 NRD=56.1253 NRS=24.6053 M=1 R=6.66667
+ SA=75001.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_516_297#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=1.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_516_297#_M1005_d N_A2_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.29 AS=0.135 PD=2.58 PS=1.27 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__a2111o_1.pxi.spice"
*
.ends
*
*

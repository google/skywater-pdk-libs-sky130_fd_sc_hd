* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_16.pxi.spice
* Created: Tue Sep  1 19:11:02 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%A N_A_M1000_g N_A_M1001_g
+ N_A_M1002_g N_A_M1003_g N_A_M1004_g N_A_M1005_g N_A_M1007_g N_A_M1006_g
+ N_A_M1008_g N_A_M1009_g N_A_M1011_g N_A_M1010_g N_A_M1016_g N_A_M1012_g
+ N_A_M1017_g N_A_M1013_g N_A_M1018_g N_A_M1014_g N_A_c_125_n N_A_c_126_n
+ N_A_M1021_g N_A_M1015_g N_A_M1023_g N_A_M1019_g N_A_M1024_g N_A_M1020_g
+ N_A_M1026_g N_A_M1022_g N_A_M1032_g N_A_M1025_g N_A_M1033_g N_A_M1027_g
+ N_A_M1035_g N_A_M1028_g N_A_M1036_g N_A_M1029_g N_A_M1037_g N_A_M1030_g
+ N_A_M1031_g N_A_M1034_g N_A_M1038_g N_A_M1039_g A N_A_c_229_p N_A_c_235_p
+ N_A_c_243_p N_A_c_309_p N_A_c_320_p N_A_c_137_n N_A_c_138_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%KAPWR N_KAPWR_M1000_d
+ N_KAPWR_M1001_d N_KAPWR_M1003_d N_KAPWR_M1006_d N_KAPWR_M1010_d
+ N_KAPWR_M1013_d N_KAPWR_M1015_d N_KAPWR_M1020_d N_KAPWR_M1025_d
+ N_KAPWR_M1028_d N_KAPWR_M1030_d N_KAPWR_M1034_d N_KAPWR_M1039_d
+ N_KAPWR_c_473_n N_KAPWR_c_479_n N_KAPWR_c_481_n N_KAPWR_c_482_n
+ N_KAPWR_c_557_p N_KAPWR_c_484_n N_KAPWR_c_562_p N_KAPWR_c_486_n
+ N_KAPWR_c_488_n N_KAPWR_c_490_n N_KAPWR_c_491_n N_KAPWR_c_493_n
+ N_KAPWR_c_495_n N_KAPWR_c_496_n N_KAPWR_c_498_n N_KAPWR_c_499_n
+ N_KAPWR_c_501_n N_KAPWR_c_502_n N_KAPWR_c_504_n N_KAPWR_c_505_n
+ N_KAPWR_c_587_p N_KAPWR_c_507_n N_KAPWR_c_592_p N_KAPWR_c_509_n
+ N_KAPWR_c_598_p KAPWR N_KAPWR_c_474_n N_KAPWR_c_513_n N_KAPWR_c_515_n
+ N_KAPWR_c_517_n N_KAPWR_c_519_n N_KAPWR_c_521_n N_KAPWR_c_523_n
+ N_KAPWR_c_525_n N_KAPWR_c_527_n N_KAPWR_c_529_n N_KAPWR_c_475_n
+ N_KAPWR_c_476_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%Y N_Y_M1004_s N_Y_M1008_s
+ N_Y_M1016_s N_Y_M1018_s N_Y_M1023_s N_Y_M1026_s N_Y_M1033_s N_Y_M1036_s
+ N_Y_M1000_s N_Y_M1002_s N_Y_M1005_s N_Y_M1009_s N_Y_M1012_s N_Y_M1014_s
+ N_Y_M1019_s N_Y_M1022_s N_Y_M1027_s N_Y_M1029_s N_Y_M1031_s N_Y_M1038_s
+ N_Y_c_726_n N_Y_c_898_n N_Y_c_727_n N_Y_c_728_n N_Y_c_718_n N_Y_c_730_n
+ N_Y_c_719_n N_Y_c_732_n N_Y_c_720_n N_Y_c_734_n N_Y_c_721_n N_Y_c_722_n
+ N_Y_c_737_n N_Y_c_723_n N_Y_c_739_n N_Y_c_724_n N_Y_c_741_n N_Y_c_725_n
+ N_Y_c_743_n N_Y_c_744_n N_Y_c_745_n N_Y_c_746_n N_Y_c_859_n N_Y_c_861_n
+ N_Y_c_747_n N_Y_c_867_n N_Y_c_869_n N_Y_c_871_n N_Y_c_748_n N_Y_c_749_n
+ N_Y_c_750_n Y Y PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%Y
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%VGND N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_M1011_d N_VGND_M1017_d N_VGND_M1021_d N_VGND_M1024_d N_VGND_M1032_d
+ N_VGND_M1035_d N_VGND_M1037_d N_VGND_c_1072_n N_VGND_c_1073_n N_VGND_c_1074_n
+ N_VGND_c_1075_n N_VGND_c_1076_n N_VGND_c_1077_n N_VGND_c_1078_n
+ N_VGND_c_1079_n N_VGND_c_1080_n N_VGND_c_1081_n N_VGND_c_1082_n
+ N_VGND_c_1083_n N_VGND_c_1084_n N_VGND_c_1085_n N_VGND_c_1086_n
+ N_VGND_c_1087_n N_VGND_c_1088_n N_VGND_c_1089_n N_VGND_c_1090_n
+ N_VGND_c_1091_n N_VGND_c_1092_n N_VGND_c_1093_n N_VGND_c_1094_n
+ N_VGND_c_1095_n N_VGND_c_1096_n N_VGND_c_1097_n VGND N_VGND_c_1098_n
+ N_VGND_c_1099_n N_VGND_c_1100_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%VPWR VPWR N_VPWR_c_1194_n
+ N_VPWR_c_1193_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16%VPWR
cc_1 VNB N_A_M1004_g 0.0383659f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=0.445
cc_2 VNB N_A_M1007_g 0.0275203f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=0.445
cc_3 VNB N_A_M1008_g 0.0275198f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=0.445
cc_4 VNB N_A_M1011_g 0.0275203f $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=0.445
cc_5 VNB N_A_M1016_g 0.0275198f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.445
cc_6 VNB N_A_M1017_g 0.028174f $X=-0.19 $Y=-0.24 $X2=4.355 $Y2=0.445
cc_7 VNB N_A_M1018_g 0.0306683f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=0.445
cc_8 VNB N_A_c_125_n 0.0217642f $X=-0.19 $Y=-0.24 $X2=5.33 $Y2=1.17
cc_9 VNB N_A_c_126_n 0.226899f $X=-0.19 $Y=-0.24 $X2=4.895 $Y2=1.17
cc_10 VNB N_A_M1021_g 0.0300266f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=0.445
cc_11 VNB N_A_M1023_g 0.0275268f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=0.445
cc_12 VNB N_A_M1024_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=6.265 $Y2=0.445
cc_13 VNB N_A_M1026_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=0.445
cc_14 VNB N_A_M1032_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=7.125 $Y2=0.445
cc_15 VNB N_A_M1033_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=7.555 $Y2=0.445
cc_16 VNB N_A_M1035_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=0.445
cc_17 VNB N_A_M1036_g 0.0275204f $X=-0.19 $Y=-0.24 $X2=8.415 $Y2=0.445
cc_18 VNB N_A_M1037_g 0.037667f $X=-0.19 $Y=-0.24 $X2=8.845 $Y2=0.445
cc_19 VNB A 0.0766144f $X=-0.19 $Y=-0.24 $X2=1.985 $Y2=1.105
cc_20 VNB N_A_c_137_n 0.0775076f $X=-0.19 $Y=-0.24 $X2=10.46 $Y2=1.16
cc_21 VNB N_A_c_138_n 0.259413f $X=-0.19 $Y=-0.24 $X2=10.565 $Y2=1.17
cc_22 VNB N_Y_c_718_n 0.00675515f $X=-0.19 $Y=-0.24 $X2=5.33 $Y2=1.17
cc_23 VNB N_Y_c_719_n 0.00687652f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=1.985
cc_24 VNB N_Y_c_720_n 0.00689469f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=1.985
cc_25 VNB N_Y_c_721_n 0.00770315f $X=-0.19 $Y=-0.24 $X2=6.265 $Y2=1.985
cc_26 VNB N_Y_c_722_n 0.00700409f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=1.35
cc_27 VNB N_Y_c_723_n 0.00687169f $X=-0.19 $Y=-0.24 $X2=7.125 $Y2=1.35
cc_28 VNB N_Y_c_724_n 0.00687169f $X=-0.19 $Y=-0.24 $X2=7.555 $Y2=1.35
cc_29 VNB N_Y_c_725_n 0.00696467f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=1.35
cc_30 VNB N_VGND_c_1072_n 0.01839f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=1.985
cc_31 VNB N_VGND_c_1073_n 0.00402504f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=0.445
cc_32 VNB N_VGND_c_1074_n 0.00405516f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=1.985
cc_33 VNB N_VGND_c_1075_n 0.00466861f $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=0.445
cc_34 VNB N_VGND_c_1076_n 0.00463719f $X=-0.19 $Y=-0.24 $X2=3.495 $Y2=1.985
cc_35 VNB N_VGND_c_1077_n 0.00385357f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.445
cc_36 VNB N_VGND_c_1078_n 0.00407253f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=1.985
cc_37 VNB N_VGND_c_1079_n 0.00402504f $X=-0.19 $Y=-0.24 $X2=4.355 $Y2=0.445
cc_38 VNB N_VGND_c_1080_n 0.0165974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_1081_n 0.0183325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_1082_n 0.0611731f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=0.445
cc_41 VNB N_VGND_c_1083_n 0.00516809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_1084_n 0.0168213f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=1.985
cc_43 VNB N_VGND_c_1085_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=4.82 $Y2=1.985
cc_44 VNB N_VGND_c_1086_n 0.0165526f $X=-0.19 $Y=-0.24 $X2=5.33 $Y2=1.17
cc_45 VNB N_VGND_c_1087_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=4.895 $Y2=1.17
cc_46 VNB N_VGND_c_1088_n 0.0174825f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=0.445
cc_47 VNB N_VGND_c_1089_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=0.445
cc_48 VNB N_VGND_c_1090_n 0.0210033f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=1.35
cc_49 VNB N_VGND_c_1091_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=5.405 $Y2=1.985
cc_50 VNB N_VGND_c_1092_n 0.0165974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1093_n 0.00430243f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=0.99
cc_52 VNB N_VGND_c_1094_n 0.0179215f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=0.445
cc_53 VNB N_VGND_c_1095_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1096_n 0.0165974f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=1.35
cc_55 VNB N_VGND_c_1097_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=5.835 $Y2=1.985
cc_56 VNB N_VGND_c_1098_n 0.0608549f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=0.445
cc_57 VNB N_VGND_c_1099_n 0.649101f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=0.445
cc_58 VNB N_VGND_c_1100_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=7.985 $Y2=1.985
cc_59 VNB N_VPWR_c_1193_n 0.459507f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.35
cc_60 VPB N_A_M1000_g 0.0240838f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_61 VPB N_A_M1001_g 0.0171919f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.985
cc_62 VPB N_A_M1002_g 0.0171919f $X=-0.19 $Y=1.305 $X2=1.345 $Y2=1.985
cc_63 VPB N_A_M1003_g 0.0171696f $X=-0.19 $Y=1.305 $X2=1.775 $Y2=1.985
cc_64 VPB N_A_M1005_g 0.0171412f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=1.985
cc_65 VPB N_A_M1006_g 0.0167979f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=1.985
cc_66 VPB N_A_M1009_g 0.0167978f $X=-0.19 $Y=1.305 $X2=3.065 $Y2=1.985
cc_67 VPB N_A_M1010_g 0.0167979f $X=-0.19 $Y=1.305 $X2=3.495 $Y2=1.985
cc_68 VPB N_A_M1012_g 0.0167978f $X=-0.19 $Y=1.305 $X2=3.925 $Y2=1.985
cc_69 VPB N_A_M1013_g 0.0171663f $X=-0.19 $Y=1.305 $X2=4.355 $Y2=1.985
cc_70 VPB N_A_M1014_g 0.0185867f $X=-0.19 $Y=1.305 $X2=4.82 $Y2=1.985
cc_71 VPB N_A_c_125_n 0.00935665f $X=-0.19 $Y=1.305 $X2=5.33 $Y2=1.17
cc_72 VPB N_A_c_126_n 0.049742f $X=-0.19 $Y=1.305 $X2=4.895 $Y2=1.17
cc_73 VPB N_A_M1015_g 0.0182207f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=1.985
cc_74 VPB N_A_M1019_g 0.0167992f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=1.985
cc_75 VPB N_A_M1020_g 0.016798f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=1.985
cc_76 VPB N_A_M1022_g 0.016798f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=1.985
cc_77 VPB N_A_M1025_g 0.016798f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=1.985
cc_78 VPB N_A_M1027_g 0.016798f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=1.985
cc_79 VPB N_A_M1028_g 0.016798f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=1.985
cc_80 VPB N_A_M1029_g 0.016798f $X=-0.19 $Y=1.305 $X2=8.415 $Y2=1.985
cc_81 VPB N_A_M1030_g 0.0171405f $X=-0.19 $Y=1.305 $X2=8.845 $Y2=1.985
cc_82 VPB N_A_M1031_g 0.0171685f $X=-0.19 $Y=1.305 $X2=9.275 $Y2=1.985
cc_83 VPB N_A_M1034_g 0.0171919f $X=-0.19 $Y=1.305 $X2=9.705 $Y2=1.985
cc_84 VPB N_A_M1038_g 0.0171919f $X=-0.19 $Y=1.305 $X2=10.135 $Y2=1.985
cc_85 VPB N_A_M1039_g 0.0240835f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.985
cc_86 VPB N_A_c_138_n 0.0580561f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.17
cc_87 VPB N_KAPWR_c_473_n 0.0116666f $X=-0.19 $Y=1.305 $X2=4.355 $Y2=1.985
cc_88 VPB N_KAPWR_c_474_n 0.0318208f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=0.445
cc_89 VPB N_KAPWR_c_475_n 0.0195476f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=1.17
cc_90 VPB N_KAPWR_c_476_n 0.0121012f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=1.17
cc_91 VPB N_Y_c_726_n 0.0016373f $X=-0.19 $Y=1.305 $X2=4.355 $Y2=1.35
cc_92 VPB N_Y_c_727_n 0.00328873f $X=-0.19 $Y=1.305 $X2=4.82 $Y2=0.99
cc_93 VPB N_Y_c_728_n 0.00275521f $X=-0.19 $Y=1.305 $X2=4.82 $Y2=1.35
cc_94 VPB N_Y_c_718_n 0.00112034f $X=-0.19 $Y=1.305 $X2=5.33 $Y2=1.17
cc_95 VPB N_Y_c_730_n 0.00261217f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=0.445
cc_96 VPB N_Y_c_719_n 0.00104035f $X=-0.19 $Y=1.305 $X2=5.405 $Y2=1.985
cc_97 VPB N_Y_c_732_n 0.00261217f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=0.445
cc_98 VPB N_Y_c_720_n 0.0010602f $X=-0.19 $Y=1.305 $X2=5.835 $Y2=1.985
cc_99 VPB N_Y_c_734_n 0.00283159f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=0.445
cc_100 VPB N_Y_c_721_n 0.00109244f $X=-0.19 $Y=1.305 $X2=6.265 $Y2=1.985
cc_101 VPB N_Y_c_722_n 0.00107025f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=1.35
cc_102 VPB N_Y_c_737_n 0.00266908f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=0.99
cc_103 VPB N_Y_c_723_n 0.00104488f $X=-0.19 $Y=1.305 $X2=7.125 $Y2=1.35
cc_104 VPB N_Y_c_739_n 0.00266908f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=0.99
cc_105 VPB N_Y_c_724_n 0.00104488f $X=-0.19 $Y=1.305 $X2=7.555 $Y2=1.35
cc_106 VPB N_Y_c_741_n 0.00266908f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=0.99
cc_107 VPB N_Y_c_725_n 0.00112789f $X=-0.19 $Y=1.305 $X2=7.985 $Y2=1.35
cc_108 VPB N_Y_c_743_n 0.00248501f $X=-0.19 $Y=1.305 $X2=8.415 $Y2=0.99
cc_109 VPB N_Y_c_744_n 0.00279943f $X=-0.19 $Y=1.305 $X2=8.415 $Y2=1.35
cc_110 VPB N_Y_c_745_n 0.00102678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_Y_c_746_n 4.29584e-19 $X=-0.19 $Y=1.305 $X2=8.845 $Y2=1.985
cc_112 VPB N_Y_c_747_n 0.00335197f $X=-0.19 $Y=1.305 $X2=9.275 $Y2=1.985
cc_113 VPB N_Y_c_748_n 4.27809e-19 $X=-0.19 $Y=1.305 $X2=10.135 $Y2=1.985
cc_114 VPB N_Y_c_749_n 0.00102678f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.35
cc_115 VPB N_Y_c_750_n 0.0021101f $X=-0.19 $Y=1.305 $X2=10.565 $Y2=1.985
cc_116 VPB N_VPWR_c_1194_n 0.293856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_1193_n 0.0436453f $X=-0.19 $Y=1.305 $X2=1.345 $Y2=1.35
cc_118 N_A_M1038_g N_KAPWR_c_473_n 0.00240782f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1039_g N_KAPWR_c_473_n 0.00580645f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_M1000_g N_KAPWR_c_479_n 0.00580645f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_M1001_g N_KAPWR_c_479_n 0.00169511f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_M1001_g N_KAPWR_c_481_n 0.00113476f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_M1002_g N_KAPWR_c_482_n 0.00238856f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_M1003_g N_KAPWR_c_482_n 0.00240782f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_M1005_g N_KAPWR_c_484_n 0.00240782f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_M1006_g N_KAPWR_c_484_n 0.00240782f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_M1010_g N_KAPWR_c_486_n 0.0064105f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_M1012_g N_KAPWR_c_486_n 0.0062148f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1009_g N_KAPWR_c_488_n 0.00240782f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_M1010_g N_KAPWR_c_488_n 0.00238856f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_M1012_g N_KAPWR_c_490_n 0.0013166f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_M1013_g N_KAPWR_c_491_n 0.00527887f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1014_g N_KAPWR_c_491_n 0.00723471f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1012_g N_KAPWR_c_493_n 0.00150248f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1013_g N_KAPWR_c_493_n 0.00277381f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1014_g N_KAPWR_c_495_n 0.00104387f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1014_g N_KAPWR_c_496_n 0.00431712f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1015_g N_KAPWR_c_496_n 0.00111723f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1015_g N_KAPWR_c_498_n 0.00159783f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1019_g N_KAPWR_c_499_n 0.00248487f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1020_g N_KAPWR_c_499_n 0.00227298f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1020_g N_KAPWR_c_501_n 6.09479e-19 $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1022_g N_KAPWR_c_502_n 0.00240782f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1025_g N_KAPWR_c_502_n 0.00227298f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1025_g N_KAPWR_c_504_n 6.09479e-19 $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1027_g N_KAPWR_c_505_n 0.00240782f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1028_g N_KAPWR_c_505_n 0.00240782f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1029_g N_KAPWR_c_507_n 0.00240782f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1030_g N_KAPWR_c_507_n 0.00240782f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1031_g N_KAPWR_c_509_n 0.00240782f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1034_g N_KAPWR_c_509_n 0.00240782f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1000_g N_KAPWR_c_474_n 0.0102684f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_153 A N_KAPWR_c_474_n 0.0044789f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A_M1001_g N_KAPWR_c_513_n 0.00621593f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_KAPWR_c_513_n 0.00641148f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1003_g N_KAPWR_c_515_n 0.00636143f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1005_g N_KAPWR_c_515_n 0.00637716f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_M1006_g N_KAPWR_c_517_n 0.00637772f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1009_g N_KAPWR_c_517_n 0.00636195f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1015_g N_KAPWR_c_519_n 0.00688381f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_M1019_g N_KAPWR_c_519_n 0.00615138f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_M1020_g N_KAPWR_c_521_n 0.00616537f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_M1022_g N_KAPWR_c_521_n 0.00637711f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1025_g N_KAPWR_c_523_n 0.00618171f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_M1027_g N_KAPWR_c_523_n 0.00637772f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_M1028_g N_KAPWR_c_525_n 0.00637785f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_M1029_g N_KAPWR_c_525_n 0.00637728f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_M1030_g N_KAPWR_c_527_n 0.00637728f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_M1031_g N_KAPWR_c_527_n 0.00637728f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_M1034_g N_KAPWR_c_529_n 0.0063773f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_M1038_g N_KAPWR_c_529_n 0.00637893f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_M1039_g N_KAPWR_c_475_n 0.0070151f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_c_137_n N_KAPWR_c_475_n 0.0023947f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_M1000_g N_Y_c_726_n 9.2188e-19 $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_c_126_n N_Y_c_726_n 0.00258307f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_176 A N_Y_c_726_n 0.0138667f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_177 N_A_M1001_g N_Y_c_727_n 0.0108326f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_M1002_g N_Y_c_727_n 0.0109021f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_c_126_n N_Y_c_727_n 0.00249109f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_180 A N_Y_c_727_n 0.0496576f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A_c_229_p N_Y_c_727_n 2.42369e-19 $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_182 N_A_M1003_g N_Y_c_728_n 0.0108201f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1005_g N_Y_c_728_n 0.0111822f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_c_126_n N_Y_c_728_n 0.00249109f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_185 A N_Y_c_728_n 0.030024f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A_c_229_p N_Y_c_728_n 0.0149363f $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_187 N_A_c_235_p N_Y_c_728_n 0.00428581f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_188 N_A_M1004_g N_Y_c_718_n 0.00687088f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_M1005_g N_Y_c_718_n 0.00163185f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_M1007_g N_Y_c_718_n 0.00479472f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A_M1006_g N_Y_c_718_n 9.05456e-19 $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_c_126_n N_Y_c_718_n 0.026551f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_193 A N_Y_c_718_n 0.0270465f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_194 N_A_c_235_p N_Y_c_718_n 0.0315188f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_195 N_A_c_243_p N_Y_c_718_n 0.00339471f $X=2.215 $Y=1.19 $X2=0 $Y2=0
cc_196 N_A_M1006_g N_Y_c_730_n 0.0127237f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_M1009_g N_Y_c_730_n 0.0128168f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_c_126_n N_Y_c_730_n 0.00443815f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_199 N_A_c_235_p N_Y_c_730_n 0.0255685f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_200 N_A_M1008_g N_Y_c_719_n 0.00483858f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_201 N_A_M1009_g N_Y_c_719_n 9.14001e-19 $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_M1011_g N_Y_c_719_n 0.00488763f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A_M1010_g N_Y_c_719_n 9.2326e-19 $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_c_126_n N_Y_c_719_n 0.0306427f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_205 N_A_c_235_p N_Y_c_719_n 0.0369292f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_206 N_A_M1010_g N_Y_c_732_n 0.0128203f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_M1012_g N_Y_c_732_n 0.0127594f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_c_126_n N_Y_c_732_n 0.00443815f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_209 N_A_c_235_p N_Y_c_732_n 0.0255685f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_210 N_A_M1016_g N_Y_c_720_n 0.0047937f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A_M1012_g N_Y_c_720_n 9.05401e-19 $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_M1017_g N_Y_c_720_n 0.00486847f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A_M1013_g N_Y_c_720_n 9.20002e-19 $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_c_126_n N_Y_c_720_n 0.0304611f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_215 N_A_c_235_p N_Y_c_720_n 0.0352566f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_216 N_A_M1013_g N_Y_c_734_n 0.013299f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_M1014_g N_Y_c_734_n 0.0165644f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_c_126_n N_Y_c_734_n 0.0059915f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_219 N_A_c_235_p N_Y_c_734_n 0.027541f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_220 N_A_M1018_g N_Y_c_721_n 0.00605274f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_221 N_A_M1014_g N_Y_c_721_n 0.00114052f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A_c_125_n N_Y_c_721_n 0.0417629f $X=5.33 $Y=1.17 $X2=0 $Y2=0
cc_223 N_A_M1021_g N_Y_c_721_n 0.00937526f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_224 N_A_M1015_g N_Y_c_721_n 0.0010184f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_c_235_p N_Y_c_721_n 0.0483297f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_226 N_A_M1023_g N_Y_c_722_n 0.00507366f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_M1019_g N_Y_c_722_n 9.59045e-19 $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_M1024_g N_Y_c_722_n 0.00484361f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_M1020_g N_Y_c_722_n 9.14964e-19 $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_c_235_p N_Y_c_722_n 0.0364786f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_231 N_A_c_138_n N_Y_c_722_n 0.0309751f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_232 N_A_M1020_g N_Y_c_737_n 0.012819f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A_M1022_g N_Y_c_737_n 0.0128281f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_c_235_p N_Y_c_737_n 0.0257897f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_235 N_A_c_138_n N_Y_c_737_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_236 N_A_M1026_g N_Y_c_723_n 0.00484361f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A_M1022_g N_Y_c_723_n 9.14964e-19 $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A_M1032_g N_Y_c_723_n 0.00484361f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A_M1025_g N_Y_c_723_n 9.14964e-19 $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_c_235_p N_Y_c_723_n 0.0363628f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_241 N_A_c_138_n N_Y_c_723_n 0.0305483f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_242 N_A_M1025_g N_Y_c_739_n 0.012819f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_M1027_g N_Y_c_739_n 0.0128281f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_c_235_p N_Y_c_739_n 0.0257897f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_245 N_A_c_138_n N_Y_c_739_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_246 N_A_M1033_g N_Y_c_724_n 0.00484361f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_247 N_A_M1027_g N_Y_c_724_n 9.14964e-19 $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_M1035_g N_Y_c_724_n 0.00484361f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_249 N_A_M1028_g N_Y_c_724_n 9.14964e-19 $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_c_235_p N_Y_c_724_n 0.0363628f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_251 N_A_c_138_n N_Y_c_724_n 0.0305483f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_252 N_A_M1028_g N_Y_c_741_n 0.0128173f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_M1029_g N_Y_c_741_n 0.012689f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A_c_235_p N_Y_c_741_n 0.0257897f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_255 N_A_c_138_n N_Y_c_741_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_256 N_A_M1036_g N_Y_c_725_n 0.00484361f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_257 N_A_M1029_g N_Y_c_725_n 9.14964e-19 $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_M1037_g N_Y_c_725_n 0.00730344f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_M1030_g N_Y_c_725_n 0.00172986f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_c_235_p N_Y_c_725_n 0.0345046f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_261 N_A_c_309_p N_Y_c_725_n 0.00117738f $X=9.4 $Y=1.19 $X2=0 $Y2=0
cc_262 N_A_c_137_n N_Y_c_725_n 0.0277667f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_c_138_n N_Y_c_725_n 0.0278283f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_264 N_A_M1030_g N_Y_c_743_n 0.0112371f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_M1031_g N_Y_c_743_n 0.0108839f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_c_235_p N_Y_c_743_n 0.00932131f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_267 N_A_c_309_p N_Y_c_743_n 0.0028903f $X=9.4 $Y=1.19 $X2=0 $Y2=0
cc_268 N_A_c_137_n N_Y_c_743_n 0.0303464f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_c_138_n N_Y_c_743_n 0.00249109f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_270 N_A_M1034_g N_Y_c_744_n 0.0107624f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_M1038_g N_Y_c_744_n 0.01091f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_c_320_p N_Y_c_744_n 0.0112216f $X=9.89 $Y=1.19 $X2=0 $Y2=0
cc_273 N_A_c_137_n N_Y_c_744_n 0.0434858f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_c_138_n N_Y_c_744_n 0.00249109f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_275 N_A_M1002_g N_Y_c_745_n 0.00140497f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_M1003_g N_Y_c_745_n 0.00140623f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_c_126_n N_Y_c_745_n 0.00258307f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_278 A N_Y_c_745_n 0.0112313f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_279 N_A_c_229_p N_Y_c_745_n 0.00432607f $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_280 N_A_M1005_g N_Y_c_746_n 0.00268766f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_M1006_g N_Y_c_746_n 0.00140623f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A_M1009_g N_Y_c_859_n 0.00140623f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A_M1010_g N_Y_c_859_n 0.00140497f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_M1012_g N_Y_c_861_n 0.00140497f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A_M1013_g N_Y_c_861_n 0.00142997f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A_M1015_g N_Y_c_747_n 0.0130118f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A_M1019_g N_Y_c_747_n 0.012864f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A_c_235_p N_Y_c_747_n 0.0284261f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_289 N_A_c_138_n N_Y_c_747_n 0.00443815f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_290 N_A_M1019_g N_Y_c_867_n 0.00141126f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_M1020_g N_Y_c_867_n 0.00140623f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A_M1022_g N_Y_c_869_n 0.00140623f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_293 N_A_M1025_g N_Y_c_869_n 0.00140623f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A_M1027_g N_Y_c_871_n 0.00140623f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A_M1028_g N_Y_c_871_n 0.00140623f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A_M1029_g N_Y_c_748_n 0.00140623f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A_M1030_g N_Y_c_748_n 0.00273624f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A_M1031_g N_Y_c_749_n 0.00140623f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_M1034_g N_Y_c_749_n 0.00140623f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A_c_320_p N_Y_c_749_n 0.00432607f $X=9.89 $Y=1.19 $X2=0 $Y2=0
cc_301 N_A_c_137_n N_Y_c_749_n 0.0112313f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_c_138_n N_Y_c_749_n 0.00258307f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_303 N_A_M1038_g N_Y_c_750_n 0.00140623f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A_M1039_g N_Y_c_750_n 0.00237484f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A_c_137_n N_Y_c_750_n 0.0172117f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_c_138_n N_Y_c_750_n 0.00258307f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_307 N_A_M1014_g Y 0.00874672f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_M1015_g Y 0.00668472f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_M1004_g N_VGND_c_1072_n 0.00372544f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_310 N_A_c_126_n N_VGND_c_1072_n 0.00146648f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_311 A N_VGND_c_1072_n 0.0131993f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A_c_229_p N_VGND_c_1072_n 0.00160784f $X=2.1 $Y=1.19 $X2=0 $Y2=0
cc_313 N_A_M1007_g N_VGND_c_1073_n 0.00167629f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_314 N_A_M1008_g N_VGND_c_1073_n 0.00169877f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_315 N_A_c_126_n N_VGND_c_1073_n 0.00357354f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_316 N_A_c_235_p N_VGND_c_1073_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_317 N_A_M1011_g N_VGND_c_1074_n 0.00167629f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_318 N_A_M1016_g N_VGND_c_1074_n 0.00173246f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_319 N_A_c_126_n N_VGND_c_1074_n 0.00357354f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_320 N_A_c_235_p N_VGND_c_1074_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_321 N_A_M1017_g N_VGND_c_1075_n 0.00166077f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_322 N_A_M1018_g N_VGND_c_1075_n 0.00315583f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_323 N_A_c_126_n N_VGND_c_1075_n 0.00482428f $X=4.895 $Y=1.17 $X2=0 $Y2=0
cc_324 N_A_c_235_p N_VGND_c_1075_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_325 N_A_M1021_g N_VGND_c_1076_n 0.00312236f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_326 N_A_M1023_g N_VGND_c_1076_n 0.00169877f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_327 N_A_c_235_p N_VGND_c_1076_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_328 N_A_c_138_n N_VGND_c_1076_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_329 N_A_M1024_g N_VGND_c_1077_n 0.00165467f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_330 N_A_M1026_g N_VGND_c_1077_n 0.0015561f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_331 N_A_c_235_p N_VGND_c_1077_n 0.00775425f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_332 N_A_c_138_n N_VGND_c_1077_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_333 N_A_M1032_g N_VGND_c_1078_n 0.00172922f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_334 N_A_M1033_g N_VGND_c_1078_n 0.00169877f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_335 N_A_c_235_p N_VGND_c_1078_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_336 N_A_c_138_n N_VGND_c_1078_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_337 N_A_M1035_g N_VGND_c_1079_n 0.00167629f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_338 N_A_M1036_g N_VGND_c_1079_n 0.00169877f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_339 N_A_c_235_p N_VGND_c_1079_n 0.00914515f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_340 N_A_c_138_n N_VGND_c_1079_n 0.00357354f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_341 N_A_M1036_g N_VGND_c_1080_n 0.00585385f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_342 N_A_M1037_g N_VGND_c_1080_n 0.00585385f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_343 N_A_M1037_g N_VGND_c_1081_n 0.00368624f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_344 N_A_c_235_p N_VGND_c_1081_n 0.00148989f $X=9.285 $Y=1.19 $X2=0 $Y2=0
cc_345 N_A_c_137_n N_VGND_c_1081_n 0.0131863f $X=10.46 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A_c_138_n N_VGND_c_1081_n 0.00145246f $X=10.565 $Y=1.17 $X2=0 $Y2=0
cc_347 N_A_M1004_g N_VGND_c_1084_n 0.00585385f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_348 N_A_M1007_g N_VGND_c_1084_n 0.00585385f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_349 N_A_M1008_g N_VGND_c_1086_n 0.00585385f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_350 N_A_M1011_g N_VGND_c_1086_n 0.00585385f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_351 N_A_M1016_g N_VGND_c_1088_n 0.00585385f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_352 N_A_M1017_g N_VGND_c_1088_n 0.00585385f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_353 N_A_M1018_g N_VGND_c_1090_n 0.00585385f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_354 N_A_M1021_g N_VGND_c_1090_n 0.00585385f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_355 N_A_M1023_g N_VGND_c_1092_n 0.00585385f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_356 N_A_M1024_g N_VGND_c_1092_n 0.00585385f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_357 N_A_M1026_g N_VGND_c_1094_n 0.00585385f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_358 N_A_M1032_g N_VGND_c_1094_n 0.00585385f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_359 N_A_M1033_g N_VGND_c_1096_n 0.00585385f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_360 N_A_M1035_g N_VGND_c_1096_n 0.00585385f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_361 N_A_M1004_g N_VGND_c_1099_n 0.0119802f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_362 N_A_M1007_g N_VGND_c_1099_n 0.010643f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_363 N_A_M1008_g N_VGND_c_1099_n 0.0106305f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_364 N_A_M1011_g N_VGND_c_1099_n 0.010643f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_365 N_A_M1016_g N_VGND_c_1099_n 0.0106305f $X=3.925 $Y=0.445 $X2=0 $Y2=0
cc_366 N_A_M1017_g N_VGND_c_1099_n 0.0107976f $X=4.355 $Y=0.445 $X2=0 $Y2=0
cc_367 N_A_M1018_g N_VGND_c_1099_n 0.0111111f $X=4.82 $Y=0.445 $X2=0 $Y2=0
cc_368 N_A_M1021_g N_VGND_c_1099_n 0.0110068f $X=5.405 $Y=0.445 $X2=0 $Y2=0
cc_369 N_A_M1023_g N_VGND_c_1099_n 0.0106305f $X=5.835 $Y=0.445 $X2=0 $Y2=0
cc_370 N_A_M1024_g N_VGND_c_1099_n 0.010643f $X=6.265 $Y=0.445 $X2=0 $Y2=0
cc_371 N_A_M1026_g N_VGND_c_1099_n 0.0107309f $X=6.695 $Y=0.445 $X2=0 $Y2=0
cc_372 N_A_M1032_g N_VGND_c_1099_n 0.010643f $X=7.125 $Y=0.445 $X2=0 $Y2=0
cc_373 N_A_M1033_g N_VGND_c_1099_n 0.0106305f $X=7.555 $Y=0.445 $X2=0 $Y2=0
cc_374 N_A_M1035_g N_VGND_c_1099_n 0.010643f $X=7.985 $Y=0.445 $X2=0 $Y2=0
cc_375 N_A_M1036_g N_VGND_c_1099_n 0.0106305f $X=8.415 $Y=0.445 $X2=0 $Y2=0
cc_376 N_A_M1037_g N_VGND_c_1099_n 0.0119927f $X=8.845 $Y=0.445 $X2=0 $Y2=0
cc_377 N_A_M1000_g N_VPWR_c_1194_n 0.00541359f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_378 N_A_M1001_g N_VPWR_c_1194_n 0.00547467f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A_M1002_g N_VPWR_c_1194_n 0.00547467f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A_M1003_g N_VPWR_c_1194_n 0.0054895f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A_M1005_g N_VPWR_c_1194_n 0.0054895f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_382 N_A_M1006_g N_VPWR_c_1194_n 0.0054895f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_383 N_A_M1009_g N_VPWR_c_1194_n 0.0054895f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_384 N_A_M1010_g N_VPWR_c_1194_n 0.00547467f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_385 N_A_M1012_g N_VPWR_c_1194_n 0.00547467f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_386 N_A_M1013_g N_VPWR_c_1194_n 0.00577801f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_387 N_A_M1014_g N_VPWR_c_1194_n 0.00570217f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_388 N_A_M1015_g N_VPWR_c_1194_n 0.00539883f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_389 N_A_M1019_g N_VPWR_c_1194_n 0.0055505f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_390 N_A_M1020_g N_VPWR_c_1194_n 0.0054895f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A_M1022_g N_VPWR_c_1194_n 0.0054895f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A_M1025_g N_VPWR_c_1194_n 0.0054895f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A_M1027_g N_VPWR_c_1194_n 0.0054895f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A_M1028_g N_VPWR_c_1194_n 0.0054895f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_395 N_A_M1029_g N_VPWR_c_1194_n 0.0054895f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_396 N_A_M1030_g N_VPWR_c_1194_n 0.0054895f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A_M1031_g N_VPWR_c_1194_n 0.0054895f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_398 N_A_M1034_g N_VPWR_c_1194_n 0.0054895f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_399 N_A_M1038_g N_VPWR_c_1194_n 0.0054895f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A_M1039_g N_VPWR_c_1194_n 0.00541359f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A_M1000_g N_VPWR_c_1193_n 0.00604751f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A_M1001_g N_VPWR_c_1193_n 0.00512084f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_403 N_A_M1002_g N_VPWR_c_1193_n 0.00515166f $X=1.345 $Y=1.985 $X2=0 $Y2=0
cc_404 N_A_M1003_g N_VPWR_c_1193_n 0.00515546f $X=1.775 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A_M1005_g N_VPWR_c_1193_n 0.00515546f $X=2.205 $Y=1.985 $X2=0 $Y2=0
cc_406 N_A_M1006_g N_VPWR_c_1193_n 0.00515546f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_407 N_A_M1009_g N_VPWR_c_1193_n 0.00515546f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A_M1010_g N_VPWR_c_1193_n 0.00515166f $X=3.495 $Y=1.985 $X2=0 $Y2=0
cc_409 N_A_M1012_g N_VPWR_c_1193_n 0.00515166f $X=3.925 $Y=1.985 $X2=0 $Y2=0
cc_410 N_A_M1013_g N_VPWR_c_1193_n 0.00529604f $X=4.355 $Y=1.985 $X2=0 $Y2=0
cc_411 N_A_M1014_g N_VPWR_c_1193_n 0.00566991f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_412 N_A_M1015_g N_VPWR_c_1193_n 0.0054963f $X=5.405 $Y=1.985 $X2=0 $Y2=0
cc_413 N_A_M1019_g N_VPWR_c_1193_n 0.00517073f $X=5.835 $Y=1.985 $X2=0 $Y2=0
cc_414 N_A_M1020_g N_VPWR_c_1193_n 0.00515546f $X=6.265 $Y=1.985 $X2=0 $Y2=0
cc_415 N_A_M1022_g N_VPWR_c_1193_n 0.00515546f $X=6.695 $Y=1.985 $X2=0 $Y2=0
cc_416 N_A_M1025_g N_VPWR_c_1193_n 0.00515546f $X=7.125 $Y=1.985 $X2=0 $Y2=0
cc_417 N_A_M1027_g N_VPWR_c_1193_n 0.00515546f $X=7.555 $Y=1.985 $X2=0 $Y2=0
cc_418 N_A_M1028_g N_VPWR_c_1193_n 0.00515546f $X=7.985 $Y=1.985 $X2=0 $Y2=0
cc_419 N_A_M1029_g N_VPWR_c_1193_n 0.00515546f $X=8.415 $Y=1.985 $X2=0 $Y2=0
cc_420 N_A_M1030_g N_VPWR_c_1193_n 0.00515546f $X=8.845 $Y=1.985 $X2=0 $Y2=0
cc_421 N_A_M1031_g N_VPWR_c_1193_n 0.00515546f $X=9.275 $Y=1.985 $X2=0 $Y2=0
cc_422 N_A_M1034_g N_VPWR_c_1193_n 0.00515546f $X=9.705 $Y=1.985 $X2=0 $Y2=0
cc_423 N_A_M1038_g N_VPWR_c_1193_n 0.00515546f $X=10.135 $Y=1.985 $X2=0 $Y2=0
cc_424 N_A_M1039_g N_VPWR_c_1193_n 0.006069f $X=10.565 $Y=1.985 $X2=0 $Y2=0
cc_425 N_KAPWR_c_479_n N_Y_M1000_s 0.00322826f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_426 N_KAPWR_c_482_n N_Y_M1002_s 0.00177005f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_427 N_KAPWR_c_484_n N_Y_M1005_s 0.00176933f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_428 N_KAPWR_c_488_n N_Y_M1009_s 0.00176892f $X=3.63 $Y=2.21 $X2=0 $Y2=0
cc_429 N_KAPWR_c_493_n N_Y_M1012_s 0.00176912f $X=4.49 $Y=2.21 $X2=0 $Y2=0
cc_430 N_KAPWR_c_496_n N_Y_M1014_s 0.00441571f $X=5.39 $Y=2.21 $X2=0 $Y2=0
cc_431 N_KAPWR_c_499_n N_Y_M1019_s 0.00176899f $X=6.31 $Y=2.21 $X2=0 $Y2=0
cc_432 N_KAPWR_c_502_n N_Y_M1022_s 0.00176899f $X=7.17 $Y=2.21 $X2=0 $Y2=0
cc_433 N_KAPWR_c_505_n N_Y_M1027_s 0.00176899f $X=8.07 $Y=2.21 $X2=0 $Y2=0
cc_434 N_KAPWR_c_507_n N_Y_M1029_s 0.00176899f $X=8.9 $Y=2.21 $X2=0 $Y2=0
cc_435 N_KAPWR_c_509_n N_Y_M1031_s 0.00177005f $X=9.76 $Y=2.21 $X2=0 $Y2=0
cc_436 N_KAPWR_c_473_n N_Y_M1038_s 0.00201707f $X=10.66 $Y=2.24 $X2=0 $Y2=0
cc_437 N_KAPWR_c_479_n N_Y_c_898_n 0.018488f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_438 N_KAPWR_c_481_n N_Y_c_898_n 0.00154073f $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_439 N_KAPWR_c_474_n N_Y_c_898_n 0.0315662f $X=0.275 $Y=1.66 $X2=0 $Y2=0
cc_440 N_KAPWR_c_513_n N_Y_c_898_n 0.024621f $X=1.13 $Y=2 $X2=0 $Y2=0
cc_441 N_KAPWR_c_476_n N_Y_c_898_n 3.6717e-19 $X=0.36 $Y=2.21 $X2=0 $Y2=0
cc_442 N_KAPWR_M1001_d N_Y_c_727_n 0.00171895f $X=0.99 $Y=1.485 $X2=0 $Y2=0
cc_443 N_KAPWR_c_479_n N_Y_c_727_n 0.00443585f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_444 N_KAPWR_c_481_n N_Y_c_727_n 0.00223607f $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_445 N_KAPWR_c_482_n N_Y_c_727_n 0.00574928f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_446 N_KAPWR_c_513_n N_Y_c_727_n 0.0165472f $X=1.13 $Y=2 $X2=0 $Y2=0
cc_447 N_KAPWR_M1003_d N_Y_c_728_n 0.00171493f $X=1.85 $Y=1.485 $X2=0 $Y2=0
cc_448 N_KAPWR_c_482_n N_Y_c_728_n 0.00548259f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_449 N_KAPWR_c_557_p N_Y_c_728_n 0.00128894f $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_450 N_KAPWR_c_484_n N_Y_c_728_n 0.00527026f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_451 N_KAPWR_c_515_n N_Y_c_728_n 0.0159201f $X=1.99 $Y=2 $X2=0 $Y2=0
cc_452 N_KAPWR_M1006_d N_Y_c_730_n 0.00172416f $X=2.71 $Y=1.485 $X2=0 $Y2=0
cc_453 N_KAPWR_c_484_n N_Y_c_730_n 0.00405284f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_454 N_KAPWR_c_562_p N_Y_c_730_n 0.00131231f $X=3 $Y=2.21 $X2=0 $Y2=0
cc_455 N_KAPWR_c_488_n N_Y_c_730_n 0.00419718f $X=3.63 $Y=2.21 $X2=0 $Y2=0
cc_456 N_KAPWR_c_517_n N_Y_c_730_n 0.0161977f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_457 N_KAPWR_M1010_d N_Y_c_732_n 0.00169697f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_458 N_KAPWR_c_486_n N_Y_c_732_n 0.0162415f $X=3.775 $Y=2.21 $X2=0 $Y2=0
cc_459 N_KAPWR_c_488_n N_Y_c_732_n 0.00427651f $X=3.63 $Y=2.21 $X2=0 $Y2=0
cc_460 N_KAPWR_c_490_n N_Y_c_732_n 0.00254989f $X=3.92 $Y=2.21 $X2=0 $Y2=0
cc_461 N_KAPWR_c_493_n N_Y_c_732_n 0.00278719f $X=4.49 $Y=2.21 $X2=0 $Y2=0
cc_462 N_KAPWR_M1013_d N_Y_c_734_n 0.00206135f $X=4.43 $Y=1.485 $X2=0 $Y2=0
cc_463 N_KAPWR_c_491_n N_Y_c_734_n 0.0163991f $X=4.635 $Y=2.21 $X2=0 $Y2=0
cc_464 N_KAPWR_c_493_n N_Y_c_734_n 0.005332f $X=4.49 $Y=2.21 $X2=0 $Y2=0
cc_465 N_KAPWR_c_495_n N_Y_c_734_n 0.00200446f $X=4.78 $Y=2.21 $X2=0 $Y2=0
cc_466 N_KAPWR_c_496_n N_Y_c_734_n 0.00369414f $X=5.39 $Y=2.21 $X2=0 $Y2=0
cc_467 N_KAPWR_M1020_d N_Y_c_737_n 0.00172416f $X=6.34 $Y=1.485 $X2=0 $Y2=0
cc_468 N_KAPWR_c_499_n N_Y_c_737_n 0.00395683f $X=6.31 $Y=2.21 $X2=0 $Y2=0
cc_469 N_KAPWR_c_501_n N_Y_c_737_n 0.00147241f $X=6.6 $Y=2.21 $X2=0 $Y2=0
cc_470 N_KAPWR_c_502_n N_Y_c_737_n 0.00431776f $X=7.17 $Y=2.21 $X2=0 $Y2=0
cc_471 N_KAPWR_c_521_n N_Y_c_737_n 0.0161887f $X=6.48 $Y=2 $X2=0 $Y2=0
cc_472 N_KAPWR_M1025_d N_Y_c_739_n 0.00172416f $X=7.2 $Y=1.485 $X2=0 $Y2=0
cc_473 N_KAPWR_c_502_n N_Y_c_739_n 0.00395683f $X=7.17 $Y=2.21 $X2=0 $Y2=0
cc_474 N_KAPWR_c_504_n N_Y_c_739_n 0.00147241f $X=7.46 $Y=2.21 $X2=0 $Y2=0
cc_475 N_KAPWR_c_505_n N_Y_c_739_n 0.00431776f $X=8.07 $Y=2.21 $X2=0 $Y2=0
cc_476 N_KAPWR_c_523_n N_Y_c_739_n 0.0161887f $X=7.34 $Y=2 $X2=0 $Y2=0
cc_477 N_KAPWR_M1028_d N_Y_c_741_n 0.00172416f $X=8.06 $Y=1.485 $X2=0 $Y2=0
cc_478 N_KAPWR_c_505_n N_Y_c_741_n 0.00427637f $X=8.07 $Y=2.21 $X2=0 $Y2=0
cc_479 N_KAPWR_c_587_p N_Y_c_741_n 0.00130852f $X=8.36 $Y=2.21 $X2=0 $Y2=0
cc_480 N_KAPWR_c_507_n N_Y_c_741_n 0.00414655f $X=8.9 $Y=2.21 $X2=0 $Y2=0
cc_481 N_KAPWR_c_525_n N_Y_c_741_n 0.0162022f $X=8.2 $Y=2 $X2=0 $Y2=0
cc_482 N_KAPWR_M1030_d N_Y_c_743_n 0.00171493f $X=8.92 $Y=1.485 $X2=0 $Y2=0
cc_483 N_KAPWR_c_507_n N_Y_c_743_n 0.00406824f $X=8.9 $Y=2.21 $X2=0 $Y2=0
cc_484 N_KAPWR_c_592_p N_Y_c_743_n 0.00128894f $X=9.19 $Y=2.21 $X2=0 $Y2=0
cc_485 N_KAPWR_c_509_n N_Y_c_743_n 0.00561047f $X=9.76 $Y=2.21 $X2=0 $Y2=0
cc_486 N_KAPWR_c_527_n N_Y_c_743_n 0.0160103f $X=9.06 $Y=2 $X2=0 $Y2=0
cc_487 N_KAPWR_M1034_d N_Y_c_744_n 0.00171493f $X=9.78 $Y=1.485 $X2=0 $Y2=0
cc_488 N_KAPWR_c_473_n N_Y_c_744_n 0.00561047f $X=10.66 $Y=2.24 $X2=0 $Y2=0
cc_489 N_KAPWR_c_509_n N_Y_c_744_n 0.00548259f $X=9.76 $Y=2.21 $X2=0 $Y2=0
cc_490 N_KAPWR_c_598_p N_Y_c_744_n 0.00128894f $X=10.05 $Y=2.21 $X2=0 $Y2=0
cc_491 N_KAPWR_c_529_n N_Y_c_744_n 0.0159801f $X=9.92 $Y=2 $X2=0 $Y2=0
cc_492 N_KAPWR_c_481_n N_Y_c_745_n 3.7042e-19 $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_493 N_KAPWR_c_482_n N_Y_c_745_n 0.0185366f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_494 N_KAPWR_c_557_p N_Y_c_745_n 4.44943e-19 $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_495 N_KAPWR_c_513_n N_Y_c_745_n 0.0247795f $X=1.13 $Y=2 $X2=0 $Y2=0
cc_496 N_KAPWR_c_515_n N_Y_c_745_n 0.024745f $X=1.99 $Y=2 $X2=0 $Y2=0
cc_497 N_KAPWR_c_557_p N_Y_c_746_n 4.09742e-19 $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_498 N_KAPWR_c_484_n N_Y_c_746_n 0.0207379f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_499 N_KAPWR_c_562_p N_Y_c_746_n 4.20762e-19 $X=3 $Y=2.21 $X2=0 $Y2=0
cc_500 N_KAPWR_c_515_n N_Y_c_746_n 0.0247213f $X=1.99 $Y=2 $X2=0 $Y2=0
cc_501 N_KAPWR_c_517_n N_Y_c_746_n 0.0247263f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_502 N_KAPWR_c_562_p N_Y_c_859_n 4.32468e-19 $X=3 $Y=2.21 $X2=0 $Y2=0
cc_503 N_KAPWR_c_486_n N_Y_c_859_n 0.0247849f $X=3.775 $Y=2.21 $X2=0 $Y2=0
cc_504 N_KAPWR_c_488_n N_Y_c_859_n 0.0219432f $X=3.63 $Y=2.21 $X2=0 $Y2=0
cc_505 N_KAPWR_c_490_n N_Y_c_859_n 3.61953e-19 $X=3.92 $Y=2.21 $X2=0 $Y2=0
cc_506 N_KAPWR_c_517_n N_Y_c_859_n 0.0247494f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_507 N_KAPWR_c_486_n N_Y_c_861_n 0.024621f $X=3.775 $Y=2.21 $X2=0 $Y2=0
cc_508 N_KAPWR_c_490_n N_Y_c_861_n 0.00156049f $X=3.92 $Y=2.21 $X2=0 $Y2=0
cc_509 N_KAPWR_c_491_n N_Y_c_861_n 0.0224648f $X=4.635 $Y=2.21 $X2=0 $Y2=0
cc_510 N_KAPWR_c_493_n N_Y_c_861_n 0.0215158f $X=4.49 $Y=2.21 $X2=0 $Y2=0
cc_511 N_KAPWR_c_495_n N_Y_c_861_n 3.77781e-19 $X=4.78 $Y=2.21 $X2=0 $Y2=0
cc_512 N_KAPWR_M1015_d N_Y_c_747_n 0.00173041f $X=5.48 $Y=1.485 $X2=0 $Y2=0
cc_513 N_KAPWR_c_496_n N_Y_c_747_n 0.00438817f $X=5.39 $Y=2.21 $X2=0 $Y2=0
cc_514 N_KAPWR_c_498_n N_Y_c_747_n 0.00296134f $X=5.68 $Y=2.21 $X2=0 $Y2=0
cc_515 N_KAPWR_c_499_n N_Y_c_747_n 0.00466889f $X=6.31 $Y=2.21 $X2=0 $Y2=0
cc_516 N_KAPWR_c_519_n N_Y_c_747_n 0.0162521f $X=5.615 $Y=2 $X2=0 $Y2=0
cc_517 N_KAPWR_c_498_n N_Y_c_867_n 3.49974e-19 $X=5.68 $Y=2.21 $X2=0 $Y2=0
cc_518 N_KAPWR_c_499_n N_Y_c_867_n 0.0217888f $X=6.31 $Y=2.21 $X2=0 $Y2=0
cc_519 N_KAPWR_c_501_n N_Y_c_867_n 0.00148428f $X=6.6 $Y=2.21 $X2=0 $Y2=0
cc_520 N_KAPWR_c_519_n N_Y_c_867_n 0.024157f $X=5.615 $Y=2 $X2=0 $Y2=0
cc_521 N_KAPWR_c_521_n N_Y_c_867_n 0.0245532f $X=6.48 $Y=2 $X2=0 $Y2=0
cc_522 N_KAPWR_c_501_n N_Y_c_869_n 3.99336e-19 $X=6.6 $Y=2.21 $X2=0 $Y2=0
cc_523 N_KAPWR_c_502_n N_Y_c_869_n 0.0217503f $X=7.17 $Y=2.21 $X2=0 $Y2=0
cc_524 N_KAPWR_c_504_n N_Y_c_869_n 0.00148428f $X=7.46 $Y=2.21 $X2=0 $Y2=0
cc_525 N_KAPWR_c_521_n N_Y_c_869_n 0.0247052f $X=6.48 $Y=2 $X2=0 $Y2=0
cc_526 N_KAPWR_c_523_n N_Y_c_869_n 0.0245532f $X=7.34 $Y=2 $X2=0 $Y2=0
cc_527 N_KAPWR_c_504_n N_Y_c_871_n 3.99336e-19 $X=7.46 $Y=2.21 $X2=0 $Y2=0
cc_528 N_KAPWR_c_505_n N_Y_c_871_n 0.0217503f $X=8.07 $Y=2.21 $X2=0 $Y2=0
cc_529 N_KAPWR_c_587_p N_Y_c_871_n 4.09742e-19 $X=8.36 $Y=2.21 $X2=0 $Y2=0
cc_530 N_KAPWR_c_523_n N_Y_c_871_n 0.0247263f $X=7.34 $Y=2 $X2=0 $Y2=0
cc_531 N_KAPWR_c_525_n N_Y_c_871_n 0.0247312f $X=8.2 $Y=2 $X2=0 $Y2=0
cc_532 N_KAPWR_c_587_p N_Y_c_748_n 2.70415e-19 $X=8.36 $Y=2.21 $X2=0 $Y2=0
cc_533 N_KAPWR_c_507_n N_Y_c_748_n 0.0217503f $X=8.9 $Y=2.21 $X2=0 $Y2=0
cc_534 N_KAPWR_c_592_p N_Y_c_748_n 2.70415e-19 $X=9.19 $Y=2.21 $X2=0 $Y2=0
cc_535 N_KAPWR_c_525_n N_Y_c_748_n 0.0247107f $X=8.2 $Y=2 $X2=0 $Y2=0
cc_536 N_KAPWR_c_527_n N_Y_c_748_n 0.0247107f $X=9.06 $Y=2 $X2=0 $Y2=0
cc_537 N_KAPWR_c_592_p N_Y_c_749_n 4.09742e-19 $X=9.19 $Y=2.21 $X2=0 $Y2=0
cc_538 N_KAPWR_c_509_n N_Y_c_749_n 0.0185462f $X=9.76 $Y=2.21 $X2=0 $Y2=0
cc_539 N_KAPWR_c_598_p N_Y_c_749_n 4.44943e-19 $X=10.05 $Y=2.21 $X2=0 $Y2=0
cc_540 N_KAPWR_c_527_n N_Y_c_749_n 0.0247107f $X=9.06 $Y=2 $X2=0 $Y2=0
cc_541 N_KAPWR_c_529_n N_Y_c_749_n 0.0247263f $X=9.92 $Y=2 $X2=0 $Y2=0
cc_542 N_KAPWR_c_473_n N_Y_c_750_n 0.0204891f $X=10.66 $Y=2.24 $X2=0 $Y2=0
cc_543 N_KAPWR_c_598_p N_Y_c_750_n 4.09742e-19 $X=10.05 $Y=2.21 $X2=0 $Y2=0
cc_544 N_KAPWR_c_529_n N_Y_c_750_n 0.0247312f $X=9.92 $Y=2 $X2=0 $Y2=0
cc_545 N_KAPWR_c_475_n N_Y_c_750_n 0.0253725f $X=10.775 $Y=2 $X2=0 $Y2=0
cc_546 N_KAPWR_c_491_n Y 0.0249171f $X=4.635 $Y=2.21 $X2=0 $Y2=0
cc_547 N_KAPWR_c_495_n Y 0.00137507f $X=4.78 $Y=2.21 $X2=0 $Y2=0
cc_548 N_KAPWR_c_496_n Y 0.0270411f $X=5.39 $Y=2.21 $X2=0 $Y2=0
cc_549 N_KAPWR_c_498_n Y 0.00157041f $X=5.68 $Y=2.21 $X2=0 $Y2=0
cc_550 N_KAPWR_c_519_n Y 0.0384994f $X=5.615 $Y=2 $X2=0 $Y2=0
cc_551 N_KAPWR_c_473_n N_VPWR_c_1194_n 0.00231062f $X=10.66 $Y=2.24 $X2=0 $Y2=0
cc_552 N_KAPWR_c_479_n N_VPWR_c_1194_n 0.00191865f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_553 N_KAPWR_c_481_n N_VPWR_c_1194_n 2.25071e-19 $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_554 N_KAPWR_c_482_n N_VPWR_c_1194_n 0.00216428f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_555 N_KAPWR_c_484_n N_VPWR_c_1194_n 0.00216924f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_556 N_KAPWR_c_486_n N_VPWR_c_1194_n 0.0188556f $X=3.775 $Y=2.21 $X2=0 $Y2=0
cc_557 N_KAPWR_c_488_n N_VPWR_c_1194_n 0.00216689f $X=3.63 $Y=2.21 $X2=0 $Y2=0
cc_558 N_KAPWR_c_490_n N_VPWR_c_1194_n 9.13511e-19 $X=3.92 $Y=2.21 $X2=0 $Y2=0
cc_559 N_KAPWR_c_491_n N_VPWR_c_1194_n 0.0189299f $X=4.635 $Y=2.21 $X2=0 $Y2=0
cc_560 N_KAPWR_c_493_n N_VPWR_c_1194_n 0.00135031f $X=4.49 $Y=2.21 $X2=0 $Y2=0
cc_561 N_KAPWR_c_495_n N_VPWR_c_1194_n 0.00168435f $X=4.78 $Y=2.21 $X2=0 $Y2=0
cc_562 N_KAPWR_c_496_n N_VPWR_c_1194_n 0.00114201f $X=5.39 $Y=2.21 $X2=0 $Y2=0
cc_563 N_KAPWR_c_498_n N_VPWR_c_1194_n 2.25213e-19 $X=5.68 $Y=2.21 $X2=0 $Y2=0
cc_564 N_KAPWR_c_499_n N_VPWR_c_1194_n 0.00196555f $X=6.31 $Y=2.21 $X2=0 $Y2=0
cc_565 N_KAPWR_c_501_n N_VPWR_c_1194_n 2.22852e-19 $X=6.6 $Y=2.21 $X2=0 $Y2=0
cc_566 N_KAPWR_c_502_n N_VPWR_c_1194_n 0.00194568f $X=7.17 $Y=2.21 $X2=0 $Y2=0
cc_567 N_KAPWR_c_504_n N_VPWR_c_1194_n 2.22852e-19 $X=7.46 $Y=2.21 $X2=0 $Y2=0
cc_568 N_KAPWR_c_505_n N_VPWR_c_1194_n 0.00216924f $X=8.07 $Y=2.21 $X2=0 $Y2=0
cc_569 N_KAPWR_c_507_n N_VPWR_c_1194_n 0.00216924f $X=8.9 $Y=2.21 $X2=0 $Y2=0
cc_570 N_KAPWR_c_509_n N_VPWR_c_1194_n 0.00216924f $X=9.76 $Y=2.21 $X2=0 $Y2=0
cc_571 N_KAPWR_c_474_n N_VPWR_c_1194_n 0.0210175f $X=0.275 $Y=1.66 $X2=0 $Y2=0
cc_572 N_KAPWR_c_513_n N_VPWR_c_1194_n 0.0188556f $X=1.13 $Y=2 $X2=0 $Y2=0
cc_573 N_KAPWR_c_515_n N_VPWR_c_1194_n 0.0188428f $X=1.99 $Y=2 $X2=0 $Y2=0
cc_574 N_KAPWR_c_517_n N_VPWR_c_1194_n 0.0188428f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_575 N_KAPWR_c_519_n N_VPWR_c_1194_n 0.0188556f $X=5.615 $Y=2 $X2=0 $Y2=0
cc_576 N_KAPWR_c_521_n N_VPWR_c_1194_n 0.0188428f $X=6.48 $Y=2 $X2=0 $Y2=0
cc_577 N_KAPWR_c_523_n N_VPWR_c_1194_n 0.0188428f $X=7.34 $Y=2 $X2=0 $Y2=0
cc_578 N_KAPWR_c_525_n N_VPWR_c_1194_n 0.0188428f $X=8.2 $Y=2 $X2=0 $Y2=0
cc_579 N_KAPWR_c_527_n N_VPWR_c_1194_n 0.0188428f $X=9.06 $Y=2 $X2=0 $Y2=0
cc_580 N_KAPWR_c_529_n N_VPWR_c_1194_n 0.0188428f $X=9.92 $Y=2 $X2=0 $Y2=0
cc_581 N_KAPWR_c_475_n N_VPWR_c_1194_n 0.020925f $X=10.775 $Y=2 $X2=0 $Y2=0
cc_582 N_KAPWR_c_476_n N_VPWR_c_1194_n 4.45124e-19 $X=0.36 $Y=2.21 $X2=0 $Y2=0
cc_583 N_KAPWR_M1000_d N_VPWR_c_1193_n 0.00113413f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_584 N_KAPWR_M1001_d N_VPWR_c_1193_n 0.00113459f $X=0.99 $Y=1.485 $X2=0 $Y2=0
cc_585 N_KAPWR_M1003_d N_VPWR_c_1193_n 0.00113449f $X=1.85 $Y=1.485 $X2=0 $Y2=0
cc_586 N_KAPWR_M1006_d N_VPWR_c_1193_n 0.00113449f $X=2.71 $Y=1.485 $X2=0 $Y2=0
cc_587 N_KAPWR_M1010_d N_VPWR_c_1193_n 0.00113459f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_588 N_KAPWR_M1013_d N_VPWR_c_1193_n 0.00127744f $X=4.43 $Y=1.485 $X2=0 $Y2=0
cc_589 N_KAPWR_M1015_d N_VPWR_c_1193_n 0.00113459f $X=5.48 $Y=1.485 $X2=0 $Y2=0
cc_590 N_KAPWR_M1020_d N_VPWR_c_1193_n 0.00113449f $X=6.34 $Y=1.485 $X2=0 $Y2=0
cc_591 N_KAPWR_M1025_d N_VPWR_c_1193_n 0.00113449f $X=7.2 $Y=1.485 $X2=0 $Y2=0
cc_592 N_KAPWR_M1028_d N_VPWR_c_1193_n 0.00113449f $X=8.06 $Y=1.485 $X2=0 $Y2=0
cc_593 N_KAPWR_M1030_d N_VPWR_c_1193_n 0.00113449f $X=8.92 $Y=1.485 $X2=0 $Y2=0
cc_594 N_KAPWR_M1034_d N_VPWR_c_1193_n 0.00113449f $X=9.78 $Y=1.485 $X2=0 $Y2=0
cc_595 N_KAPWR_M1039_d N_VPWR_c_1193_n 0.00109164f $X=10.64 $Y=1.485 $X2=0 $Y2=0
cc_596 N_KAPWR_c_486_n N_VPWR_c_1193_n 0.0029506f $X=3.775 $Y=2.21 $X2=0 $Y2=0
cc_597 N_KAPWR_c_491_n N_VPWR_c_1193_n 0.00298824f $X=4.635 $Y=2.21 $X2=0 $Y2=0
cc_598 N_KAPWR_c_474_n N_VPWR_c_1193_n 0.00299564f $X=0.275 $Y=1.66 $X2=0 $Y2=0
cc_599 N_KAPWR_c_513_n N_VPWR_c_1193_n 0.0029506f $X=1.13 $Y=2 $X2=0 $Y2=0
cc_600 N_KAPWR_c_515_n N_VPWR_c_1193_n 0.00293281f $X=1.99 $Y=2 $X2=0 $Y2=0
cc_601 N_KAPWR_c_517_n N_VPWR_c_1193_n 0.00293281f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_602 N_KAPWR_c_519_n N_VPWR_c_1193_n 0.0029506f $X=5.615 $Y=2 $X2=0 $Y2=0
cc_603 N_KAPWR_c_521_n N_VPWR_c_1193_n 0.00293281f $X=6.48 $Y=2 $X2=0 $Y2=0
cc_604 N_KAPWR_c_523_n N_VPWR_c_1193_n 0.00293281f $X=7.34 $Y=2 $X2=0 $Y2=0
cc_605 N_KAPWR_c_525_n N_VPWR_c_1193_n 0.00293281f $X=8.2 $Y=2 $X2=0 $Y2=0
cc_606 N_KAPWR_c_527_n N_VPWR_c_1193_n 0.00293281f $X=9.06 $Y=2 $X2=0 $Y2=0
cc_607 N_KAPWR_c_529_n N_VPWR_c_1193_n 0.00293281f $X=9.92 $Y=2 $X2=0 $Y2=0
cc_608 N_KAPWR_c_475_n N_VPWR_c_1193_n 0.00297054f $X=10.775 $Y=2 $X2=0 $Y2=0
cc_609 N_KAPWR_c_476_n N_VPWR_c_1193_n 1.11967f $X=0.36 $Y=2.21 $X2=0 $Y2=0
cc_610 N_Y_c_725_n N_VGND_c_1080_n 0.0125932f $X=8.63 $Y=0.445 $X2=0 $Y2=0
cc_611 N_Y_c_718_n N_VGND_c_1084_n 0.0118195f $X=2.42 $Y=0.445 $X2=0 $Y2=0
cc_612 N_Y_c_719_n N_VGND_c_1086_n 0.012748f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_613 N_Y_c_720_n N_VGND_c_1088_n 0.0122837f $X=4.14 $Y=0.445 $X2=0 $Y2=0
cc_614 N_Y_c_721_n N_VGND_c_1090_n 0.0197173f $X=5.065 $Y=0.445 $X2=0 $Y2=0
cc_615 N_Y_c_722_n N_VGND_c_1092_n 0.0125932f $X=6.05 $Y=0.445 $X2=0 $Y2=0
cc_616 N_Y_c_723_n N_VGND_c_1094_n 0.0125932f $X=6.91 $Y=0.445 $X2=0 $Y2=0
cc_617 N_Y_c_724_n N_VGND_c_1096_n 0.0125932f $X=7.77 $Y=0.445 $X2=0 $Y2=0
cc_618 N_Y_M1004_s N_VGND_c_1099_n 0.00423669f $X=2.28 $Y=0.235 $X2=0 $Y2=0
cc_619 N_Y_M1008_s N_VGND_c_1099_n 0.0031965f $X=3.14 $Y=0.235 $X2=0 $Y2=0
cc_620 N_Y_M1016_s N_VGND_c_1099_n 0.0037166f $X=4 $Y=0.235 $X2=0 $Y2=0
cc_621 N_Y_M1018_s N_VGND_c_1099_n 0.00654074f $X=4.895 $Y=0.235 $X2=0 $Y2=0
cc_622 N_Y_M1023_s N_VGND_c_1099_n 0.00336987f $X=5.91 $Y=0.235 $X2=0 $Y2=0
cc_623 N_Y_M1026_s N_VGND_c_1099_n 0.00336987f $X=6.77 $Y=0.235 $X2=0 $Y2=0
cc_624 N_Y_M1033_s N_VGND_c_1099_n 0.00336987f $X=7.63 $Y=0.235 $X2=0 $Y2=0
cc_625 N_Y_M1036_s N_VGND_c_1099_n 0.00336987f $X=8.49 $Y=0.235 $X2=0 $Y2=0
cc_626 N_Y_c_718_n N_VGND_c_1099_n 0.00848423f $X=2.42 $Y=0.445 $X2=0 $Y2=0
cc_627 N_Y_c_719_n N_VGND_c_1099_n 0.00962561f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_628 N_Y_c_720_n N_VGND_c_1099_n 0.00905492f $X=4.14 $Y=0.445 $X2=0 $Y2=0
cc_629 N_Y_c_721_n N_VGND_c_1099_n 0.01324f $X=5.065 $Y=0.445 $X2=0 $Y2=0
cc_630 N_Y_c_722_n N_VGND_c_1099_n 0.00943538f $X=6.05 $Y=0.445 $X2=0 $Y2=0
cc_631 N_Y_c_723_n N_VGND_c_1099_n 0.00943538f $X=6.91 $Y=0.445 $X2=0 $Y2=0
cc_632 N_Y_c_724_n N_VGND_c_1099_n 0.00943538f $X=7.77 $Y=0.445 $X2=0 $Y2=0
cc_633 N_Y_c_725_n N_VGND_c_1099_n 0.00943538f $X=8.63 $Y=0.445 $X2=0 $Y2=0
cc_634 N_Y_c_898_n N_VPWR_c_1194_n 0.0117442f $X=0.7 $Y=2.3 $X2=0 $Y2=0
cc_635 N_Y_c_745_n N_VPWR_c_1194_n 0.0117442f $X=1.56 $Y=1.62 $X2=0 $Y2=0
cc_636 N_Y_c_746_n N_VPWR_c_1194_n 0.0117442f $X=2.42 $Y=1.62 $X2=0 $Y2=0
cc_637 N_Y_c_859_n N_VPWR_c_1194_n 0.0117442f $X=3.28 $Y=1.62 $X2=0 $Y2=0
cc_638 N_Y_c_861_n N_VPWR_c_1194_n 0.0117442f $X=4.14 $Y=1.62 $X2=0 $Y2=0
cc_639 N_Y_c_867_n N_VPWR_c_1194_n 0.0117442f $X=6.05 $Y=1.62 $X2=0 $Y2=0
cc_640 N_Y_c_869_n N_VPWR_c_1194_n 0.0117442f $X=6.91 $Y=1.62 $X2=0 $Y2=0
cc_641 N_Y_c_871_n N_VPWR_c_1194_n 0.0117442f $X=7.77 $Y=1.62 $X2=0 $Y2=0
cc_642 N_Y_c_748_n N_VPWR_c_1194_n 0.0117442f $X=8.63 $Y=1.62 $X2=0 $Y2=0
cc_643 N_Y_c_749_n N_VPWR_c_1194_n 0.0117442f $X=9.49 $Y=1.62 $X2=0 $Y2=0
cc_644 N_Y_c_750_n N_VPWR_c_1194_n 0.0117442f $X=10.35 $Y=1.62 $X2=0 $Y2=0
cc_645 Y N_VPWR_c_1194_n 0.0118139f $X=5.205 $Y=1.445 $X2=0 $Y2=0
cc_646 N_Y_M1000_s N_VPWR_c_1193_n 0.00157789f $X=0.56 $Y=1.485 $X2=0 $Y2=0
cc_647 N_Y_M1002_s N_VPWR_c_1193_n 0.00157789f $X=1.42 $Y=1.485 $X2=0 $Y2=0
cc_648 N_Y_M1005_s N_VPWR_c_1193_n 0.00157789f $X=2.28 $Y=1.485 $X2=0 $Y2=0
cc_649 N_Y_M1009_s N_VPWR_c_1193_n 0.00157789f $X=3.14 $Y=1.485 $X2=0 $Y2=0
cc_650 N_Y_M1012_s N_VPWR_c_1193_n 0.00157789f $X=4 $Y=1.485 $X2=0 $Y2=0
cc_651 N_Y_M1014_s N_VPWR_c_1193_n 0.00285594f $X=4.895 $Y=1.485 $X2=0 $Y2=0
cc_652 N_Y_M1019_s N_VPWR_c_1193_n 0.00157789f $X=5.91 $Y=1.485 $X2=0 $Y2=0
cc_653 N_Y_M1022_s N_VPWR_c_1193_n 0.00157789f $X=6.77 $Y=1.485 $X2=0 $Y2=0
cc_654 N_Y_M1027_s N_VPWR_c_1193_n 0.00157789f $X=7.63 $Y=1.485 $X2=0 $Y2=0
cc_655 N_Y_M1029_s N_VPWR_c_1193_n 0.00157789f $X=8.49 $Y=1.485 $X2=0 $Y2=0
cc_656 N_Y_M1031_s N_VPWR_c_1193_n 0.00157789f $X=9.35 $Y=1.485 $X2=0 $Y2=0
cc_657 N_Y_M1038_s N_VPWR_c_1193_n 0.00157789f $X=10.21 $Y=1.485 $X2=0 $Y2=0
cc_658 N_Y_c_898_n N_VPWR_c_1193_n 0.00154881f $X=0.7 $Y=2.3 $X2=0 $Y2=0
cc_659 N_Y_c_745_n N_VPWR_c_1193_n 0.00154881f $X=1.56 $Y=1.62 $X2=0 $Y2=0
cc_660 N_Y_c_746_n N_VPWR_c_1193_n 0.00154881f $X=2.42 $Y=1.62 $X2=0 $Y2=0
cc_661 N_Y_c_859_n N_VPWR_c_1193_n 0.00154881f $X=3.28 $Y=1.62 $X2=0 $Y2=0
cc_662 N_Y_c_861_n N_VPWR_c_1193_n 0.00154881f $X=4.14 $Y=1.62 $X2=0 $Y2=0
cc_663 N_Y_c_867_n N_VPWR_c_1193_n 0.00154881f $X=6.05 $Y=1.62 $X2=0 $Y2=0
cc_664 N_Y_c_869_n N_VPWR_c_1193_n 0.00154881f $X=6.91 $Y=1.62 $X2=0 $Y2=0
cc_665 N_Y_c_871_n N_VPWR_c_1193_n 0.00154881f $X=7.77 $Y=1.62 $X2=0 $Y2=0
cc_666 N_Y_c_748_n N_VPWR_c_1193_n 0.00154881f $X=8.63 $Y=1.62 $X2=0 $Y2=0
cc_667 N_Y_c_749_n N_VPWR_c_1193_n 0.00154881f $X=9.49 $Y=1.62 $X2=0 $Y2=0
cc_668 N_Y_c_750_n N_VPWR_c_1193_n 0.00154881f $X=10.35 $Y=1.62 $X2=0 $Y2=0
cc_669 Y N_VPWR_c_1193_n 0.00155926f $X=5.205 $Y=1.445 $X2=0 $Y2=0

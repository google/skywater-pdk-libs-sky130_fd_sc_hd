* NGSPICE file created from sky130_fd_sc_hd__o311ai_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A2 a_138_47# VNB nshort w=420000u l=150000u
+  ad=2.31e+11p pd=2.78e+06u as=3.696e+11p ps=3.44e+06u
M1001 a_222_369# A2 a_138_369# VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=1.728e+11p ps=1.82e+06u
M1002 VPWR B1 Y VPB phighvt w=640000u l=150000u
+  ad=4.16e+11p pd=3.86e+06u as=4.864e+11p ps=4.08e+06u
M1003 Y C1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_138_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_138_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 a_458_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1007 a_458_47# B1 a_138_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_138_369# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A3 a_222_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_4.pxi.spice
* Created: Tue Sep  1 19:11:20 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%A N_A_M1000_g N_A_M1002_g N_A_M1001_g
+ N_A_c_68_n N_A_M1003_g N_A_M1004_g N_A_c_71_n N_A_M1008_g N_A_M1005_g
+ N_A_c_74_n N_A_M1009_g N_A_M1006_g N_A_M1007_g N_A_c_78_n N_A_c_79_n
+ N_A_c_80_n N_A_c_81_n N_A_c_82_n N_A_c_83_n N_A_c_84_n A A A A A
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%KAPWR N_KAPWR_M1000_s N_KAPWR_M1001_s
+ N_KAPWR_M1005_s N_KAPWR_M1007_s N_KAPWR_c_177_n N_KAPWR_c_178_n
+ N_KAPWR_c_181_n N_KAPWR_c_183_n N_KAPWR_c_184_n N_KAPWR_c_186_n KAPWR
+ N_KAPWR_c_187_n N_KAPWR_c_188_n N_KAPWR_c_190_n N_KAPWR_c_192_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%Y N_Y_M1002_s N_Y_M1008_s N_Y_M1000_d
+ N_Y_M1004_d N_Y_M1006_d N_Y_c_251_n N_Y_c_252_n N_Y_c_253_n N_Y_c_263_n
+ N_Y_c_264_n N_Y_c_281_n N_Y_c_265_n N_Y_c_254_n N_Y_c_255_n N_Y_c_293_n
+ N_Y_c_266_n N_Y_c_256_n N_Y_c_257_n N_Y_c_304_n N_Y_c_267_n N_Y_c_268_n
+ N_Y_c_258_n N_Y_c_269_n N_Y_c_259_n N_Y_c_270_n Y Y Y N_Y_c_261_n N_Y_c_272_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%Y
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%VGND N_VGND_M1002_d N_VGND_M1003_d
+ N_VGND_M1009_d N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n VGND
+ N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n
+ N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%VPWR VPWR N_VPWR_c_438_n
+ N_VPWR_c_437_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4%VPWR
cc_1 VNB N_A_M1000_g 5.00591e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_2 VNB N_A_M1002_g 0.0369233f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.445
cc_3 VNB N_A_M1001_g 4.57532e-19 $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.985
cc_4 VNB N_A_c_68_n 0.0126448f $X=-0.19 $Y=-0.24 $X2=1.3 $Y2=1.16
cc_5 VNB N_A_M1003_g 0.0279614f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.445
cc_6 VNB N_A_M1004_g 4.57707e-19 $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.985
cc_7 VNB N_A_c_71_n 0.0126445f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_8 VNB N_A_M1008_g 0.0279614f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.445
cc_9 VNB N_A_M1005_g 4.57707e-19 $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.985
cc_10 VNB N_A_c_74_n 0.0126448f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.16
cc_11 VNB N_A_M1009_g 0.0367478f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=0.445
cc_12 VNB N_A_M1006_g 4.57415e-19 $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.985
cc_13 VNB N_A_M1007_g 4.94191e-19 $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.985
cc_14 VNB N_A_c_78_n 0.0151897f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_15 VNB N_A_c_79_n 0.0172072f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.16
cc_16 VNB N_A_c_80_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.16
cc_17 VNB N_A_c_81_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.16
cc_18 VNB N_A_c_82_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_19 VNB N_A_c_83_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.16
cc_20 VNB N_A_c_84_n 0.0321714f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.16
cc_21 VNB N_Y_c_251_n 0.0201292f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.445
cc_22 VNB N_Y_c_252_n 0.0142122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_253_n 0.0104981f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.295
cc_24 VNB N_Y_c_254_n 0.00119645f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.985
cc_25 VNB N_Y_c_255_n 0.00514362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_256_n 0.00119511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_257_n 0.0120925f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.985
cc_28 VNB N_Y_c_258_n 0.00208412f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.16
cc_29 VNB N_Y_c_259_n 0.00203725f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_30 VNB Y 0.0231444f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.105
cc_31 VNB N_Y_c_261_n 0.0132357f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_32 VNB N_VGND_c_392_n 0.00482504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_393_n 0.00400382f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.445
cc_34 VNB N_VGND_c_394_n 0.00484653f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.985
cc_35 VNB N_VGND_c_395_n 0.0184172f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.16
cc_36 VNB N_VGND_c_396_n 0.0154375f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.295
cc_37 VNB N_VGND_c_397_n 0.0152868f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_38 VNB N_VGND_c_398_n 0.0194663f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.985
cc_39 VNB N_VGND_c_399_n 0.191074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_400_n 0.00564654f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.985
cc_41 VNB N_VGND_c_401_n 0.00497354f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.16
cc_42 VNB N_VGND_c_402_n 0.00574268f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_43 VNB N_VPWR_c_437_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.295
cc_44 VPB N_A_M1000_g 0.0232949f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_45 VPB N_A_M1001_g 0.0195526f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.985
cc_46 VPB N_A_M1004_g 0.0195731f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_47 VPB N_A_M1005_g 0.0195731f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_48 VPB N_A_M1006_g 0.0195506f $X=-0.19 $Y=1.305 $X2=2.235 $Y2=1.985
cc_49 VPB N_A_M1007_g 0.0231846f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.985
cc_50 VPB N_KAPWR_c_177_n 0.0122581f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.16
cc_51 VPB N_KAPWR_c_178_n 0.00948585f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=0.445
cc_52 VPB N_Y_c_251_n 0.00764075f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=0.445
cc_53 VPB N_Y_c_263_n 0.00273171f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_54 VPB N_Y_c_264_n 0.00777503f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_55 VPB N_Y_c_265_n 0.00324518f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=0.445
cc_56 VPB N_Y_c_266_n 0.00324518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_Y_c_267_n 0.00177748f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.16
cc_58 VPB N_Y_c_268_n 0.00126996f $X=-0.19 $Y=1.305 $X2=2.31 $Y2=1.16
cc_59 VPB N_Y_c_269_n 0.00126996f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.16
cc_60 VPB N_Y_c_270_n 0.00126996f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_61 VPB Y 0.00841183f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.105
cc_62 VPB N_Y_c_272_n 0.00831511f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_63 VPB N_VPWR_c_438_n 0.0892897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_437_n 0.0427359f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.295
cc_65 N_A_M1006_g N_KAPWR_c_178_n 0.00243525f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1007_g N_KAPWR_c_178_n 0.00247485f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_KAPWR_c_181_n 0.00247485f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_M1001_g N_KAPWR_c_181_n 0.00243525f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_M1001_g N_KAPWR_c_183_n 5.00343e-19 $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A_M1004_g N_KAPWR_c_184_n 0.00247485f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_KAPWR_c_184_n 0.00247485f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_M1006_g N_KAPWR_c_186_n 5.00343e-19 $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_KAPWR_c_187_n 0.00689624f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_M1001_g N_KAPWR_c_188_n 0.00675868f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_KAPWR_c_188_n 0.00695476f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1005_g N_KAPWR_c_190_n 0.00695476f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_KAPWR_c_190_n 0.00675868f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1007_g N_KAPWR_c_192_n 0.00695417f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_Y_c_251_n 0.00284045f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_c_78_n N_Y_c_251_n 0.0135164f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_81 A N_Y_c_251_n 0.0178211f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_Y_c_252_n 0.0142819f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_c_78_n N_Y_c_252_n 0.01134f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_84 A N_Y_c_252_n 0.042008f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A_M1000_g N_Y_c_263_n 0.0130871f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_86 A N_Y_c_263_n 0.0139884f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_M1000_g N_Y_c_281_n 4.8033e-19 $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1001_g N_Y_c_281_n 4.8033e-19 $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1001_g N_Y_c_265_n 0.011554f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_c_68_n N_Y_c_265_n 0.00216422f $X=1.3 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_M1004_g N_Y_c_265_n 0.0115772f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_92 A N_Y_c_265_n 0.0490463f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_M1002_g N_Y_c_254_n 0.00194229f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_M1003_g N_Y_c_254_n 0.00105846f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_M1003_g N_Y_c_255_n 0.0122413f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_c_71_n N_Y_c_255_n 0.00225558f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_M1008_g N_Y_c_255_n 0.0122413f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_98 A N_Y_c_255_n 0.0424729f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_99 N_A_M1004_g N_Y_c_293_n 4.8033e-19 $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_M1005_g N_Y_c_293_n 4.8033e-19 $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_M1005_g N_Y_c_266_n 0.0115772f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_c_74_n N_Y_c_266_n 0.00216422f $X=2.16 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_M1006_g N_Y_c_266_n 0.011554f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_104 A N_Y_c_266_n 0.0490463f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_105 N_A_M1008_g N_Y_c_256_n 0.00105549f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_M1009_g N_Y_c_256_n 0.00192273f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_Y_c_257_n 0.0142819f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_c_84_n N_Y_c_257_n 0.0116658f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_109 A N_Y_c_257_n 0.0368972f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_110 N_A_M1006_g N_Y_c_304_n 4.8033e-19 $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_M1007_g N_Y_c_304_n 4.8033e-19 $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_M1007_g N_Y_c_267_n 0.0139395f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_113 A N_Y_c_267_n 0.00879289f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_114 N_A_c_79_n N_Y_c_268_n 0.00225251f $X=0.87 $Y=1.16 $X2=0 $Y2=0
cc_115 A N_Y_c_268_n 0.0139725f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A_c_68_n N_Y_c_258_n 0.00233861f $X=1.3 $Y=1.16 $X2=0 $Y2=0
cc_117 A N_Y_c_258_n 0.02119f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_c_71_n N_Y_c_269_n 0.00225251f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_119 A N_Y_c_269_n 0.0139725f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A_c_74_n N_Y_c_259_n 0.00233861f $X=2.16 $Y=1.16 $X2=0 $Y2=0
cc_121 A N_Y_c_259_n 0.0207824f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_c_84_n N_Y_c_270_n 0.00225251f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_123 A N_Y_c_270_n 0.0139725f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_M1009_g Y 0.00326216f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_c_84_n Y 0.0152731f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_126 A Y 0.0181732f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A_M1002_g N_VGND_c_392_n 0.00341694f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_M1003_g N_VGND_c_393_n 0.00161372f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A_M1008_g N_VGND_c_393_n 0.00160701f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_M1009_g N_VGND_c_394_n 0.00344739f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_M1002_g N_VGND_c_396_n 0.00437852f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_M1003_g N_VGND_c_396_n 0.00437852f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_M1008_g N_VGND_c_397_n 0.00437852f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A_M1009_g N_VGND_c_397_n 0.00437852f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_M1002_g N_VGND_c_399_n 0.00718425f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_M1003_g N_VGND_c_399_n 0.00588456f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_M1008_g N_VGND_c_399_n 0.00588456f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_M1009_g N_VGND_c_399_n 0.00717171f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_VPWR_c_438_n 0.0054895f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1001_g N_VPWR_c_438_n 0.0054895f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1004_g N_VPWR_c_438_n 0.0054895f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1005_g N_VPWR_c_438_n 0.0054895f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1006_g N_VPWR_c_438_n 0.0054895f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1007_g N_VPWR_c_438_n 0.0054895f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_VPWR_c_437_n 0.00613268f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1001_g N_VPWR_c_437_n 0.00516436f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1004_g N_VPWR_c_437_n 0.00516436f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_VPWR_c_437_n 0.00516436f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_VPWR_c_437_n 0.00516436f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_VPWR_c_437_n 0.00616432f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_151 N_KAPWR_c_181_n N_Y_M1000_d 0.00182099f $X=0.995 $Y=2.21 $X2=0 $Y2=0
cc_152 N_KAPWR_c_184_n N_Y_M1004_d 0.00182099f $X=1.895 $Y=2.21 $X2=0 $Y2=0
cc_153 N_KAPWR_c_178_n N_Y_M1006_d 0.00182099f $X=2.775 $Y=2.24 $X2=0 $Y2=0
cc_154 N_KAPWR_M1000_s N_Y_c_263_n 0.00110444f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_155 N_KAPWR_c_177_n N_Y_c_263_n 6.18045e-19 $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_156 N_KAPWR_c_181_n N_Y_c_263_n 0.00534243f $X=0.995 $Y=2.21 $X2=0 $Y2=0
cc_157 N_KAPWR_c_187_n N_Y_c_263_n 0.0101368f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_158 N_KAPWR_M1000_s N_Y_c_264_n 0.00249672f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_159 N_KAPWR_c_177_n N_Y_c_264_n 0.00180545f $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_160 N_KAPWR_c_187_n N_Y_c_264_n 0.0119953f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_161 N_KAPWR_c_177_n N_Y_c_281_n 4.04466e-19 $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_162 N_KAPWR_c_181_n N_Y_c_281_n 0.0183847f $X=0.995 $Y=2.21 $X2=0 $Y2=0
cc_163 N_KAPWR_c_183_n N_Y_c_281_n 0.00147497f $X=1.285 $Y=2.21 $X2=0 $Y2=0
cc_164 N_KAPWR_c_187_n N_Y_c_281_n 0.0248872f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_165 N_KAPWR_c_188_n N_Y_c_281_n 0.0247324f $X=1.16 $Y=1.965 $X2=0 $Y2=0
cc_166 N_KAPWR_M1001_s N_Y_c_265_n 0.00171343f $X=1.02 $Y=1.485 $X2=0 $Y2=0
cc_167 N_KAPWR_c_181_n N_Y_c_265_n 0.00516424f $X=0.995 $Y=2.21 $X2=0 $Y2=0
cc_168 N_KAPWR_c_183_n N_Y_c_265_n 0.00118572f $X=1.285 $Y=2.21 $X2=0 $Y2=0
cc_169 N_KAPWR_c_184_n N_Y_c_265_n 0.00534243f $X=1.895 $Y=2.21 $X2=0 $Y2=0
cc_170 N_KAPWR_c_188_n N_Y_c_265_n 0.0164188f $X=1.16 $Y=1.965 $X2=0 $Y2=0
cc_171 N_KAPWR_c_183_n N_Y_c_293_n 4.04466e-19 $X=1.285 $Y=2.21 $X2=0 $Y2=0
cc_172 N_KAPWR_c_184_n N_Y_c_293_n 0.0183847f $X=1.895 $Y=2.21 $X2=0 $Y2=0
cc_173 N_KAPWR_c_186_n N_Y_c_293_n 4.04466e-19 $X=2.185 $Y=2.21 $X2=0 $Y2=0
cc_174 N_KAPWR_c_188_n N_Y_c_293_n 0.024908f $X=1.16 $Y=1.965 $X2=0 $Y2=0
cc_175 N_KAPWR_c_190_n N_Y_c_293_n 0.024908f $X=2.02 $Y=1.965 $X2=0 $Y2=0
cc_176 N_KAPWR_M1005_s N_Y_c_266_n 0.00171343f $X=1.88 $Y=1.485 $X2=0 $Y2=0
cc_177 N_KAPWR_c_178_n N_Y_c_266_n 0.00516424f $X=2.775 $Y=2.24 $X2=0 $Y2=0
cc_178 N_KAPWR_c_184_n N_Y_c_266_n 0.00534243f $X=1.895 $Y=2.21 $X2=0 $Y2=0
cc_179 N_KAPWR_c_186_n N_Y_c_266_n 0.00118572f $X=2.185 $Y=2.21 $X2=0 $Y2=0
cc_180 N_KAPWR_c_190_n N_Y_c_266_n 0.0164188f $X=2.02 $Y=1.965 $X2=0 $Y2=0
cc_181 N_KAPWR_c_178_n N_Y_c_304_n 0.0187695f $X=2.775 $Y=2.24 $X2=0 $Y2=0
cc_182 N_KAPWR_c_186_n N_Y_c_304_n 0.00147497f $X=2.185 $Y=2.21 $X2=0 $Y2=0
cc_183 N_KAPWR_c_190_n N_Y_c_304_n 0.0247324f $X=2.02 $Y=1.965 $X2=0 $Y2=0
cc_184 N_KAPWR_c_192_n N_Y_c_304_n 0.0248872f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_185 N_KAPWR_M1007_s N_Y_c_267_n 3.8191e-19 $X=2.74 $Y=1.485 $X2=0 $Y2=0
cc_186 N_KAPWR_c_178_n N_Y_c_267_n 0.00566427f $X=2.775 $Y=2.24 $X2=0 $Y2=0
cc_187 N_KAPWR_c_192_n N_Y_c_267_n 0.00466491f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_188 N_KAPWR_M1007_s N_Y_c_272_n 0.00444506f $X=2.74 $Y=1.485 $X2=0 $Y2=0
cc_189 N_KAPWR_c_178_n N_Y_c_272_n 0.00459252f $X=2.775 $Y=2.24 $X2=0 $Y2=0
cc_190 N_KAPWR_c_192_n N_Y_c_272_n 0.018036f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_191 N_KAPWR_c_177_n N_VPWR_c_438_n 5.71511e-19 $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_192 N_KAPWR_c_178_n N_VPWR_c_438_n 0.00274212f $X=2.775 $Y=2.24 $X2=0 $Y2=0
cc_193 N_KAPWR_c_181_n N_VPWR_c_438_n 0.00195383f $X=0.995 $Y=2.21 $X2=0 $Y2=0
cc_194 N_KAPWR_c_183_n N_VPWR_c_438_n 2.22823e-19 $X=1.285 $Y=2.21 $X2=0 $Y2=0
cc_195 N_KAPWR_c_184_n N_VPWR_c_438_n 0.00217991f $X=1.895 $Y=2.21 $X2=0 $Y2=0
cc_196 N_KAPWR_c_187_n N_VPWR_c_438_n 0.0209643f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_197 N_KAPWR_c_188_n N_VPWR_c_438_n 0.0189011f $X=1.16 $Y=1.965 $X2=0 $Y2=0
cc_198 N_KAPWR_c_190_n N_VPWR_c_438_n 0.0189011f $X=2.02 $Y=1.965 $X2=0 $Y2=0
cc_199 N_KAPWR_c_192_n N_VPWR_c_438_n 0.0209643f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_200 N_KAPWR_M1000_s N_VPWR_c_437_n 0.00125752f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_201 N_KAPWR_M1001_s N_VPWR_c_437_n 0.00113449f $X=1.02 $Y=1.485 $X2=0 $Y2=0
cc_202 N_KAPWR_M1005_s N_VPWR_c_437_n 0.00113449f $X=1.88 $Y=1.485 $X2=0 $Y2=0
cc_203 N_KAPWR_M1007_s N_VPWR_c_437_n 0.00159683f $X=2.74 $Y=1.485 $X2=0 $Y2=0
cc_204 N_KAPWR_c_177_n N_VPWR_c_437_n 0.31744f $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_205 N_KAPWR_c_187_n N_VPWR_c_437_n 0.00299364f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_206 N_KAPWR_c_188_n N_VPWR_c_437_n 0.00295042f $X=1.16 $Y=1.965 $X2=0 $Y2=0
cc_207 N_KAPWR_c_190_n N_VPWR_c_437_n 0.00295042f $X=2.02 $Y=1.965 $X2=0 $Y2=0
cc_208 N_KAPWR_c_192_n N_VPWR_c_437_n 0.00299364f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_209 N_Y_c_252_n N_VGND_c_392_n 0.0212491f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_210 N_Y_c_255_n N_VGND_c_393_n 0.0164203f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_211 N_Y_c_257_n N_VGND_c_394_n 0.0214243f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_212 N_Y_c_252_n N_VGND_c_395_n 0.00440462f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_213 N_Y_c_253_n N_VGND_c_395_n 0.00289403f $X=0.275 $Y=0.81 $X2=0 $Y2=0
cc_214 N_Y_c_252_n N_VGND_c_396_n 0.0022979f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_215 N_Y_c_254_n N_VGND_c_396_n 0.01283f $X=1.16 $Y=0.445 $X2=0 $Y2=0
cc_216 N_Y_c_255_n N_VGND_c_396_n 0.0022979f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_217 N_Y_c_255_n N_VGND_c_397_n 0.0022979f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_218 N_Y_c_256_n N_VGND_c_397_n 0.0126752f $X=2.02 $Y=0.445 $X2=0 $Y2=0
cc_219 N_Y_c_257_n N_VGND_c_397_n 0.0022979f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_220 N_Y_c_257_n N_VGND_c_398_n 0.00333776f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_221 N_Y_c_261_n N_VGND_c_398_n 0.00510712f $X=2.985 $Y=0.895 $X2=0 $Y2=0
cc_222 N_Y_M1002_s N_VGND_c_399_n 0.00234276f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_223 N_Y_M1008_s N_VGND_c_399_n 0.0023674f $X=1.88 $Y=0.235 $X2=0 $Y2=0
cc_224 N_Y_c_252_n N_VGND_c_399_n 0.0125077f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_225 N_Y_c_253_n N_VGND_c_399_n 0.00478629f $X=0.275 $Y=0.81 $X2=0 $Y2=0
cc_226 N_Y_c_254_n N_VGND_c_399_n 0.00978777f $X=1.16 $Y=0.445 $X2=0 $Y2=0
cc_227 N_Y_c_255_n N_VGND_c_399_n 0.00837675f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_228 N_Y_c_256_n N_VGND_c_399_n 0.00959809f $X=2.02 $Y=0.445 $X2=0 $Y2=0
cc_229 N_Y_c_257_n N_VGND_c_399_n 0.0106771f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_230 N_Y_c_261_n N_VGND_c_399_n 0.0084464f $X=2.985 $Y=0.895 $X2=0 $Y2=0
cc_231 N_Y_c_281_n N_VPWR_c_438_n 0.0098434f $X=0.73 $Y=1.83 $X2=0 $Y2=0
cc_232 N_Y_c_293_n N_VPWR_c_438_n 0.0098434f $X=1.59 $Y=1.83 $X2=0 $Y2=0
cc_233 N_Y_c_304_n N_VPWR_c_438_n 0.0098434f $X=2.45 $Y=1.83 $X2=0 $Y2=0
cc_234 N_Y_M1000_d N_VPWR_c_437_n 0.00159777f $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_235 N_Y_M1004_d N_VPWR_c_437_n 0.00159777f $X=1.45 $Y=1.485 $X2=0 $Y2=0
cc_236 N_Y_M1006_d N_VPWR_c_437_n 0.00159777f $X=2.31 $Y=1.485 $X2=0 $Y2=0
cc_237 N_Y_c_281_n N_VPWR_c_437_n 0.00158462f $X=0.73 $Y=1.83 $X2=0 $Y2=0
cc_238 N_Y_c_293_n N_VPWR_c_437_n 0.00158462f $X=1.59 $Y=1.83 $X2=0 $Y2=0
cc_239 N_Y_c_304_n N_VPWR_c_437_n 0.00158462f $X=2.45 $Y=1.83 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dlymetal6s6s_1.spice
* Created: Tue Sep  1 19:07:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlymetal6s6s_1.pex.spice"
.subckt sky130_fd_sc_hd__dlymetal6s6s_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_63_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_240_47#_M1006_d N_A_63_47#_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=4.608 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A_240_47#_M1000_g N_A_346_47#_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_523_47#_M1005_d N_A_346_47#_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=4.608 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_523_47#_M1003_g N_A_629_47#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_629_47#_M1008_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=4.608 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_A_63_47#_M1011_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=11.7215 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_240_47#_M1009_d N_A_63_47#_M1009_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.198239 PD=2.52 PS=1.8662 NRD=0 NRS=3.9203 M=1 R=6.66667
+ SA=75000.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_240_47#_M1010_g N_A_346_47#_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=11.7215 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_523_47#_M1007_d N_A_346_47#_M1007_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.198239 PD=2.52 PS=1.8662 NRD=0 NRS=3.9203 M=1 R=6.66667
+ SA=75000.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_523_47#_M1001_g N_A_629_47#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=11.7215 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_629_47#_M1004_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.198239 PD=2.52 PS=1.8662 NRD=0 NRS=3.9203 M=1 R=6.66667
+ SA=75000.4 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_90 VPB 0 3.72505e-19 $X=0.125 $Y=2.635
*
.include "sky130_fd_sc_hd__dlymetal6s6s_1.pxi.spice"
*
.ends
*
*

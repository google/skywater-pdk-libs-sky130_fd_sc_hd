* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 a_1061_369# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=2.755e+11p pd=2.33e+06u as=1.505e+12p ps=1.348e+07u
M1001 a_193_369# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.947e+11p pd=1.94e+06u as=0p ps=0u
M1002 VPWR A3 a_373_413# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.29e+11p ps=2.66e+06u
M1003 VGND a_789_316# X VNB nshort w=650000u l=150000u
+  ad=1.04515e+12p pd=1.034e+07u as=3.51e+11p ps=3.68e+06u
M1004 VPWR a_789_316# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1005 X a_789_316# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_288_47# a_27_47# a_193_47# VNB nshort w=360000u l=150000u
+  ad=2.532e+11p pd=2.88e+06u as=1.32e+11p ps=1.49e+06u
M1007 a_873_316# a_601_345# a_789_316# VNB nshort w=420000u l=150000u
+  ad=2.532e+11p pd=2.88e+06u as=1.155e+11p ps=1.39e+06u
M1008 VPWR a_789_316# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_601_345# S1 VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1010 a_873_316# S0 a_1065_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.572e+11p ps=1.61e+06u
M1011 VGND a_789_316# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_789_316# S1 a_288_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_873_316# S1 a_789_316# VPB phighvt w=540000u l=150000u
+  ad=2.538e+11p pd=2.98e+06u as=1.458e+11p ps=1.62e+06u
M1014 X a_789_316# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_789_316# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1280_413# S0 a_873_316# VPB phighvt w=420000u l=150000u
+  ad=2.107e+11p pd=1.99e+06u as=0p ps=0u
M1017 a_373_413# a_27_47# a_288_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.538e+11p ps=2.98e+06u
M1018 a_193_47# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_789_316# a_601_345# a_288_47# VPB phighvt w=540000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A0 a_1282_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1021 VPWR S0 a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1022 VPWR A0 a_1280_413# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_873_316# a_27_47# a_1061_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1065_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_288_47# S0 a_193_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_398_47# S0 a_288_47# VNB nshort w=360000u l=150000u
+  ad=1.341e+11p pd=1.5e+06u as=0p ps=0u
M1027 a_601_345# S1 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1028 a_1282_47# a_27_47# a_873_316# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND S0 a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1030 VGND A3 a_398_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 X a_789_316# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__xor2_1.pex.spice
* Created: Tue Sep  1 19:33:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XOR2_1%B 1 3 6 8 10 13 16 20 21 23 24 29 30 34
c84 29 0 5.71701e-20 $X=0.51 $Y=1.16
c85 21 0 3.51517e-19 $X=1.77 $Y=1.16
c86 16 0 7.82759e-20 $X=1.645 $Y=1.445
r87 32 34 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.67 $Y=1.53 $X2=0.69
+ $Y2=1.53
r88 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r89 24 32 4.20453 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.547 $Y=1.53
+ $X2=0.67 $Y2=1.53
r90 24 30 11.134 $w=3.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.547 $Y=1.445
+ $X2=0.547 $Y2=1.16
r91 24 34 2.0877 $w=1.68e-07 $l=3.2e-08 $layer=LI1_cond $X=0.722 $Y=1.53
+ $X2=0.69 $Y2=1.53
r92 23 24 54.6717 $w=1.68e-07 $l=8.38e-07 $layer=LI1_cond $X=1.56 $Y=1.53
+ $X2=0.722 $Y2=1.53
r93 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r94 17 20 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.645 $Y=1.16
+ $X2=1.77 $Y2=1.16
r95 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=1.445
+ $X2=1.56 $Y2=1.53
r96 15 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.245
+ $X2=1.645 $Y2=1.16
r97 15 16 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.645 $Y=1.245
+ $X2=1.645 $Y2=1.445
r98 11 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.16
r99 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.985
r100 8 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=0.995
+ $X2=1.77 $Y2=1.16
r101 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.77 $Y=0.995
+ $X2=1.77 $Y2=0.56
r102 4 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.325
+ $X2=0.51 $Y2=1.16
r103 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.51 $Y=1.325
+ $X2=0.51 $Y2=1.985
r104 1 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=1.16
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_1%A 1 3 6 8 10 13 15 22
c44 15 0 1.99162e-19 $X=1.15 $Y=1.19
r45 20 22 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.095 $Y=1.16
+ $X2=1.35 $Y2=1.16
r46 17 20 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=1.095 $Y2=1.16
r47 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.16 $X2=1.095 $Y2=1.16
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.985
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=0.56
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.93 $Y=1.325 $X2=0.93
+ $Y2=1.985
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.93 $Y=0.995 $X2=0.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_1%A_35_297# 1 2 7 9 12 14 15 18 20 22 23 26 28
+ 32 35 36
c86 36 0 5.71701e-20 $X=0.72 $Y=0.74
c87 14 0 7.82759e-20 $X=2.615 $Y=1.16
r88 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r89 30 32 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.22 $Y=0.825
+ $X2=2.22 $Y2=1.16
r90 29 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.74
+ $X2=0.72 $Y2=0.74
r91 28 30 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.105 $Y=0.74
+ $X2=2.22 $Y2=0.825
r92 28 29 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=2.105 $Y=0.74
+ $X2=0.805 $Y2=0.74
r93 24 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.655
+ $X2=0.72 $Y2=0.74
r94 24 26 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.72 $Y=0.655
+ $X2=0.72 $Y2=0.5
r95 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=0.74
+ $X2=0.72 $Y2=0.74
r96 22 23 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.635 $Y=0.74
+ $X2=0.255 $Y2=0.74
r97 18 35 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=0.275 $Y=1.975
+ $X2=0.275 $Y2=1.785
r98 18 20 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.275 $Y=1.975
+ $X2=0.275 $Y2=2
r99 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.255 $Y2=0.74
r100 16 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.785
r101 14 33 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.615 $Y=1.16
+ $X2=2.25 $Y2=1.16
r102 14 15 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.16
+ $X2=2.615 $Y2=0.995
r103 10 15 37.0704 $w=1.5e-07 $l=3.745e-07 $layer=POLY_cond $X=2.71 $Y=1.325
+ $X2=2.615 $Y2=0.995
r104 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.71 $Y=1.325
+ $X2=2.71 $Y2=1.985
r105 7 15 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.69 $Y=0.995
+ $X2=2.615 $Y2=0.995
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.69 $Y=0.995
+ $X2=2.69 $Y2=0.56
r107 2 20 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.175
+ $Y=1.485 $X2=0.3 $Y2=2
r108 1 26 182 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.235 $X2=0.72 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_1%VPWR 1 2 9 13 16 17 19 20 21 34 35
r42 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 31 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 25 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 19 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.98 $Y2=2.72
r53 18 31 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.98 $Y2=2.72
r55 16 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=1.14 $Y2=2.72
r57 15 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.225 $Y=2.72
+ $X2=1.61 $Y2=2.72
r58 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.72
+ $X2=1.14 $Y2=2.72
r59 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.72
r60 11 13 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.29
r61 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635 $X2=1.14
+ $Y2=2.72
r62 7 9 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=1.95
r63 2 13 600 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.485 $X2=1.98 $Y2=2.29
r64 1 9 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=1.485 $X2=1.14 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_1%A_285_297# 1 2 9 14 16
c27 14 0 1.52356e-19 $X=1.56 $Y=1.95
r28 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.87
+ $X2=1.56 $Y2=1.87
r29 9 16 5.87433 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.235 $Y=1.87 $X2=2.435
+ $Y2=1.87
r30 9 10 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.235 $Y=1.87
+ $X2=1.725 $Y2=1.87
r31 2 16 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=2.375
+ $Y=1.485 $X2=2.5 $Y2=1.95
r32 1 14 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.425
+ $Y=1.485 $X2=1.56 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_1%X 1 2 7 12 13
r33 16 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.975 $Y=1.45
+ $X2=2.59 $Y2=1.45
r34 13 16 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.99 $Y=1.45
+ $X2=2.975 $Y2=1.45
r35 13 20 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=2.975 $Y=1.575
+ $X2=2.975 $Y2=2.3
r36 13 16 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=2.975 $Y=1.575
+ $X2=2.975 $Y2=1.535
r37 12 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=1.365
+ $X2=2.59 $Y2=1.45
r38 11 12 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.59 $Y=0.485
+ $X2=2.59 $Y2=1.365
r39 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=0.4
+ $X2=2.59 $Y2=0.485
r40 7 9 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.505 $Y=0.4 $X2=2.48
+ $Y2=0.4
r41 2 20 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.485 $X2=2.92 $Y2=2.3
r42 2 13 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.485 $X2=2.92 $Y2=1.62
r43 1 9 91 $w=1.7e-07 $l=7.12741e-07 $layer=licon1_NDIFF $count=2 $X=1.845
+ $Y=0.235 $X2=2.48 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_1%VGND 1 2 3 10 12 16 18 20 22 24 29 41 45
r51 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r54 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r55 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r56 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r57 32 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r58 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r59 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r60 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.61
+ $Y2=0
r61 29 44 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=3.032
+ $Y2=0
r62 29 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.53
+ $Y2=0
r63 28 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r64 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r65 25 38 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.232
+ $Y2=0
r66 25 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.69
+ $Y2=0
r67 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r68 24 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.69
+ $Y2=0
r69 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r70 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 18 44 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=3.032 $Y2=0
r72 18 20 13.114 $w=2.88e-07 $l=3.3e-07 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0.415
r73 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r74 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.39
r75 10 38 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.232 $Y2=0
r76 10 12 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.3 $Y2=0.39
r77 3 20 91 $w=1.7e-07 $l=2.49199e-07 $layer=licon1_NDIFF $count=2 $X=2.765
+ $Y=0.235 $X2=2.93 $Y2=0.415
r78 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.39
r79 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__sdfsbp_2.pex.spice
* Created: Thu Aug 27 14:46:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%SCD 1 2 3 5 6 8 11 13 14
r32 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r33 14 19 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.53
+ $X2=0.212 $Y2=1.16
r34 13 19 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r35 9 11 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.315 $Y=1.695
+ $X2=0.47 $Y2=1.695
r36 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=1.695
r37 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=2.165
r38 3 18 87.63 $w=2.63e-07 $l=4.97242e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.325 $Y2=1.16
r39 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r40 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.315 $Y=1.62
+ $X2=0.315 $Y2=1.695
r41 1 18 39.0634 $w=2.63e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.325 $Y2=1.16
r42 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.315 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%SCE 3 5 7 11 15 17 19 20 26 27 33
c106 27 0 1.45056e-19 $X=2.53 $Y=1.19
c107 26 0 9.29321e-20 $X=2.53 $Y=1.19
r108 33 36 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.16
+ $X2=2.585 $Y2=1.325
r109 33 35 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.16
+ $X2=2.585 $Y2=0.995
r110 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.16 $X2=2.57 $Y2=1.16
r111 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r112 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.19
+ $X2=0.69 $Y2=1.19
r113 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r114 19 20 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.835 $Y2=1.19
r115 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.735
+ $Y=1.25 $X2=0.735 $Y2=1.25
r116 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.19
+ $X2=0.69 $Y2=1.19
r117 15 36 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.66 $Y=2.165
+ $X2=2.66 $Y2=1.325
r118 11 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.655 $Y=0.445
+ $X2=2.655 $Y2=0.995
r119 5 30 38.6139 $w=3.32e-07 $l=2.12238e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.782 $Y2=1.25
r120 5 7 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.89 $Y2=2.165
r121 1 30 38.6139 $w=3.32e-07 $l=1.8747e-07 $layer=POLY_cond $X=0.83 $Y=1.085
+ $X2=0.782 $Y2=1.25
r122 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.83 $Y=1.085 $X2=0.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%D 1 3 6 8 9 13
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=0.93 $X2=1.25 $Y2=0.93
r44 9 14 24.262 $w=2.83e-07 $l=6e-07 $layer=LI1_cond $X=1.192 $Y=1.53 $X2=1.192
+ $Y2=0.93
r45 8 14 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=1.192 $Y=0.85 $X2=1.192
+ $Y2=0.93
r46 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.095
+ $X2=1.25 $Y2=0.93
r47 4 6 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.25 $Y=1.095 $X2=1.25
+ $Y2=2.165
r48 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.765
+ $X2=1.25 $Y2=0.93
r49 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.25 $Y=0.765 $X2=1.25
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_328_21# 1 2 9 13 18 19 20 22 32 34
r79 36 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.715 $Y=1.16
+ $X2=1.73 $Y2=1.16
r80 32 34 1.59569 $w=3.23e-07 $l=4.5e-08 $layer=LI1_cond $X=2.405 $Y=1.922
+ $X2=2.45 $Y2=1.922
r81 20 22 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.395 $Y=0.715
+ $X2=2.395 $Y2=0.44
r82 19 38 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=2.065 $Y=1.16
+ $X2=1.73 $Y2=1.16
r83 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.065
+ $Y=1.16 $X2=2.065 $Y2=1.16
r84 16 32 10.567 $w=3.23e-07 $l=2.98e-07 $layer=LI1_cond $X=2.107 $Y=1.922
+ $X2=2.405 $Y2=1.922
r85 16 18 27.1163 $w=2.53e-07 $l=6e-07 $layer=LI1_cond $X=2.107 $Y=1.76
+ $X2=2.107 $Y2=1.16
r86 15 20 16.8115 $w=1.88e-07 $l=2.88e-07 $layer=LI1_cond $X=2.107 $Y=0.81
+ $X2=2.395 $Y2=0.81
r87 15 18 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=2.107 $Y=0.905
+ $X2=2.107 $Y2=1.16
r88 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r89 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=2.165
r90 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=0.995
+ $X2=1.715 $Y2=1.16
r91 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.715 $Y=0.995
+ $X2=1.715 $Y2=0.445
r92 2 34 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.845 $X2=2.45 $Y2=1.99
r93 1 22 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.235 $X2=2.445 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%CLK 4 5 7 8 10 13 17 19 20 21 22 28 30
c78 30 0 8.82473e-21 $X=3.43 $Y=1.09
c79 22 0 1.05862e-19 $X=3.45 $Y=1.19
c80 13 0 1.07468e-19 $X=3.595 $Y=0.805
c81 4 0 2.11828e-19 $X=3.49 $Y=1.62
r82 36 43 7.01796 $w=1.95e-07 $l=2.8e-07 $layer=LI1_cond $X=3.002 $Y=1.615
+ $X2=3.002 $Y2=1.335
r83 32 43 7.01796 $w=1.95e-07 $l=2.8e-07 $layer=LI1_cond $X=3.002 $Y=1.055
+ $X2=3.002 $Y2=1.335
r84 28 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.42
r85 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.09
r86 22 43 9.14146 $w=5.58e-07 $l=4.28e-07 $layer=LI1_cond $X=3.43 $Y=1.335
+ $X2=3.002 $Y2=1.335
r87 22 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.255 $X2=3.43 $Y2=1.255
r88 21 36 14.5035 $w=1.93e-07 $l=2.55e-07 $layer=LI1_cond $X=3.002 $Y=1.87
+ $X2=3.002 $Y2=1.615
r89 20 43 0.256303 $w=5.58e-07 $l=1.2e-08 $layer=LI1_cond $X=2.99 $Y=1.335
+ $X2=3.002 $Y2=1.335
r90 19 32 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.002 $Y=0.85
+ $X2=3.002 $Y2=1.055
r91 15 17 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=3.49 $Y=1.695
+ $X2=3.6 $Y2=1.695
r92 11 13 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=3.49 $Y=0.805
+ $X2=3.595 $Y2=0.805
r93 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.6 $Y=1.77 $X2=3.6
+ $Y2=1.695
r94 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.6 $Y=1.77 $X2=3.6
+ $Y2=2.165
r95 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=0.73
+ $X2=3.595 $Y2=0.805
r96 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.595 $Y=0.73 $X2=3.595
+ $Y2=0.445
r97 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=1.62 $X2=3.49
+ $Y2=1.695
r98 4 31 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.49 $Y=1.62 $X2=3.49
+ $Y2=1.42
r99 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=0.805
r100 1 30 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.49 $Y=0.88
+ $X2=3.49 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_652_47# 1 2 8 9 11 12 14 16 18 20 23 27
+ 31 33 36 40 42 43 44 45 47 49 54 55 56 57 60 61 63 64 65 66 67 76 81 82
c288 81 0 1.18775e-19 $X=5.38 $Y=1.74
c289 76 0 2.10875e-19 $X=7.645 $Y=1.87
c290 64 0 1.51716e-19 $X=5.2 $Y=1.87
c291 61 0 9.42889e-20 $X=8.93 $Y=1.1
c292 60 0 3.15377e-19 $X=8.93 $Y=1.1
c293 49 0 7.55977e-20 $X=3.91 $Y=1.255
c294 12 0 1.20946e-19 $X=4.02 $Y=1.68
c295 8 0 3.22574e-20 $X=3.985 $Y=1.09
r296 81 84 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.74
+ $X2=5.38 $Y2=1.905
r297 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.38
+ $Y=1.74 $X2=5.38 $Y2=1.74
r298 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.645 $Y=1.87
+ $X2=7.645 $Y2=1.87
r299 73 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.345 $Y=1.87
+ $X2=5.345 $Y2=1.87
r300 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=1.87
+ $X2=3.91 $Y2=1.87
r301 67 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.49 $Y=1.87
+ $X2=5.345 $Y2=1.87
r302 66 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.5 $Y=1.87
+ $X2=7.645 $Y2=1.87
r303 66 67 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=7.5 $Y=1.87
+ $X2=5.49 $Y2=1.87
r304 65 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=1.87
+ $X2=3.91 $Y2=1.87
r305 64 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.2 $Y=1.87
+ $X2=5.345 $Y2=1.87
r306 64 65 1.41708 $w=1.4e-07 $l=1.145e-06 $layer=MET1_cond $X=5.2 $Y=1.87
+ $X2=4.055 $Y2=1.87
r307 63 77 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=7.885 $Y=1.83
+ $X2=7.645 $Y2=1.83
r308 61 89 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.93 $Y=1.1
+ $X2=8.93 $Y2=0.935
r309 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.93
+ $Y=1.1 $X2=8.93 $Y2=1.1
r310 58 60 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=8.957 $Y=0.895
+ $X2=8.957 $Y2=1.1
r311 56 58 6.94684 $w=2e-07 $l=1.69791e-07 $layer=LI1_cond $X=8.83 $Y=0.795
+ $X2=8.957 $Y2=0.895
r312 56 57 42.9773 $w=1.98e-07 $l=7.75e-07 $layer=LI1_cond $X=8.83 $Y=0.795
+ $X2=8.055 $Y2=0.795
r313 55 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.97 $Y=1.16
+ $X2=7.97 $Y2=1.325
r314 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.16 $X2=7.97 $Y2=1.16
r315 52 63 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.97 $Y=1.705
+ $X2=7.885 $Y2=1.83
r316 52 54 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.97 $Y=1.705
+ $X2=7.97 $Y2=1.16
r317 51 57 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.97 $Y=0.895
+ $X2=8.055 $Y2=0.795
r318 51 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.97 $Y=0.895
+ $X2=7.97 $Y2=1.16
r319 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=1.255 $X2=3.91 $Y2=1.255
r320 47 70 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=1.83
+ $X2=3.865 $Y2=1.915
r321 47 49 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.865 $Y=1.83
+ $X2=3.865 $Y2=1.255
r322 46 49 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.865 $Y=0.885
+ $X2=3.865 $Y2=1.255
r323 44 70 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.735 $Y=1.915
+ $X2=3.865 $Y2=1.915
r324 44 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.735 $Y=1.915
+ $X2=3.475 $Y2=1.915
r325 42 46 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.865 $Y2=0.885
r326 42 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.47 $Y2=0.8
r327 38 45 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=3.372 $Y=2
+ $X2=3.475 $Y2=1.915
r328 38 40 8.65632 $w=2.03e-07 $l=1.6e-07 $layer=LI1_cond $X=3.372 $Y=2
+ $X2=3.372 $Y2=2.16
r329 34 43 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.37 $Y=0.715
+ $X2=3.47 $Y2=0.8
r330 34 36 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.37 $Y=0.715
+ $X2=3.37 $Y2=0.44
r331 31 89 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.99 $Y=0.445
+ $X2=8.99 $Y2=0.935
r332 27 87 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.91 $Y=2.065
+ $X2=7.91 $Y2=1.325
r333 23 84 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.435 $Y=2.275
+ $X2=5.435 $Y2=1.905
r334 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.955 $Y=0.73
+ $X2=4.955 $Y2=0.445
r335 17 33 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.09 $Y=0.805 $X2=4
+ $Y2=0.805
r336 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.88 $Y=0.805
+ $X2=4.955 $Y2=0.73
r337 16 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.88 $Y=0.805
+ $X2=4.09 $Y2=0.805
r338 12 50 91.0612 $w=2.44e-07 $l=4.65564e-07 $layer=POLY_cond $X=4.02 $Y=1.68
+ $X2=3.935 $Y2=1.255
r339 12 14 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.02 $Y=1.68
+ $X2=4.02 $Y2=2.165
r340 9 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=4.015 $Y=0.73
+ $X2=4 $Y2=0.805
r341 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.015 $Y=0.73
+ $X2=4.015 $Y2=0.445
r342 8 50 39.7006 $w=2.44e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.985 $Y=1.09
+ $X2=3.935 $Y2=1.255
r343 7 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=4 $Y2=0.805
r344 7 8 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.985 $Y2=1.09
r345 2 40 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.845 $X2=3.39 $Y2=2.16
r346 1 36 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.26
+ $Y=0.235 $X2=3.385 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_818_47# 1 2 8 9 11 13 15 18 21 23 25 29
+ 31 32 38 42 43 45 46 49 52 53 60 69
c194 69 0 8.03561e-20 $X=4.327 $Y=1.09
c195 49 0 3.35674e-20 $X=4.37 $Y=1.19
c196 32 0 2.4546e-19 $X=5.345 $Y=0.86
c197 31 0 1.78833e-19 $X=5.345 $Y=0.73
c198 23 0 5.6211e-20 $X=8.54 $Y=1.905
c199 9 0 1.51716e-19 $X=5.24 $Y=1.165
r200 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.56
+ $Y=1.74 $X2=8.56 $Y2=1.74
r201 59 60 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.255
+ $X2=4.745 $Y2=1.255
r202 56 59 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=4.405 $Y=1.255
+ $X2=4.67 $Y2=1.255
r203 53 63 27.5584 $w=2.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.535 $Y=1.19
+ $X2=8.535 $Y2=1.74
r204 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.565 $Y=1.19
+ $X2=8.565 $Y2=1.19
r205 49 70 8.46186 $w=3.23e-07 $l=2.3e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.42
r206 49 69 6.15528 $w=3.23e-07 $l=1e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.09
r207 49 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.255 $X2=4.405 $Y2=1.255
r208 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.19
r209 46 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=1.19
+ $X2=4.37 $Y2=1.19
r210 45 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.42 $Y=1.19
+ $X2=8.565 $Y2=1.19
r211 45 46 4.83291 $w=1.4e-07 $l=3.905e-06 $layer=MET1_cond $X=8.42 $Y=1.19
+ $X2=4.515 $Y2=1.19
r212 43 70 29.9635 $w=2.73e-07 $l=7.15e-07 $layer=LI1_cond $X=4.302 $Y=2.135
+ $X2=4.302 $Y2=1.42
r213 42 43 6.5155 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=4.292 $Y=2.3
+ $X2=4.292 $Y2=2.135
r214 40 69 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.25 $Y=0.585
+ $X2=4.25 $Y2=1.09
r215 38 40 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=4.222 $Y=0.42
+ $X2=4.222 $Y2=0.585
r216 31 32 60.6369 $w=1.6e-07 $l=1.3e-07 $layer=POLY_cond $X=5.345 $Y=0.73
+ $X2=5.345 $Y2=0.86
r217 27 29 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.67 $Y=1.915
+ $X2=4.96 $Y2=1.915
r218 23 62 38.5495 $w=3.2e-07 $l=1.81659e-07 $layer=POLY_cond $X=8.54 $Y=1.905
+ $X2=8.505 $Y2=1.74
r219 23 25 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.54 $Y=1.905
+ $X2=8.54 $Y2=2.275
r220 19 62 38.5495 $w=3.2e-07 $l=2.14942e-07 $layer=POLY_cond $X=8.39 $Y=1.575
+ $X2=8.505 $Y2=1.74
r221 19 21 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=8.39 $Y=1.575
+ $X2=8.39 $Y2=0.555
r222 18 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.375 $Y=0.445
+ $X2=5.375 $Y2=0.73
r223 15 32 106.596 $w=1.6e-07 $l=2.3e-07 $layer=POLY_cond $X=5.32 $Y=1.09
+ $X2=5.32 $Y2=0.86
r224 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.96 $Y=1.99
+ $X2=4.96 $Y2=1.915
r225 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.96 $Y=1.99
+ $X2=4.96 $Y2=2.275
r226 9 15 26.9672 $w=1.5e-07 $l=1.11355e-07 $layer=POLY_cond $X=5.24 $Y=1.165
+ $X2=5.32 $Y2=1.09
r227 9 60 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.24 $Y=1.165
+ $X2=4.745 $Y2=1.165
r228 8 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.84
+ $X2=4.67 $Y2=1.915
r229 7 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=1.42
+ $X2=4.67 $Y2=1.255
r230 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.67 $Y=1.42 $X2=4.67
+ $Y2=1.84
r231 2 42 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=1.845 $X2=4.23 $Y2=2.3
r232 1 38 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.235 $X2=4.225 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_1132_21# 1 2 9 11 14 18 19 21 23 24 27 31
+ 33 37 40
c101 40 0 1.41649e-19 $X=5.81 $Y=0.765
c102 37 0 1.35477e-19 $X=5.795 $Y=0.93
c103 33 0 1.39478e-19 $X=5.817 $Y=0.72
c104 21 0 4.57149e-20 $X=6.335 $Y=0.72
c105 19 0 8.87939e-20 $X=6.06 $Y=1.74
r106 37 41 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=1.095
r107 37 40 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=0.765
r108 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.795
+ $Y=0.93 $X2=5.795 $Y2=0.93
r109 33 36 6.12691 $w=3.93e-07 $l=2.1e-07 $layer=LI1_cond $X=5.817 $Y=0.72
+ $X2=5.817 $Y2=0.93
r110 29 31 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=6.712 $Y=2.105
+ $X2=6.712 $Y2=2.285
r111 25 27 6.70025 $w=2.13e-07 $l=1.25e-07 $layer=LI1_cond $X=6.442 $Y=0.635
+ $X2=6.442 $Y2=0.51
r112 23 29 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.712 $Y2=2.105
r113 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.145 $Y2=2.02
r114 22 33 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=6.015 $Y=0.72
+ $X2=5.817 $Y2=0.72
r115 21 25 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.335 $Y=0.72
+ $X2=6.442 $Y2=0.635
r116 21 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.335 $Y=0.72
+ $X2=6.015 $Y2=0.72
r117 19 42 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.06 $Y=1.74
+ $X2=5.885 $Y2=1.74
r118 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.06
+ $Y=1.74 $X2=6.06 $Y2=1.74
r119 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.06 $Y=1.935
+ $X2=6.145 $Y2=2.02
r120 16 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.06 $Y=1.935
+ $X2=6.06 $Y2=1.74
r121 12 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.905
+ $X2=5.885 $Y2=1.74
r122 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.885 $Y=1.905
+ $X2=5.885 $Y2=2.275
r123 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.575
+ $X2=5.885 $Y2=1.74
r124 11 41 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.885 $Y=1.575
+ $X2=5.885 $Y2=1.095
r125 9 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.735 $Y=0.445
+ $X2=5.735 $Y2=0.765
r126 2 31 600 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_PDIFF $count=1 $X=6.555
+ $Y=2.065 $X2=6.715 $Y2=2.285
r127 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.465 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_1006_47# 1 2 11 13 15 18 21 25 29 31 35
+ 36 38 43 46 47 48 50 51 52 55 58
c158 55 0 1.39478e-19 $X=6.39 $Y=1.095
c159 47 0 1.35477e-19 $X=6.305 $Y=1.185
r160 51 59 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=7.472 $Y=1.16
+ $X2=7.472 $Y2=1.325
r161 51 58 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=7.472 $Y=1.16
+ $X2=7.472 $Y2=0.995
r162 50 52 3.56026 $w=3.48e-07 $l=1e-07 $layer=LI1_cond $X=7.455 $Y=1.15
+ $X2=7.355 $Y2=1.15
r163 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.455
+ $Y=1.16 $X2=7.455 $Y2=1.16
r164 48 52 33.805 $w=2.98e-07 $l=8.8e-07 $layer=LI1_cond $X=6.475 $Y=1.125
+ $X2=7.355 $Y2=1.125
r165 46 56 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.39 $Y=1.23
+ $X2=6.39 $Y2=1.365
r166 46 55 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.39 $Y=1.23
+ $X2=6.39 $Y2=1.095
r167 45 48 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.475 $Y2=1.185
r168 45 47 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.305 $Y2=1.185
r169 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.39
+ $Y=1.23 $X2=6.39 $Y2=1.23
r170 40 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=1.31
+ $X2=5.72 $Y2=1.31
r171 40 47 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.805 $Y=1.31
+ $X2=6.305 $Y2=1.31
r172 37 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=1.395
+ $X2=5.72 $Y2=1.31
r173 37 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.72 $Y=1.395
+ $X2=5.72 $Y2=2.135
r174 35 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=1.31
+ $X2=5.72 $Y2=1.31
r175 35 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.635 $Y=1.31
+ $X2=5.45 $Y2=1.31
r176 31 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.635 $Y=2.3
+ $X2=5.72 $Y2=2.135
r177 31 33 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.635 $Y=2.3
+ $X2=5.225 $Y2=2.3
r178 27 36 22.8143 $w=1.03e-07 $l=2.36715e-07 $layer=LI1_cond $X=5.252 $Y=1.225
+ $X2=5.45 $Y2=1.31
r179 27 29 23.4865 $w=3.93e-07 $l=8.05e-07 $layer=LI1_cond $X=5.252 $Y=1.225
+ $X2=5.252 $Y2=0.42
r180 23 25 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.48 $Y=0.805
+ $X2=6.675 $Y2=0.805
r181 21 59 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.55 $Y=2.065
+ $X2=7.55 $Y2=1.325
r182 18 58 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.51 $Y=0.555
+ $X2=7.51 $Y2=0.995
r183 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.675 $Y=0.73
+ $X2=6.675 $Y2=0.805
r184 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.675 $Y=0.73
+ $X2=6.675 $Y2=0.445
r185 11 56 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=6.48 $Y=2.275
+ $X2=6.48 $Y2=1.365
r186 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.48 $Y=0.88
+ $X2=6.48 $Y2=0.805
r187 7 55 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.48 $Y=0.88
+ $X2=6.48 $Y2=1.095
r188 2 33 600 $w=1.7e-07 $l=3.1603e-07 $layer=licon1_PDIFF $count=1 $X=5.035
+ $Y=2.065 $X2=5.225 $Y2=2.3
r189 1 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.235 $X2=5.165 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%SET_B 5 9 11 13 16 19 23 25 29 30 32 34 35
+ 41 46 47 48 57
c136 47 0 5.67121e-20 $X=6.9 $Y=1.68
c137 29 0 8.40823e-20 $X=9.77 $Y=1.64
c138 23 0 1.13886e-19 $X=9.78 $Y=1.835
c139 9 0 4.57149e-20 $X=7.035 $Y=0.445
c140 5 0 1.54163e-19 $X=6.97 $Y=2.275
r141 46 49 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.845
r142 46 48 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.515
r143 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.9
+ $Y=1.68 $X2=6.9 $Y2=1.68
r144 42 57 4.69647 $w=2.88e-07 $l=9e-08 $layer=LI1_cond $X=9.025 $Y=1.58
+ $X2=9.115 $Y2=1.58
r145 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.025 $Y=1.53
+ $X2=9.025 $Y2=1.53
r146 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.87 $Y=1.53
+ $X2=6.725 $Y2=1.53
r147 34 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.88 $Y=1.53
+ $X2=9.025 $Y2=1.53
r148 34 35 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=8.88 $Y=1.53
+ $X2=6.87 $Y2=1.53
r149 32 47 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=6.725 $Y=1.605
+ $X2=6.9 $Y2=1.605
r150 32 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.725 $Y=1.53
+ $X2=6.725 $Y2=1.53
r151 29 57 36.3227 $w=1.98e-07 $l=6.55e-07 $layer=LI1_cond $X=9.77 $Y=1.625
+ $X2=9.115 $Y2=1.625
r152 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.77
+ $Y=1.64 $X2=9.77 $Y2=1.64
r153 25 30 4.13703 $w=2.9e-07 $l=2e-08 $layer=POLY_cond $X=9.78 $Y=1.62 $X2=9.78
+ $Y2=1.64
r154 25 26 43.9218 $w=2.9e-07 $l=1.45e-07 $layer=POLY_cond $X=9.78 $Y=1.62
+ $X2=9.78 $Y2=1.475
r155 23 30 40.336 $w=2.9e-07 $l=1.95e-07 $layer=POLY_cond $X=9.78 $Y=1.835
+ $X2=9.78 $Y2=1.64
r156 20 23 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=9.535 $Y=1.91
+ $X2=9.78 $Y2=1.91
r157 19 48 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.97 $Y=1.365
+ $X2=6.97 $Y2=1.515
r158 18 19 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=7.002 $Y=1.215
+ $X2=7.002 $Y2=1.365
r159 16 26 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=9.85 $Y=0.445
+ $X2=9.85 $Y2=1.475
r160 11 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.535 $Y=1.985
+ $X2=9.535 $Y2=1.91
r161 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.535 $Y=1.985
+ $X2=9.535 $Y2=2.275
r162 9 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.035 $Y=0.445
+ $X2=7.035 $Y2=1.215
r163 5 49 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.97 $Y=2.275
+ $X2=6.97 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_1781_295# 1 2 9 11 12 15 18 21 22 24 25
+ 28 31 35 37
c103 25 0 9.42889e-20 $X=9.515 $Y=1.27
c104 15 0 1.08286e-19 $X=9.35 $Y=0.445
c105 12 0 1.81319e-19 $X=9.055 $Y=1.55
c106 11 0 1.34058e-19 $X=9.275 $Y=1.55
r107 33 35 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=10.55 $Y=0.42
+ $X2=10.82 $Y2=0.42
r108 31 37 4.27425 $w=2.12e-07 $l=1.12916e-07 $layer=LI1_cond $X=10.82 $Y=1.185
+ $X2=10.755 $Y2=1.27
r109 30 35 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.82 $Y=0.585
+ $X2=10.82 $Y2=0.42
r110 30 31 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=10.82 $Y=0.585
+ $X2=10.82 $Y2=1.185
r111 26 37 4.27425 $w=2.12e-07 $l=1.0015e-07 $layer=LI1_cond $X=10.722 $Y=1.355
+ $X2=10.755 $Y2=1.27
r112 26 28 43.7458 $w=2.43e-07 $l=9.3e-07 $layer=LI1_cond $X=10.722 $Y=1.355
+ $X2=10.722 $Y2=2.285
r113 24 37 2.15711 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=10.6 $Y=1.27
+ $X2=10.755 $Y2=1.27
r114 24 25 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=10.6 $Y=1.27
+ $X2=9.515 $Y2=1.27
r115 22 40 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=9.42 $Y=1.02
+ $X2=9.42 $Y2=1.185
r116 22 39 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=9.42 $Y=1.02
+ $X2=9.42 $Y2=0.855
r117 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.43
+ $Y=1.02 $X2=9.43 $Y2=1.02
r118 19 25 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.4 $Y=1.185
+ $X2=9.515 $Y2=1.27
r119 19 21 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.4 $Y=1.185
+ $X2=9.4 $Y2=1.02
r120 18 40 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.35 $Y=1.475
+ $X2=9.35 $Y2=1.185
r121 15 39 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.35 $Y=0.445
+ $X2=9.35 $Y2=0.855
r122 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.275 $Y=1.55
+ $X2=9.35 $Y2=1.475
r123 11 12 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=9.275 $Y=1.55
+ $X2=9.055 $Y2=1.55
r124 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.98 $Y=1.625
+ $X2=9.055 $Y2=1.55
r125 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=8.98 $Y=1.625
+ $X2=8.98 $Y2=2.275
r126 2 28 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=10.55
+ $Y=2.065 $X2=10.685 $Y2=2.285
r127 1 33 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=10.41
+ $Y=0.235 $X2=10.55 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_1597_329# 1 2 3 10 12 13 17 19 21 23 26
+ 28 30 33 35 36 39 43 47 48 52 56 60 63 64 66 69 73 74 76 80 82
c180 82 0 8.40823e-20 $X=10.342 $Y=1.555
c181 76 0 1.44514e-19 $X=8.905 $Y=1.98
c182 64 0 1.08286e-19 $X=9.855 $Y=0.93
c183 47 0 1.25776e-19 $X=12.84 $Y=1.16
r184 74 83 42.008 $w=4.15e-07 $l=1.35e-07 $layer=POLY_cond $X=10.342 $Y=1.69
+ $X2=10.342 $Y2=1.825
r185 74 82 23.1986 $w=4.15e-07 $l=1.35e-07 $layer=POLY_cond $X=10.342 $Y=1.69
+ $X2=10.342 $Y2=1.555
r186 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.3
+ $Y=1.69 $X2=10.3 $Y2=1.69
r187 71 73 7.26926 $w=3.23e-07 $l=2.05e-07 $layer=LI1_cond $X=10.267 $Y=1.895
+ $X2=10.267 $Y2=1.69
r188 70 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.93 $Y=1.98
+ $X2=9.795 $Y2=1.98
r189 69 71 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=10.105 $Y=1.98
+ $X2=10.267 $Y2=1.895
r190 69 70 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.105 $Y=1.98
+ $X2=9.93 $Y2=1.98
r191 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.395
+ $Y=0.93 $X2=10.395 $Y2=0.93
r192 64 66 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=9.855 $Y=0.93
+ $X2=10.395 $Y2=0.93
r193 63 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.77 $Y=0.845
+ $X2=9.855 $Y2=0.93
r194 62 63 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.77 $Y=0.515
+ $X2=9.77 $Y2=0.845
r195 58 80 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=2.065
+ $X2=9.795 $Y2=1.98
r196 58 60 9.39028 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.795 $Y=2.065
+ $X2=9.795 $Y2=2.285
r197 57 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=1.98
+ $X2=8.905 $Y2=1.98
r198 56 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.66 $Y=1.98
+ $X2=9.795 $Y2=1.98
r199 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.66 $Y=1.98
+ $X2=8.99 $Y2=1.98
r200 52 62 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=9.685 $Y=0.395
+ $X2=9.77 $Y2=0.515
r201 52 54 50.6595 $w=2.38e-07 $l=1.055e-06 $layer=LI1_cond $X=9.685 $Y=0.395
+ $X2=8.63 $Y2=0.395
r202 48 76 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=8.905 $Y=2.292
+ $X2=8.905 $Y2=1.98
r203 48 50 18.9207 $w=3.33e-07 $l=5.5e-07 $layer=LI1_cond $X=8.82 $Y=2.292
+ $X2=8.27 $Y2=2.292
r204 45 46 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.415 $Y=1.16
+ $X2=11.835 $Y2=1.16
r205 41 47 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.84 $Y=1.325
+ $X2=12.84 $Y2=1.16
r206 41 43 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=12.84 $Y=1.325
+ $X2=12.84 $Y2=2.1
r207 37 47 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.84 $Y=0.995
+ $X2=12.84 $Y2=1.16
r208 37 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=12.84 $Y=0.995
+ $X2=12.84 $Y2=0.445
r209 36 46 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.91 $Y=1.16
+ $X2=11.835 $Y2=1.16
r210 35 47 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.765 $Y=1.16
+ $X2=12.84 $Y2=1.16
r211 35 36 149.506 $w=3.3e-07 $l=8.55e-07 $layer=POLY_cond $X=12.765 $Y=1.16
+ $X2=11.91 $Y2=1.16
r212 31 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.835 $Y=1.325
+ $X2=11.835 $Y2=1.16
r213 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.835 $Y=1.325
+ $X2=11.835 $Y2=1.985
r214 28 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.835 $Y=0.995
+ $X2=11.835 $Y2=1.16
r215 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.835 $Y=0.995
+ $X2=11.835 $Y2=0.56
r216 24 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.415 $Y=1.325
+ $X2=11.415 $Y2=1.16
r217 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.415 $Y=1.325
+ $X2=11.415 $Y2=1.985
r218 21 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.415 $Y=0.995
+ $X2=11.415 $Y2=1.16
r219 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.415 $Y=0.995
+ $X2=11.415 $Y2=0.56
r220 20 67 39.452 $w=2.81e-07 $l=2.3e-07 $layer=POLY_cond $X=10.405 $Y=1.16
+ $X2=10.405 $Y2=0.93
r221 19 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.34 $Y=1.16
+ $X2=11.415 $Y2=1.16
r222 19 20 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=11.34 $Y=1.16
+ $X2=10.55 $Y2=1.16
r223 17 83 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=10.475 $Y=2.275
+ $X2=10.475 $Y2=1.825
r224 13 20 27.4241 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=10.405 $Y=1.325
+ $X2=10.405 $Y2=1.16
r225 13 82 47.5758 $w=2.9e-07 $l=2.3e-07 $layer=POLY_cond $X=10.405 $Y=1.325
+ $X2=10.405 $Y2=1.555
r226 10 67 38.716 $w=2.81e-07 $l=1.96914e-07 $layer=POLY_cond $X=10.335 $Y=0.765
+ $X2=10.405 $Y2=0.93
r227 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.335 $Y=0.765
+ $X2=10.335 $Y2=0.445
r228 3 60 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=9.61
+ $Y=2.065 $X2=9.745 $Y2=2.285
r229 2 50 600 $w=1.7e-07 $l=7.745e-07 $layer=licon1_PDIFF $count=1 $X=7.985
+ $Y=1.645 $X2=8.27 $Y2=2.29
r230 1 54 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=0.235 $X2=8.63 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_2501_47# 1 2 7 9 12 14 16 19 23 27 31 34
+ 38
r60 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=13.315 $Y=1.16
+ $X2=13.735 $Y2=1.16
r61 32 37 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=13.26 $Y=1.16
+ $X2=13.315 $Y2=1.16
r62 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.26
+ $Y=1.16 $X2=13.26 $Y2=1.16
r63 29 34 0.63164 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=12.715 $Y=1.16
+ $X2=12.622 $Y2=1.16
r64 29 31 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=12.715 $Y=1.16
+ $X2=13.26 $Y2=1.16
r65 25 34 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.622 $Y=1.325
+ $X2=12.622 $Y2=1.16
r66 25 27 36.57 $w=1.83e-07 $l=6.1e-07 $layer=LI1_cond $X=12.622 $Y=1.325
+ $X2=12.622 $Y2=1.935
r67 21 34 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.622 $Y=0.995
+ $X2=12.622 $Y2=1.16
r68 21 23 33.2727 $w=1.83e-07 $l=5.55e-07 $layer=LI1_cond $X=12.622 $Y=0.995
+ $X2=12.622 $Y2=0.44
r69 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.735 $Y=1.325
+ $X2=13.735 $Y2=1.16
r70 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.735 $Y=1.325
+ $X2=13.735 $Y2=1.985
r71 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.735 $Y=0.995
+ $X2=13.735 $Y2=1.16
r72 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.735 $Y=0.995
+ $X2=13.735 $Y2=0.56
r73 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.315 $Y=1.325
+ $X2=13.315 $Y2=1.16
r74 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.315 $Y=1.325
+ $X2=13.315 $Y2=1.985
r75 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.315 $Y=0.995
+ $X2=13.315 $Y2=1.16
r76 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.315 $Y=0.995
+ $X2=13.315 $Y2=0.56
r77 2 27 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=12.505
+ $Y=1.78 $X2=12.63 $Y2=1.935
r78 1 23 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=12.505
+ $Y=0.235 $X2=12.63 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_27_369# 1 2 9 12 13 15 18
r41 13 15 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=1.185 $Y=2.36
+ $X2=1.94 $Y2=2.36
r42 12 13 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.1 $Y=2.255
+ $X2=1.185 $Y2=2.36
r43 11 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.1 $Y=2.075 $X2=1.1
+ $Y2=2.255
r44 10 18 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.96
+ $X2=0.215 $Y2=1.96
r45 9 11 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.015 $Y=1.96
+ $X2=1.1 $Y2=2.075
r46 9 10 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=1.96
+ $X2=0.345 $Y2=1.96
r47 2 15 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.845 $X2=1.94 $Y2=2.34
r48 1 18 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48 54
+ 58 62 68 74 76 78 83 84 86 87 89 90 91 93 98 106 111 129 133 138 144 147 150
+ 153 158 164 166 169 173
c219 173 0 1.14377e-19 $X=14.03 $Y=2.72
c220 44 0 1.20946e-19 $X=3.81 $Y=2.36
c221 40 0 3.22446e-20 $X=2.87 $Y=2.34
r222 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r223 169 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r224 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r225 162 164 15.2496 $w=6.78e-07 $l=4.25e-07 $layer=LI1_cond $X=7.59 $Y=2.465
+ $X2=8.015 $Y2=2.465
r226 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r227 160 162 6.42013 $w=6.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.225 $Y=2.465
+ $X2=7.59 $Y2=2.465
r228 157 163 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r229 156 160 1.67099 $w=6.78e-07 $l=9.5e-08 $layer=LI1_cond $X=7.13 $Y=2.465
+ $X2=7.225 $Y2=2.465
r230 156 158 9.00537 $w=6.78e-07 $l=7e-08 $layer=LI1_cond $X=7.13 $Y=2.465
+ $X2=7.06 $Y2=2.465
r231 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r232 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r233 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r234 150 151 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r235 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r236 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r237 142 173 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.03 $Y2=2.72
r238 142 170 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=13.11 $Y2=2.72
r239 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r240 139 169 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=13.24 $Y=2.72
+ $X2=13.062 $Y2=2.72
r241 139 141 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=13.24 $Y=2.72
+ $X2=13.57 $Y2=2.72
r242 138 172 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=13.91 $Y=2.72
+ $X2=14.085 $Y2=2.72
r243 138 141 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.91 $Y=2.72
+ $X2=13.57 $Y2=2.72
r244 137 170 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r245 137 167 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r246 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r247 134 166 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.315 $Y=2.72
+ $X2=12.17 $Y2=2.72
r248 134 136 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.315 $Y=2.72
+ $X2=12.65 $Y2=2.72
r249 133 169 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=12.885 $Y=2.72
+ $X2=13.062 $Y2=2.72
r250 133 136 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=12.885 $Y=2.72
+ $X2=12.65 $Y2=2.72
r251 132 167 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r252 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r253 129 166 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=12.17 $Y2=2.72
r254 129 131 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=11.73 $Y2=2.72
r255 128 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r256 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r257 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r258 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r259 122 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r260 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r261 119 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r262 119 163 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r263 118 121 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r264 118 164 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.015 $Y2=2.72
r265 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r266 115 154 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r267 115 151 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r268 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r269 112 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=3.81 $Y2=2.72
r270 112 114 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=5.75 $Y2=2.72
r271 111 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=2.72
+ $X2=6.165 $Y2=2.72
r272 111 114 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6 $Y=2.72
+ $X2=5.75 $Y2=2.72
r273 110 151 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r274 110 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r275 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r276 107 147 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.1 $Y=2.72
+ $X2=2.902 $Y2=2.72
r277 107 109 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.1 $Y=2.72
+ $X2=3.45 $Y2=2.72
r278 106 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=2.72
+ $X2=3.81 $Y2=2.72
r279 106 109 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.645 $Y=2.72
+ $X2=3.45 $Y2=2.72
r280 105 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r281 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r282 102 105 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r283 102 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r284 101 104 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r285 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r286 99 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r287 99 101 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r288 98 147 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.902 $Y2=2.72
r289 98 104 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.53 $Y2=2.72
r290 93 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r291 93 95 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r292 91 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r293 91 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r294 89 127 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.08 $Y=2.72
+ $X2=10.81 $Y2=2.72
r295 89 90 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.08 $Y=2.72
+ $X2=11.185 $Y2=2.72
r296 88 131 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=11.29 $Y=2.72
+ $X2=11.73 $Y2=2.72
r297 88 90 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.29 $Y=2.72
+ $X2=11.185 $Y2=2.72
r298 86 124 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=10.1 $Y=2.72
+ $X2=9.89 $Y2=2.72
r299 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.1 $Y=2.72
+ $X2=10.265 $Y2=2.72
r300 85 127 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.43 $Y=2.72
+ $X2=10.81 $Y2=2.72
r301 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.43 $Y=2.72
+ $X2=10.265 $Y2=2.72
r302 83 121 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.16 $Y=2.72
+ $X2=8.97 $Y2=2.72
r303 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=2.72
+ $X2=9.325 $Y2=2.72
r304 82 124 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.89 $Y2=2.72
r305 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.325 $Y2=2.72
r306 78 81 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=14.042 $Y=1.66
+ $X2=14.042 $Y2=2.34
r307 76 172 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=14.042
+ $Y=2.635 $X2=14.085 $Y2=2.72
r308 76 81 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=14.042 $Y=2.635
+ $X2=14.042 $Y2=2.34
r309 72 169 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=13.062 $Y=2.635
+ $X2=13.062 $Y2=2.72
r310 72 74 22.7242 $w=3.53e-07 $l=7e-07 $layer=LI1_cond $X=13.062 $Y=2.635
+ $X2=13.062 $Y2=1.935
r311 68 71 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=12.17 $Y=1.66
+ $X2=12.17 $Y2=2.34
r312 66 166 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.17 $Y=2.635
+ $X2=12.17 $Y2=2.72
r313 66 71 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=12.17 $Y=2.635
+ $X2=12.17 $Y2=2.34
r314 62 65 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=11.185 $Y=1.66
+ $X2=11.185 $Y2=2.34
r315 60 90 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=2.635
+ $X2=11.185 $Y2=2.72
r316 60 65 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=11.185 $Y=2.635
+ $X2=11.185 $Y2=2.34
r317 56 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=2.635
+ $X2=10.265 $Y2=2.72
r318 56 58 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.265 $Y=2.635
+ $X2=10.265 $Y2=2.34
r319 52 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=2.635
+ $X2=9.325 $Y2=2.72
r320 52 54 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.325 $Y=2.635
+ $X2=9.325 $Y2=2.36
r321 51 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=6.165 $Y2=2.72
r322 51 158 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=7.06 $Y2=2.72
r323 46 153 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.165 $Y=2.635
+ $X2=6.165 $Y2=2.72
r324 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.165 $Y=2.635
+ $X2=6.165 $Y2=2.36
r325 42 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=2.635
+ $X2=3.81 $Y2=2.72
r326 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.81 $Y=2.635
+ $X2=3.81 $Y2=2.36
r327 38 147 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.902 $Y=2.635
+ $X2=2.902 $Y2=2.72
r328 38 40 8.60685 $w=3.93e-07 $l=2.95e-07 $layer=LI1_cond $X=2.902 $Y=2.635
+ $X2=2.902 $Y2=2.34
r329 34 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r330 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.36
r331 11 81 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=13.81
+ $Y=1.485 $X2=13.995 $Y2=2.34
r332 11 78 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=13.81
+ $Y=1.485 $X2=13.995 $Y2=1.66
r333 10 74 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=12.915
+ $Y=1.78 $X2=13.1 $Y2=1.935
r334 9 71 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=11.91
+ $Y=1.485 $X2=12.11 $Y2=2.34
r335 9 68 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=11.91
+ $Y=1.485 $X2=12.11 $Y2=1.66
r336 8 65 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=11.08
+ $Y=1.485 $X2=11.205 $Y2=2.34
r337 8 62 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=11.08
+ $Y=1.485 $X2=11.205 $Y2=1.66
r338 7 58 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=2.065 $X2=10.265 $Y2=2.34
r339 6 54 600 $w=1.7e-07 $l=4.08258e-07 $layer=licon1_PDIFF $count=1 $X=9.055
+ $Y=2.065 $X2=9.325 $Y2=2.36
r340 5 160 600 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=2.065 $X2=7.225 $Y2=2.36
r341 4 48 600 $w=1.7e-07 $l=3.84057e-07 $layer=licon1_PDIFF $count=1 $X=5.96
+ $Y=2.065 $X2=6.165 $Y2=2.36
r342 3 44 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.845 $X2=3.81 $Y2=2.36
r343 2 40 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=1.845 $X2=2.87 $Y2=2.34
r344 1 36 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%A_181_47# 1 2 3 4 13 19 21 23 26 30 34 35
+ 36 39 42
c124 42 0 3.35674e-20 $X=4.885 $Y=1.53
c125 34 0 1.07774e-19 $X=4.695 $Y=0.92
c126 21 0 1.18775e-19 $X=4.777 $Y=1.615
c127 19 0 1.78833e-19 $X=4.745 $Y=0.42
r128 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.885 $Y=1.53
+ $X2=4.885 $Y2=1.53
r129 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.53
+ $X2=1.61 $Y2=1.53
r130 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.53
+ $X2=1.61 $Y2=1.53
r131 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.74 $Y=1.53
+ $X2=4.885 $Y2=1.53
r132 35 36 3.6943 $w=1.4e-07 $l=2.985e-06 $layer=MET1_cond $X=4.74 $Y=1.53
+ $X2=1.755 $Y2=1.53
r133 33 39 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.6 $Y=0.72 $X2=1.6
+ $Y2=1.53
r134 31 39 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.6 $Y=1.845
+ $X2=1.6 $Y2=1.53
r135 30 31 2.10789 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=1.6 $Y=1.965 $X2=1.6
+ $Y2=1.845
r136 28 30 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=1.52 $Y=1.965 $X2=1.6
+ $Y2=1.965
r137 26 43 5.45986 $w=2.62e-07 $l=9.31128e-08 $layer=LI1_cond $X=4.8 $Y=1.445
+ $X2=4.817 $Y2=1.53
r138 26 34 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.8 $Y=1.445
+ $X2=4.8 $Y2=0.92
r139 21 43 4.23541 $w=2.62e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.777 $Y=1.615
+ $X2=4.817 $Y2=1.53
r140 21 23 35.0855 $w=2.23e-07 $l=6.85e-07 $layer=LI1_cond $X=4.777 $Y=1.615
+ $X2=4.777 $Y2=2.3
r141 17 34 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=4.695 $Y=0.73
+ $X2=4.695 $Y2=0.92
r142 17 19 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=4.695 $Y=0.73
+ $X2=4.695 $Y2=0.42
r143 13 33 3.63177 $w=5.51e-07 $l=3.43511e-07 $layer=LI1_cond $X=1.495 $Y=0.425
+ $X2=1.6 $Y2=0.72
r144 13 15 15.4224 $w=3.38e-07 $l=4.55e-07 $layer=LI1_cond $X=1.495 $Y=0.425
+ $X2=1.04 $Y2=0.425
r145 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=2.065 $X2=4.75 $Y2=2.3
r146 3 28 600 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=1.845 $X2=1.52 $Y2=1.97
r147 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.62
+ $Y=0.235 $X2=4.745 $Y2=0.42
r148 1 15 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=0.905
+ $Y=0.235 $X2=1.04 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%Q_N 1 2 7 8 9 10 11 12 20
r19 12 37 3.64697 $w=3.93e-07 $l=1.25e-07 $layer=LI1_cond $X=11.657 $Y=2.21
+ $X2=11.657 $Y2=2.335
r20 11 12 9.91976 $w=3.93e-07 $l=3.4e-07 $layer=LI1_cond $X=11.657 $Y=1.87
+ $X2=11.657 $Y2=2.21
r21 11 31 6.27279 $w=3.93e-07 $l=2.15e-07 $layer=LI1_cond $X=11.657 $Y=1.87
+ $X2=11.657 $Y2=1.655
r22 10 31 3.64697 $w=3.93e-07 $l=1.25e-07 $layer=LI1_cond $X=11.657 $Y=1.53
+ $X2=11.657 $Y2=1.655
r23 9 10 9.91976 $w=3.93e-07 $l=3.4e-07 $layer=LI1_cond $X=11.657 $Y=1.19
+ $X2=11.657 $Y2=1.53
r24 8 9 9.91976 $w=3.93e-07 $l=3.4e-07 $layer=LI1_cond $X=11.657 $Y=0.85
+ $X2=11.657 $Y2=1.19
r25 7 8 9.91976 $w=3.93e-07 $l=3.4e-07 $layer=LI1_cond $X=11.657 $Y=0.51
+ $X2=11.657 $Y2=0.85
r26 7 20 3.79285 $w=3.93e-07 $l=1.3e-07 $layer=LI1_cond $X=11.657 $Y=0.51
+ $X2=11.657 $Y2=0.38
r27 2 37 400 $w=1.7e-07 $l=9.15014e-07 $layer=licon1_PDIFF $count=1 $X=11.49
+ $Y=1.485 $X2=11.625 $Y2=2.335
r28 2 31 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=11.49
+ $Y=1.485 $X2=11.625 $Y2=1.655
r29 1 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=11.49
+ $Y=0.235 $X2=11.625 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%Q 1 2 7 8 9 10 11 12 23 30 46
c22 30 0 1.25776e-19 $X=13.63 $Y=0.85
r23 46 47 2.39662 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=13.575 $Y=1.53
+ $X2=13.575 $Y2=1.495
r24 30 44 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=13.627 $Y=0.85
+ $X2=13.627 $Y2=0.825
r25 12 39 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=13.575 $Y=2.21
+ $X2=13.575 $Y2=1.945
r26 11 39 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=13.575 $Y=1.87
+ $X2=13.575 $Y2=1.945
r27 11 35 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=13.575 $Y=1.87
+ $X2=13.575 $Y2=1.66
r28 10 35 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=13.575 $Y=1.555
+ $X2=13.575 $Y2=1.66
r29 10 46 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=13.575 $Y=1.555
+ $X2=13.575 $Y2=1.53
r30 10 47 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=13.627 $Y=1.47
+ $X2=13.627 $Y2=1.495
r31 9 10 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=13.627 $Y=1.19
+ $X2=13.627 $Y2=1.47
r32 8 44 2.22201 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=13.575 $Y=0.795
+ $X2=13.575 $Y2=0.825
r33 8 21 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=13.575 $Y=0.795
+ $X2=13.575 $Y2=0.66
r34 8 9 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=13.627 $Y=0.88
+ $X2=13.627 $Y2=1.19
r35 8 30 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=13.627 $Y=0.88
+ $X2=13.627 $Y2=0.85
r36 7 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=13.575 $Y=0.51
+ $X2=13.575 $Y2=0.66
r37 7 23 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=13.575 $Y=0.51
+ $X2=13.575 $Y2=0.44
r38 2 39 300 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_PDIFF $count=2 $X=13.39
+ $Y=1.485 $X2=13.525 $Y2=1.945
r39 1 23 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=13.39
+ $Y=0.235 $X2=13.525 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_2%VGND 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48 52
+ 56 58 61 63 66 67 69 70 72 73 74 80 84 89 109 113 118 124 131 134 138 145 149
+ 151 154 158
c204 158 0 2.71124e-20 $X=14.03 $Y=0
c205 89 0 2.79334e-19 $X=5.665 $Y=0
c206 40 0 4.13602e-20 $X=2.865 $Y=0.38
r207 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r208 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r209 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r210 147 149 11.5282 $w=8.88e-07 $l=1.15e-07 $layer=LI1_cond $X=7.59 $Y=0.36
+ $X2=7.705 $Y2=0.36
r211 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r212 144 147 4.72921 $w=8.88e-07 $l=3.45e-07 $layer=LI1_cond $X=7.245 $Y=0.36
+ $X2=7.59 $Y2=0.36
r213 144 145 17.1485 $w=8.88e-07 $l=5.25e-07 $layer=LI1_cond $X=7.245 $Y=0.36
+ $X2=6.72 $Y2=0.36
r214 138 141 9.0902 $w=4.98e-07 $l=3.8e-07 $layer=LI1_cond $X=5.915 $Y=0
+ $X2=5.915 $Y2=0.38
r215 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r216 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r217 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r218 124 129 8.24843 $w=6.36e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=0
+ $X2=0.35 $Y2=0.43
r219 124 127 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r220 122 158 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r221 122 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=13.11 $Y2=0
r222 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r223 119 154 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=13.24 $Y=0
+ $X2=13.062 $Y2=0
r224 119 121 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=13.24 $Y=0
+ $X2=13.57 $Y2=0
r225 118 157 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=13.91 $Y=0
+ $X2=14.085 $Y2=0
r226 118 121 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.91 $Y=0
+ $X2=13.57 $Y2=0
r227 117 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r228 117 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r229 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r230 114 151 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.315 $Y=0
+ $X2=12.17 $Y2=0
r231 114 116 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.315 $Y=0
+ $X2=12.65 $Y2=0
r232 113 154 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=12.885 $Y=0
+ $X2=13.062 $Y2=0
r233 113 116 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=12.885 $Y=0
+ $X2=12.65 $Y2=0
r234 112 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r235 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r236 109 151 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.025 $Y=0
+ $X2=12.17 $Y2=0
r237 109 111 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=0
+ $X2=11.73 $Y2=0
r238 108 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r239 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r240 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r241 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r242 102 105 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.89 $Y2=0
r243 102 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r244 101 104 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=9.89 $Y2=0
r245 101 149 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=7.705 $Y2=0
r246 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r247 98 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r248 98 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=5.75 $Y2=0
r249 97 145 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.72
+ $Y2=0
r250 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r251 95 138 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.165 $Y=0
+ $X2=5.915 $Y2=0
r252 95 97 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.165 $Y=0
+ $X2=6.67 $Y2=0
r253 93 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r254 93 135 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=3.91 $Y2=0
r255 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r256 90 134 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=3.79
+ $Y2=0
r257 90 92 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.94 $Y=0 $X2=5.29
+ $Y2=0
r258 89 138 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=5.665 $Y=0
+ $X2=5.915 $Y2=0
r259 89 92 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.665 $Y=0
+ $X2=5.29 $Y2=0
r260 88 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r261 88 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.99 $Y2=0
r262 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r263 85 131 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.9
+ $Y2=0
r264 85 87 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.45
+ $Y2=0
r265 84 134 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.79
+ $Y2=0
r266 84 87 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.45
+ $Y2=0
r267 83 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r268 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r269 80 131 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.9
+ $Y2=0
r270 80 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.53
+ $Y2=0
r271 79 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r272 79 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r273 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r274 76 124 8.69404 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=0.7 $Y=0 $X2=0.35
+ $Y2=0
r275 76 78 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.7 $Y=0 $X2=1.61
+ $Y2=0
r276 74 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r277 74 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r278 72 107 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=10.81 $Y2=0
r279 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=11.205 $Y2=0
r280 71 111 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=11.29 $Y=0
+ $X2=11.73 $Y2=0
r281 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.29 $Y=0
+ $X2=11.205 $Y2=0
r282 69 104 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.035 $Y=0
+ $X2=9.89 $Y2=0
r283 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.035 $Y=0
+ $X2=10.16 $Y2=0
r284 68 107 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=10.285 $Y=0
+ $X2=10.81 $Y2=0
r285 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.285 $Y=0
+ $X2=10.16 $Y2=0
r286 66 78 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.61
+ $Y2=0
r287 66 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.965
+ $Y2=0
r288 65 82 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.53
+ $Y2=0
r289 65 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.965
+ $Y2=0
r290 61 157 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=14.042
+ $Y=0.085 $X2=14.085 $Y2=0
r291 61 63 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=14.042 $Y=0.085
+ $X2=14.042 $Y2=0.38
r292 58 154 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=13.062 $Y=0.085
+ $X2=13.062 $Y2=0
r293 58 60 9.4507 $w=3.55e-07 $l=2.75e-07 $layer=LI1_cond $X=13.062 $Y=0.085
+ $X2=13.062 $Y2=0.36
r294 54 151 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.17 $Y=0.085
+ $X2=12.17 $Y2=0
r295 54 56 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=12.17 $Y=0.085
+ $X2=12.17 $Y2=0.38
r296 50 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=0.085
+ $X2=11.205 $Y2=0
r297 50 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.205 $Y=0.085
+ $X2=11.205 $Y2=0.38
r298 46 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.16 $Y=0.085
+ $X2=10.16 $Y2=0
r299 46 48 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=10.16 $Y=0.085
+ $X2=10.16 $Y2=0.36
r300 42 134 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r301 42 44 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.36
r302 38 131 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0
r303 38 40 8.49927 $w=3.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.9 $Y=0.085
+ $X2=2.9 $Y2=0.38
r304 34 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=0.085
+ $X2=1.965 $Y2=0
r305 34 36 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.965 $Y=0.085
+ $X2=1.965 $Y2=0.38
r306 11 63 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=13.81
+ $Y=0.235 $X2=13.995 $Y2=0.38
r307 10 60 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=12.915
+ $Y=0.235 $X2=13.075 $Y2=0.36
r308 9 56 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=11.91
+ $Y=0.235 $X2=12.11 $Y2=0.38
r309 8 52 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=11.08
+ $Y=0.235 $X2=11.205 $Y2=0.38
r310 7 48 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=9.925
+ $Y=0.235 $X2=10.12 $Y2=0.36
r311 6 144 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.11
+ $Y=0.235 $X2=7.245 $Y2=0.36
r312 5 141 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.81
+ $Y=0.235 $X2=5.945 $Y2=0.38
r313 4 44 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.235 $X2=3.805 $Y2=0.36
r314 3 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.235 $X2=2.865 $Y2=0.38
r315 2 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.235 $X2=1.925 $Y2=0.38
r316 1 129 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends


* NGSPICE file created from sky130_fd_sc_hd__o21ba_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VGND A2 a_448_47# VNB nshort w=650000u l=150000u
+  ad=3.76e+11p pd=3.81e+06u as=3.8675e+11p ps=3.79e+06u
M1001 a_544_297# A2 a_79_199# VPB phighvt w=1e+06u l=150000u
+  ad=2.1e+11p pd=2.42e+06u as=3.3e+11p ps=2.66e+06u
M1002 a_222_93# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1003 a_222_93# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=9.515e+11p ps=7.99e+06u
M1004 a_79_199# a_222_93# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_79_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1006 VPWR a_79_199# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1007 VPWR A1 a_544_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_448_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_448_47# a_222_93# a_79_199# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
.ends


* File: sky130_fd_sc_hd__bufinv_8.pxi.spice
* Created: Thu Aug 27 14:10:34 2020
* 
x_PM_SKY130_FD_SC_HD__BUFINV_8%A N_A_c_127_n N_A_M1023_g N_A_M1017_g A
+ N_A_c_129_n PM_SKY130_FD_SC_HD__BUFINV_8%A
x_PM_SKY130_FD_SC_HD__BUFINV_8%A_109_47# N_A_109_47#_M1023_d N_A_109_47#_M1017_d
+ N_A_109_47#_M1002_g N_A_109_47#_M1001_g N_A_109_47#_M1003_g
+ N_A_109_47#_M1019_g N_A_109_47#_M1005_g N_A_109_47#_M1020_g
+ N_A_109_47#_c_157_n N_A_109_47#_c_167_n N_A_109_47#_c_158_n
+ N_A_109_47#_c_159_n N_A_109_47#_c_160_n N_A_109_47#_c_168_n
+ N_A_109_47#_c_161_n N_A_109_47#_c_162_n N_A_109_47#_c_163_n
+ PM_SKY130_FD_SC_HD__BUFINV_8%A_109_47#
x_PM_SKY130_FD_SC_HD__BUFINV_8%A_215_47# N_A_215_47#_M1002_d N_A_215_47#_M1003_d
+ N_A_215_47#_M1001_s N_A_215_47#_M1019_s N_A_215_47#_M1004_g
+ N_A_215_47#_M1000_g N_A_215_47#_M1006_g N_A_215_47#_M1007_g
+ N_A_215_47#_M1009_g N_A_215_47#_M1008_g N_A_215_47#_M1011_g
+ N_A_215_47#_M1010_g N_A_215_47#_M1012_g N_A_215_47#_M1014_g
+ N_A_215_47#_M1013_g N_A_215_47#_M1015_g N_A_215_47#_M1016_g
+ N_A_215_47#_M1021_g N_A_215_47#_M1018_g N_A_215_47#_M1022_g
+ N_A_215_47#_c_261_n N_A_215_47#_c_278_n N_A_215_47#_c_262_n
+ N_A_215_47#_c_263_n N_A_215_47#_c_279_n N_A_215_47#_c_280_n
+ N_A_215_47#_c_306_n N_A_215_47#_c_309_n N_A_215_47#_c_264_n
+ N_A_215_47#_c_265_n N_A_215_47#_c_266_n N_A_215_47#_c_267_n
+ N_A_215_47#_c_282_n N_A_215_47#_c_268_n N_A_215_47#_c_269_n
+ PM_SKY130_FD_SC_HD__BUFINV_8%A_215_47#
x_PM_SKY130_FD_SC_HD__BUFINV_8%VPWR N_VPWR_M1017_s N_VPWR_M1001_d N_VPWR_M1020_d
+ N_VPWR_M1007_s N_VPWR_M1010_s N_VPWR_M1015_s N_VPWR_M1022_s N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n
+ N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n
+ N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n
+ N_VPWR_c_507_n VPWR N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_490_n
+ N_VPWR_c_511_n N_VPWR_c_512_n PM_SKY130_FD_SC_HD__BUFINV_8%VPWR
x_PM_SKY130_FD_SC_HD__BUFINV_8%Y N_Y_M1004_s N_Y_M1009_s N_Y_M1012_s N_Y_M1016_s
+ N_Y_M1000_d N_Y_M1008_d N_Y_M1014_d N_Y_M1021_d N_Y_c_604_n N_Y_c_605_n
+ N_Y_c_585_n N_Y_c_586_n N_Y_c_594_n N_Y_c_595_n N_Y_c_632_n N_Y_c_636_n
+ N_Y_c_587_n N_Y_c_596_n N_Y_c_648_n N_Y_c_652_n N_Y_c_588_n N_Y_c_597_n
+ N_Y_c_664_n N_Y_c_667_n N_Y_c_589_n N_Y_c_598_n N_Y_c_590_n N_Y_c_599_n
+ N_Y_c_591_n N_Y_c_600_n N_Y_c_592_n N_Y_c_601_n Y Y
+ PM_SKY130_FD_SC_HD__BUFINV_8%Y
x_PM_SKY130_FD_SC_HD__BUFINV_8%VGND N_VGND_M1023_s N_VGND_M1002_s N_VGND_M1005_s
+ N_VGND_M1006_d N_VGND_M1011_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_c_753_n
+ N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n N_VGND_c_763_n
+ N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n N_VGND_c_767_n N_VGND_c_768_n
+ N_VGND_c_769_n VGND N_VGND_c_770_n N_VGND_c_771_n N_VGND_c_772_n
+ N_VGND_c_773_n N_VGND_c_774_n PM_SKY130_FD_SC_HD__BUFINV_8%VGND
cc_1 VNB N_A_c_127_n 0.0247926f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A 0.00900655f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_129_n 0.0437109f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_109_47#_M1002_g 0.0216102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_109_47#_M1001_g 5.49071e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_109_47#_M1003_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_109_47#_M1019_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_109_47#_M1005_g 0.0175122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_109_47#_M1020_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_109_47#_c_157_n 0.00452528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_109_47#_c_158_n 0.00444855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_109_47#_c_159_n 0.0210275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_109_47#_c_160_n 0.00344329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_109_47#_c_161_n 8.10809e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_109_47#_c_162_n 0.00236261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_109_47#_c_163_n 0.0499058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_215_47#_M1004_g 0.0176384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_215_47#_M1000_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_215_47#_M1006_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_215_47#_M1007_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_215_47#_M1009_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_215_47#_M1008_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_215_47#_M1011_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_215_47#_M1010_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_215_47#_M1012_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_215_47#_M1014_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_215_47#_M1013_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_215_47#_M1015_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_215_47#_M1016_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_215_47#_M1021_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_215_47#_M1018_g 0.0211059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_215_47#_M1022_g 5.13413e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_215_47#_c_261_n 0.00451034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_215_47#_c_262_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_215_47#_c_263_n 0.004399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_215_47#_c_264_n 0.00354558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_215_47#_c_265_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_215_47#_c_266_n 0.00682104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_215_47#_c_267_n 0.00345692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_215_47#_c_268_n 0.0013705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_215_47#_c_269_n 0.12942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_490_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_585_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_586_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_587_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_588_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_Y_c_589_n 0.0190968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_Y_c_590_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_Y_c_591_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_592_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB Y 0.0245101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_753_n 0.0110515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_754_n 0.00654843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_755_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_756_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_757_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_758_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_759_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_760_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_761_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_762_n 0.0168651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_763_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_764_n 0.0174747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_765_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_766_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_767_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_768_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_769_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_770_n 0.0309534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_771_n 0.0175311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_772_n 0.328612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_773_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_774_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_A_M1017_g 0.0284139f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_75 VPB N_A_c_129_n 0.0126558f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_76 VPB N_A_109_47#_M1001_g 0.0240397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_109_47#_M1019_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_109_47#_M1020_g 0.0194268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_109_47#_c_167_n 0.00700329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_109_47#_c_168_n 0.00146952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_109_47#_c_161_n 0.00508712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_215_47#_M1000_g 0.0196632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_215_47#_M1007_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_215_47#_M1008_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_215_47#_M1010_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_215_47#_M1014_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_215_47#_M1015_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_215_47#_M1021_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_215_47#_M1022_g 0.0234522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_215_47#_c_278_n 0.00784989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_215_47#_c_279_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_215_47#_c_280_n 0.00447011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_215_47#_c_265_n 0.00301948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_215_47#_c_282_n 0.00360324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_491_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_492_n 0.00753549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_493_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_494_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_495_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_496_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_497_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_498_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_499_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_500_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_501_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_502_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_503_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_504_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_505_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_506_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_507_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_508_n 0.0313815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_509_n 0.0191681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_490_n 0.0705489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_511_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_512_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_Y_c_594_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_595_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_596_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_Y_c_597_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_Y_c_598_n 0.00454525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_Y_c_599_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_Y_c_600_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_Y_c_601_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB Y 0.00886484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB Y 0.0249431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 N_A_c_127_n N_A_109_47#_c_157_n 0.00551285f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_M1017_g N_A_109_47#_c_167_n 0.00853007f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_c_127_n N_A_109_47#_c_158_n 0.0064171f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_127_n N_A_109_47#_c_160_n 0.00300034f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_M1017_g N_A_109_47#_c_168_n 0.00258868f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_c_129_n N_A_109_47#_c_161_n 0.00742031f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_133 A N_A_109_47#_c_162_n 0.0170591f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_c_129_n N_A_109_47#_c_162_n 0.00521701f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_127_n N_A_215_47#_c_263_n 3.65437e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_M1017_g N_VPWR_c_492_n 0.0053541f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_137 A N_VPWR_c_492_n 0.0136987f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_c_129_n N_VPWR_c_492_n 0.00415776f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_M1017_g N_VPWR_c_508_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1017_g N_VPWR_c_490_n 0.0117818f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_c_127_n N_VGND_c_754_n 0.00482486f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_142 A N_VGND_c_754_n 0.0136981f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_c_129_n N_VGND_c_754_n 0.00431355f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_c_127_n N_VGND_c_770_n 0.00541562f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_127_n N_VGND_c_772_n 0.011782f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_109_47#_M1005_g N_A_215_47#_M1004_g 0.021435f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_147 N_A_109_47#_M1020_g N_A_215_47#_M1000_g 0.021435f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_109_47#_M1002_g N_A_215_47#_c_261_n 0.00636826f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_149 N_A_109_47#_M1003_g N_A_215_47#_c_261_n 5.23702e-19 $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_150 N_A_109_47#_c_157_n N_A_215_47#_c_261_n 0.0365376f $X=0.68 $Y=0.4 $X2=0
+ $Y2=0
cc_151 N_A_109_47#_M1001_g N_A_215_47#_c_278_n 0.0102729f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_109_47#_M1019_g N_A_215_47#_c_278_n 6.98608e-19 $X=1.83 $Y=1.985
+ $X2=0 $Y2=0
cc_153 N_A_109_47#_c_168_n N_A_215_47#_c_278_n 0.0653749f $X=0.68 $Y=1.63 $X2=0
+ $Y2=0
cc_154 N_A_109_47#_M1002_g N_A_215_47#_c_262_n 0.00850187f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_155 N_A_109_47#_M1003_g N_A_215_47#_c_262_n 0.00850187f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_156 N_A_109_47#_c_159_n N_A_215_47#_c_262_n 0.0596152f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A_109_47#_c_163_n N_A_215_47#_c_262_n 0.00205431f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_109_47#_M1002_g N_A_215_47#_c_263_n 0.00126794f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_159 N_A_109_47#_c_157_n N_A_215_47#_c_263_n 0.0138613f $X=0.68 $Y=0.4 $X2=0
+ $Y2=0
cc_160 N_A_109_47#_c_159_n N_A_215_47#_c_263_n 0.0278128f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_109_47#_M1001_g N_A_215_47#_c_279_n 0.0107189f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_109_47#_M1019_g N_A_215_47#_c_279_n 0.0107189f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_109_47#_c_159_n N_A_215_47#_c_279_n 0.0596157f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_109_47#_c_163_n N_A_215_47#_c_279_n 0.00198252f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_109_47#_M1001_g N_A_215_47#_c_280_n 0.00168781f $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_166 N_A_109_47#_c_159_n N_A_215_47#_c_280_n 0.0279329f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_109_47#_c_161_n N_A_215_47#_c_280_n 0.0134952f $X=0.68 $Y=1.545 $X2=0
+ $Y2=0
cc_168 N_A_109_47#_M1002_g N_A_215_47#_c_306_n 5.24491e-19 $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_169 N_A_109_47#_M1003_g N_A_215_47#_c_306_n 0.00647394f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_170 N_A_109_47#_M1005_g N_A_215_47#_c_306_n 0.00647394f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_171 N_A_109_47#_M1001_g N_A_215_47#_c_309_n 6.99397e-19 $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_172 N_A_109_47#_M1019_g N_A_215_47#_c_309_n 0.0103785f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_109_47#_M1020_g N_A_215_47#_c_309_n 0.0103785f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_109_47#_M1005_g N_A_215_47#_c_264_n 0.00412488f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_175 N_A_109_47#_c_163_n N_A_215_47#_c_265_n 0.00407173f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_A_109_47#_M1003_g N_A_215_47#_c_267_n 0.00123754f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_177 N_A_109_47#_M1005_g N_A_215_47#_c_267_n 0.0107176f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_178 N_A_109_47#_c_163_n N_A_215_47#_c_267_n 0.00205431f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_109_47#_M1019_g N_A_215_47#_c_282_n 0.00139111f $X=1.83 $Y=1.985
+ $X2=0 $Y2=0
cc_180 N_A_109_47#_M1020_g N_A_215_47#_c_282_n 0.0131306f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_109_47#_c_163_n N_A_215_47#_c_282_n 0.00198252f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A_109_47#_c_159_n N_A_215_47#_c_268_n 0.0176501f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_183 N_A_109_47#_c_163_n N_A_215_47#_c_268_n 0.00200384f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_109_47#_c_163_n N_A_215_47#_c_269_n 0.021435f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_109_47#_c_161_n N_VPWR_c_492_n 0.00318841f $X=0.68 $Y=1.545 $X2=0
+ $Y2=0
cc_186 N_A_109_47#_M1001_g N_VPWR_c_493_n 0.0027696f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_109_47#_M1019_g N_VPWR_c_493_n 0.00154685f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_109_47#_M1020_g N_VPWR_c_494_n 0.00154685f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_109_47#_M1019_g N_VPWR_c_500_n 0.00541359f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_109_47#_M1020_g N_VPWR_c_500_n 0.00541359f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_109_47#_M1001_g N_VPWR_c_508_n 0.00541359f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_109_47#_c_167_n N_VPWR_c_508_n 0.0210382f $X=0.68 $Y=2.31 $X2=0 $Y2=0
cc_193 N_A_109_47#_M1017_d N_VPWR_c_490_n 0.00209319f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_194 N_A_109_47#_M1001_g N_VPWR_c_490_n 0.0108276f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_109_47#_M1019_g N_VPWR_c_490_n 0.00950154f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_109_47#_M1020_g N_VPWR_c_490_n 0.00952874f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_109_47#_c_167_n N_VPWR_c_490_n 0.0124268f $X=0.68 $Y=2.31 $X2=0 $Y2=0
cc_198 N_A_109_47#_M1005_g N_Y_c_604_n 5.23702e-19 $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_109_47#_M1020_g N_Y_c_605_n 6.98608e-19 $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_109_47#_c_157_n N_VGND_c_754_n 0.0248793f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_201 N_A_109_47#_M1002_g N_VGND_c_755_n 0.00268723f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_A_109_47#_M1003_g N_VGND_c_755_n 0.00146448f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_A_109_47#_M1005_g N_VGND_c_756_n 0.00146448f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_109_47#_M1003_g N_VGND_c_762_n 0.00423644f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_205 N_A_109_47#_M1005_g N_VGND_c_762_n 0.00423644f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_206 N_A_109_47#_M1002_g N_VGND_c_770_n 0.00424619f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_109_47#_c_157_n N_VGND_c_770_n 0.020363f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_208 N_A_109_47#_M1023_d N_VGND_c_772_n 0.0020946f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_209 N_A_109_47#_M1002_g N_VGND_c_772_n 0.00706231f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_210 N_A_109_47#_M1003_g N_VGND_c_772_n 0.00575105f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_A_109_47#_M1005_g N_VGND_c_772_n 0.00577825f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_212 N_A_109_47#_c_157_n N_VGND_c_772_n 0.0123884f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_213 N_A_215_47#_c_279_n N_VPWR_M1001_d 0.00165831f $X=1.875 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_215_47#_c_282_n N_VPWR_M1020_d 0.00187252f $X=2.46 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_215_47#_c_279_n N_VPWR_c_493_n 0.0126919f $X=1.875 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_215_47#_M1000_g N_VPWR_c_494_n 0.00154685f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_215_47#_c_282_n N_VPWR_c_494_n 0.0126919f $X=2.46 $Y=1.53 $X2=0 $Y2=0
cc_218 N_A_215_47#_M1007_g N_VPWR_c_495_n 0.00146448f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_215_47#_M1008_g N_VPWR_c_495_n 0.00146448f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_215_47#_M1010_g N_VPWR_c_496_n 0.00146448f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_215_47#_M1014_g N_VPWR_c_496_n 0.00146448f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_215_47#_M1015_g N_VPWR_c_497_n 0.00146448f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_215_47#_M1021_g N_VPWR_c_497_n 0.00146448f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_215_47#_M1021_g N_VPWR_c_498_n 0.00541359f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_215_47#_M1022_g N_VPWR_c_498_n 0.00541359f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_215_47#_M1022_g N_VPWR_c_499_n 0.00316354f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_215_47#_c_309_n N_VPWR_c_500_n 0.0189039f $X=2.04 $Y=1.63 $X2=0 $Y2=0
cc_228 N_A_215_47#_M1000_g N_VPWR_c_502_n 0.00541359f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_215_47#_M1007_g N_VPWR_c_502_n 0.00541359f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_215_47#_M1008_g N_VPWR_c_504_n 0.00541359f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_215_47#_M1010_g N_VPWR_c_504_n 0.00541359f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_215_47#_M1014_g N_VPWR_c_506_n 0.00541359f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_215_47#_M1015_g N_VPWR_c_506_n 0.00541359f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_215_47#_c_278_n N_VPWR_c_508_n 0.0210382f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_235 N_A_215_47#_M1001_s N_VPWR_c_490_n 0.00209319f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_236 N_A_215_47#_M1019_s N_VPWR_c_490_n 0.00215201f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_237 N_A_215_47#_M1000_g N_VPWR_c_490_n 0.00952874f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_215_47#_M1007_g N_VPWR_c_490_n 0.00950154f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A_215_47#_M1008_g N_VPWR_c_490_n 0.00950154f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_215_47#_M1010_g N_VPWR_c_490_n 0.00950154f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_215_47#_M1014_g N_VPWR_c_490_n 0.00950154f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_215_47#_M1015_g N_VPWR_c_490_n 0.00950154f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_215_47#_M1021_g N_VPWR_c_490_n 0.00950154f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_A_215_47#_M1022_g N_VPWR_c_490_n 0.0108276f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_A_215_47#_c_278_n N_VPWR_c_490_n 0.0124268f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_246 N_A_215_47#_c_309_n N_VPWR_c_490_n 0.0122217f $X=2.04 $Y=1.63 $X2=0 $Y2=0
cc_247 N_A_215_47#_M1004_g N_Y_c_604_n 0.00636826f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_215_47#_M1006_g N_Y_c_604_n 0.00636826f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A_215_47#_M1009_g N_Y_c_604_n 5.23702e-19 $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A_215_47#_c_306_n N_Y_c_604_n 0.00518536f $X=2.04 $Y=0.4 $X2=0 $Y2=0
cc_251 N_A_215_47#_M1000_g N_Y_c_605_n 0.0102729f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_215_47#_M1007_g N_Y_c_605_n 0.0106215f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_215_47#_M1008_g N_Y_c_605_n 7.66249e-19 $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A_215_47#_c_309_n N_Y_c_605_n 0.00518536f $X=2.04 $Y=1.63 $X2=0 $Y2=0
cc_255 N_A_215_47#_M1006_g N_Y_c_585_n 0.00850187f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A_215_47#_M1009_g N_Y_c_585_n 0.00850187f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_257 N_A_215_47#_c_266_n N_Y_c_585_n 0.0359512f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_215_47#_c_269_n N_Y_c_585_n 0.00205431f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_215_47#_M1004_g N_Y_c_586_n 0.00240257f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_215_47#_M1006_g N_Y_c_586_n 0.00109384f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_215_47#_c_266_n N_Y_c_586_n 0.0265235f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_215_47#_c_267_n N_Y_c_586_n 0.00795337f $X=2.46 $Y=0.82 $X2=0 $Y2=0
cc_263 N_A_215_47#_c_269_n N_Y_c_586_n 0.00213376f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_215_47#_M1007_g N_Y_c_594_n 0.0107189f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_215_47#_M1008_g N_Y_c_594_n 0.0107189f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_215_47#_c_266_n N_Y_c_594_n 0.0359514f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_215_47#_c_269_n N_Y_c_594_n 0.00198252f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_215_47#_M1000_g N_Y_c_595_n 0.00265135f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_215_47#_M1007_g N_Y_c_595_n 0.00134262f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_215_47#_c_266_n N_Y_c_595_n 0.026643f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_215_47#_c_282_n N_Y_c_595_n 0.0088897f $X=2.46 $Y=1.53 $X2=0 $Y2=0
cc_272 N_A_215_47#_c_269_n N_Y_c_595_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_215_47#_M1006_g N_Y_c_632_n 5.23702e-19 $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A_215_47#_M1009_g N_Y_c_632_n 0.00636826f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_275 N_A_215_47#_M1011_g N_Y_c_632_n 0.00636826f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A_215_47#_M1012_g N_Y_c_632_n 5.23702e-19 $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A_215_47#_M1007_g N_Y_c_636_n 7.66249e-19 $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A_215_47#_M1008_g N_Y_c_636_n 0.0106215f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A_215_47#_M1010_g N_Y_c_636_n 0.0106215f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A_215_47#_M1014_g N_Y_c_636_n 7.66249e-19 $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_215_47#_M1011_g N_Y_c_587_n 0.00850187f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_215_47#_M1012_g N_Y_c_587_n 0.00850187f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_215_47#_c_266_n N_Y_c_587_n 0.0359512f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_215_47#_c_269_n N_Y_c_587_n 0.00205431f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_215_47#_M1010_g N_Y_c_596_n 0.0107189f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A_215_47#_M1014_g N_Y_c_596_n 0.0107189f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A_215_47#_c_266_n N_Y_c_596_n 0.0359514f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_215_47#_c_269_n N_Y_c_596_n 0.00198252f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A_215_47#_M1011_g N_Y_c_648_n 5.23702e-19 $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_215_47#_M1012_g N_Y_c_648_n 0.00636826f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_215_47#_M1013_g N_Y_c_648_n 0.00636826f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A_215_47#_M1016_g N_Y_c_648_n 5.23702e-19 $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_215_47#_M1010_g N_Y_c_652_n 7.66249e-19 $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A_215_47#_M1014_g N_Y_c_652_n 0.0106215f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A_215_47#_M1015_g N_Y_c_652_n 0.0106215f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A_215_47#_M1021_g N_Y_c_652_n 7.66249e-19 $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A_215_47#_M1013_g N_Y_c_588_n 0.00850187f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A_215_47#_M1016_g N_Y_c_588_n 0.00850187f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A_215_47#_c_266_n N_Y_c_588_n 0.0359512f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_215_47#_c_269_n N_Y_c_588_n 0.00205431f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A_215_47#_M1015_g N_Y_c_597_n 0.0107189f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_302 N_A_215_47#_M1021_g N_Y_c_597_n 0.0107189f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A_215_47#_c_266_n N_Y_c_597_n 0.0359514f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A_215_47#_c_269_n N_Y_c_597_n 0.00198252f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_305 N_A_215_47#_M1013_g N_Y_c_664_n 5.23702e-19 $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A_215_47#_M1016_g N_Y_c_664_n 0.00636826f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_215_47#_M1018_g N_Y_c_664_n 0.0109928f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A_215_47#_M1015_g N_Y_c_667_n 7.66249e-19 $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_215_47#_M1021_g N_Y_c_667_n 0.0106215f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_215_47#_M1022_g N_Y_c_667_n 0.0167471f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A_215_47#_M1018_g N_Y_c_589_n 0.0105322f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_312 N_A_215_47#_c_266_n N_Y_c_589_n 0.0139209f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_215_47#_M1022_g N_Y_c_598_n 0.0127492f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A_215_47#_c_266_n N_Y_c_598_n 0.0139209f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_215_47#_M1009_g N_Y_c_590_n 0.00110541f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A_215_47#_M1011_g N_Y_c_590_n 0.00110541f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A_215_47#_c_266_n N_Y_c_590_n 0.0265235f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_215_47#_c_269_n N_Y_c_590_n 0.00213376f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_215_47#_M1008_g N_Y_c_599_n 0.00135419f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_215_47#_M1010_g N_Y_c_599_n 0.00135419f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A_215_47#_c_266_n N_Y_c_599_n 0.026643f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_215_47#_c_269_n N_Y_c_599_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_215_47#_M1012_g N_Y_c_591_n 0.00110541f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_324 N_A_215_47#_M1013_g N_Y_c_591_n 0.00110541f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A_215_47#_c_266_n N_Y_c_591_n 0.0265235f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_215_47#_c_269_n N_Y_c_591_n 0.00213376f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_215_47#_M1014_g N_Y_c_600_n 0.00135419f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_215_47#_M1015_g N_Y_c_600_n 0.00135419f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_215_47#_c_266_n N_Y_c_600_n 0.026643f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_215_47#_c_269_n N_Y_c_600_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_215_47#_M1016_g N_Y_c_592_n 0.00110541f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_332 N_A_215_47#_M1018_g N_Y_c_592_n 0.00110541f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_333 N_A_215_47#_c_266_n N_Y_c_592_n 0.0265235f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_215_47#_c_269_n N_Y_c_592_n 0.00213376f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_215_47#_M1021_g N_Y_c_601_n 0.00135419f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_215_47#_M1022_g N_Y_c_601_n 0.00135419f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_215_47#_c_266_n N_Y_c_601_n 0.026643f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_215_47#_c_269_n N_Y_c_601_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A_215_47#_M1018_g Y 0.00601334f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A_215_47#_c_266_n Y 0.015258f $X=5.52 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_215_47#_c_269_n Y 0.00701084f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_342 N_A_215_47#_c_262_n N_VGND_M1002_s 0.00162006f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_343 N_A_215_47#_c_267_n N_VGND_M1005_s 0.00186748f $X=2.46 $Y=0.82 $X2=0
+ $Y2=0
cc_344 N_A_215_47#_c_262_n N_VGND_c_755_n 0.0122414f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_345 N_A_215_47#_M1004_g N_VGND_c_756_n 0.00146448f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_346 N_A_215_47#_c_267_n N_VGND_c_756_n 0.0122414f $X=2.46 $Y=0.82 $X2=0 $Y2=0
cc_347 N_A_215_47#_M1006_g N_VGND_c_757_n 0.00146448f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_348 N_A_215_47#_M1009_g N_VGND_c_757_n 0.00146448f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_349 N_A_215_47#_M1011_g N_VGND_c_758_n 0.00146448f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_215_47#_M1012_g N_VGND_c_758_n 0.00146448f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_351 N_A_215_47#_M1013_g N_VGND_c_759_n 0.00146448f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_352 N_A_215_47#_M1016_g N_VGND_c_759_n 0.00146448f $X=5.19 $Y=0.56 $X2=0
+ $Y2=0
cc_353 N_A_215_47#_M1016_g N_VGND_c_760_n 0.00424619f $X=5.19 $Y=0.56 $X2=0
+ $Y2=0
cc_354 N_A_215_47#_M1018_g N_VGND_c_760_n 0.00424619f $X=5.61 $Y=0.56 $X2=0
+ $Y2=0
cc_355 N_A_215_47#_M1018_g N_VGND_c_761_n 0.00316354f $X=5.61 $Y=0.56 $X2=0
+ $Y2=0
cc_356 N_A_215_47#_c_262_n N_VGND_c_762_n 0.00390702f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_357 N_A_215_47#_c_306_n N_VGND_c_762_n 0.0179571f $X=2.04 $Y=0.4 $X2=0 $Y2=0
cc_358 N_A_215_47#_M1004_g N_VGND_c_764_n 0.00541562f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_359 N_A_215_47#_M1006_g N_VGND_c_764_n 0.00424619f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_215_47#_M1009_g N_VGND_c_766_n 0.00424619f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_361 N_A_215_47#_M1011_g N_VGND_c_766_n 0.00424619f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_215_47#_M1012_g N_VGND_c_768_n 0.00424619f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_363 N_A_215_47#_M1013_g N_VGND_c_768_n 0.00424619f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_364 N_A_215_47#_c_261_n N_VGND_c_770_n 0.020318f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_365 N_A_215_47#_c_262_n N_VGND_c_770_n 0.00193763f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_366 N_A_215_47#_M1002_d N_VGND_c_772_n 0.0020946f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_215_47#_M1003_d N_VGND_c_772_n 0.00215347f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_215_47#_M1004_g N_VGND_c_772_n 0.00952891f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_369 N_A_215_47#_M1006_g N_VGND_c_772_n 0.00573624f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_370 N_A_215_47#_M1009_g N_VGND_c_772_n 0.00573624f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_371 N_A_215_47#_M1011_g N_VGND_c_772_n 0.00573624f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_372 N_A_215_47#_M1012_g N_VGND_c_772_n 0.00573624f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_373 N_A_215_47#_M1013_g N_VGND_c_772_n 0.00573624f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_374 N_A_215_47#_M1016_g N_VGND_c_772_n 0.00573624f $X=5.19 $Y=0.56 $X2=0
+ $Y2=0
cc_375 N_A_215_47#_M1018_g N_VGND_c_772_n 0.00706231f $X=5.61 $Y=0.56 $X2=0
+ $Y2=0
cc_376 N_A_215_47#_c_261_n N_VGND_c_772_n 0.0123792f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_377 N_A_215_47#_c_262_n N_VGND_c_772_n 0.012122f $X=1.875 $Y=0.82 $X2=0 $Y2=0
cc_378 N_A_215_47#_c_306_n N_VGND_c_772_n 0.0120759f $X=2.04 $Y=0.4 $X2=0 $Y2=0
cc_379 N_A_215_47#_c_267_n N_VGND_c_772_n 6.28727e-19 $X=2.46 $Y=0.82 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_490_n N_Y_M1000_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_490_n N_Y_M1008_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_490_n N_Y_M1014_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_490_n N_Y_M1021_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_502_n N_Y_c_605_n 0.0189039f $X=3.215 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_490_n N_Y_c_605_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_M1007_s N_Y_c_594_n 0.00185611f $X=3.165 $Y=1.485 $X2=0 $Y2=0
cc_387 N_VPWR_c_495_n N_Y_c_594_n 0.0104788f $X=3.3 $Y=2 $X2=0 $Y2=0
cc_388 N_VPWR_c_504_n N_Y_c_636_n 0.0189039f $X=4.055 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_490_n N_Y_c_636_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_M1010_s N_Y_c_596_n 0.00185611f $X=4.005 $Y=1.485 $X2=0 $Y2=0
cc_391 N_VPWR_c_496_n N_Y_c_596_n 0.0104788f $X=4.14 $Y=2 $X2=0 $Y2=0
cc_392 N_VPWR_c_506_n N_Y_c_652_n 0.0189039f $X=4.895 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_490_n N_Y_c_652_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_M1015_s N_Y_c_597_n 0.00185611f $X=4.845 $Y=1.485 $X2=0 $Y2=0
cc_395 N_VPWR_c_497_n N_Y_c_597_n 0.0104788f $X=4.98 $Y=2 $X2=0 $Y2=0
cc_396 N_VPWR_c_498_n N_Y_c_667_n 0.0189039f $X=5.735 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_490_n N_Y_c_667_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_M1022_s N_Y_c_598_n 0.00406309f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_399 N_VPWR_c_499_n N_Y_c_598_n 0.0108818f $X=5.82 $Y=2 $X2=0 $Y2=0
cc_400 N_Y_c_585_n N_VGND_M1006_d 0.00162006f $X=3.555 $Y=0.82 $X2=0 $Y2=0
cc_401 N_Y_c_587_n N_VGND_M1011_d 0.00162006f $X=4.395 $Y=0.82 $X2=0 $Y2=0
cc_402 N_Y_c_588_n N_VGND_M1013_d 0.00162006f $X=5.235 $Y=0.82 $X2=0 $Y2=0
cc_403 N_Y_c_589_n N_VGND_M1018_d 0.0031176f $X=5.97 $Y=0.82 $X2=0 $Y2=0
cc_404 N_Y_c_585_n N_VGND_c_757_n 0.0122414f $X=3.555 $Y=0.82 $X2=0 $Y2=0
cc_405 N_Y_c_587_n N_VGND_c_758_n 0.0122414f $X=4.395 $Y=0.82 $X2=0 $Y2=0
cc_406 N_Y_c_588_n N_VGND_c_759_n 0.0122414f $X=5.235 $Y=0.82 $X2=0 $Y2=0
cc_407 N_Y_c_588_n N_VGND_c_760_n 0.00193763f $X=5.235 $Y=0.82 $X2=0 $Y2=0
cc_408 N_Y_c_664_n N_VGND_c_760_n 0.0182681f $X=5.4 $Y=0.4 $X2=0 $Y2=0
cc_409 N_Y_c_589_n N_VGND_c_760_n 0.00193763f $X=5.97 $Y=0.82 $X2=0 $Y2=0
cc_410 N_Y_c_589_n N_VGND_c_761_n 0.0127122f $X=5.97 $Y=0.82 $X2=0 $Y2=0
cc_411 N_Y_c_604_n N_VGND_c_764_n 0.0182681f $X=2.88 $Y=0.4 $X2=0 $Y2=0
cc_412 N_Y_c_585_n N_VGND_c_764_n 0.00193763f $X=3.555 $Y=0.82 $X2=0 $Y2=0
cc_413 N_Y_c_585_n N_VGND_c_766_n 0.00193763f $X=3.555 $Y=0.82 $X2=0 $Y2=0
cc_414 N_Y_c_632_n N_VGND_c_766_n 0.0182681f $X=3.72 $Y=0.4 $X2=0 $Y2=0
cc_415 N_Y_c_587_n N_VGND_c_766_n 0.00193763f $X=4.395 $Y=0.82 $X2=0 $Y2=0
cc_416 N_Y_c_587_n N_VGND_c_768_n 0.00193763f $X=4.395 $Y=0.82 $X2=0 $Y2=0
cc_417 N_Y_c_648_n N_VGND_c_768_n 0.0182681f $X=4.56 $Y=0.4 $X2=0 $Y2=0
cc_418 N_Y_c_588_n N_VGND_c_768_n 0.00193763f $X=5.235 $Y=0.82 $X2=0 $Y2=0
cc_419 N_Y_c_589_n N_VGND_c_771_n 0.00736076f $X=5.97 $Y=0.82 $X2=0 $Y2=0
cc_420 N_Y_M1004_s N_VGND_c_772_n 0.00215347f $X=2.745 $Y=0.235 $X2=0 $Y2=0
cc_421 N_Y_M1009_s N_VGND_c_772_n 0.00215347f $X=3.585 $Y=0.235 $X2=0 $Y2=0
cc_422 N_Y_M1012_s N_VGND_c_772_n 0.00215347f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_423 N_Y_M1016_s N_VGND_c_772_n 0.00215347f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_424 N_Y_c_604_n N_VGND_c_772_n 0.0121741f $X=2.88 $Y=0.4 $X2=0 $Y2=0
cc_425 N_Y_c_585_n N_VGND_c_772_n 0.00825759f $X=3.555 $Y=0.82 $X2=0 $Y2=0
cc_426 N_Y_c_632_n N_VGND_c_772_n 0.0121741f $X=3.72 $Y=0.4 $X2=0 $Y2=0
cc_427 N_Y_c_587_n N_VGND_c_772_n 0.00825759f $X=4.395 $Y=0.82 $X2=0 $Y2=0
cc_428 N_Y_c_648_n N_VGND_c_772_n 0.0121741f $X=4.56 $Y=0.4 $X2=0 $Y2=0
cc_429 N_Y_c_588_n N_VGND_c_772_n 0.00825759f $X=5.235 $Y=0.82 $X2=0 $Y2=0
cc_430 N_Y_c_664_n N_VGND_c_772_n 0.0121741f $X=5.4 $Y=0.4 $X2=0 $Y2=0
cc_431 N_Y_c_589_n N_VGND_c_772_n 0.0169393f $X=5.97 $Y=0.82 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkinv_4.pxi.spice
* Created: Thu Aug 27 14:12:42 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINV_4%A N_A_M1000_g N_A_M1002_g N_A_M1001_g N_A_c_76_n
+ N_A_M1003_g N_A_M1004_g N_A_c_79_n N_A_M1008_g N_A_M1005_g N_A_c_82_n
+ N_A_M1009_g N_A_M1006_g N_A_M1007_g N_A_c_86_n N_A_c_87_n N_A_c_88_n
+ N_A_c_89_n N_A_c_90_n N_A_c_91_n N_A_c_92_n A A A A A
+ PM_SKY130_FD_SC_HD__CLKINV_4%A
x_PM_SKY130_FD_SC_HD__CLKINV_4%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_M1005_s
+ N_VPWR_M1007_s N_VPWR_c_172_n N_VPWR_c_173_n N_VPWR_c_174_n N_VPWR_c_175_n
+ N_VPWR_c_176_n N_VPWR_c_177_n N_VPWR_c_178_n N_VPWR_c_179_n VPWR
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_182_n N_VPWR_c_171_n
+ PM_SKY130_FD_SC_HD__CLKINV_4%VPWR
x_PM_SKY130_FD_SC_HD__CLKINV_4%Y N_Y_M1002_s N_Y_M1008_s N_Y_M1000_d N_Y_M1004_d
+ N_Y_M1006_d N_Y_c_223_n N_Y_c_224_n N_Y_c_225_n N_Y_c_235_n N_Y_c_236_n
+ N_Y_c_294_n N_Y_c_237_n N_Y_c_226_n N_Y_c_227_n N_Y_c_298_n N_Y_c_238_n
+ N_Y_c_228_n N_Y_c_229_n N_Y_c_302_n N_Y_c_239_n N_Y_c_240_n N_Y_c_230_n
+ N_Y_c_241_n N_Y_c_231_n N_Y_c_242_n Y Y Y N_Y_c_233_n N_Y_c_244_n
+ PM_SKY130_FD_SC_HD__CLKINV_4%Y
x_PM_SKY130_FD_SC_HD__CLKINV_4%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_M1009_d
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n VGND N_VGND_c_333_n
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n
+ N_VGND_c_339_n N_VGND_c_340_n PM_SKY130_FD_SC_HD__CLKINV_4%VGND
cc_1 VNB N_A_M1000_g 5.00591e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_2 VNB N_A_M1002_g 0.0369233f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.445
cc_3 VNB N_A_M1001_g 4.57532e-19 $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.985
cc_4 VNB N_A_c_76_n 0.0126448f $X=-0.19 $Y=-0.24 $X2=1.3 $Y2=1.16
cc_5 VNB N_A_M1003_g 0.0279614f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.445
cc_6 VNB N_A_M1004_g 4.57707e-19 $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.985
cc_7 VNB N_A_c_79_n 0.0126445f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_8 VNB N_A_M1008_g 0.0279614f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=0.445
cc_9 VNB N_A_M1005_g 4.57707e-19 $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.985
cc_10 VNB N_A_c_82_n 0.0126448f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.16
cc_11 VNB N_A_M1009_g 0.0367478f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=0.445
cc_12 VNB N_A_M1006_g 4.57415e-19 $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.985
cc_13 VNB N_A_M1007_g 4.94191e-19 $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.985
cc_14 VNB N_A_c_86_n 0.0151897f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_15 VNB N_A_c_87_n 0.0172072f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.16
cc_16 VNB N_A_c_88_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.16
cc_17 VNB N_A_c_89_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.16
cc_18 VNB N_A_c_90_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_19 VNB N_A_c_91_n 0.00429822f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.16
cc_20 VNB N_A_c_92_n 0.0321714f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.16
cc_21 VNB N_VPWR_c_171_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_22 VNB N_Y_c_223_n 0.0201292f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.445
cc_23 VNB N_Y_c_224_n 0.0142122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_225_n 0.0104981f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.295
cc_25 VNB N_Y_c_226_n 0.00119645f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.985
cc_26 VNB N_Y_c_227_n 0.00514362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_228_n 0.00119511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_229_n 0.0120925f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.985
cc_29 VNB N_Y_c_230_n 0.00208412f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.16
cc_30 VNB N_Y_c_231_n 0.00203725f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_31 VNB Y 0.0231444f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.105
cc_32 VNB N_Y_c_233_n 0.0132357f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_33 VNB N_VGND_c_330_n 0.00482504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_331_n 0.00400382f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.445
cc_35 VNB N_VGND_c_332_n 0.00484653f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=1.985
cc_36 VNB N_VGND_c_333_n 0.0184172f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.16
cc_37 VNB N_VGND_c_334_n 0.0154375f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.295
cc_38 VNB N_VGND_c_335_n 0.0152868f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_39 VNB N_VGND_c_336_n 0.0194663f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=1.985
cc_40 VNB N_VGND_c_337_n 0.191074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_338_n 0.00564654f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.985
cc_42 VNB N_VGND_c_339_n 0.00497354f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.16
cc_43 VNB N_VGND_c_340_n 0.00574268f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_44 VPB N_A_M1000_g 0.0232949f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_45 VPB N_A_M1001_g 0.0195526f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.985
cc_46 VPB N_A_M1004_g 0.0195731f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_47 VPB N_A_M1005_g 0.0195731f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_48 VPB N_A_M1006_g 0.0195506f $X=-0.19 $Y=1.305 $X2=2.235 $Y2=1.985
cc_49 VPB N_A_M1007_g 0.0231846f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.985
cc_50 VPB N_VPWR_c_172_n 0.0115225f $X=-0.19 $Y=1.305 $X2=1.3 $Y2=1.16
cc_51 VPB N_VPWR_c_173_n 0.0329354f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.025
cc_52 VPB N_VPWR_c_174_n 0.00400996f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.295
cc_53 VPB N_VPWR_c_175_n 0.00400996f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_54 VPB N_VPWR_c_176_n 0.0122918f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.025
cc_55 VPB N_VPWR_c_177_n 0.0329156f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=0.445
cc_56 VPB N_VPWR_c_178_n 0.0167849f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_57 VPB N_VPWR_c_179_n 0.00497514f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.985
cc_58 VPB N_VPWR_c_180_n 0.0167849f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_59 VPB N_VPWR_c_181_n 0.0167406f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.295
cc_60 VPB N_VPWR_c_182_n 0.00497514f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.16
cc_61 VPB N_VPWR_c_171_n 0.0422076f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_62 VPB N_Y_c_223_n 0.00764075f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=0.445
cc_63 VPB N_Y_c_235_n 0.00236425f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_64 VPB N_Y_c_236_n 0.00749967f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_65 VPB N_Y_c_237_n 0.00246432f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=0.445
cc_66 VPB N_Y_c_238_n 0.00241839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_Y_c_239_n 0.00136408f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.16
cc_68 VPB N_Y_c_240_n 0.00206815f $X=-0.19 $Y=1.305 $X2=2.31 $Y2=1.16
cc_69 VPB N_Y_c_241_n 0.00206815f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.16
cc_70 VPB N_Y_c_242_n 0.0021151f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_71 VPB Y 0.00841183f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.105
cc_72 VPB N_Y_c_244_n 0.00784985f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_73 N_A_M1000_g N_VPWR_c_173_n 0.00343841f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_M1001_g N_VPWR_c_174_n 0.00161372f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_VPWR_c_174_n 0.00161372f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1005_g N_VPWR_c_175_n 0.00161372f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_VPWR_c_175_n 0.00161372f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1007_g N_VPWR_c_177_n 0.0034537f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1004_g N_VPWR_c_178_n 0.00585385f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_M1005_g N_VPWR_c_178_n 0.00585385f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_VPWR_c_180_n 0.00585385f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_M1001_g N_VPWR_c_180_n 0.00585385f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_VPWR_c_181_n 0.00585385f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1007_g N_VPWR_c_181_n 0.00585385f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1000_g N_VPWR_c_171_n 0.0115347f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_VPWR_c_171_n 0.0105664f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_VPWR_c_171_n 0.0105664f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1005_g N_VPWR_c_171_n 0.0105664f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_VPWR_c_171_n 0.0105664f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_M1007_g N_VPWR_c_171_n 0.0115663f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_Y_c_223_n 0.00284045f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_c_86_n N_Y_c_223_n 0.0135164f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_93 A N_Y_c_223_n 0.0178211f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A_M1002_g N_Y_c_224_n 0.0142819f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_c_86_n N_Y_c_224_n 0.01134f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_96 A N_Y_c_224_n 0.042008f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A_M1000_g N_Y_c_235_n 0.0165836f $X=0.515 $Y=1.985 $X2=0 $Y2=0
cc_98 A N_Y_c_235_n 0.011067f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_99 N_A_M1001_g N_Y_c_237_n 0.0150738f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_c_76_n N_Y_c_237_n 0.00216422f $X=1.3 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_M1004_g N_Y_c_237_n 0.0150738f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_102 A N_Y_c_237_n 0.0428385f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_Y_c_226_n 0.00194229f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_M1003_g N_Y_c_226_n 0.00105846f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_M1003_g N_Y_c_227_n 0.0122413f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_c_79_n N_Y_c_227_n 0.00225558f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_M1008_g N_Y_c_227_n 0.0122413f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_108 A N_Y_c_227_n 0.0424729f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_109 N_A_M1005_g N_Y_c_238_n 0.0150738f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_c_82_n N_Y_c_238_n 0.00216422f $X=2.16 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_M1006_g N_Y_c_238_n 0.0150738f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_112 A N_Y_c_238_n 0.0424733f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_113 N_A_M1008_g N_Y_c_228_n 0.00105549f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_M1009_g N_Y_c_228_n 0.00192273f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_M1009_g N_Y_c_229_n 0.0142819f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_c_92_n N_Y_c_229_n 0.0116658f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_117 A N_Y_c_229_n 0.0368972f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_M1007_g N_Y_c_239_n 0.0174361f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_119 A N_Y_c_239_n 0.0055064f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A_c_87_n N_Y_c_240_n 0.00225251f $X=0.87 $Y=1.16 $X2=0 $Y2=0
cc_121 A N_Y_c_240_n 0.0209598f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_c_76_n N_Y_c_230_n 0.00233861f $X=1.3 $Y=1.16 $X2=0 $Y2=0
cc_123 A N_Y_c_230_n 0.02119f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_c_79_n N_Y_c_241_n 0.00225251f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_125 A N_Y_c_241_n 0.0209598f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_126 N_A_c_82_n N_Y_c_231_n 0.00233861f $X=2.16 $Y=1.16 $X2=0 $Y2=0
cc_127 A N_Y_c_231_n 0.0207824f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A_c_92_n N_Y_c_242_n 0.00225251f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_129 A N_Y_c_242_n 0.0213708f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A_M1009_g Y 0.00326216f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_c_92_n Y 0.0152731f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_132 A Y 0.0181732f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_133 N_A_M1002_g N_VGND_c_330_n 0.00341694f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A_M1003_g N_VGND_c_331_n 0.00161372f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_M1008_g N_VGND_c_331_n 0.00160701f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_M1009_g N_VGND_c_332_n 0.00344739f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_M1002_g N_VGND_c_334_n 0.00437852f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_VGND_c_334_n 0.00437852f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_M1008_g N_VGND_c_335_n 0.00437852f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_M1009_g N_VGND_c_335_n 0.00437852f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_M1002_g N_VGND_c_337_n 0.00718425f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_VGND_c_337_n 0.00588456f $X=1.375 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_M1008_g N_VGND_c_337_n 0.00588456f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_M1009_g N_VGND_c_337_n 0.00717171f $X=2.235 $Y=0.445 $X2=0 $Y2=0
cc_145 N_VPWR_c_171_n N_Y_M1000_d 0.00319983f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_146 N_VPWR_c_171_n N_Y_M1004_d 0.00319983f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_147 N_VPWR_c_171_n N_Y_M1006_d 0.00302653f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_148 N_VPWR_M1000_s N_Y_c_235_n 0.00113743f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_149 N_VPWR_c_173_n N_Y_c_235_n 0.00875025f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_150 N_VPWR_M1000_s N_Y_c_236_n 0.0025525f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_151 N_VPWR_c_173_n N_Y_c_236_n 0.0153867f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_152 N_VPWR_c_180_n N_Y_c_294_n 0.0124093f $X=1.03 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_171_n N_Y_c_294_n 0.00960102f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_M1001_s N_Y_c_237_n 0.00176461f $X=1.02 $Y=1.485 $X2=0 $Y2=0
cc_155 N_VPWR_c_174_n N_Y_c_237_n 0.0135055f $X=1.16 $Y=1.965 $X2=0 $Y2=0
cc_156 N_VPWR_c_178_n N_Y_c_298_n 0.0124093f $X=1.89 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_171_n N_Y_c_298_n 0.00960102f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_M1005_s N_Y_c_238_n 0.00176461f $X=1.88 $Y=1.485 $X2=0 $Y2=0
cc_159 N_VPWR_c_175_n N_Y_c_238_n 0.0135055f $X=2.02 $Y=1.965 $X2=0 $Y2=0
cc_160 N_VPWR_c_181_n N_Y_c_302_n 0.0125603f $X=2.75 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_171_n N_Y_c_302_n 0.00979076f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_162 N_VPWR_M1007_s N_Y_c_239_n 3.93317e-19 $X=2.74 $Y=1.485 $X2=0 $Y2=0
cc_163 N_VPWR_c_177_n N_Y_c_239_n 0.00305515f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_164 N_VPWR_M1007_s N_Y_c_244_n 0.00409082f $X=2.74 $Y=1.485 $X2=0 $Y2=0
cc_165 N_VPWR_c_177_n N_Y_c_244_n 0.0271316f $X=2.88 $Y=1.965 $X2=0 $Y2=0
cc_166 N_Y_c_224_n N_VGND_c_330_n 0.0212491f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_167 N_Y_c_227_n N_VGND_c_331_n 0.0164203f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_168 N_Y_c_229_n N_VGND_c_332_n 0.0214243f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_169 N_Y_c_224_n N_VGND_c_333_n 0.00440462f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_170 N_Y_c_225_n N_VGND_c_333_n 0.00289403f $X=0.275 $Y=0.81 $X2=0 $Y2=0
cc_171 N_Y_c_224_n N_VGND_c_334_n 0.0022979f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_172 N_Y_c_226_n N_VGND_c_334_n 0.01283f $X=1.16 $Y=0.445 $X2=0 $Y2=0
cc_173 N_Y_c_227_n N_VGND_c_334_n 0.0022979f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_174 N_Y_c_227_n N_VGND_c_335_n 0.0022979f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_175 N_Y_c_228_n N_VGND_c_335_n 0.0126752f $X=2.02 $Y=0.445 $X2=0 $Y2=0
cc_176 N_Y_c_229_n N_VGND_c_335_n 0.0022979f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_177 N_Y_c_229_n N_VGND_c_336_n 0.00333776f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_178 N_Y_c_233_n N_VGND_c_336_n 0.00510712f $X=2.985 $Y=0.895 $X2=0 $Y2=0
cc_179 N_Y_M1002_s N_VGND_c_337_n 0.00234276f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_180 N_Y_M1008_s N_VGND_c_337_n 0.0023674f $X=1.88 $Y=0.235 $X2=0 $Y2=0
cc_181 N_Y_c_224_n N_VGND_c_337_n 0.0125077f $X=1.03 $Y=0.81 $X2=0 $Y2=0
cc_182 N_Y_c_225_n N_VGND_c_337_n 0.00478629f $X=0.275 $Y=0.81 $X2=0 $Y2=0
cc_183 N_Y_c_226_n N_VGND_c_337_n 0.00978777f $X=1.16 $Y=0.445 $X2=0 $Y2=0
cc_184 N_Y_c_227_n N_VGND_c_337_n 0.00837675f $X=1.89 $Y=0.81 $X2=0 $Y2=0
cc_185 N_Y_c_228_n N_VGND_c_337_n 0.00959809f $X=2.02 $Y=0.445 $X2=0 $Y2=0
cc_186 N_Y_c_229_n N_VGND_c_337_n 0.0106771f $X=2.835 $Y=0.81 $X2=0 $Y2=0
cc_187 N_Y_c_233_n N_VGND_c_337_n 0.0084464f $X=2.985 $Y=0.895 $X2=0 $Y2=0

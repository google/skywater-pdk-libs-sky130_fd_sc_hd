# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__o41ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.170000 1.075000 7.940000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 1.075000 5.980000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.075000 4.020000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.700000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 2.160000 0.905000 ;
        RECT 0.515000 1.445000 3.885000 1.615000 ;
        RECT 0.515000 1.615000 0.845000 2.465000 ;
        RECT 1.355000 1.615000 1.685000 2.465000 ;
        RECT 1.870000 0.905000 2.160000 1.445000 ;
        RECT 2.715000 1.615000 3.045000 2.125000 ;
        RECT 3.555000 1.615000 3.885000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  2.625000 0.465000 ;
      RECT 0.085000  0.465000  0.345000 0.905000 ;
      RECT 0.085000  1.445000  0.345000 2.635000 ;
      RECT 1.015000  1.835000  1.185000 2.635000 ;
      RECT 1.855000  1.835000  2.105000 2.635000 ;
      RECT 2.295000  1.785000  2.545000 2.295000 ;
      RECT 2.295000  2.295000  4.225000 2.465000 ;
      RECT 2.350000  0.465000  2.625000 0.735000 ;
      RECT 2.350000  0.735000  9.865000 0.905000 ;
      RECT 2.795000  0.085000  2.965000 0.545000 ;
      RECT 3.135000  0.255000  3.465000 0.735000 ;
      RECT 3.215000  1.785000  3.385000 2.295000 ;
      RECT 3.635000  0.085000  3.805000 0.545000 ;
      RECT 3.975000  0.255000  4.305000 0.735000 ;
      RECT 4.055000  1.445000  5.985000 1.615000 ;
      RECT 4.055000  1.615000  4.225000 2.295000 ;
      RECT 4.395000  1.785000  4.645000 2.295000 ;
      RECT 4.395000  2.295000  7.685000 2.465000 ;
      RECT 4.475000  0.085000  4.645000 0.545000 ;
      RECT 4.815000  0.255000  5.145000 0.735000 ;
      RECT 4.815000  1.615000  5.145000 2.125000 ;
      RECT 5.315000  0.085000  5.485000 0.545000 ;
      RECT 5.315000  1.785000  5.485000 2.295000 ;
      RECT 5.655000  0.255000  5.985000 0.735000 ;
      RECT 5.655000  1.615000  5.985000 2.125000 ;
      RECT 6.175000  0.260000  6.505000 0.735000 ;
      RECT 6.175000  1.445000  9.865000 1.615000 ;
      RECT 6.175000  1.615000  6.505000 2.125000 ;
      RECT 6.675000  0.085000  6.845000 0.545000 ;
      RECT 6.675000  1.785000  6.845000 2.295000 ;
      RECT 7.015000  0.260000  7.345000 0.735000 ;
      RECT 7.015000  1.615000  7.345000 2.125000 ;
      RECT 7.515000  0.085000  7.685000 0.545000 ;
      RECT 7.515000  1.785000  7.685000 2.295000 ;
      RECT 7.855000  0.260000  8.185000 0.735000 ;
      RECT 7.855000  1.615000  8.185000 2.465000 ;
      RECT 8.355000  0.085000  8.525000 0.545000 ;
      RECT 8.355000  1.835000  8.525000 2.635000 ;
      RECT 8.695000  0.260000  9.025000 0.735000 ;
      RECT 8.695000  1.615000  9.025000 2.465000 ;
      RECT 9.195000  0.085000  9.365000 0.545000 ;
      RECT 9.195000  1.835000  9.365000 2.635000 ;
      RECT 9.535000  0.260000  9.865000 0.735000 ;
      RECT 9.535000  1.615000  9.865000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_4
END LIBRARY

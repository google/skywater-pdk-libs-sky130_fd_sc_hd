* File: sky130_fd_sc_hd__einvp_2.spice
* Created: Thu Aug 27 14:20:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__einvp_2.pex.spice"
.subckt sky130_fd_sc_hd__einvp_2  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_TE_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=7.14 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1008_d N_TE_M1000_g N_A_204_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.08775 PD=1.18458 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_TE_M1009_g N_A_204_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_204_47#_M1006_d N_A_M1006_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_204_47#_M1007_d N_A_M1007_g N_Z_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_TE_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1664 AS=0.1664 PD=1.8 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_215_309#_M1001_d N_A_27_47#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.2444 AS=0.1269 PD=2.4 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75000.2
+ SB=75001.5 A=0.141 P=2.18 MULT=1
MM1003 N_A_215_309#_M1003_d N_A_27_47#_M1003_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.155294 AS=0.1269 PD=1.28402 PS=1.21 NRD=5.2205 NRS=0 M=1 R=6.26667
+ SA=75000.6 SB=75001.1 A=0.141 P=2.18 MULT=1
MM1002 N_A_215_309#_M1003_d N_A_M1002_g N_Z_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165206 AS=0.135 PD=1.36598 PS=1.27 NRD=3.9203 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_215_309#_M1005_d N_A_M1005_g N_Z_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_58 VPB 0 1.1096e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__einvp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__buf_2.spice.SKY130_FD_SC_HD__BUF_2.pxi
* Created: Thu Aug 27 14:09:44 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_2%A N_A_M1004_g N_A_M1001_g A N_A_c_41_n
+ PM_SKY130_FD_SC_HD__BUF_2%A
x_PM_SKY130_FD_SC_HD__BUF_2%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_70_n N_A_27_47#_M1003_g N_A_27_47#_M1000_g N_A_27_47#_c_71_n
+ N_A_27_47#_M1005_g N_A_27_47#_M1002_g N_A_27_47#_c_139_p N_A_27_47#_c_79_n
+ N_A_27_47#_c_72_n N_A_27_47#_c_73_n N_A_27_47#_c_80_n N_A_27_47#_c_81_n
+ N_A_27_47#_c_82_n N_A_27_47#_c_74_n N_A_27_47#_c_75_n N_A_27_47#_c_76_n
+ PM_SKY130_FD_SC_HD__BUF_2%A_27_47#
x_PM_SKY130_FD_SC_HD__BUF_2%VPWR N_VPWR_M1001_d N_VPWR_M1002_d N_VPWR_c_149_n
+ N_VPWR_c_150_n N_VPWR_c_151_n VPWR VPWR N_VPWR_c_152_n N_VPWR_c_153_n
+ N_VPWR_c_154_n N_VPWR_c_148_n PM_SKY130_FD_SC_HD__BUF_2%VPWR
x_PM_SKY130_FD_SC_HD__BUF_2%X N_X_M1003_s N_X_M1000_s N_X_c_179_n N_X_c_181_n
+ N_X_c_177_n X X X PM_SKY130_FD_SC_HD__BUF_2%X
x_PM_SKY130_FD_SC_HD__BUF_2%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_c_201_n
+ N_VGND_c_202_n N_VGND_c_203_n VGND VGND N_VGND_c_204_n N_VGND_c_205_n
+ N_VGND_c_206_n N_VGND_c_207_n PM_SKY130_FD_SC_HD__BUF_2%VGND
cc_1 VNB N_A_M1004_g 0.0381123f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.0174906f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A_c_41_n 0.0349516f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_c_70_n 0.0158658f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.125
cc_5 VNB N_A_27_47#_c_71_n 0.0204757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_72_n 0.00287879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_73_n 0.00742394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_74_n 0.00221485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_75_n 0.00102941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_76_n 0.0484055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_VPWR_c_148_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_X_c_177_n 7.39732e-19 $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_13 VNB N_VGND_c_201_n 0.00278085f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_14 VNB N_VGND_c_202_n 0.0100714f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_15 VNB N_VGND_c_203_n 0.0352119f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_16 VNB N_VGND_c_204_n 0.0174195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_205_n 0.0154765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_206_n 0.00513086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_207_n 0.124444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VPB N_A_M1001_g 0.0465559f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.125
cc_21 VPB A 0.00733067f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_22 VPB N_A_c_41_n 0.00920847f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_23 VPB N_A_27_47#_M1000_g 0.0187981f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_24 VPB N_A_27_47#_M1002_g 0.0253024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A_27_47#_c_79_n 0.00658534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_47#_c_80_n 0.00565572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_27_47#_c_81_n 0.00830017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_c_82_n 0.00146014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_27_47#_c_76_n 0.00846909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_149_n 0.00321136f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_31 VPB N_VPWR_c_150_n 0.0100455f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_32 VPB N_VPWR_c_151_n 0.0463009f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_33 VPB N_VPWR_c_152_n 0.0183831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_153_n 0.0154765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_154_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_148_n 0.0499797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_X_c_177_n 0.00107597f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_38 N_A_M1004_g N_A_27_47#_c_70_n 0.0198678f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_39 N_A_M1001_g N_A_27_47#_M1000_g 0.0202342f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_40 N_A_M1001_g N_A_27_47#_c_79_n 0.0043143f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_41 N_A_M1004_g N_A_27_47#_c_72_n 0.0163494f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_42 A N_A_27_47#_c_72_n 0.00690379f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_43 N_A_c_41_n N_A_27_47#_c_72_n 3.36787e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_44 A N_A_27_47#_c_73_n 0.0143207f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_45 N_A_c_41_n N_A_27_47#_c_73_n 0.00127129f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_46 N_A_M1001_g N_A_27_47#_c_80_n 0.0196498f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_47 A N_A_27_47#_c_80_n 0.00690389f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_48 N_A_c_41_n N_A_27_47#_c_80_n 3.19113e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_49 A N_A_27_47#_c_81_n 0.0145573f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A_c_41_n N_A_27_47#_c_81_n 0.00123585f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_M1001_g N_A_27_47#_c_82_n 0.00337476f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_52 N_A_c_41_n N_A_27_47#_c_74_n 0.00337476f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_M1004_g N_A_27_47#_c_75_n 0.00337476f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_54 A N_A_27_47#_c_75_n 0.0196676f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_55 A N_A_27_47#_c_76_n 3.3412e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_c_41_n N_A_27_47#_c_76_n 0.0210574f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_M1001_g N_VPWR_c_149_n 0.00291026f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_58 N_A_M1001_g N_VPWR_c_152_n 0.00545548f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_148_n 0.0109879f $X=0.47 $Y=2.125 $X2=0 $Y2=0
cc_60 N_A_M1004_g N_VGND_c_201_n 0.00316741f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_VGND_c_204_n 0.00425094f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_62 N_A_M1004_g N_VGND_c_207_n 0.00677097f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_63 N_A_27_47#_c_80_n N_VPWR_M1001_d 0.00584788f $X=0.72 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_64 N_A_27_47#_c_82_n N_VPWR_M1001_d 5.70224e-19 $X=0.805 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_27_47#_M1000_g N_VPWR_c_149_n 0.0103255f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_27_47#_M1002_g N_VPWR_c_149_n 7.08894e-19 $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_67 N_A_27_47#_c_79_n N_VPWR_c_149_n 0.00127645f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_68 N_A_27_47#_c_80_n N_VPWR_c_149_n 0.0210439f $X=0.72 $Y=1.62 $X2=0 $Y2=0
cc_69 N_A_27_47#_c_76_n N_VPWR_c_149_n 3.28752e-19 $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_27_47#_M1002_g N_VPWR_c_151_n 0.00313486f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_71 N_A_27_47#_c_79_n N_VPWR_c_152_n 0.0120448f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_72 N_A_27_47#_M1000_g N_VPWR_c_153_n 0.00505556f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_73 N_A_27_47#_M1002_g N_VPWR_c_153_n 0.0054895f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_27_47#_M1000_g N_VPWR_c_148_n 0.00858194f $X=0.945 $Y=1.985 $X2=0
+ $Y2=0
cc_75 N_A_27_47#_M1002_g N_VPWR_c_148_n 0.0106843f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_79_n N_VPWR_c_148_n 0.00646998f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_71_n N_X_c_179_n 0.00231511f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_76_n N_X_c_179_n 0.0015213f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_27_47#_M1002_g N_X_c_181_n 0.00190975f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_76_n N_X_c_181_n 0.00145049f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_70_n N_X_c_177_n 0.00114857f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_27_47#_M1000_g N_X_c_177_n 0.00163853f $X=0.945 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_71_n N_X_c_177_n 0.0049544f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_27_47#_M1002_g N_X_c_177_n 0.00886214f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_80_n N_X_c_177_n 0.00141452f $X=0.72 $Y=1.62 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_82_n N_X_c_177_n 0.0109809f $X=0.805 $Y=1.535 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_74_n N_X_c_177_n 0.0230865f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_75_n N_X_c_177_n 0.00859268f $X=0.847 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_76_n N_X_c_177_n 0.0248224f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_71_n X 0.00574565f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_27_47#_M1002_g X 0.00916849f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_72_n N_VGND_M1004_d 0.00596397f $X=0.72 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_27_47#_c_75_n N_VGND_M1004_d 9.19341e-19 $X=0.847 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_27_47#_c_70_n N_VGND_c_201_n 0.00627222f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_71_n N_VGND_c_201_n 6.06599e-19 $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_72_n N_VGND_c_201_n 0.0182694f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_76_n N_VGND_c_201_n 3.34628e-19 $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_71_n N_VGND_c_203_n 0.00402932f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_139_p N_VGND_c_204_n 0.01143f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_72_n N_VGND_c_204_n 0.00307419f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_70_n N_VGND_c_205_n 0.00505556f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_71_n N_VGND_c_205_n 0.0054895f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_27_47#_M1004_s N_VGND_c_207_n 0.00369894f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_70_n N_VGND_c_207_n 0.00858194f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_71_n N_VGND_c_207_n 0.0106843f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_139_p N_VGND_c_207_n 0.00643448f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_72_n N_VGND_c_207_n 0.00682895f $X=0.72 $Y=0.72 $X2=0 $Y2=0
cc_108 N_VPWR_c_148_n N_X_M1000_s 0.00359141f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_109 N_VPWR_c_153_n X 0.0151965f $X=1.49 $Y=2.72 $X2=0 $Y2=0
cc_110 N_VPWR_c_148_n X 0.00963372f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_111 N_VPWR_c_151_n N_VGND_c_203_n 0.00998951f $X=1.575 $Y=1.66 $X2=0 $Y2=0
cc_112 X N_VGND_c_203_n 0.0248733f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_113 X N_VGND_c_205_n 0.0151383f $X=1.06 $Y=0.425 $X2=0 $Y2=0
cc_114 N_X_M1003_s N_VGND_c_207_n 0.00359141f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_115 X N_VGND_c_207_n 0.00961963f $X=1.06 $Y=0.425 $X2=0 $Y2=0

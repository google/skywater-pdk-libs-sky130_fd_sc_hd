* File: sky130_fd_sc_hd__or4bb_4.pxi.spice
* Created: Tue Sep  1 19:29:12 2020
* 
x_PM_SKY130_FD_SC_HD__OR4BB_4%C_N N_C_N_M1017_g N_C_N_M1014_g C_N C_N
+ N_C_N_c_112_n N_C_N_c_113_n N_C_N_c_114_n PM_SKY130_FD_SC_HD__OR4BB_4%C_N
x_PM_SKY130_FD_SC_HD__OR4BB_4%D_N N_D_N_M1016_g N_D_N_M1018_g D_N N_D_N_c_146_n
+ N_D_N_c_147_n PM_SKY130_FD_SC_HD__OR4BB_4%D_N
x_PM_SKY130_FD_SC_HD__OR4BB_4%A_205_93# N_A_205_93#_M1016_d N_A_205_93#_M1018_d
+ N_A_205_93#_c_179_n N_A_205_93#_M1004_g N_A_205_93#_M1002_g
+ N_A_205_93#_c_180_n N_A_205_93#_c_181_n N_A_205_93#_c_188_n
+ N_A_205_93#_c_189_n N_A_205_93#_c_182_n N_A_205_93#_c_183_n
+ N_A_205_93#_c_184_n PM_SKY130_FD_SC_HD__OR4BB_4%A_205_93#
x_PM_SKY130_FD_SC_HD__OR4BB_4%A_27_410# N_A_27_410#_M1014_s N_A_27_410#_M1017_s
+ N_A_27_410#_M1007_g N_A_27_410#_M1003_g N_A_27_410#_c_245_n
+ N_A_27_410#_c_252_n N_A_27_410#_c_253_n N_A_27_410#_c_254_n
+ N_A_27_410#_c_255_n N_A_27_410#_c_256_n N_A_27_410#_c_246_n
+ N_A_27_410#_c_247_n N_A_27_410#_c_248_n N_A_27_410#_c_259_n
+ N_A_27_410#_c_249_n PM_SKY130_FD_SC_HD__OR4BB_4%A_27_410#
x_PM_SKY130_FD_SC_HD__OR4BB_4%B N_B_c_332_n N_B_M1005_g N_B_M1000_g N_B_c_333_n
+ N_B_c_334_n B B B PM_SKY130_FD_SC_HD__OR4BB_4%B
x_PM_SKY130_FD_SC_HD__OR4BB_4%A N_A_M1011_g N_A_M1019_g A N_A_c_371_n
+ N_A_c_372_n N_A_c_373_n PM_SKY130_FD_SC_HD__OR4BB_4%A
x_PM_SKY130_FD_SC_HD__OR4BB_4%A_315_380# N_A_315_380#_M1004_d
+ N_A_315_380#_M1005_d N_A_315_380#_M1002_s N_A_315_380#_c_412_n
+ N_A_315_380#_M1008_g N_A_315_380#_M1001_g N_A_315_380#_c_413_n
+ N_A_315_380#_M1009_g N_A_315_380#_M1006_g N_A_315_380#_c_414_n
+ N_A_315_380#_M1012_g N_A_315_380#_M1010_g N_A_315_380#_c_415_n
+ N_A_315_380#_M1015_g N_A_315_380#_M1013_g N_A_315_380#_c_424_n
+ N_A_315_380#_c_416_n N_A_315_380#_c_441_n N_A_315_380#_c_455_n
+ N_A_315_380#_c_442_n N_A_315_380#_c_544_p N_A_315_380#_c_467_n
+ N_A_315_380#_c_417_n N_A_315_380#_c_418_n N_A_315_380#_c_495_p
+ N_A_315_380#_c_462_n N_A_315_380#_c_419_n
+ PM_SKY130_FD_SC_HD__OR4BB_4%A_315_380#
x_PM_SKY130_FD_SC_HD__OR4BB_4%VPWR N_VPWR_M1017_d N_VPWR_M1019_d N_VPWR_M1006_s
+ N_VPWR_M1013_s N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n VPWR N_VPWR_c_566_n N_VPWR_c_567_n
+ N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_559_n
+ PM_SKY130_FD_SC_HD__OR4BB_4%VPWR
x_PM_SKY130_FD_SC_HD__OR4BB_4%X N_X_M1008_d N_X_M1012_d N_X_M1001_d N_X_M1010_d
+ N_X_c_646_n N_X_c_687_n N_X_c_655_n N_X_c_647_n N_X_c_640_n N_X_c_641_n
+ N_X_c_670_n N_X_c_691_n N_X_c_648_n N_X_c_642_n N_X_c_643_n N_X_c_649_n X
+ N_X_c_645_n PM_SKY130_FD_SC_HD__OR4BB_4%X
x_PM_SKY130_FD_SC_HD__OR4BB_4%VGND N_VGND_M1014_d N_VGND_M1004_s N_VGND_M1007_d
+ N_VGND_M1011_d N_VGND_M1009_s N_VGND_M1015_s N_VGND_c_714_n N_VGND_c_715_n
+ N_VGND_c_716_n N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n N_VGND_c_720_n
+ N_VGND_c_721_n N_VGND_c_722_n VGND N_VGND_c_723_n N_VGND_c_724_n
+ N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n
+ N_VGND_c_730_n N_VGND_c_731_n PM_SKY130_FD_SC_HD__OR4BB_4%VGND
cc_1 VNB N_C_N_c_112_n 0.023245f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_2 VNB N_C_N_c_113_n 0.00603475f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_C_N_c_114_n 0.0208027f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_4 VNB D_N 0.0023067f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_5 VNB N_D_N_c_146_n 0.026211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_D_N_c_147_n 0.0189641f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_7 VNB N_A_205_93#_c_179_n 0.0190119f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=0.675
cc_8 VNB N_A_205_93#_c_180_n 0.0252082f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_9 VNB N_A_205_93#_c_181_n 0.00975485f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_10 VNB N_A_205_93#_c_182_n 0.0111553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_205_93#_c_183_n 0.00338114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_205_93#_c_184_n 0.00280828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_c_245_n 0.0222773f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_14 VNB N_A_27_410#_c_246_n 6.47944e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_410#_c_247_n 0.022675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_410#_c_248_n 0.0186165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_410#_c_249_n 0.0171358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_332_n 0.0162189f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_19 VNB N_B_c_333_n 0.00583329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_c_334_n 0.0186258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_c_371_n 0.0229306f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_22 VNB N_A_c_372_n 6.43385e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_23 VNB N_A_c_373_n 0.0174079f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_24 VNB N_A_315_380#_c_412_n 0.0163299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_315_380#_c_413_n 0.0157937f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_26 VNB N_A_315_380#_c_414_n 0.0157971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_315_380#_c_415_n 0.0191578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_315_380#_c_416_n 0.00293881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_315_380#_c_417_n 0.00157854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_315_380#_c_418_n 0.00376665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_315_380#_c_419_n 0.0647168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_559_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_640_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_641_n 0.00187124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_642_n 0.00105843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_643_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB X 0.0199442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_645_n 0.00846039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_714_n 0.0151127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_715_n 0.00882935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_716_n 0.0145978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_717_n 3.29237e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_718_n 0.00239633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_719_n 0.0148447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_720_n 0.0035091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_721_n 0.0106873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_722_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_723_n 0.0196515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_724_n 0.0135943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_725_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_726_n 0.0242387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_727_n 0.00507259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_728_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_729_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_730_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_731_n 0.296148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VPB N_C_N_M1017_g 0.0560403f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.26
cc_58 VPB N_C_N_c_112_n 0.00472379f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_59 VPB N_C_N_c_113_n 0.0023481f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_60 VPB N_D_N_M1018_g 0.0229391f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.675
cc_61 VPB D_N 5.12388e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_62 VPB N_D_N_c_146_n 0.00583771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_205_93#_M1002_g 0.022559f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_64 VPB N_A_205_93#_c_180_n 0.0112048f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_65 VPB N_A_205_93#_c_181_n 0.00131448f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_66 VPB N_A_205_93#_c_188_n 0.00888098f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.325
cc_67 VPB N_A_205_93#_c_189_n 0.00354994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_205_93#_c_183_n 0.00175284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_410#_M1003_g 0.0191524f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_70 VPB N_A_27_410#_c_245_n 0.026212f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_71 VPB N_A_27_410#_c_252_n 0.016454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_410#_c_253_n 0.00753281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_410#_c_254_n 0.00711414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_410#_c_255_n 0.00769888f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_410#_c_256_n 0.00384172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_410#_c_246_n 0.00102304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_410#_c_247_n 0.00583162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_410#_c_259_n 0.0113037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_B_M1000_g 0.0174072f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.675
cc_80 VPB N_B_c_333_n 0.00536776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_B_c_334_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB B 2.2639e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_83 VPB N_A_M1019_g 0.0193215f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.675
cc_84 VPB A 0.00385897f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_85 VPB N_A_c_371_n 0.00445127f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_86 VPB N_A_c_372_n 0.00148828f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_87 VPB N_A_315_380#_M1001_g 0.0199018f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_88 VPB N_A_315_380#_M1006_g 0.0182214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_315_380#_M1010_g 0.0182002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_315_380#_M1013_g 0.0219116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_315_380#_c_424_n 0.00301662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_315_380#_c_416_n 0.00111305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_315_380#_c_419_n 0.0102664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_560_n 0.00735188f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_95 VPB N_VPWR_c_561_n 0.00463796f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.19
cc_96 VPB N_VPWR_c_562_n 0.0181285f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.53
cc_97 VPB N_VPWR_c_563_n 0.00399514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_564_n 0.0112901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_565_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_566_n 0.0145108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_567_n 0.0649032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_568_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_569_n 0.00519112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_570_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_571_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_559_n 0.0544428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_X_c_646_n 0.00246856f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_108 VPB N_X_c_647_n 0.00252706f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.53
cc_109 VPB N_X_c_648_n 0.01047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_X_c_649_n 0.00220075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB X 0.00743877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 N_C_N_M1017_g N_D_N_M1018_g 0.0243394f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_113 N_C_N_c_113_n N_D_N_M1018_g 0.00410692f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_114 N_C_N_c_112_n D_N 2.85663e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C_N_c_113_n D_N 0.0259635f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_N_c_112_n N_D_N_c_146_n 0.019221f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_117 N_C_N_c_113_n N_D_N_c_146_n 0.00225922f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C_N_c_114_n N_D_N_c_147_n 0.0104665f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_119 N_C_N_c_113_n N_A_205_93#_c_188_n 0.011488f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C_N_c_113_n N_A_205_93#_c_183_n 0.00634775f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C_N_M1017_g N_A_27_410#_c_245_n 0.0132977f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_122 N_C_N_c_112_n N_A_27_410#_c_245_n 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_123 N_C_N_c_113_n N_A_27_410#_c_245_n 0.0528067f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C_N_c_114_n N_A_27_410#_c_245_n 0.0052679f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_125 N_C_N_M1017_g N_A_27_410#_c_252_n 0.00143901f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_126 N_C_N_M1017_g N_A_27_410#_c_253_n 0.0143338f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_127 N_C_N_c_112_n N_A_27_410#_c_253_n 8.32653e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_128 N_C_N_c_113_n N_A_27_410#_c_253_n 0.0279958f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_129 N_C_N_M1017_g N_A_27_410#_c_254_n 0.00257483f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_130 N_C_N_c_114_n N_A_27_410#_c_248_n 3.39179e-19 $X=0.51 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_C_N_c_113_n N_VPWR_M1017_d 0.00432228f $X=0.51 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_132 N_C_N_M1017_g N_VPWR_c_560_n 0.0100087f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_133 N_C_N_M1017_g N_VPWR_c_566_n 0.00334979f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_134 N_C_N_M1017_g N_VPWR_c_559_n 0.0048928f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_135 N_C_N_c_113_n N_VGND_c_714_n 0.0108718f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_136 N_C_N_c_114_n N_VGND_c_714_n 0.00422719f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_137 N_C_N_c_114_n N_VGND_c_726_n 0.00510437f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_138 N_C_N_c_114_n N_VGND_c_731_n 0.00512902f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_139 D_N N_A_205_93#_c_180_n 9.47065e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_140 N_D_N_c_146_n N_A_205_93#_c_180_n 0.0150223f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_141 N_D_N_M1018_g N_A_205_93#_c_188_n 0.00312367f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_142 D_N N_A_205_93#_c_188_n 0.0141649f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_143 N_D_N_c_146_n N_A_205_93#_c_188_n 0.00349053f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_144 N_D_N_M1018_g N_A_205_93#_c_189_n 0.00312224f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_145 D_N N_A_205_93#_c_182_n 0.012483f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_146 N_D_N_c_146_n N_A_205_93#_c_182_n 0.00272654f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_147 N_D_N_c_147_n N_A_205_93#_c_182_n 3.44947e-19 $X=1.03 $Y=0.995 $X2=0
+ $Y2=0
cc_148 D_N N_A_205_93#_c_183_n 0.0269017f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_149 N_D_N_c_146_n N_A_205_93#_c_183_n 0.00101647f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_150 N_D_N_c_147_n N_A_205_93#_c_184_n 0.0042717f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_151 N_D_N_M1018_g N_A_27_410#_c_253_n 0.0147166f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_152 D_N N_A_27_410#_c_253_n 0.00124584f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_153 N_D_N_M1018_g N_A_315_380#_c_424_n 3.47028e-19 $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_154 N_D_N_M1018_g N_VPWR_c_567_n 0.00259183f $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_155 N_D_N_M1018_g N_VPWR_c_559_n 0.00417489f $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_156 N_D_N_c_147_n N_VGND_c_714_n 0.00290717f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_157 N_D_N_c_147_n N_VGND_c_715_n 0.00311391f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_158 N_D_N_c_147_n N_VGND_c_723_n 0.00510437f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_159 N_D_N_c_147_n N_VGND_c_731_n 0.00512902f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_205_93#_M1002_g N_A_27_410#_M1003_g 0.0419995f $X=1.91 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_205_93#_M1018_d N_A_27_410#_c_253_n 0.00214482f $X=1.03 $Y=1.485
+ $X2=0 $Y2=0
cc_162 N_A_205_93#_c_188_n N_A_27_410#_c_253_n 0.0191176f $X=1.405 $Y=1.61 $X2=0
+ $Y2=0
cc_163 N_A_205_93#_M1002_g N_A_27_410#_c_254_n 0.00269181f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_164 N_A_205_93#_M1002_g N_A_27_410#_c_255_n 0.0120949f $X=1.91 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_205_93#_c_188_n N_A_27_410#_c_255_n 0.0070528f $X=1.405 $Y=1.61 $X2=0
+ $Y2=0
cc_166 N_A_205_93#_M1002_g N_A_27_410#_c_246_n 0.00516899f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_167 N_A_205_93#_c_181_n N_A_27_410#_c_246_n 3.09204e-19 $X=1.9 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_205_93#_c_181_n N_A_27_410#_c_247_n 0.017052f $X=1.9 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_A_205_93#_c_179_n N_A_27_410#_c_249_n 0.019656f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_205_93#_c_188_n N_A_315_380#_M1002_s 0.00232997f $X=1.405 $Y=1.61
+ $X2=0 $Y2=0
cc_171 N_A_205_93#_c_189_n N_A_315_380#_M1002_s 4.62701e-19 $X=1.5 $Y=1.525
+ $X2=0 $Y2=0
cc_172 N_A_205_93#_M1002_g N_A_315_380#_c_424_n 0.0101303f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_173 N_A_205_93#_c_180_n N_A_315_380#_c_424_n 0.00348139f $X=1.815 $Y=1.16
+ $X2=0 $Y2=0
cc_174 N_A_205_93#_c_188_n N_A_315_380#_c_424_n 0.0052433f $X=1.405 $Y=1.61
+ $X2=0 $Y2=0
cc_175 N_A_205_93#_c_183_n N_A_315_380#_c_424_n 0.00260172f $X=1.61 $Y=1.16
+ $X2=0 $Y2=0
cc_176 N_A_205_93#_c_179_n N_A_315_380#_c_416_n 0.00427172f $X=1.89 $Y=0.995
+ $X2=0 $Y2=0
cc_177 N_A_205_93#_M1002_g N_A_315_380#_c_416_n 0.0207589f $X=1.91 $Y=1.985
+ $X2=0 $Y2=0
cc_178 N_A_205_93#_c_181_n N_A_315_380#_c_416_n 0.00916997f $X=1.9 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_205_93#_c_188_n N_A_315_380#_c_416_n 0.00780797f $X=1.405 $Y=1.61
+ $X2=0 $Y2=0
cc_180 N_A_205_93#_c_189_n N_A_315_380#_c_416_n 0.00849713f $X=1.5 $Y=1.525
+ $X2=0 $Y2=0
cc_181 N_A_205_93#_c_183_n N_A_315_380#_c_416_n 0.0177065f $X=1.61 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A_205_93#_c_184_n N_A_315_380#_c_416_n 0.0071734f $X=1.55 $Y=0.995
+ $X2=0 $Y2=0
cc_183 N_A_205_93#_c_179_n N_A_315_380#_c_441_n 0.00541038f $X=1.89 $Y=0.995
+ $X2=0 $Y2=0
cc_184 N_A_205_93#_c_179_n N_A_315_380#_c_442_n 0.00588026f $X=1.89 $Y=0.995
+ $X2=0 $Y2=0
cc_185 N_A_205_93#_c_182_n N_A_315_380#_c_442_n 0.00841187f $X=1.16 $Y=0.66
+ $X2=0 $Y2=0
cc_186 N_A_205_93#_M1002_g N_VPWR_c_567_n 0.00357877f $X=1.91 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_205_93#_M1002_g N_VPWR_c_559_n 0.00688262f $X=1.91 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_205_93#_c_182_n N_VGND_M1004_s 0.00275812f $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_189 N_A_205_93#_c_184_n N_VGND_M1004_s 6.72012e-19 $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_205_93#_c_182_n N_VGND_c_714_n 8.07382e-19 $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_191 N_A_205_93#_c_179_n N_VGND_c_715_n 0.01001f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_205_93#_c_180_n N_VGND_c_715_n 0.00364602f $X=1.815 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_A_205_93#_c_182_n N_VGND_c_715_n 0.00836503f $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_194 N_A_205_93#_c_183_n N_VGND_c_715_n 0.00340568f $X=1.61 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_205_93#_c_179_n N_VGND_c_716_n 0.00435058f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_205_93#_c_179_n N_VGND_c_717_n 6.75279e-19 $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_205_93#_c_182_n N_VGND_c_723_n 0.0100997f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_198 N_A_205_93#_c_179_n N_VGND_c_731_n 0.00726129f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_205_93#_c_182_n N_VGND_c_731_n 0.0138693f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_200 N_A_27_410#_c_249_n N_B_c_332_n 0.0251622f $X=2.36 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_201 N_A_27_410#_M1003_g N_B_M1000_g 0.0548318f $X=2.42 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_27_410#_c_255_n N_B_M1000_g 7.55916e-19 $X=2.275 $Y=2.38 $X2=0 $Y2=0
cc_203 N_A_27_410#_c_246_n N_B_M1000_g 0.00278336f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_27_410#_c_246_n N_B_c_333_n 0.0274089f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_27_410#_c_247_n N_B_c_333_n 0.00284781f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_27_410#_c_246_n N_B_c_334_n 3.68507e-19 $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_27_410#_c_247_n N_B_c_334_n 0.0203414f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_27_410#_M1003_g B 0.00302042f $X=2.42 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_27_410#_c_255_n B 0.0035615f $X=2.275 $Y=2.38 $X2=0 $Y2=0
cc_210 N_A_27_410#_c_246_n B 0.0332087f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_27_410#_c_255_n N_A_315_380#_M1002_s 0.00480304f $X=2.275 $Y=2.38
+ $X2=0 $Y2=0
cc_212 N_A_27_410#_M1003_g N_A_315_380#_c_424_n 5.92223e-19 $X=2.42 $Y=1.985
+ $X2=0 $Y2=0
cc_213 N_A_27_410#_c_253_n N_A_315_380#_c_424_n 0.00620564f $X=1.125 $Y=1.95
+ $X2=0 $Y2=0
cc_214 N_A_27_410#_c_254_n N_A_315_380#_c_424_n 0.00626935f $X=1.21 $Y=2.295
+ $X2=0 $Y2=0
cc_215 N_A_27_410#_c_255_n N_A_315_380#_c_424_n 0.0331132f $X=2.275 $Y=2.38
+ $X2=0 $Y2=0
cc_216 N_A_27_410#_c_246_n N_A_315_380#_c_424_n 0.0136829f $X=2.36 $Y=1.16 $X2=0
+ $Y2=0
cc_217 N_A_27_410#_M1003_g N_A_315_380#_c_416_n 0.00179169f $X=2.42 $Y=1.985
+ $X2=0 $Y2=0
cc_218 N_A_27_410#_c_253_n N_A_315_380#_c_416_n 0.00266088f $X=1.125 $Y=1.95
+ $X2=0 $Y2=0
cc_219 N_A_27_410#_c_246_n N_A_315_380#_c_416_n 0.0697478f $X=2.36 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_A_27_410#_c_247_n N_A_315_380#_c_416_n 0.00201257f $X=2.36 $Y=1.16
+ $X2=0 $Y2=0
cc_221 N_A_27_410#_c_249_n N_A_315_380#_c_416_n 0.00338056f $X=2.36 $Y=0.995
+ $X2=0 $Y2=0
cc_222 N_A_27_410#_c_246_n N_A_315_380#_c_455_n 0.0108856f $X=2.36 $Y=1.16 $X2=0
+ $Y2=0
cc_223 N_A_27_410#_c_247_n N_A_315_380#_c_455_n 3.62043e-19 $X=2.36 $Y=1.16
+ $X2=0 $Y2=0
cc_224 N_A_27_410#_c_249_n N_A_315_380#_c_455_n 0.0131138f $X=2.36 $Y=0.995
+ $X2=0 $Y2=0
cc_225 N_A_27_410#_c_247_n N_A_315_380#_c_442_n 0.00189854f $X=2.36 $Y=1.16
+ $X2=0 $Y2=0
cc_226 N_A_27_410#_c_253_n N_VPWR_M1017_d 0.00538813f $X=1.125 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_227 N_A_27_410#_c_253_n N_VPWR_c_560_n 0.0229102f $X=1.125 $Y=1.95 $X2=0
+ $Y2=0
cc_228 N_A_27_410#_c_254_n N_VPWR_c_560_n 0.00501924f $X=1.21 $Y=2.295 $X2=0
+ $Y2=0
cc_229 N_A_27_410#_c_256_n N_VPWR_c_560_n 0.0106159f $X=1.295 $Y=2.38 $X2=0
+ $Y2=0
cc_230 N_A_27_410#_c_252_n N_VPWR_c_566_n 0.0168632f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_231 N_A_27_410#_c_253_n N_VPWR_c_566_n 0.00256078f $X=1.125 $Y=1.95 $X2=0
+ $Y2=0
cc_232 N_A_27_410#_M1003_g N_VPWR_c_567_n 0.00433573f $X=2.42 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_27_410#_c_253_n N_VPWR_c_567_n 0.00431784f $X=1.125 $Y=1.95 $X2=0
+ $Y2=0
cc_234 N_A_27_410#_c_255_n N_VPWR_c_567_n 0.0685563f $X=2.275 $Y=2.38 $X2=0
+ $Y2=0
cc_235 N_A_27_410#_c_256_n N_VPWR_c_567_n 0.0120734f $X=1.295 $Y=2.38 $X2=0
+ $Y2=0
cc_236 N_A_27_410#_M1003_g N_VPWR_c_559_n 0.00738288f $X=2.42 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_27_410#_c_252_n N_VPWR_c_559_n 0.00987599f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_238 N_A_27_410#_c_253_n N_VPWR_c_559_n 0.0128853f $X=1.125 $Y=1.95 $X2=0
+ $Y2=0
cc_239 N_A_27_410#_c_255_n N_VPWR_c_559_n 0.0418903f $X=2.275 $Y=2.38 $X2=0
+ $Y2=0
cc_240 N_A_27_410#_c_256_n N_VPWR_c_559_n 0.00652563f $X=1.295 $Y=2.38 $X2=0
+ $Y2=0
cc_241 N_A_27_410#_c_255_n A_397_297# 0.00940368f $X=2.275 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_242 N_A_27_410#_c_246_n A_397_297# 0.00775786f $X=2.36 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_27_410#_c_248_n N_VGND_c_714_n 0.0104991f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_244 N_A_27_410#_c_249_n N_VGND_c_715_n 6.60171e-19 $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_27_410#_c_249_n N_VGND_c_716_n 0.00341689f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_27_410#_c_249_n N_VGND_c_717_n 0.00770433f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_27_410#_c_248_n N_VGND_c_726_n 0.00957361f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_248 N_A_27_410#_c_248_n N_VGND_c_731_n 0.0105585f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_249 N_A_27_410#_c_249_n N_VGND_c_731_n 0.00431054f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_B_M1000_g N_A_M1019_g 0.0564998f $X=2.84 $Y=1.985 $X2=0 $Y2=0
cc_251 B N_A_M1019_g 0.00915664f $X=2.925 $Y=1.785 $X2=0 $Y2=0
cc_252 N_B_c_333_n A 0.0102741f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_253 N_B_c_333_n N_A_c_371_n 0.00373575f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B_c_334_n N_A_c_371_n 0.0203414f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B_c_333_n N_A_c_372_n 0.0271074f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B_c_334_n N_A_c_372_n 3.68507e-19 $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B_c_332_n N_A_c_373_n 0.0243955f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B_c_332_n N_A_315_380#_c_455_n 0.0110728f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_259 N_B_c_333_n N_A_315_380#_c_455_n 0.018276f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B_c_334_n N_A_315_380#_c_455_n 2.98597e-19 $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B_c_333_n N_A_315_380#_c_462_n 0.00316818f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_262 B N_VPWR_c_561_n 0.031049f $X=2.925 $Y=1.785 $X2=0 $Y2=0
cc_263 N_B_M1000_g N_VPWR_c_567_n 0.00419108f $X=2.84 $Y=1.985 $X2=0 $Y2=0
cc_264 B N_VPWR_c_567_n 0.0126498f $X=2.925 $Y=1.785 $X2=0 $Y2=0
cc_265 N_B_M1000_g N_VPWR_c_559_n 0.00651073f $X=2.84 $Y=1.985 $X2=0 $Y2=0
cc_266 B N_VPWR_c_559_n 0.0110804f $X=2.925 $Y=1.785 $X2=0 $Y2=0
cc_267 B A_583_297# 0.0164072f $X=2.925 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_268 N_B_c_332_n N_VGND_c_717_n 0.00732663f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B_c_332_n N_VGND_c_724_n 0.00341689f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B_c_332_n N_VGND_c_731_n 0.00405445f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_c_373_n N_A_315_380#_c_412_n 0.0200495f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_M1019_g N_A_315_380#_M1001_g 0.0173803f $X=3.26 $Y=1.985 $X2=0 $Y2=0
cc_273 A N_A_315_380#_M1001_g 0.00128363f $X=3.385 $Y=1.445 $X2=0 $Y2=0
cc_274 N_A_c_372_n N_A_315_380#_M1001_g 0.00219223f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_275 A N_A_315_380#_c_467_n 0.00495213f $X=3.385 $Y=1.445 $X2=0 $Y2=0
cc_276 N_A_c_371_n N_A_315_380#_c_467_n 0.00173573f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_c_372_n N_A_315_380#_c_467_n 0.0104547f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_278 N_A_c_373_n N_A_315_380#_c_467_n 0.0134819f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_c_371_n N_A_315_380#_c_417_n 5.07416e-19 $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_c_372_n N_A_315_380#_c_417_n 0.00568393f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_281 N_A_c_373_n N_A_315_380#_c_417_n 0.00336447f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_282 A N_A_315_380#_c_418_n 0.00707041f $X=3.385 $Y=1.445 $X2=0 $Y2=0
cc_283 N_A_c_371_n N_A_315_380#_c_418_n 0.00124527f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_c_372_n N_A_315_380#_c_418_n 0.0137152f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_c_371_n N_A_315_380#_c_419_n 0.0161964f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_c_372_n N_A_315_380#_c_419_n 7.74805e-19 $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_287 A N_VPWR_M1019_d 0.00433176f $X=3.385 $Y=1.445 $X2=0 $Y2=0
cc_288 N_A_M1019_g N_VPWR_c_561_n 0.00789297f $X=3.26 $Y=1.985 $X2=0 $Y2=0
cc_289 A N_VPWR_c_561_n 0.0193325f $X=3.385 $Y=1.445 $X2=0 $Y2=0
cc_290 N_A_M1019_g N_VPWR_c_567_n 0.00585385f $X=3.26 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_M1019_g N_VPWR_c_559_n 0.0109527f $X=3.26 $Y=1.985 $X2=0 $Y2=0
cc_292 A N_X_c_646_n 0.00229946f $X=3.385 $Y=1.445 $X2=0 $Y2=0
cc_293 N_A_c_373_n N_VGND_c_717_n 6.8876e-19 $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_c_373_n N_VGND_c_718_n 0.00318791f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_c_373_n N_VGND_c_724_n 0.00428022f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_c_373_n N_VGND_c_731_n 0.00603983f $X=3.32 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A_315_380#_M1001_g N_VPWR_c_561_n 0.00430866f $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_315_380#_M1001_g N_VPWR_c_562_n 0.00585385f $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_315_380#_M1006_g N_VPWR_c_562_n 0.00585385f $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A_315_380#_M1006_g N_VPWR_c_563_n 0.00165046f $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A_315_380#_M1010_g N_VPWR_c_563_n 0.00157837f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A_315_380#_M1013_g N_VPWR_c_565_n 0.00338128f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_315_380#_M1010_g N_VPWR_c_568_n 0.00585385f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A_315_380#_M1013_g N_VPWR_c_568_n 0.00585385f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_A_315_380#_M1002_s N_VPWR_c_559_n 0.00210147f $X=1.575 $Y=1.9 $X2=0
+ $Y2=0
cc_306 N_A_315_380#_M1001_g N_VPWR_c_559_n 0.0108486f $X=3.79 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_A_315_380#_M1006_g N_VPWR_c_559_n 0.0104367f $X=4.21 $Y=1.985 $X2=0
+ $Y2=0
cc_308 N_A_315_380#_M1010_g N_VPWR_c_559_n 0.0104367f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_315_380#_M1013_g N_VPWR_c_559_n 0.011391f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_315_380#_c_424_n A_397_297# 0.00215179f $X=1.935 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_311 N_A_315_380#_c_416_n A_397_297# 0.00402758f $X=2.02 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_312 N_A_315_380#_M1001_g N_X_c_646_n 2.80238e-19 $X=3.79 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A_315_380#_c_495_p N_X_c_646_n 0.0172286f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_315_380#_c_419_n N_X_c_646_n 0.00226413f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_315_380#_c_413_n N_X_c_655_n 0.00701434f $X=4.21 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A_315_380#_c_414_n N_X_c_655_n 5.23786e-19 $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_315_380#_M1006_g N_X_c_647_n 0.0134538f $X=4.21 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A_315_380#_M1010_g N_X_c_647_n 0.013468f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A_315_380#_c_495_p N_X_c_647_n 0.03482f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_315_380#_c_419_n N_X_c_647_n 0.00216069f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_315_380#_c_413_n N_X_c_640_n 0.00870364f $X=4.21 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_315_380#_c_414_n N_X_c_640_n 0.00865686f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_315_380#_c_495_p N_X_c_640_n 0.0356734f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A_315_380#_c_419_n N_X_c_640_n 0.00222133f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_315_380#_c_412_n N_X_c_641_n 8.16938e-19 $X=3.79 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_315_380#_c_413_n N_X_c_641_n 0.00250064f $X=4.21 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_315_380#_c_417_n N_X_c_641_n 0.00357582f $X=3.66 $Y=1.075 $X2=0 $Y2=0
cc_328 N_A_315_380#_c_495_p N_X_c_641_n 0.01996f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_315_380#_c_419_n N_X_c_641_n 0.00230339f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_315_380#_c_413_n N_X_c_670_n 5.22228e-19 $X=4.21 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_315_380#_c_414_n N_X_c_670_n 0.00630972f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_315_380#_c_415_n N_X_c_670_n 0.0109314f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_315_380#_M1013_g N_X_c_648_n 0.0158823f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A_315_380#_c_495_p N_X_c_648_n 0.00401279f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_315_380#_c_415_n N_X_c_642_n 0.0113022f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A_315_380#_c_495_p N_X_c_642_n 0.00200821f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_315_380#_c_414_n N_X_c_643_n 0.00113286f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_315_380#_c_415_n N_X_c_643_n 0.00113286f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_315_380#_c_495_p N_X_c_643_n 0.026256f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_315_380#_c_419_n N_X_c_643_n 0.00230339f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_315_380#_c_495_p N_X_c_649_n 0.0172286f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_342 N_A_315_380#_c_419_n N_X_c_649_n 0.00226413f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_315_380#_c_415_n X 0.0211223f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A_315_380#_c_495_p X 0.0137227f $X=4.87 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A_315_380#_c_455_n N_VGND_M1007_d 0.00664072f $X=2.965 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_315_380#_c_467_n N_VGND_M1011_d 0.00616911f $X=3.575 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A_315_380#_c_417_n N_VGND_M1011_d 7.20909e-19 $X=3.66 $Y=1.075 $X2=0
+ $Y2=0
cc_348 N_A_315_380#_c_441_n N_VGND_c_715_n 0.00960696f $X=2.18 $Y=0.49 $X2=0
+ $Y2=0
cc_349 N_A_315_380#_c_441_n N_VGND_c_716_n 0.00852533f $X=2.18 $Y=0.49 $X2=0
+ $Y2=0
cc_350 N_A_315_380#_c_442_n N_VGND_c_716_n 0.00502163f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_351 N_A_315_380#_c_441_n N_VGND_c_717_n 0.0117247f $X=2.18 $Y=0.49 $X2=0
+ $Y2=0
cc_352 N_A_315_380#_c_455_n N_VGND_c_717_n 0.0160613f $X=2.965 $Y=0.74 $X2=0
+ $Y2=0
cc_353 N_A_315_380#_c_412_n N_VGND_c_718_n 0.00675761f $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_315_380#_c_413_n N_VGND_c_718_n 5.99174e-19 $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A_315_380#_c_467_n N_VGND_c_718_n 0.0224385f $X=3.575 $Y=0.74 $X2=0
+ $Y2=0
cc_356 N_A_315_380#_c_412_n N_VGND_c_719_n 0.00496106f $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_315_380#_c_413_n N_VGND_c_719_n 0.00423334f $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_315_380#_c_413_n N_VGND_c_720_n 0.00138579f $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_359 N_A_315_380#_c_414_n N_VGND_c_720_n 0.00146448f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_360 N_A_315_380#_c_415_n N_VGND_c_722_n 0.00316354f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_315_380#_c_455_n N_VGND_c_724_n 0.00232396f $X=2.965 $Y=0.74 $X2=0
+ $Y2=0
cc_362 N_A_315_380#_c_544_p N_VGND_c_724_n 0.00846569f $X=3.05 $Y=0.49 $X2=0
+ $Y2=0
cc_363 N_A_315_380#_c_467_n N_VGND_c_724_n 0.0029785f $X=3.575 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_315_380#_c_414_n N_VGND_c_725_n 0.00423334f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_365 N_A_315_380#_c_415_n N_VGND_c_725_n 0.00423334f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_315_380#_M1004_d N_VGND_c_731_n 0.00390697f $X=1.965 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_315_380#_M1005_d N_VGND_c_731_n 0.00256656f $X=2.915 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_315_380#_c_412_n N_VGND_c_731_n 0.00822344f $X=3.79 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_315_380#_c_413_n N_VGND_c_731_n 0.00575518f $X=4.21 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_315_380#_c_414_n N_VGND_c_731_n 0.0057163f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A_315_380#_c_415_n N_VGND_c_731_n 0.00667051f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A_315_380#_c_441_n N_VGND_c_731_n 0.00618681f $X=2.18 $Y=0.49 $X2=0
+ $Y2=0
cc_373 N_A_315_380#_c_455_n N_VGND_c_731_n 0.00554474f $X=2.965 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_315_380#_c_442_n N_VGND_c_731_n 0.00936859f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_375 N_A_315_380#_c_544_p N_VGND_c_731_n 0.00625722f $X=3.05 $Y=0.49 $X2=0
+ $Y2=0
cc_376 N_A_315_380#_c_467_n N_VGND_c_731_n 0.00734097f $X=3.575 $Y=0.74 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_559_n A_397_297# 0.00289104f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_378 N_VPWR_c_559_n A_499_297# 0.0115413f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_379 N_VPWR_c_559_n A_583_297# 0.0046981f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_380 N_VPWR_c_559_n N_X_M1001_d 0.00284632f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_559_n N_X_M1010_d 0.00284632f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_562_n N_X_c_687_n 0.0142343f $X=4.295 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_559_n N_X_c_687_n 0.00955092f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_M1006_s N_X_c_647_n 0.00165831f $X=4.285 $Y=1.485 $X2=0 $Y2=0
cc_385 N_VPWR_c_563_n N_X_c_647_n 0.0126919f $X=4.42 $Y=1.96 $X2=0 $Y2=0
cc_386 N_VPWR_c_568_n N_X_c_691_n 0.0142343f $X=5.135 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_559_n N_X_c_691_n 0.00955092f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_M1013_s N_X_c_648_n 0.00283464f $X=5.125 $Y=1.485 $X2=0 $Y2=0
cc_389 N_VPWR_c_565_n N_X_c_648_n 0.0179737f $X=5.26 $Y=1.96 $X2=0 $Y2=0
cc_390 N_X_c_640_n N_VGND_M1009_s 0.00162089f $X=4.675 $Y=0.815 $X2=0 $Y2=0
cc_391 N_X_c_642_n N_VGND_M1015_s 2.28588e-19 $X=5.205 $Y=0.815 $X2=0 $Y2=0
cc_392 N_X_c_645_n N_VGND_M1015_s 0.0030148f $X=5.32 $Y=0.905 $X2=0 $Y2=0
cc_393 N_X_c_655_n N_VGND_c_719_n 0.0151398f $X=4 $Y=0.485 $X2=0 $Y2=0
cc_394 N_X_c_640_n N_VGND_c_719_n 0.00198695f $X=4.675 $Y=0.815 $X2=0 $Y2=0
cc_395 N_X_c_640_n N_VGND_c_720_n 0.0122559f $X=4.675 $Y=0.815 $X2=0 $Y2=0
cc_396 N_X_c_645_n N_VGND_c_721_n 0.00149748f $X=5.32 $Y=0.905 $X2=0 $Y2=0
cc_397 N_X_c_642_n N_VGND_c_722_n 0.00177288f $X=5.205 $Y=0.815 $X2=0 $Y2=0
cc_398 N_X_c_645_n N_VGND_c_722_n 0.0120207f $X=5.32 $Y=0.905 $X2=0 $Y2=0
cc_399 N_X_c_640_n N_VGND_c_725_n 0.00198695f $X=4.675 $Y=0.815 $X2=0 $Y2=0
cc_400 N_X_c_670_n N_VGND_c_725_n 0.0188551f $X=4.84 $Y=0.39 $X2=0 $Y2=0
cc_401 N_X_c_642_n N_VGND_c_725_n 0.00198695f $X=5.205 $Y=0.815 $X2=0 $Y2=0
cc_402 N_X_M1008_d N_VGND_c_731_n 0.00393857f $X=3.865 $Y=0.235 $X2=0 $Y2=0
cc_403 N_X_M1012_d N_VGND_c_731_n 0.00215201f $X=4.705 $Y=0.235 $X2=0 $Y2=0
cc_404 N_X_c_655_n N_VGND_c_731_n 0.00940698f $X=4 $Y=0.485 $X2=0 $Y2=0
cc_405 N_X_c_640_n N_VGND_c_731_n 0.00835832f $X=4.675 $Y=0.815 $X2=0 $Y2=0
cc_406 N_X_c_670_n N_VGND_c_731_n 0.0122069f $X=4.84 $Y=0.39 $X2=0 $Y2=0
cc_407 N_X_c_642_n N_VGND_c_731_n 0.00396723f $X=5.205 $Y=0.815 $X2=0 $Y2=0
cc_408 N_X_c_645_n N_VGND_c_731_n 0.00317702f $X=5.32 $Y=0.905 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__xnor3_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__xnor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425000 1.075000 8.835000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.605000 0.995000 7.775000 1.445000 ;
        RECT 7.605000 1.445000 8.185000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 1.075000 3.560000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.375000 0.875000 0.995000 ;
        RECT 0.625000 0.995000 1.710000 1.325000 ;
        RECT 0.625000 1.325000 0.955000 2.425000 ;
        RECT 1.465000 0.350000 1.725000 0.925000 ;
        RECT 1.465000 0.925000 1.710000 0.995000 ;
        RECT 1.465000 1.325000 1.710000 1.440000 ;
        RECT 1.465000 1.440000 1.745000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.285000  0.085000 0.455000 0.735000 ;
        RECT 1.125000  0.085000 1.295000 0.735000 ;
        RECT 1.895000  0.085000 2.145000 0.525000 ;
        RECT 4.855000  0.085000 5.025000 0.865000 ;
        RECT 8.855000  0.085000 9.025000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.285000 1.490000 0.455000 2.635000 ;
        RECT 1.125000 1.495000 1.295000 2.635000 ;
        RECT 1.915000 2.215000 2.250000 2.635000 ;
        RECT 4.605000 2.235000 4.935000 2.635000 ;
        RECT 8.775000 2.275000 9.110000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.880000 0.995000 2.085000 1.325000 ;
      RECT 1.910000 0.695000 2.485000 0.865000 ;
      RECT 1.910000 0.865000 2.085000 0.995000 ;
      RECT 1.915000 1.325000 2.085000 1.875000 ;
      RECT 1.915000 1.875000 2.600000 2.045000 ;
      RECT 2.315000 0.255000 3.885000 0.425000 ;
      RECT 2.315000 0.425000 2.485000 0.695000 ;
      RECT 2.315000 1.535000 3.900000 1.705000 ;
      RECT 2.430000 2.045000 2.600000 2.235000 ;
      RECT 2.430000 2.235000 3.900000 2.405000 ;
      RECT 2.655000 0.595000 2.825000 1.535000 ;
      RECT 2.940000 1.895000 5.440000 2.065000 ;
      RECT 3.125000 0.625000 4.345000 0.795000 ;
      RECT 3.125000 0.795000 3.505000 0.905000 ;
      RECT 3.450000 0.425000 3.885000 0.455000 ;
      RECT 3.730000 0.995000 4.005000 1.325000 ;
      RECT 3.730000 1.325000 3.900000 1.535000 ;
      RECT 4.055000 0.285000 4.685000 0.455000 ;
      RECT 4.070000 1.525000 4.455000 1.695000 ;
      RECT 4.175000 0.795000 4.345000 1.375000 ;
      RECT 4.175000 1.375000 4.455000 1.525000 ;
      RECT 4.515000 0.455000 4.685000 1.035000 ;
      RECT 4.515000 1.035000 4.795000 1.205000 ;
      RECT 4.625000 1.205000 4.795000 1.895000 ;
      RECT 5.025000 1.445000 5.445000 1.715000 ;
      RECT 5.205000 0.415000 5.445000 1.445000 ;
      RECT 5.270000 2.065000 5.440000 2.275000 ;
      RECT 5.270000 2.275000 8.365000 2.445000 ;
      RECT 5.625000 0.265000 6.035000 0.485000 ;
      RECT 5.625000 0.485000 5.835000 0.595000 ;
      RECT 5.625000 0.595000 5.795000 2.105000 ;
      RECT 5.965000 0.720000 6.375000 0.825000 ;
      RECT 5.965000 0.825000 6.175000 0.890000 ;
      RECT 5.965000 0.890000 6.135000 2.275000 ;
      RECT 6.005000 0.655000 6.375000 0.720000 ;
      RECT 6.205000 0.320000 6.375000 0.655000 ;
      RECT 6.315000 1.445000 7.095000 1.615000 ;
      RECT 6.315000 1.615000 6.730000 2.045000 ;
      RECT 6.330000 0.995000 6.755000 1.270000 ;
      RECT 6.545000 0.630000 6.755000 0.995000 ;
      RECT 6.925000 0.255000 8.070000 0.425000 ;
      RECT 6.925000 0.425000 7.095000 1.445000 ;
      RECT 7.265000 0.595000 7.435000 1.935000 ;
      RECT 7.265000 1.935000 9.575000 2.105000 ;
      RECT 7.605000 0.425000 8.070000 0.465000 ;
      RECT 7.945000 0.730000 8.150000 0.945000 ;
      RECT 7.945000 0.945000 8.255000 1.275000 ;
      RECT 8.355000 1.495000 9.175000 1.705000 ;
      RECT 8.395000 0.295000 8.685000 0.735000 ;
      RECT 8.395000 0.735000 9.175000 0.750000 ;
      RECT 8.435000 0.750000 9.175000 0.905000 ;
      RECT 9.005000 0.905000 9.175000 0.995000 ;
      RECT 9.005000 0.995000 9.235000 1.325000 ;
      RECT 9.005000 1.325000 9.175000 1.495000 ;
      RECT 9.090000 1.875000 9.575000 1.935000 ;
      RECT 9.275000 0.255000 9.575000 0.585000 ;
      RECT 9.280000 2.105000 9.575000 2.465000 ;
      RECT 9.405000 0.585000 9.575000 1.875000 ;
    LAYER mcon ;
      RECT 4.285000 1.445000 4.455000 1.615000 ;
      RECT 5.205000 0.765000 5.375000 0.935000 ;
      RECT 5.665000 0.425000 5.835000 0.595000 ;
      RECT 6.585000 0.765000 6.755000 0.935000 ;
      RECT 6.585000 1.445000 6.755000 1.615000 ;
      RECT 7.965000 0.765000 8.135000 0.935000 ;
      RECT 8.425000 0.425000 8.595000 0.595000 ;
    LAYER met1 ;
      RECT 4.225000 1.415000 4.515000 1.460000 ;
      RECT 4.225000 1.460000 6.815000 1.600000 ;
      RECT 4.225000 1.600000 4.515000 1.645000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.780000 8.195000 0.920000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.605000 0.395000 5.895000 0.440000 ;
      RECT 5.605000 0.440000 8.655000 0.580000 ;
      RECT 5.605000 0.580000 5.895000 0.625000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
      RECT 6.525000 1.415000 6.815000 1.460000 ;
      RECT 6.525000 1.600000 6.815000 1.645000 ;
      RECT 7.905000 0.735000 8.195000 0.780000 ;
      RECT 7.905000 0.920000 8.195000 0.965000 ;
      RECT 8.365000 0.395000 8.655000 0.440000 ;
      RECT 8.365000 0.580000 8.655000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_4

* File: sky130_fd_sc_hd__o311a_1.spice.pex
* Created: Thu Aug 27 14:38:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311A_1%A_81_21# 1 2 3 10 12 15 19 20 22 23 25 26 27
+ 29 31 32 33 35 36 38 43
c99 19 0 1.79971e-19 $X=0.69 $Y=1.16
r100 43 45 15.3743 $w=5.83e-07 $l=4.25e-07 $layer=LI1_cond $X=3.302 $Y=0.4
+ $X2=3.302 $Y2=0.825
r101 36 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.45 $Y=1.58
+ $X2=3.095 $Y2=1.58
r102 36 38 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=1.665
+ $X2=3.45 $Y2=1.815
r103 35 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=1.495
+ $X2=3.095 $Y2=1.58
r104 35 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.095 $Y=1.495
+ $X2=3.095 $Y2=0.825
r105 32 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=1.58
+ $X2=3.095 $Y2=1.58
r106 32 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.01 $Y=1.58
+ $X2=2.715 $Y2=1.58
r107 29 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=2.295
+ $X2=2.55 $Y2=2.38
r108 29 31 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.55 $Y=2.295
+ $X2=2.55 $Y2=1.68
r109 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.55 $Y=1.665
+ $X2=2.715 $Y2=1.58
r110 28 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=1.68
r111 26 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=2.38
+ $X2=2.55 $Y2=2.38
r112 26 27 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.385 $Y=2.38
+ $X2=1.35 $Y2=2.38
r113 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.265 $Y=2.295
+ $X2=1.35 $Y2=2.38
r114 24 25 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.265 $Y=1.665
+ $X2=1.265 $Y2=2.295
r115 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=1.58
+ $X2=1.265 $Y2=1.665
r116 22 23 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.18 $Y=1.58
+ $X2=0.775 $Y2=1.58
r117 20 49 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.69 $Y=1.16
+ $X2=0.48 $Y2=1.16
r118 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.16 $X2=0.69 $Y2=1.16
r119 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=1.495
+ $X2=0.775 $Y2=1.58
r120 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=1.495
+ $X2=0.69 $Y2=1.16
r121 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r122 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.985
r123 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r124 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=0.56
r125 3 38 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.815
r126 2 41 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.485 $X2=2.55 $Y2=2.36
r127 2 31 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.485 $X2=2.55 $Y2=1.68
r128 1 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%A1 3 6 8 11 13
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.16
+ $X2=1.195 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.16
+ $X2=1.195 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.16 $X2=1.195 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.255 $Y=1.985
+ $X2=1.255 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.255 $Y=0.56
+ $X2=1.255 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%A2 3 6 8 9 10 15 16 17
c36 16 0 5.26758e-20 $X=1.705 $Y=1.16
r37 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.16
+ $X2=1.705 $Y2=1.325
r38 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.16
+ $X2=1.705 $Y2=0.995
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.705
+ $Y=1.16 $X2=1.705 $Y2=1.16
r40 9 10 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.655 $Y=1.53
+ $X2=1.655 $Y2=1.87
r41 9 29 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.655 $Y=1.53
+ $X2=1.655 $Y2=1.325
r42 8 29 5.09704 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.62 $Y=1.19
+ $X2=1.62 $Y2=1.325
r43 8 16 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=1.62 $Y=1.19 $X2=1.62
+ $Y2=1.16
r44 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.985
+ $X2=1.765 $Y2=1.325
r45 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.765 $Y=0.56
+ $X2=1.765 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%A3 3 6 8 9 10 15 16 17
r35 15 18 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=1.325
r36 15 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=0.995
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.185
+ $Y=1.16 $X2=2.185 $Y2=1.16
r38 9 10 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.097 $Y=1.53
+ $X2=2.097 $Y2=1.87
r39 9 29 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=2.097 $Y=1.53
+ $X2=2.097 $Y2=1.325
r40 8 29 5.81314 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.125 $Y=1.19
+ $X2=2.125 $Y2=1.325
r41 8 16 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=2.125 $Y=1.19 $X2=2.125
+ $Y2=1.16
r42 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.335 $Y=1.985
+ $X2=2.335 $Y2=1.325
r43 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.335 $Y=0.56
+ $X2=2.335 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%B1 3 7 8 11 12 13
r35 11 14 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.772 $Y=1.16
+ $X2=2.772 $Y2=1.325
r36 11 13 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.772 $Y=1.16
+ $X2=2.772 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.16 $X2=2.755 $Y2=1.16
r38 8 12 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.525 $Y=1.16
+ $X2=2.755 $Y2=1.16
r39 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.85 $Y=0.56 $X2=2.85
+ $Y2=0.995
r40 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.76 $Y=1.985
+ $X2=2.76 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%C1 1 3 6 8 13
r26 10 13 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.435 $Y2=1.16
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.435
+ $Y=1.16 $X2=3.435 $Y2=1.16
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r29 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.325 $X2=3.21
+ $Y2=1.985
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995 $X2=3.21
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%X 1 2 7 8 9 10 11 12 43
r14 27 43 1.81098 $w=3.48e-07 $l=5.5e-08 $layer=LI1_cond $X=0.26 $Y=1.245
+ $X2=0.26 $Y2=1.19
r15 12 38 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.21 $X2=0.26
+ $Y2=2.34
r16 11 12 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.87
+ $X2=0.26 $Y2=2.21
r17 11 32 6.91466 $w=3.48e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=1.87
+ $X2=0.26 $Y2=1.66
r18 10 32 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=1.53 $X2=0.26
+ $Y2=1.66
r19 9 43 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.175
+ $X2=0.26 $Y2=1.19
r20 9 41 4.08923 $w=3.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.26 $Y=1.175
+ $X2=0.26 $Y2=1.07
r21 9 10 8.89028 $w=3.48e-07 $l=2.7e-07 $layer=LI1_cond $X=0.26 $Y=1.26 $X2=0.26
+ $Y2=1.53
r22 9 27 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.26
+ $X2=0.26 $Y2=1.245
r23 8 41 9.39028 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.22 $Y=0.85 $X2=0.22
+ $Y2=1.07
r24 7 8 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=0.51 $X2=0.22
+ $Y2=0.85
r25 2 38 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.34
r26 2 32 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.66
r27 1 7 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%VPWR 1 2 9 13 15 17 22 32 33 36 39 44
c53 1 0 1.27295e-19 $X=0.555 $Y=1.485
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 37 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 30 39 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.017 $Y2=2.72
r60 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r63 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r66 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 23 36 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=1.01 $Y=2.72
+ $X2=0.807 $Y2=2.72
r68 23 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.01 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 22 39 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.9 $Y=2.72
+ $X2=3.017 $Y2=2.72
r70 22 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.9 $Y=2.72 $X2=2.53
+ $Y2=2.72
r71 19 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 17 36 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.807 $Y2=2.72
r73 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 15 44 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r75 11 39 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.017 $Y=2.635
+ $X2=3.017 $Y2=2.72
r76 11 13 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=3.017 $Y=2.635
+ $X2=3.017 $Y2=2
r77 7 36 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.807 $Y=2.635
+ $X2=0.807 $Y2=2.72
r78 7 9 17.5001 $w=4.03e-07 $l=6.15e-07 $layer=LI1_cond $X=0.807 $Y=2.635
+ $X2=0.807 $Y2=2.02
r79 2 13 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.835
+ $Y=1.485 $X2=2.985 $Y2=2
r80 1 9 300 $w=1.7e-07 $l=6.56258e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.825 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%VGND 1 2 9 13 15 17 22 32 33 36 39 44
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r49 37 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r50 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r52 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r53 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r54 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r55 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r56 27 39 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.027
+ $Y2=0
r57 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.53
+ $Y2=0
r58 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r59 26 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r60 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r61 23 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=0.86
+ $Y2=0
r62 23 25 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.61
+ $Y2=0
r63 22 39 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=2.027
+ $Y2=0
r64 22 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.61
+ $Y2=0
r65 19 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 17 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.86
+ $Y2=0
r67 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r68 15 44 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r69 11 39 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.027 $Y=0.085
+ $X2=2.027 $Y2=0
r70 11 13 8.45125 $w=3.73e-07 $l=2.75e-07 $layer=LI1_cond $X=2.027 $Y=0.085
+ $X2=2.027 $Y2=0.36
r71 7 36 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=0.085 $X2=0.86
+ $Y2=0
r72 7 9 4.90928 $w=6.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0.36
r73 2 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=2.05 $Y2=0.36
r74 1 9 45.5 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_NDIFF $count=4 $X=0.555
+ $Y=0.235 $X2=1.03 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_1%A_266_47# 1 2 9 11 12 13 15
r21 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.655
+ $X2=2.595 $Y2=0.74
r22 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.595 $Y=0.655
+ $X2=2.595 $Y2=0.4
r23 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=0.74
+ $X2=2.595 $Y2=0.74
r24 11 12 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.43 $Y=0.74
+ $X2=1.66 $Y2=0.74
r25 7 12 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.512 $Y=0.655
+ $X2=1.66 $Y2=0.74
r26 7 9 3.71126 $w=2.93e-07 $l=9.5e-08 $layer=LI1_cond $X=1.512 $Y=0.655
+ $X2=1.512 $Y2=0.56
r27 2 18 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.235 $X2=2.595 $Y2=0.74
r28 2 15 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.235 $X2=2.595 $Y2=0.4
r29 1 9 182 $w=1.7e-07 $l=4.05123e-07 $layer=licon1_NDIFF $count=1 $X=1.33
+ $Y=0.235 $X2=1.51 $Y2=0.56
.ends


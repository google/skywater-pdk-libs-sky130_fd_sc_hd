* File: sky130_fd_sc_hd__nor4b_1.pex.spice
* Created: Tue Sep  1 19:19:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4B_1%A_91_199# 1 2 9 12 16 17 19 20 24 26 29
c63 19 0 1.48372e-19 $X=2.965 $Y=1.9
r64 26 27 14.3668 $w=2.59e-07 $l=3.05e-07 $layer=LI1_cond $X=2.745 $Y=0.655
+ $X2=3.05 $Y2=0.655
r65 23 27 3.20129 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.05 $Y=0.825
+ $X2=3.05 $Y2=0.655
r66 23 24 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=3.05 $Y=0.825
+ $X2=3.05 $Y2=1.795
r67 20 22 105.628 $w=2.08e-07 $l=2e-06 $layer=LI1_cond $X=0.745 $Y=1.9 $X2=2.745
+ $Y2=1.9
r68 19 24 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.965 $Y=1.9
+ $X2=3.05 $Y2=1.795
r69 19 22 11.619 $w=2.08e-07 $l=2.2e-07 $layer=LI1_cond $X=2.965 $Y=1.9
+ $X2=2.745 $Y2=1.9
r70 17 30 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.16
+ $X2=0.63 $Y2=1.325
r71 17 29 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.16
+ $X2=0.63 $Y2=0.995
r72 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r73 14 20 6.82129 $w=2.1e-07 $l=1.53786e-07 $layer=LI1_cond $X=0.635 $Y=1.795
+ $X2=0.745 $Y2=1.9
r74 14 16 33.2637 $w=2.18e-07 $l=6.35e-07 $layer=LI1_cond $X=0.635 $Y=1.795
+ $X2=0.635 $Y2=1.16
r75 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=1.325
r76 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.73 $Y=0.56 $X2=0.73
+ $Y2=0.995
r77 2 22 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.68 $X2=2.745 $Y2=1.9
r78 1 26 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=2.61
+ $Y=0.465 $X2=2.745 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%C 1 3 6 8 11
c36 11 0 1.48372e-19 $X=1.15 $Y=1.16
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.16 $X2=1.15 $Y2=1.16
r38 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.325
+ $X2=1.15 $Y2=1.16
r39 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.15 $Y=1.325 $X2=1.15
+ $Y2=1.985
r40 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=0.995
+ $X2=1.15 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.15 $Y=0.995 $X2=1.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%B 1 3 6 8 11
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.16 $X2=1.63 $Y2=1.16
r37 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.325
+ $X2=1.63 $Y2=1.16
r38 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.63 $Y=1.325 $X2=1.63
+ $Y2=1.985
r39 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=0.995
+ $X2=1.63 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.63 $Y=0.995 $X2=1.63
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%A 3 6 8 11 13
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.16
+ $X2=2.11 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.16
+ $X2=2.11 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.16 $X2=2.11 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.05 $Y=1.985
+ $X2=2.05 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.05 $Y=0.56 $X2=2.05
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%D_N 3 6 8 11 13
r30 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.59 $Y2=1.325
r31 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.59 $Y2=0.995
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.16 $X2=2.59 $Y2=1.16
r33 6 14 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.535 $Y=1.89
+ $X2=2.535 $Y2=1.325
r34 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.535 $Y=0.675
+ $X2=2.535 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%Y 1 2 3 10 11 14 16 20 23 24
c42 10 0 1.57721e-19 $X=0.855 $Y=0.74
r43 22 24 46.3193 $w=2.58e-07 $l=1.045e-06 $layer=LI1_cond $X=0.215 $Y=0.825
+ $X2=0.215 $Y2=1.87
r44 18 20 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=1.825 $Y=0.655
+ $X2=1.825 $Y2=0.495
r45 17 23 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.055 $Y=0.74 $X2=0.955
+ $Y2=0.74
r46 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.725 $Y=0.74
+ $X2=1.825 $Y2=0.655
r47 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.725 $Y=0.74
+ $X2=1.055 $Y2=0.74
r48 12 23 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=0.655
+ $X2=0.955 $Y2=0.74
r49 12 14 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=0.955 $Y=0.655
+ $X2=0.955 $Y2=0.495
r50 11 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.215 $Y2=0.825
r51 10 23 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.855 $Y=0.74 $X2=0.955
+ $Y2=0.74
r52 10 11 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.855 $Y=0.74
+ $X2=0.345 $Y2=0.74
r53 3 24 300 $w=1.7e-07 $l=5.18748e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.945
r54 2 20 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.235 $X2=1.84 $Y2=0.495
r55 1 14 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=0.805
+ $Y=0.235 $X2=0.94 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%VPWR 1 6 9 10 11 21 22
r33 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r34 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r35 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 14 18 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 11 19 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 11 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r39 9 18 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.095 $Y=2.72
+ $X2=2.07 $Y2=2.72
r40 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=2.72
+ $X2=2.26 $Y2=2.72
r41 8 21 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.425 $Y=2.72
+ $X2=2.99 $Y2=2.72
r42 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.72
+ $X2=2.26 $Y2=2.72
r43 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=2.635 $X2=2.26
+ $Y2=2.72
r44 4 6 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.26 $Y=2.635
+ $X2=2.26 $Y2=2.27
r45 1 6 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.485 $X2=2.26 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_1%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 44
+ 45
c50 23 0 1.57721e-19 $X=0.355 $Y=0
r51 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r53 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r54 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r55 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r56 31 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r57 31 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 29 41 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.07
+ $Y2=0
r59 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.26
+ $Y2=0
r60 28 44 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.99
+ $Y2=0
r61 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.26
+ $Y2=0
r62 26 38 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.15
+ $Y2=0
r63 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.39
+ $Y2=0
r64 25 41 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=2.07
+ $Y2=0
r65 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.39
+ $Y2=0
r66 23 34 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.23
+ $Y2=0
r67 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.52
+ $Y2=0
r68 22 38 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.685 $Y=0 $X2=1.15
+ $Y2=0
r69 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=0 $X2=0.52
+ $Y2=0
r70 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0
r71 18 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0.39
r72 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=0.085
+ $X2=1.39 $Y2=0
r73 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.39 $Y=0.085
+ $X2=1.39 $Y2=0.39
r74 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0
r75 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0.36
r76 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.125
+ $Y=0.235 $X2=2.26 $Y2=0.39
r77 2 16 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.235 $X2=1.39 $Y2=0.39
r78 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.375
+ $Y=0.235 $X2=0.52 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__a211o_2.pxi.spice
* Created: Tue Sep  1 18:50:52 2020
* 
x_PM_SKY130_FD_SC_HD__A211O_2%A_79_21# N_A_79_21#_M1008_d N_A_79_21#_M1006_d
+ N_A_79_21#_M1000_d N_A_79_21#_c_57_n N_A_79_21#_M1010_g N_A_79_21#_M1002_g
+ N_A_79_21#_M1005_g N_A_79_21#_c_58_n N_A_79_21#_M1011_g N_A_79_21#_c_59_n
+ N_A_79_21#_c_72_p N_A_79_21#_c_136_p N_A_79_21#_c_66_n N_A_79_21#_c_67_n
+ N_A_79_21#_c_73_p N_A_79_21#_c_60_n N_A_79_21#_c_61_n N_A_79_21#_c_68_n
+ N_A_79_21#_c_86_p N_A_79_21#_c_62_n PM_SKY130_FD_SC_HD__A211O_2%A_79_21#
x_PM_SKY130_FD_SC_HD__A211O_2%A2 N_A2_c_162_n N_A2_M1001_g N_A2_M1007_g A2
+ N_A2_c_164_n PM_SKY130_FD_SC_HD__A211O_2%A2
x_PM_SKY130_FD_SC_HD__A211O_2%A1 N_A1_M1008_g N_A1_M1003_g A1 N_A1_c_193_n
+ N_A1_c_194_n N_A1_c_195_n PM_SKY130_FD_SC_HD__A211O_2%A1
x_PM_SKY130_FD_SC_HD__A211O_2%B1 N_B1_M1004_g N_B1_M1009_g B1 N_B1_c_227_n
+ N_B1_c_228_n PM_SKY130_FD_SC_HD__A211O_2%B1
x_PM_SKY130_FD_SC_HD__A211O_2%C1 N_C1_c_256_n N_C1_M1006_g N_C1_M1000_g C1
+ N_C1_c_258_n PM_SKY130_FD_SC_HD__A211O_2%C1
x_PM_SKY130_FD_SC_HD__A211O_2%VPWR N_VPWR_M1002_d N_VPWR_M1005_d N_VPWR_M1007_d
+ N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n VPWR
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_280_n N_VPWR_c_289_n
+ N_VPWR_c_290_n PM_SKY130_FD_SC_HD__A211O_2%VPWR
x_PM_SKY130_FD_SC_HD__A211O_2%X N_X_M1010_d N_X_M1002_s N_X_c_345_p N_X_c_346_p
+ X N_X_c_332_n PM_SKY130_FD_SC_HD__A211O_2%X
x_PM_SKY130_FD_SC_HD__A211O_2%A_299_297# N_A_299_297#_M1007_s
+ N_A_299_297#_M1003_d N_A_299_297#_c_351_n N_A_299_297#_c_348_n
+ N_A_299_297#_c_353_n PM_SKY130_FD_SC_HD__A211O_2%A_299_297#
x_PM_SKY130_FD_SC_HD__A211O_2%VGND N_VGND_M1010_s N_VGND_M1011_s N_VGND_M1004_d
+ N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n VGND N_VGND_c_378_n
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n
+ PM_SKY130_FD_SC_HD__A211O_2%VGND
cc_1 VNB N_A_79_21#_c_57_n 0.0216709f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_2 VNB N_A_79_21#_c_58_n 0.0182902f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_3 VNB N_A_79_21#_c_59_n 0.00419078f $X=-0.19 $Y=-0.24 $X2=1.085 $Y2=1.16
cc_4 VNB N_A_79_21#_c_60_n 0.00784647f $X=-0.19 $Y=-0.24 $X2=3.255 $Y2=0.785
cc_5 VNB N_A_79_21#_c_61_n 0.0165135f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.4
cc_6 VNB N_A_79_21#_c_62_n 0.0580499f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_7 VNB N_A2_c_162_n 0.0186394f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=0.235
cc_8 VNB A2 0.00202517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A2_c_164_n 0.0298244f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_10 VNB N_A1_c_193_n 0.0212772f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_11 VNB N_A1_c_194_n 0.00612773f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_12 VNB N_A1_c_195_n 0.0183415f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_13 VNB B1 0.00624789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B1_c_227_n 0.0193163f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB N_B1_c_228_n 0.0177911f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_16 VNB N_C1_c_256_n 0.0227688f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=0.235
cc_17 VNB C1 0.00942206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_C1_c_258_n 0.0372638f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_19 VNB N_VPWR_c_280_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_332_n 0.00171134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_375_n 0.0107461f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_22 VNB N_VGND_c_376_n 0.035393f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_23 VNB N_VGND_c_377_n 0.00526585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_378_n 0.0257853f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.49
cc_25 VNB N_VGND_c_379_n 0.0174308f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.575
cc_26 VNB N_VGND_c_380_n 0.199451f $X=-0.19 $Y=-0.24 $X2=2.44 $Y2=0.695
cc_27 VNB N_VGND_c_381_n 0.0146003f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.4
cc_28 VNB N_VGND_c_382_n 0.0162868f $X=-0.19 $Y=-0.24 $X2=2.44 $Y2=0.785
cc_29 VNB N_VGND_c_383_n 0.00526062f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_30 VPB N_A_79_21#_M1002_g 0.025936f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_31 VPB N_A_79_21#_M1005_g 0.0218202f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_32 VPB N_A_79_21#_c_59_n 0.00336285f $X=-0.19 $Y=1.305 $X2=1.085 $Y2=1.16
cc_33 VPB N_A_79_21#_c_66_n 0.0164753f $X=-0.19 $Y=1.305 $X2=3.255 $Y2=1.575
cc_34 VPB N_A_79_21#_c_67_n 0.00299909f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.575
cc_35 VPB N_A_79_21#_c_68_n 0.0260659f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=1.755
cc_36 VPB N_A_79_21#_c_62_n 0.0138444f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_37 VPB N_A2_M1007_g 0.0243941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A2_c_164_n 0.00780582f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_39 VPB N_A1_M1003_g 0.0210736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A1_c_193_n 0.00510692f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_41 VPB N_B1_M1009_g 0.0191018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B1_c_227_n 0.00437045f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_43 VPB N_C1_M1000_g 0.0255936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_C1_c_258_n 0.00930724f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_45 VPB N_VPWR_c_281_n 0.0107202f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1
cc_46 VPB N_VPWR_c_282_n 0.0436299f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_47 VPB N_VPWR_c_283_n 0.010744f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_48 VPB N_VPWR_c_284_n 0.00527793f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_49 VPB N_VPWR_c_285_n 0.0178439f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_50 VPB N_VPWR_c_286_n 0.0183278f $X=-0.19 $Y=1.305 $X2=3.255 $Y2=1.575
cc_51 VPB N_VPWR_c_287_n 0.0418017f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=0.4
cc_52 VPB N_VPWR_c_280_n 0.0521446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_289_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_54 VPB N_VPWR_c_290_n 0.00525752f $X=-0.19 $Y=1.305 $X2=1.085 $Y2=1.16
cc_55 VPB N_X_c_332_n 0.00248033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_299_297#_c_348_n 0.00631724f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_57 N_A_79_21#_c_58_n N_A2_c_162_n 0.00848426f $X=0.9 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_58 N_A_79_21#_c_59_n N_A2_c_162_n 0.00274362f $X=1.085 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_59 N_A_79_21#_c_72_p N_A2_c_162_n 0.0132514f $X=2.275 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_60 N_A_79_21#_c_73_p N_A2_c_162_n 0.00131571f $X=2.44 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_61 N_A_79_21#_c_59_n N_A2_M1007_g 0.00451736f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_66_n N_A2_M1007_g 0.0142782f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_59_n A2 0.0189785f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_72_p A2 0.0193792f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_66_n A2 0.0180506f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_62_n A2 6.46526e-19 $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_59_n N_A2_c_164_n 0.00311755f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_72_p N_A2_c_164_n 0.0066792f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_66_n N_A2_c_164_n 0.00609418f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_62_n N_A2_c_164_n 0.0142329f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_66_n N_A1_M1003_g 0.0115751f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_66_n N_A1_c_193_n 0.00376493f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_86_p N_A1_c_193_n 0.0039881f $X=2.44 $Y=0.785 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_72_p N_A1_c_194_n 0.0195177f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_66_n N_A1_c_194_n 0.0266212f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_86_p N_A1_c_194_n 0.0113517f $X=2.44 $Y=0.785 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_72_p N_A1_c_195_n 0.00959468f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_73_p N_A1_c_195_n 0.00816096f $X=2.44 $Y=0.36 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_86_p N_A1_c_195_n 6.8073e-19 $X=2.44 $Y=0.785 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_66_n N_B1_M1009_g 0.0144697f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_68_n N_B1_M1009_g 0.00224314f $X=3.42 $Y=1.755 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_66_n B1 0.023855f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_60_n B1 0.0294284f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_66_n N_B1_c_227_n 0.00308881f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_60_n N_B1_c_227_n 0.00321658f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_60_n N_B1_c_228_n 0.0131325f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_61_n N_B1_c_228_n 5.27165e-19 $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_60_n N_C1_c_256_n 0.0114696f $X=3.255 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_79_21#_c_61_n N_C1_c_256_n 0.00626231f $X=3.42 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_79_21#_c_66_n N_C1_M1000_g 0.0143092f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_68_n N_C1_M1000_g 0.0121743f $X=3.42 $Y=1.755 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_66_n C1 0.0197603f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_60_n C1 0.023444f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_66_n N_C1_c_258_n 0.00679036f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_60_n N_C1_c_258_n 0.00694884f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_67_n N_VPWR_M1005_d 0.00398804f $X=1.31 $Y=1.575 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_66_n N_VPWR_M1007_d 0.00644456f $X=3.255 $Y=1.575 $X2=0 $Y2=0
cc_98 N_A_79_21#_M1002_g N_VPWR_c_282_n 0.0034372f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_79_21#_M1005_g N_VPWR_c_283_n 0.00324789f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_67_n N_VPWR_c_283_n 0.0210201f $X=1.31 $Y=1.575 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_62_n N_VPWR_c_283_n 8.18903e-19 $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_79_21#_M1002_g N_VPWR_c_285_n 0.00585385f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_M1005_g N_VPWR_c_285_n 0.00585385f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_79_21#_c_68_n N_VPWR_c_287_n 0.0110564f $X=3.42 $Y=1.755 $X2=0 $Y2=0
cc_105 N_A_79_21#_M1000_d N_VPWR_c_280_n 0.00228331f $X=3.285 $Y=1.485 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_M1002_g N_VPWR_c_280_n 0.0114668f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_79_21#_M1005_g N_VPWR_c_280_n 0.0119014f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_68_n N_VPWR_c_280_n 0.0115304f $X=3.42 $Y=1.755 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_57_n N_X_c_332_n 0.0026937f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_110 N_A_79_21#_M1002_g N_X_c_332_n 0.00479385f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_79_21#_M1005_g N_X_c_332_n 0.00183748f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_58_n N_X_c_332_n 9.34096e-19 $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_59_n N_X_c_332_n 0.0382115f $X=1.085 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_62_n N_X_c_332_n 0.0297275f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_66_n N_A_299_297#_M1007_s 0.00485213f $X=3.255 $Y=1.575
+ $X2=-0.19 $Y2=-0.24
cc_116 N_A_79_21#_c_66_n N_A_299_297#_M1003_d 0.00558159f $X=3.255 $Y=1.575
+ $X2=0 $Y2=0
cc_117 N_A_79_21#_c_66_n N_A_299_297#_c_351_n 0.0367882f $X=3.255 $Y=1.575 $X2=0
+ $Y2=0
cc_118 N_A_79_21#_c_66_n N_A_299_297#_c_348_n 0.0210659f $X=3.255 $Y=1.575 $X2=0
+ $Y2=0
cc_119 N_A_79_21#_c_66_n N_A_299_297#_c_353_n 0.0181279f $X=3.255 $Y=1.575 $X2=0
+ $Y2=0
cc_120 N_A_79_21#_c_68_n N_A_299_297#_c_353_n 0.0165753f $X=3.42 $Y=1.755 $X2=0
+ $Y2=0
cc_121 N_A_79_21#_c_66_n A_585_297# 0.00485323f $X=3.255 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_79_21#_c_72_p N_VGND_M1011_s 0.00711714f $X=2.275 $Y=0.785 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_c_136_p N_VGND_M1011_s 0.0053859f $X=1.31 $Y=0.785 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_60_n N_VGND_M1004_d 0.00445525f $X=3.255 $Y=0.785 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_c_57_n N_VGND_c_376_n 0.00382875f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_60_n N_VGND_c_377_n 0.0168356f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_72_p N_VGND_c_378_n 0.00684738f $X=2.275 $Y=0.785 $X2=0
+ $Y2=0
cc_128 N_A_79_21#_c_73_p N_VGND_c_378_n 0.018286f $X=2.44 $Y=0.36 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_60_n N_VGND_c_378_n 0.00260343f $X=3.255 $Y=0.785 $X2=0
+ $Y2=0
cc_130 N_A_79_21#_c_60_n N_VGND_c_379_n 0.00212534f $X=3.255 $Y=0.785 $X2=0
+ $Y2=0
cc_131 N_A_79_21#_c_61_n N_VGND_c_379_n 0.0185069f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_132 N_A_79_21#_M1008_d N_VGND_c_380_n 0.00307026f $X=2.3 $Y=0.235 $X2=0 $Y2=0
cc_133 N_A_79_21#_M1006_d N_VGND_c_380_n 0.00210124f $X=3.285 $Y=0.235 $X2=0
+ $Y2=0
cc_134 N_A_79_21#_c_57_n N_VGND_c_380_n 0.0114173f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_58_n N_VGND_c_380_n 0.00786964f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_72_p N_VGND_c_380_n 0.0146077f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_136_p N_VGND_c_380_n 0.00172085f $X=1.31 $Y=0.785 $X2=0
+ $Y2=0
cc_138 N_A_79_21#_c_73_p N_VGND_c_380_n 0.0122842f $X=2.44 $Y=0.36 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_60_n N_VGND_c_380_n 0.0098176f $X=3.255 $Y=0.785 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_61_n N_VGND_c_380_n 0.0122611f $X=3.42 $Y=0.4 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_57_n N_VGND_c_381_n 0.00585385f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_58_n N_VGND_c_381_n 0.0046653f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_57_n N_VGND_c_382_n 5.35408e-19 $X=0.47 $Y=1 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_58_n N_VGND_c_382_n 0.00866968f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_72_p N_VGND_c_382_n 0.0197185f $X=2.275 $Y=0.785 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_136_p N_VGND_c_382_n 0.0166986f $X=1.31 $Y=0.785 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_62_n N_VGND_c_382_n 8.39972e-19 $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_72_p A_348_47# 0.00998777f $X=2.275 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A2_M1007_g N_A1_M1003_g 0.0349894f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_150 A2 N_A1_c_194_n 0.0187427f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A2_c_164_n N_A1_c_194_n 0.0017831f $X=1.665 $Y=1.157 $X2=0 $Y2=0
cc_152 N_A2_c_162_n N_A1_c_195_n 0.0257368f $X=1.665 $Y=0.99 $X2=0 $Y2=0
cc_153 N_A2_c_164_n N_A1_c_195_n 0.0185886f $X=1.665 $Y=1.157 $X2=0 $Y2=0
cc_154 N_A2_M1007_g N_VPWR_c_283_n 0.00226303f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A2_M1007_g N_VPWR_c_284_n 0.00466029f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A2_M1007_g N_VPWR_c_286_n 0.00420583f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A2_M1007_g N_VPWR_c_280_n 0.00734207f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A2_M1007_g N_A_299_297#_c_351_n 0.00929228f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A2_M1007_g N_A_299_297#_c_348_n 0.00749315f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A2_c_162_n N_VGND_c_382_n 0.01516f $X=1.665 $Y=0.99 $X2=0 $Y2=0
cc_161 N_A1_M1003_g N_B1_M1009_g 0.0251746f $X=2.37 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A1_c_193_n B1 7.81088e-19 $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A1_c_194_n B1 0.0201357f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A1_c_193_n N_B1_c_227_n 0.0221726f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A1_c_194_n N_B1_c_227_n 7.32725e-19 $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_c_195_n N_B1_c_228_n 0.0186358f $X=2.297 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_M1003_g N_VPWR_c_284_n 0.00440799f $X=2.37 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A1_M1003_g N_VPWR_c_287_n 0.00434414f $X=2.37 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A1_M1003_g N_VPWR_c_280_n 0.00632473f $X=2.37 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A1_M1003_g N_A_299_297#_c_351_n 0.01096f $X=2.37 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A1_M1003_g N_A_299_297#_c_348_n 7.78734e-19 $X=2.37 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A1_c_195_n N_VGND_c_378_n 0.00423225f $X=2.297 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_195_n N_VGND_c_380_n 0.0064178f $X=2.297 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_195_n N_VGND_c_382_n 0.00254946f $X=2.297 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B1_c_228_n N_C1_c_256_n 0.0219618f $X=2.79 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_176 N_B1_M1009_g N_C1_M1000_g 0.05058f $X=2.85 $Y=1.985 $X2=0 $Y2=0
cc_177 B1 C1 0.017109f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_178 B1 N_C1_c_258_n 0.00178733f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_179 N_B1_c_227_n N_C1_c_258_n 0.05058f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_M1009_g N_VPWR_c_287_n 0.0055654f $X=2.85 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B1_M1009_g N_VPWR_c_280_n 0.0101033f $X=2.85 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B1_M1009_g N_A_299_297#_c_353_n 0.0103386f $X=2.85 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_c_228_n N_VGND_c_377_n 0.0031795f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_c_228_n N_VGND_c_378_n 0.00433717f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B1_c_228_n N_VGND_c_380_n 0.00614259f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_186 N_C1_M1000_g N_VPWR_c_287_n 0.00546688f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_187 N_C1_M1000_g N_VPWR_c_280_n 0.0106182f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_188 N_C1_M1000_g N_A_299_297#_c_353_n 0.00199801f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_C1_c_256_n N_VGND_c_377_n 0.00291251f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_190 N_C1_c_256_n N_VGND_c_379_n 0.00420829f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_191 N_C1_c_256_n N_VGND_c_380_n 0.00678018f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_192 N_VPWR_c_280_n N_X_M1002_s 0.00376664f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_285_n N_X_c_332_n 0.00738837f $X=1 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_c_280_n N_X_c_332_n 0.00816554f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_280_n N_A_299_297#_M1007_s 0.00209319f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_196 N_VPWR_c_280_n N_A_299_297#_M1003_d 0.00271317f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_197 N_VPWR_M1007_d N_A_299_297#_c_351_n 0.00612377f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_284_n N_A_299_297#_c_351_n 0.020839f $X=2.105 $Y=2.355 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_286_n N_A_299_297#_c_351_n 0.00210141f $X=1.955 $Y=2.72 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_287_n N_A_299_297#_c_351_n 0.00287255f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_280_n N_A_299_297#_c_351_n 0.0106128f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_283_n N_A_299_297#_c_348_n 0.0463287f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_203 N_VPWR_c_286_n N_A_299_297#_c_348_n 0.0209208f $X=1.955 $Y=2.72 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_280_n N_A_299_297#_c_348_n 0.0123991f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_287_n N_A_299_297#_c_353_n 0.0196507f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_280_n N_A_299_297#_c_353_n 0.0124448f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_280_n A_585_297# 0.00897657f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_208 N_VPWR_c_282_n N_VGND_c_376_n 0.0102687f $X=0.26 $Y=1.655 $X2=0 $Y2=0
cc_209 N_X_c_332_n N_VGND_c_376_n 0.00152559f $X=0.685 $Y=0.76 $X2=0 $Y2=0
cc_210 N_X_M1010_d N_VGND_c_380_n 0.00399277f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_211 N_X_c_345_p N_VGND_c_380_n 0.00839556f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_212 N_X_c_346_p N_VGND_c_380_n 2.70794e-19 $X=0.67 $Y=0.75 $X2=0 $Y2=0
cc_213 N_X_c_345_p N_VGND_c_381_n 0.0135183f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_214 N_VGND_c_380_n A_348_47# 0.00445732f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o311a_2.pxi.spice
* Created: Tue Sep  1 19:24:26 2020
* 
x_PM_SKY130_FD_SC_HD__O311A_2%A_91_21# N_A_91_21#_M1008_d N_A_91_21#_M1001_d
+ N_A_91_21#_M1003_d N_A_91_21#_c_70_n N_A_91_21#_M1009_g N_A_91_21#_M1002_g
+ N_A_91_21#_c_71_n N_A_91_21#_M1011_g N_A_91_21#_M1007_g N_A_91_21#_c_72_n
+ N_A_91_21#_c_73_n N_A_91_21#_c_85_p N_A_91_21#_c_127_p N_A_91_21#_c_86_p
+ N_A_91_21#_c_95_p N_A_91_21#_c_87_p N_A_91_21#_c_99_p N_A_91_21#_c_96_p
+ N_A_91_21#_c_105_p N_A_91_21#_c_101_p N_A_91_21#_c_74_n N_A_91_21#_c_81_n
+ N_A_91_21#_c_82_n N_A_91_21#_c_75_n PM_SKY130_FD_SC_HD__O311A_2%A_91_21#
x_PM_SKY130_FD_SC_HD__O311A_2%A1 N_A1_M1013_g N_A1_M1000_g A1 N_A1_c_181_n
+ N_A1_c_182_n PM_SKY130_FD_SC_HD__O311A_2%A1
x_PM_SKY130_FD_SC_HD__O311A_2%A2 N_A2_M1012_g N_A2_M1004_g A2 A2 A2 N_A2_c_213_n
+ N_A2_c_214_n N_A2_c_215_n PM_SKY130_FD_SC_HD__O311A_2%A2
x_PM_SKY130_FD_SC_HD__O311A_2%A3 N_A3_M1005_g N_A3_M1001_g A3 A3 A3 N_A3_c_249_n
+ N_A3_c_250_n N_A3_c_251_n PM_SKY130_FD_SC_HD__O311A_2%A3
x_PM_SKY130_FD_SC_HD__O311A_2%B1 N_B1_M1010_g N_B1_M1006_g B1 N_B1_c_284_n
+ N_B1_c_285_n N_B1_c_286_n PM_SKY130_FD_SC_HD__O311A_2%B1
x_PM_SKY130_FD_SC_HD__O311A_2%C1 N_C1_c_319_n N_C1_M1008_g N_C1_M1003_g C1
+ N_C1_c_321_n PM_SKY130_FD_SC_HD__O311A_2%C1
x_PM_SKY130_FD_SC_HD__O311A_2%VPWR N_VPWR_M1002_d N_VPWR_M1007_d N_VPWR_M1010_d
+ N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_350_n
+ VPWR N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_345_n N_VPWR_c_354_n
+ N_VPWR_c_355_n PM_SKY130_FD_SC_HD__O311A_2%VPWR
x_PM_SKY130_FD_SC_HD__O311A_2%X N_X_M1009_s N_X_M1002_s X X X X X X X
+ N_X_c_404_n PM_SKY130_FD_SC_HD__O311A_2%X
x_PM_SKY130_FD_SC_HD__O311A_2%VGND N_VGND_M1009_d N_VGND_M1011_d N_VGND_M1012_d
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n VGND
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ N_VGND_c_440_n PM_SKY130_FD_SC_HD__O311A_2%VGND
x_PM_SKY130_FD_SC_HD__O311A_2%A_360_47# N_A_360_47#_M1013_d N_A_360_47#_M1005_d
+ N_A_360_47#_c_499_n N_A_360_47#_c_487_n N_A_360_47#_c_490_n
+ N_A_360_47#_c_495_n N_A_360_47#_c_506_n PM_SKY130_FD_SC_HD__O311A_2%A_360_47#
cc_1 VNB N_A_91_21#_c_70_n 0.0215059f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_2 VNB N_A_91_21#_c_71_n 0.0184006f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_3 VNB N_A_91_21#_c_72_n 0.00157408f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=1.16
cc_4 VNB N_A_91_21#_c_73_n 0.0535018f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=1.16
cc_5 VNB N_A_91_21#_c_74_n 0.00281491f $X=-0.19 $Y=-0.24 $X2=3.555 $Y2=1.495
cc_6 VNB N_A_91_21#_c_75_n 0.0245152f $X=-0.19 $Y=-0.24 $X2=3.88 $Y2=0.4
cc_7 VNB A1 0.00290387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_181_n 0.020649f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.56
cc_9 VNB N_A1_c_182_n 0.0194735f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.325
cc_10 VNB N_A2_c_213_n 0.0208451f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.985
cc_11 VNB N_A2_c_214_n 0.00397726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_215_n 0.018451f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_13 VNB N_A3_c_249_n 0.0261176f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.985
cc_14 VNB N_A3_c_250_n 0.00452535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A3_c_251_n 0.0185884f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_16 VNB N_B1_c_284_n 0.0226542f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.56
cc_17 VNB N_B1_c_285_n 0.00347516f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.56
cc_18 VNB N_B1_c_286_n 0.0167081f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.325
cc_19 VNB N_C1_c_319_n 0.0209378f $X=-0.19 $Y=-0.24 $X2=3.745 $Y2=0.235
cc_20 VNB C1 0.0133884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_C1_c_321_n 0.0344721f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.325
cc_22 VNB N_VPWR_c_345_n 0.17485f $X=-0.19 $Y=-0.24 $X2=3.47 $Y2=1.58
cc_23 VNB X 0.00103928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_404_n 0.017348f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.985
cc_25 VNB N_VGND_c_431_n 0.0105833f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_26 VNB N_VGND_c_432_n 0.0325136f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.56
cc_27 VNB N_VGND_c_433_n 0.00180074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_434_n 0.00529728f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.325
cc_29 VNB N_VGND_c_435_n 0.0157573f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=1.495
cc_30 VNB N_VGND_c_436_n 0.0159285f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=1.58
cc_31 VNB N_VGND_c_437_n 0.0394108f $X=-0.19 $Y=-0.24 $X2=3.47 $Y2=1.58
cc_32 VNB N_VGND_c_438_n 0.217852f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=1.58
cc_33 VNB N_VGND_c_439_n 0.0104906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_440_n 0.00718038f $X=-0.19 $Y=-0.24 $X2=3.762 $Y2=0.4
cc_35 VPB N_A_91_21#_M1002_g 0.0252993f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.985
cc_36 VPB N_A_91_21#_M1007_g 0.0209812f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.985
cc_37 VPB N_A_91_21#_c_72_n 0.00280012f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.16
cc_38 VPB N_A_91_21#_c_73_n 0.0141761f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.16
cc_39 VPB N_A_91_21#_c_74_n 0.00165139f $X=-0.19 $Y=1.305 $X2=3.555 $Y2=1.495
cc_40 VPB N_A_91_21#_c_81_n 0.00763029f $X=-0.19 $Y=1.305 $X2=3.91 $Y2=1.665
cc_41 VPB N_A_91_21#_c_82_n 0.0312708f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=1.815
cc_42 VPB N_A1_M1000_g 0.0229699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB A1 0.0011816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A1_c_181_n 0.00403444f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.56
cc_45 VPB N_A2_M1004_g 0.0205099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB A2 0.00162648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A2_c_213_n 0.00452834f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.985
cc_48 VPB N_A2_c_214_n 0.00231345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A3_M1001_g 0.0206248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB A3 0.00247089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A3_c_249_n 0.00728583f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.985
cc_52 VPB N_A3_c_250_n 0.0018022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_B1_M1010_g 0.0195048f $X=-0.19 $Y=1.305 $X2=3.745 $Y2=1.485
cc_54 VPB N_B1_c_284_n 0.00509613f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.56
cc_55 VPB N_B1_c_285_n 0.00178038f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.56
cc_56 VPB N_C1_M1003_g 0.0257003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB C1 0.00297249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_C1_c_321_n 0.0096974f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.325
cc_59 VPB N_VPWR_c_346_n 0.0105574f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_60 VPB N_VPWR_c_347_n 0.0466076f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.56
cc_61 VPB N_VPWR_c_348_n 0.0185011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_349_n 0.00595031f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.325
cc_63 VPB N_VPWR_c_350_n 0.00509471f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.495
cc_64 VPB N_VPWR_c_351_n 0.0450741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_352_n 0.0167769f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.68
cc_66 VPB N_VPWR_c_345_n 0.0430844f $X=-0.19 $Y=1.305 $X2=3.47 $Y2=1.58
cc_67 VPB N_VPWR_c_354_n 0.00756851f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=1.815
cc_68 VPB N_VPWR_c_355_n 0.00449427f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=2.36
cc_69 VPB N_X_c_404_n 0.00588682f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.985
cc_70 N_A_91_21#_M1007_g N_A1_M1000_g 0.0156636f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_91_21#_c_72_n N_A1_M1000_g 0.00301901f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_91_21#_c_85_p N_A1_M1000_g 0.0105021f $X=1.64 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A_91_21#_c_86_p N_A1_M1000_g 0.0174768f $X=1.725 $Y=2.295 $X2=0 $Y2=0
cc_74 N_A_91_21#_c_87_p N_A1_M1000_g 0.00759606f $X=1.81 $Y=2.38 $X2=0 $Y2=0
cc_75 N_A_91_21#_c_72_n A1 0.024918f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_91_21#_c_73_n A1 0.00240951f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_91_21#_c_85_p A1 0.0237392f $X=1.64 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_91_21#_c_72_n N_A1_c_181_n 3.10952e-19 $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_91_21#_c_73_n N_A1_c_181_n 0.0187852f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_91_21#_c_85_p N_A1_c_181_n 0.00236315f $X=1.64 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_91_21#_c_71_n N_A1_c_182_n 0.00425898f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_91_21#_c_95_p N_A2_M1004_g 0.0124823f $X=2.845 $Y=2.38 $X2=0 $Y2=0
cc_83 N_A_91_21#_c_96_p N_A2_M1004_g 0.00110498f $X=3.01 $Y=1.68 $X2=0 $Y2=0
cc_84 N_A_91_21#_c_95_p A2 0.0121614f $X=2.845 $Y=2.38 $X2=0 $Y2=0
cc_85 N_A_91_21#_c_95_p N_A3_M1001_g 0.011169f $X=2.845 $Y=2.38 $X2=0 $Y2=0
cc_86 N_A_91_21#_c_99_p N_A3_M1001_g 5.89792e-19 $X=3.01 $Y=2.295 $X2=0 $Y2=0
cc_87 N_A_91_21#_c_96_p N_A3_M1001_g 0.00872665f $X=3.01 $Y=1.68 $X2=0 $Y2=0
cc_88 N_A_91_21#_c_101_p N_A3_M1001_g 0.00249995f $X=3.175 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_91_21#_c_95_p A3 0.0132929f $X=2.845 $Y=2.38 $X2=0 $Y2=0
cc_90 N_A_91_21#_c_99_p N_B1_M1010_g 0.00209677f $X=3.01 $Y=2.295 $X2=0 $Y2=0
cc_91 N_A_91_21#_c_96_p N_B1_M1010_g 0.00815505f $X=3.01 $Y=1.68 $X2=0 $Y2=0
cc_92 N_A_91_21#_c_105_p N_B1_M1010_g 0.0108502f $X=3.47 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A_91_21#_c_101_p N_B1_M1010_g 8.84614e-19 $X=3.175 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_91_21#_c_74_n N_B1_M1010_g 0.00352622f $X=3.555 $Y=1.495 $X2=0 $Y2=0
cc_95 N_A_91_21#_c_105_p N_B1_c_284_n 0.0027472f $X=3.47 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_91_21#_c_101_p N_B1_c_284_n 0.00134053f $X=3.175 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A_91_21#_c_74_n N_B1_c_284_n 0.00573092f $X=3.555 $Y=1.495 $X2=0 $Y2=0
cc_98 N_A_91_21#_c_105_p N_B1_c_285_n 0.00872323f $X=3.47 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A_91_21#_c_101_p N_B1_c_285_n 0.0195547f $X=3.175 $Y=1.58 $X2=0 $Y2=0
cc_100 N_A_91_21#_c_74_n N_B1_c_285_n 0.0251379f $X=3.555 $Y=1.495 $X2=0 $Y2=0
cc_101 N_A_91_21#_c_75_n N_B1_c_286_n 0.00573092f $X=3.88 $Y=0.4 $X2=0 $Y2=0
cc_102 N_A_91_21#_c_74_n N_C1_c_319_n 0.00789512f $X=3.555 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_91_21#_c_75_n N_C1_c_319_n 0.0150777f $X=3.88 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_91_21#_c_96_p N_C1_M1003_g 5.87886e-19 $X=3.01 $Y=1.68 $X2=0 $Y2=0
cc_105 N_A_91_21#_c_74_n N_C1_M1003_g 0.0084555f $X=3.555 $Y=1.495 $X2=0 $Y2=0
cc_106 N_A_91_21#_c_81_n N_C1_M1003_g 0.0166705f $X=3.91 $Y=1.665 $X2=0 $Y2=0
cc_107 N_A_91_21#_c_74_n C1 0.0230137f $X=3.555 $Y=1.495 $X2=0 $Y2=0
cc_108 N_A_91_21#_c_81_n C1 0.0181761f $X=3.91 $Y=1.665 $X2=0 $Y2=0
cc_109 N_A_91_21#_c_75_n C1 0.0200459f $X=3.88 $Y=0.4 $X2=0 $Y2=0
cc_110 N_A_91_21#_c_74_n N_C1_c_321_n 0.00752413f $X=3.555 $Y=1.495 $X2=0 $Y2=0
cc_111 N_A_91_21#_c_81_n N_C1_c_321_n 0.00297804f $X=3.91 $Y=1.665 $X2=0 $Y2=0
cc_112 N_A_91_21#_c_75_n N_C1_c_321_n 0.00315879f $X=3.88 $Y=0.4 $X2=0 $Y2=0
cc_113 N_A_91_21#_c_85_p N_VPWR_M1007_d 0.0140824f $X=1.64 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_91_21#_c_127_p N_VPWR_M1007_d 0.00321774f $X=1.245 $Y=1.58 $X2=0
+ $Y2=0
cc_115 N_A_91_21#_c_105_p N_VPWR_M1010_d 0.00507927f $X=3.47 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_91_21#_c_74_n N_VPWR_M1010_d 3.14485e-19 $X=3.555 $Y=1.495 $X2=0
+ $Y2=0
cc_117 N_A_91_21#_c_81_n N_VPWR_M1010_d 9.10335e-19 $X=3.91 $Y=1.665 $X2=0 $Y2=0
cc_118 N_A_91_21#_M1002_g N_VPWR_c_347_n 0.007691f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_91_21#_M1002_g N_VPWR_c_348_n 0.00503406f $X=0.53 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_91_21#_M1007_g N_VPWR_c_348_n 0.00541359f $X=0.95 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_91_21#_M1007_g N_VPWR_c_349_n 0.008733f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_91_21#_c_73_n N_VPWR_c_349_n 7.36359e-19 $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_91_21#_c_85_p N_VPWR_c_349_n 0.0181878f $X=1.64 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_91_21#_c_127_p N_VPWR_c_349_n 0.0146353f $X=1.245 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A_91_21#_c_99_p N_VPWR_c_350_n 0.0127992f $X=3.01 $Y=2.295 $X2=0 $Y2=0
cc_126 N_A_91_21#_c_96_p N_VPWR_c_350_n 0.032561f $X=3.01 $Y=1.68 $X2=0 $Y2=0
cc_127 N_A_91_21#_c_105_p N_VPWR_c_350_n 0.0143275f $X=3.47 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_91_21#_c_95_p N_VPWR_c_351_n 0.0589382f $X=2.845 $Y=2.38 $X2=0 $Y2=0
cc_129 N_A_91_21#_c_87_p N_VPWR_c_351_n 0.0109366f $X=1.81 $Y=2.38 $X2=0 $Y2=0
cc_130 N_A_91_21#_c_99_p N_VPWR_c_351_n 0.019051f $X=3.01 $Y=2.295 $X2=0 $Y2=0
cc_131 N_A_91_21#_c_82_n N_VPWR_c_352_n 0.0190655f $X=3.88 $Y=1.815 $X2=0 $Y2=0
cc_132 N_A_91_21#_M1001_d N_VPWR_c_345_n 0.00219216f $X=2.87 $Y=1.485 $X2=0
+ $Y2=0
cc_133 N_A_91_21#_M1003_d N_VPWR_c_345_n 0.00283025f $X=3.745 $Y=1.485 $X2=0
+ $Y2=0
cc_134 N_A_91_21#_M1002_g N_VPWR_c_345_n 0.00964666f $X=0.53 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_91_21#_M1007_g N_VPWR_c_345_n 0.0102772f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_91_21#_c_95_p N_VPWR_c_345_n 0.0372911f $X=2.845 $Y=2.38 $X2=0 $Y2=0
cc_137 N_A_91_21#_c_87_p N_VPWR_c_345_n 0.00586103f $X=1.81 $Y=2.38 $X2=0 $Y2=0
cc_138 N_A_91_21#_c_99_p N_VPWR_c_345_n 0.0123125f $X=3.01 $Y=2.295 $X2=0 $Y2=0
cc_139 N_A_91_21#_c_82_n N_VPWR_c_345_n 0.0110914f $X=3.88 $Y=1.815 $X2=0 $Y2=0
cc_140 N_A_91_21#_c_70_n X 0.0164223f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_91_21#_c_71_n X 0.00382189f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_91_21#_c_72_n X 0.0241381f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_91_21#_c_73_n X 0.0239979f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_91_21#_M1002_g X 0.0220594f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_91_21#_M1007_g X 0.0202298f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_91_21#_c_72_n X 0.0130751f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_91_21#_c_73_n X 0.00299403f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_91_21#_c_73_n N_X_c_404_n 0.0164667f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_91_21#_c_95_p A_360_297# 0.00829427f $X=2.845 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_91_21#_c_95_p A_460_297# 0.00930583f $X=2.845 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_91_21#_c_70_n N_VGND_c_432_n 0.00507496f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_91_21#_c_70_n N_VGND_c_433_n 7.95762e-19 $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_91_21#_c_71_n N_VGND_c_433_n 0.0127369f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_91_21#_c_72_n N_VGND_c_433_n 0.0143975f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_91_21#_c_73_n N_VGND_c_433_n 0.00286475f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_91_21#_c_85_p N_VGND_c_433_n 0.00488088f $X=1.64 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_91_21#_c_70_n N_VGND_c_435_n 0.00503406f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_91_21#_c_71_n N_VGND_c_435_n 0.0046653f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_91_21#_c_75_n N_VGND_c_437_n 0.0364195f $X=3.88 $Y=0.4 $X2=0 $Y2=0
cc_160 N_A_91_21#_M1008_d N_VGND_c_438_n 0.00209319f $X=3.745 $Y=0.235 $X2=0
+ $Y2=0
cc_161 N_A_91_21#_c_70_n N_VGND_c_438_n 0.00968554f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_91_21#_c_71_n N_VGND_c_438_n 0.00796766f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_91_21#_c_75_n N_VGND_c_438_n 0.0216215f $X=3.88 $Y=0.4 $X2=0 $Y2=0
cc_164 N_A_91_21#_c_101_p N_A_360_47#_c_487_n 5.79016e-19 $X=3.175 $Y=1.58 $X2=0
+ $Y2=0
cc_165 N_A_91_21#_c_74_n A_677_47# 6.54266e-19 $X=3.555 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_91_21#_c_75_n A_677_47# 0.00644001f $X=3.88 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A1_M1000_g N_A2_M1004_g 0.0429089f $X=1.725 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A1_M1000_g A2 0.0059338f $X=1.725 $Y=1.985 $X2=0 $Y2=0
cc_169 A1 N_A2_c_213_n 3.11177e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A1_c_181_n N_A2_c_213_n 0.0179535f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_171 A1 N_A2_c_214_n 0.0261113f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A1_c_181_n N_A2_c_214_n 0.0021064f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A1_c_182_n N_A2_c_215_n 0.017939f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_VPWR_c_349_n 0.00591858f $X=1.725 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A1_M1000_g N_VPWR_c_351_n 0.00357668f $X=1.725 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A1_M1000_g N_VPWR_c_345_n 0.00618337f $X=1.725 $Y=1.985 $X2=0 $Y2=0
cc_177 A1 N_VGND_c_433_n 0.0183964f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A1_c_181_n N_VGND_c_433_n 0.00262179f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A1_c_182_n N_VGND_c_433_n 0.0110619f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_182_n N_VGND_c_436_n 0.00525069f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_182_n N_VGND_c_438_n 0.00910857f $X=1.665 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_M1004_g N_A3_M1001_g 0.0302643f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A2_M1004_g A3 0.00390408f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_184 A2 A3 0.0374428f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_185 N_A2_c_213_n N_A3_c_249_n 0.0202578f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_c_214_n N_A3_c_249_n 3.33413e-19 $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A2_c_213_n N_A3_c_250_n 0.00390408f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A2_c_214_n N_A3_c_250_n 0.0374428f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_c_215_n N_A3_c_251_n 0.0235995f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_M1004_g N_VPWR_c_351_n 0.00357877f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A2_M1004_g N_VPWR_c_345_n 0.00584902f $X=2.225 $Y=1.985 $X2=0 $Y2=0
cc_192 A2 A_360_297# 0.00636701f $X=1.98 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_193 N_A2_c_215_n N_VGND_c_433_n 8.06326e-19 $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_215_n N_VGND_c_434_n 0.00364336f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_215_n N_VGND_c_436_n 0.00427293f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_215_n N_VGND_c_438_n 0.00626203f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_214_n N_A_360_47#_c_487_n 0.00880508f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A2_c_215_n N_A_360_47#_c_487_n 0.012961f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_213_n N_A_360_47#_c_490_n 6.16454e-19 $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A2_c_214_n N_A_360_47#_c_490_n 0.0160718f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A3_M1001_g N_B1_M1010_g 0.0136218f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A3_c_249_n N_B1_c_284_n 0.0204866f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A3_c_250_n N_B1_c_284_n 2.38775e-19 $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A3_c_249_n N_B1_c_285_n 0.0025442f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A3_c_250_n N_B1_c_285_n 0.0262419f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A3_c_251_n N_B1_c_286_n 0.0087356f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A3_M1001_g N_VPWR_c_351_n 0.00357842f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A3_M1001_g N_VPWR_c_345_n 0.00563013f $X=2.795 $Y=1.985 $X2=0 $Y2=0
cc_209 A3 A_460_297# 0.014726f $X=2.44 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_210 N_A3_c_251_n N_VGND_c_434_n 0.00467408f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A3_c_251_n N_VGND_c_437_n 0.00428022f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A3_c_251_n N_VGND_c_438_n 0.00635517f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A3_c_249_n N_A_360_47#_c_487_n 0.00135602f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A3_c_250_n N_A_360_47#_c_487_n 0.0206113f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A3_c_251_n N_A_360_47#_c_487_n 0.0144537f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_286_n N_C1_c_319_n 0.0368767f $X=3.232 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_217 N_B1_M1010_g N_C1_M1003_g 0.0246074f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_c_284_n N_C1_c_321_n 0.0368767f $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B1_c_285_n N_C1_c_321_n 2.80449e-19 $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B1_M1010_g N_VPWR_c_350_n 0.00510038f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B1_M1010_g N_VPWR_c_351_n 0.00539841f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_222 N_B1_M1010_g N_VPWR_c_345_n 0.00964112f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B1_c_286_n N_VGND_c_437_n 0.00585385f $X=3.232 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B1_c_286_n N_VGND_c_438_n 0.0108442f $X=3.232 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B1_c_284_n N_A_360_47#_c_495_n 0.00340725f $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_226 N_B1_c_285_n N_A_360_47#_c_495_n 0.0236139f $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_227 N_C1_M1003_g N_VPWR_c_350_n 0.00307308f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_228 N_C1_M1003_g N_VPWR_c_352_n 0.00583607f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_229 N_C1_M1003_g N_VPWR_c_345_n 0.0115712f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_230 N_C1_c_319_n N_VGND_c_437_n 0.00357668f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_231 N_C1_c_319_n N_VGND_c_438_n 0.00604465f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_232 N_VPWR_c_345_n N_X_M1002_s 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_c_347_n X 0.0758332f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_234 N_VPWR_c_348_n X 0.0206084f $X=1.075 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_345_n X 0.0130702f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_c_347_n N_X_c_404_n 0.0250529f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_237 N_VPWR_c_345_n A_360_297# 0.00281079f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_238 N_VPWR_c_345_n A_460_297# 0.00338304f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_239 X N_VGND_c_432_n 0.0478331f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_240 N_X_c_404_n N_VGND_c_432_n 0.0250529f $X=0.55 $Y=1.185 $X2=0 $Y2=0
cc_241 X N_VGND_c_435_n 0.0168871f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_242 N_X_M1009_s N_VGND_c_438_n 0.00393857f $X=0.605 $Y=0.235 $X2=0 $Y2=0
cc_243 X N_VGND_c_438_n 0.0102668f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_244 N_VGND_c_438_n N_A_360_47#_M1013_d 0.0042111f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_245 N_VGND_c_438_n N_A_360_47#_M1005_d 0.00354962f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_246 N_VGND_c_436_n N_A_360_47#_c_499_n 0.0132692f $X=2.3 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_438_n N_A_360_47#_c_499_n 0.0105075f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_M1012_d N_A_360_47#_c_487_n 0.00888498f $X=2.3 $Y=0.235 $X2=0
+ $Y2=0
cc_249 N_VGND_c_434_n N_A_360_47#_c_487_n 0.0234908f $X=2.51 $Y=0.36 $X2=0 $Y2=0
cc_250 N_VGND_c_436_n N_A_360_47#_c_487_n 0.00260706f $X=2.3 $Y=0 $X2=0 $Y2=0
cc_251 N_VGND_c_437_n N_A_360_47#_c_487_n 0.00293207f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_438_n N_A_360_47#_c_487_n 0.0110612f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_437_n N_A_360_47#_c_506_n 0.0148394f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_438_n N_A_360_47#_c_506_n 0.0121783f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_438_n A_677_47# 0.00467183f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

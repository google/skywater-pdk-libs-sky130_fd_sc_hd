# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.780000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.280000 1.275000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 1.445000 4.055000 1.625000 ;
        RECT 1.905000 1.625000 3.625000 1.765000 ;
        RECT 3.295000 0.635000 4.055000 0.855000 ;
        RECT 3.295000 1.765000 3.625000 2.125000 ;
        RECT 3.825000 0.855000 4.055000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 0.320000 1.845000 ;
      RECT 0.085000  1.845000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.850000 0.595000 ;
      RECT 0.515000  1.845000 0.950000 2.635000 ;
      RECT 1.020000  0.255000 1.730000 0.595000 ;
      RECT 1.120000  1.445000 1.735000 1.765000 ;
      RECT 1.120000  1.765000 1.410000 2.465000 ;
      RECT 1.450000  0.595000 1.730000 1.025000 ;
      RECT 1.450000  1.025000 2.965000 1.275000 ;
      RECT 1.450000  1.275000 1.735000 1.445000 ;
      RECT 1.600000  1.935000 3.125000 2.105000 ;
      RECT 1.600000  2.105000 1.810000 2.465000 ;
      RECT 1.900000  0.255000 2.170000 0.655000 ;
      RECT 1.900000  0.655000 3.125000 0.855000 ;
      RECT 1.980000  2.275000 2.310000 2.635000 ;
      RECT 2.340000  0.085000 2.670000 0.485000 ;
      RECT 2.480000  2.105000 3.125000 2.295000 ;
      RECT 2.480000  2.295000 4.055000 2.465000 ;
      RECT 2.840000  0.275000 4.050000 0.465000 ;
      RECT 2.840000  0.465000 3.125000 0.655000 ;
      RECT 3.245000  1.025000 3.655000 1.275000 ;
      RECT 3.795000  1.795000 4.055000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.105000 0.320000 1.275000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.380000  1.105000 3.550000 1.275000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 3.610000 1.260000 ;
      RECT 0.085000 1.260000 0.380000 1.305000 ;
      RECT 3.320000 1.075000 3.610000 1.120000 ;
      RECT 3.320000 1.260000 3.610000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_2
END LIBRARY

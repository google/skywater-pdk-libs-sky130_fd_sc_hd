* File: sky130_fd_sc_hd__lpflow_decapkapwr_12.pxi.spice
* Created: Tue Sep  1 19:11:33 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%VGND N_VGND_M1001_s N_VGND_M1000_g
+ N_VGND_c_22_n N_VGND_c_23_n VGND N_VGND_c_24_n N_VGND_c_25_n N_VGND_c_26_n
+ N_VGND_c_27_n PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%KAPWR N_KAPWR_M1000_s N_KAPWR_M1001_g
+ N_KAPWR_c_50_n N_KAPWR_c_55_n KAPWR N_KAPWR_c_51_n N_KAPWR_c_52_n
+ N_KAPWR_c_53_n N_KAPWR_c_57_n N_KAPWR_c_58_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%VPWR VPWR N_VPWR_c_81_n N_VPWR_c_80_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%VPWR
cc_1 VNB N_VGND_c_22_n 0.0304509f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=0.385
cc_2 VNB N_VGND_c_23_n 0.0927609f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=0.385
cc_3 VNB N_VGND_c_24_n 0.0491357f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.87
cc_4 VNB N_VGND_c_25_n 0.0241734f $X=-0.19 $Y=-0.24 $X2=2.645 $Y2=1.87
cc_5 VNB N_VGND_c_26_n 0.0439214f $X=-0.19 $Y=-0.24 $X2=5.26 $Y2=0.475
cc_6 VNB N_VGND_c_27_n 0.274429f $X=-0.19 $Y=-0.24 $X2=5.29 $Y2=0
cc_7 VNB N_KAPWR_c_50_n 0.00216151f $X=-0.19 $Y=-0.24 $X2=4.96 $Y2=0.385
cc_8 VNB N_KAPWR_c_51_n 0.173698f $X=-0.19 $Y=-0.24 $X2=2.645 $Y2=1.87
cc_9 VNB N_KAPWR_c_52_n 0.266166f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0
cc_10 VNB N_KAPWR_c_53_n 0.015517f $X=-0.19 $Y=-0.24 $X2=5.29 $Y2=0
cc_11 VNB N_VPWR_c_80_n 0.231782f $X=-0.19 $Y=-0.24 $X2=2.76 $Y2=2.05
cc_12 VPB N_VGND_c_23_n 0.00687456f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=0.385
cc_13 VPB N_VGND_c_24_n 0.139048f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.87
cc_14 VPB N_VGND_c_25_n 0.254589f $X=-0.19 $Y=1.305 $X2=2.645 $Y2=1.87
cc_15 VPB N_KAPWR_c_50_n 0.00170143f $X=-0.19 $Y=1.305 $X2=4.96 $Y2=0.385
cc_16 VPB N_KAPWR_c_55_n 0.0353425f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.87
cc_17 VPB N_KAPWR_c_53_n 0.0431548f $X=-0.19 $Y=1.305 $X2=5.29 $Y2=0
cc_18 VPB N_KAPWR_c_57_n 0.0113645f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0
cc_19 VPB N_KAPWR_c_58_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_81_n 0.128316f $X=-0.19 $Y=1.305 $X2=2.76 $Y2=2.05
cc_21 VPB N_VPWR_c_80_n 0.0425047f $X=-0.19 $Y=1.305 $X2=2.76 $Y2=2.05
cc_22 N_VGND_c_22_n N_KAPWR_c_50_n 0.178146f $X=4.96 $Y=0.385 $X2=0 $Y2=0
cc_23 N_VGND_c_23_n N_KAPWR_c_50_n 0.0326918f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_24 N_VGND_c_25_n N_KAPWR_c_50_n 0.0889517f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_25 N_VGND_c_23_n N_KAPWR_c_55_n 0.220132f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_26 N_VGND_c_24_n N_KAPWR_c_55_n 0.168296f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_27 N_VGND_c_25_n N_KAPWR_c_55_n 0.102805f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_28 N_VGND_c_22_n N_KAPWR_c_51_n 0.0203072f $X=4.96 $Y=0.385 $X2=0 $Y2=0
cc_29 N_VGND_c_23_n N_KAPWR_c_51_n 0.247023f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_30 N_VGND_c_24_n N_KAPWR_c_51_n 0.147138f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_31 N_VGND_c_25_n N_KAPWR_c_51_n 0.00421134f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_32 N_VGND_c_22_n N_KAPWR_c_52_n 0.21632f $X=4.96 $Y=0.385 $X2=0 $Y2=0
cc_33 N_VGND_c_23_n N_KAPWR_c_52_n 0.00652589f $X=2.665 $Y=0.385 $X2=0 $Y2=0
cc_34 N_VGND_c_25_n N_KAPWR_c_52_n 0.158306f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_35 N_VGND_c_26_n N_KAPWR_c_52_n 0.0242125f $X=5.26 $Y=0.475 $X2=0 $Y2=0
cc_36 N_VGND_c_25_n N_KAPWR_c_53_n 0.177935f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_37 N_VGND_c_26_n N_KAPWR_c_53_n 0.0423591f $X=5.26 $Y=0.475 $X2=0 $Y2=0
cc_38 N_VGND_c_24_n N_VPWR_c_81_n 0.112808f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_39 N_VGND_c_24_n N_VPWR_c_80_n 0.0324745f $X=1.9 $Y=1.87 $X2=0 $Y2=0
cc_40 N_VGND_c_25_n N_VPWR_c_80_n 0.0676482f $X=2.645 $Y=1.87 $X2=0 $Y2=0
cc_41 N_KAPWR_c_55_n N_VPWR_c_81_n 0.359353f $X=2.835 $Y=1.745 $X2=0 $Y2=0
cc_42 N_KAPWR_c_58_n N_VPWR_c_81_n 0.00372207f $X=0.215 $Y=2.21 $X2=0 $Y2=0
cc_43 N_KAPWR_M1000_s N_VPWR_c_80_n 0.00214099f $X=0.135 $Y=1.615 $X2=0 $Y2=0
cc_44 N_KAPWR_c_55_n N_VPWR_c_80_n 0.0445025f $X=2.835 $Y=1.745 $X2=0 $Y2=0
cc_45 N_KAPWR_c_58_n N_VPWR_c_80_n 0.549307f $X=0.215 $Y=2.21 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o2bb2a_1.pex.spice
* Created: Thu Aug 27 14:38:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%A_76_199# 1 2 9 12 16 17 20 21 22 26 29 32
+ 35 36 37 41
c98 12 0 1.14156e-19 $X=0.47 $Y=1.985
r99 37 39 2.25 $w=4.88e-07 $l=9e-08 $layer=LI1_cond $X=2.457 $Y=1.97 $X2=2.457
+ $Y2=2.06
r100 35 36 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.252 $Y=1.075
+ $X2=2.252 $Y2=1.245
r101 34 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.24 $Y=0.69
+ $X2=2.24 $Y2=1.075
r102 32 34 10.6372 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=2.2 $Y=0.485
+ $X2=2.2 $Y2=0.69
r103 27 29 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.515 $Y=1.53
+ $X2=0.74 $Y2=1.53
r104 26 37 17.3831 $w=4.88e-07 $l=5.62872e-07 $layer=LI1_cond $X=2.265 $Y=1.495
+ $X2=2.457 $Y2=1.97
r105 26 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.265 $Y=1.495
+ $X2=2.265 $Y2=1.245
r106 21 37 7.00443 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=2.18 $Y=1.97
+ $X2=2.457 $Y2=1.97
r107 21 22 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=2.18 $Y=1.97
+ $X2=0.825 $Y2=1.97
r108 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.74 $Y=1.885
+ $X2=0.825 $Y2=1.97
r109 19 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=1.615
+ $X2=0.74 $Y2=1.53
r110 19 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.74 $Y=1.615
+ $X2=0.74 $Y2=1.885
r111 17 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r112 17 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r113 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r114 14 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.515 $Y=1.445
+ $X2=0.515 $Y2=1.53
r115 14 16 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=1.445
+ $X2=0.515 $Y2=1.16
r116 12 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r117 9 41 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
r118 2 39 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.845 $X2=2.59 $Y2=2.06
r119 1 32 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.235 $X2=2.16 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%A1_N 3 7 9 12 20
c38 20 0 1.51767e-19 $X=1.155 $Y=1.19
r39 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=1.325
r40 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=0.995
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r42 9 20 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=1.135 $Y=1.175
+ $X2=1.155 $Y2=1.175
r43 9 13 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=1.135 $Y=1.175
+ $X2=0.995 $Y2=1.175
r44 7 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.955 $Y=2.055
+ $X2=0.955 $Y2=1.325
r45 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.95 $Y=0.445
+ $X2=0.95 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%A2_N 3 6 8 12 13 16
c45 12 0 1.51767e-19 $X=1.475 $Y=0.935
r46 12 17 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=1.1
r47 12 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.77
r48 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.475
+ $Y=0.935 $X2=1.475 $Y2=0.935
r49 9 13 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.18 $Y=0.735
+ $X2=1.18 $Y2=0.51
r50 8 11 15.1218 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.18 $Y=0.905
+ $X2=1.475 $Y2=0.905
r51 8 9 1.19154 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=1.18 $Y=0.905 $X2=1.18
+ $Y2=0.735
r52 6 17 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=1.505 $Y=2.055
+ $X2=1.505 $Y2=1.1
r53 3 16 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.415 $Y=0.445
+ $X2=1.415 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%A_206_369# 1 2 9 13 15 16 17 21 28 30
c70 17 0 1.14156e-19 $X=1.735 $Y=1.605
r71 28 30 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.872 $Y=1.52
+ $X2=1.872 $Y2=1.355
r72 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.52 $X2=1.925 $Y2=1.52
r73 25 30 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.82 $Y=0.565
+ $X2=1.82 $Y2=1.355
r74 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.735 $Y=0.48
+ $X2=1.82 $Y2=0.565
r75 21 23 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.735 $Y=0.48
+ $X2=1.625 $Y2=0.48
r76 17 28 3.5621 $w=2.73e-07 $l=8.5e-08 $layer=LI1_cond $X=1.872 $Y=1.605
+ $X2=1.872 $Y2=1.52
r77 17 19 26.4538 $w=2.18e-07 $l=5.05e-07 $layer=LI1_cond $X=1.735 $Y=1.605
+ $X2=1.23 $Y2=1.605
r78 15 29 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.295 $Y=1.52
+ $X2=1.925 $Y2=1.52
r79 15 16 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.52
+ $X2=2.295 $Y2=1.355
r80 11 16 37.0704 $w=1.5e-07 $l=3.70068e-07 $layer=POLY_cond $X=2.38 $Y=1.685
+ $X2=2.295 $Y2=1.355
r81 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.38 $Y=1.685
+ $X2=2.38 $Y2=2.055
r82 7 16 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.355
+ $X2=2.295 $Y2=1.355
r83 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.37 $Y=1.355 $X2=2.37
+ $Y2=0.445
r84 2 19 600 $w=1.7e-07 $l=2.98706e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.845 $X2=1.23 $Y2=1.63
r85 1 23 182 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.235 $X2=1.625 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%B2 3 7 9 12 15
r51 14 15 14.2914 $w=1.75e-07 $l=2.05e-07 $layer=LI1_cond $X=2.992 $Y=1.325
+ $X2=2.992 $Y2=1.53
r52 12 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.16
+ $X2=2.79 $Y2=1.325
r53 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.16 $X2=2.79 $Y2=1.16
r54 9 14 7.09627 $w=2.5e-07 $l=1.62788e-07 $layer=LI1_cond $X=2.905 $Y=1.2
+ $X2=2.992 $Y2=1.325
r55 9 11 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.905 $Y=1.2
+ $X2=2.79 $Y2=1.2
r56 7 18 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.85 $Y=2.055
+ $X2=2.85 $Y2=1.325
r57 1 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.995
+ $X2=2.79 $Y2=1.16
r58 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.79 $Y=0.995 $X2=2.79
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%B1 3 7 9 10 16
r27 13 16 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.415 $Y2=1.16
r28 9 10 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.422 $Y=1.16
+ $X2=3.422 $Y2=1.53
r29 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.16 $X2=3.415 $Y2=1.16
r30 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r31 5 7 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.21 $Y=1.325 $X2=3.21
+ $Y2=2.055
r32 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r33 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.21 $Y=0.995 $X2=3.21
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%X 1 2 9 13 14 15 16 19
r23 16 19 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.215 $Y=2.21
+ $X2=0.215 $Y2=1.96
r24 14 19 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.215 $Y=1.925
+ $X2=0.215 $Y2=1.96
r25 14 15 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.925
+ $X2=0.215 $Y2=1.795
r26 13 15 61.4753 $w=1.73e-07 $l=9.7e-07 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=1.795
r27 7 13 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.655
+ $X2=0.255 $Y2=0.825
r28 7 9 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.255 $Y=0.655
+ $X2=0.255 $Y2=0.38
r29 2 19 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r30 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%VPWR 1 2 3 12 14 16 18 20 25 30 36 39 47
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 39 42 11.5244 $w=3.98e-07 $l=4e-07 $layer=LI1_cond $X=1.915 $Y=2.32
+ $X2=1.915 $Y2=2.72
r54 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 34 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 31 42 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.115 $Y=2.72 $X2=1.915
+ $Y2=2.72
r59 31 33 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 30 46 4.94809 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.25 $Y=2.72
+ $X2=3.465 $Y2=2.72
r61 30 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.25 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 29 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 29 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r66 26 28 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r67 25 42 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.715 $Y=2.72 $X2=1.915
+ $Y2=2.72
r68 25 28 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.715 $Y=2.72
+ $X2=1.61 $Y2=2.72
r69 20 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r70 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 14 46 2.94584 $w=3.45e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.422 $Y=2.635
+ $X2=3.465 $Y2=2.72
r74 14 16 19.2074 $w=3.43e-07 $l=5.75e-07 $layer=LI1_cond $X=3.422 $Y=2.635
+ $X2=3.422 $Y2=2.06
r75 10 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r76 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.32
r77 3 16 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.845 $X2=3.42 $Y2=2.06
r78 2 39 600 $w=1.7e-07 $l=6.20282e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.845 $X2=1.915 $Y2=2.32
r79 1 12 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%VGND 1 2 11 15 17 19 26 27 30 33 36
r52 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r53 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 27 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r55 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0 $X2=3
+ $Y2=0
r57 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.45
+ $Y2=0
r58 23 34 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r59 23 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r60 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.705
+ $Y2=0
r62 20 22 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=1.15
+ $Y2=0
r63 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0 $X2=3
+ $Y2=0
r64 19 22 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.915 $Y=0 $X2=1.15
+ $Y2=0
r65 17 31 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r66 17 36 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r67 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0
r68 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0.39
r69 9 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r70 9 11 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.525
r71 2 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3 $Y2=0.39
r72 1 11 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.705 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_1%A_489_47# 1 2 9 11 12 15
r32 13 15 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=3.425 $Y=0.725
+ $X2=3.425 $Y2=0.435
r33 11 13 7.6914 $w=1.8e-07 $l=2.10238e-07 $layer=LI1_cond $X=3.255 $Y=0.815
+ $X2=3.425 $Y2=0.725
r34 11 12 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.255 $Y=0.815
+ $X2=2.745 $Y2=0.815
r35 7 12 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.62 $Y=0.725
+ $X2=2.745 $Y2=0.815
r36 7 9 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=2.62 $Y=0.725 $X2=2.62
+ $Y2=0.485
r37 2 15 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.435
r38 1 9 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.235 $X2=2.58 $Y2=0.485
.ends


* File: sky130_fd_sc_hd__o21a_2.spice
* Created: Thu Aug 27 14:35:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21a_2.pex.spice"
.subckt sky130_fd_sc_hd__o21a_2  VNB VPB B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_79_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.089375 PD=1.82 PS=0.925 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_79_21#_M1009_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.089375 PD=1.83 PS=0.925 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_384_47#_M1004_d N_B1_M1004_g N_A_79_21#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_384_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.091 PD=0.97 PS=0.93 NRD=3.684 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_A_384_47#_M1005_d N_A1_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.104 PD=1.83 PS=0.97 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_79_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1375 PD=2.52 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A_79_21#_M1008_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.4 AS=0.1375 PD=1.8 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1006 N_A_79_21#_M1006_d N_B1_M1006_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.4 PD=1.28 PS=1.8 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1002 A_470_297# N_A2_M1002_g N_A_79_21#_M1006_d VPB PHIGHVT L=0.15 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=20.6653 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_470_297# VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.16 PD=2.53 PS=1.32 NRD=0 NRS=20.6653 M=1 R=6.66667 SA=75002.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o21a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__dlrtn_2.spice.pex
* Created: Thu Aug 27 14:17:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRTN_2%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%A_27_47# 1 2 9 13 17 21 25 29 30 31 39 40 43
+ 46 48 53 55 57 58 61 64 65 69 79
c166 79 0 9.36962e-20 $X=3.095 $Y=1.415
c167 21 0 1.66856e-19 $X=3.15 $Y=2.275
c168 13 0 2.6965e-20 $X=0.89 $Y=2.135
c169 9 0 2.6965e-20 $X=0.89 $Y=0.445
r170 65 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.095 $Y=1.53
+ $X2=3.095 $Y2=1.415
r171 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.53
+ $X2=3.015 $Y2=1.53
r172 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r173 58 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 57 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=3.015 $Y2=1.53
r175 57 58 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=0.84 $Y2=1.53
r176 53 72 41.0874 $w=3.35e-07 $l=1.35e-07 $layer=POLY_cond $X=2.762 $Y=0.9
+ $X2=2.762 $Y2=0.765
r177 52 55 6.41701 $w=4.38e-07 $l=2.45e-07 $layer=LI1_cond $X=2.765 $Y=0.925
+ $X2=3.01 $Y2=0.925
r178 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=0.9 $X2=2.765 $Y2=0.9
r179 50 61 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r180 49 61 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r181 47 69 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r182 46 49 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r183 46 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r184 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r185 40 76 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.18 $Y2=1.875
r186 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r187 37 65 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.53
r188 37 39 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.74
r189 35 55 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.01 $Y=1.145
+ $X2=3.01 $Y2=0.925
r190 35 79 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.01 $Y=1.145
+ $X2=3.01 $Y2=1.415
r191 33 48 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r192 32 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r193 31 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r194 31 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r195 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r196 29 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r197 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r198 23 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r199 21 76 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.15 $Y=2.275
+ $X2=3.15 $Y2=1.875
r200 17 72 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.725 $Y=0.415
+ $X2=2.725 $Y2=0.765
r201 11 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r202 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r203 7 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r204 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r205 2 43 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r206 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%D 3 7 9 13 15
c40 13 0 1.09751e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%A_299_47# 1 2 7 9 12 16 18 20 21 22 23 25 32
c82 32 0 1.97325e-19 $X=2.25 $Y=0.93
r83 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=0.93 $X2=2.25 $Y2=0.93
r84 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r85 22 31 8.60998 $w=3.17e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.05 $Y=1.095
+ $X2=2.15 $Y2=0.93
r86 22 23 24.6465 $w=1.78e-07 $l=4e-07 $layer=LI1_cond $X=2.05 $Y=1.095 $X2=2.05
+ $Y2=1.495
r87 20 23 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.96 $Y=1.58
+ $X2=2.05 $Y2=1.495
r88 20 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.96 $Y=1.58
+ $X2=1.785 $Y2=1.58
r89 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r90 18 31 8.85174 $w=3.17e-07 $l=3.10805e-07 $layer=LI1_cond $X=1.96 $Y=0.7
+ $X2=2.15 $Y2=0.93
r91 18 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.96 $Y=0.7
+ $X2=1.705 $Y2=0.7
r92 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r93 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r94 10 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.095
+ $X2=2.25 $Y2=0.93
r95 10 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=1.095
+ $X2=2.25 $Y2=2.165
r96 7 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.765
+ $X2=2.25 $Y2=0.93
r97 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.765 $X2=2.25
+ $Y2=0.445
r98 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r99 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c113 38 0 1.66856e-19 $X=2.67 $Y=1.52
r114 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r115 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.612 $Y=1.87
+ $X2=2.612 $Y2=1.52
r116 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.87
+ $X2=2.555 $Y2=1.87
r117 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r119 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=2.555 $Y2=1.87
r120 26 27 1.37376 $w=1.4e-07 $l=1.11e-06 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=1.3 $Y2=1.87
r121 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r122 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r123 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r124 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r125 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r126 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r127 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.215 $Y=1.245
+ $X2=3.215 $Y2=0.415
r128 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r129 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.14 $Y=1.32
+ $X2=3.215 $Y2=1.245
r130 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.14 $Y=1.32
+ $X2=2.805 $Y2=1.32
r131 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r132 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r133 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%A_711_307# 1 2 9 13 17 19 21 22 24 27 29 32
+ 36 38 39 42 44 49 51 53 55 66
c135 66 0 5.5665e-20 $X=5.97 $Y=1.16
c136 13 0 9.36962e-20 $X=3.69 $Y=0.445
r137 65 66 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.55 $Y=1.16
+ $X2=5.97 $Y2=1.16
r138 57 59 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.63 $Y=1.7 $X2=3.69
+ $Y2=1.7
r139 54 65 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.53 $Y=1.16 $X2=5.55
+ $Y2=1.16
r140 54 62 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.53 $Y=1.16
+ $X2=5.515 $Y2=1.16
r141 53 56 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.482 $Y=1.16
+ $X2=5.482 $Y2=1.325
r142 53 55 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.482 $Y=1.16
+ $X2=5.482 $Y2=0.995
r143 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.16 $X2=5.53 $Y2=1.16
r144 49 56 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.5 $Y=1.535
+ $X2=5.5 $Y2=1.325
r145 46 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.5 $Y=0.825
+ $X2=5.5 $Y2=0.995
r146 45 51 4.08801 $w=2.5e-07 $l=1.28938e-07 $layer=LI1_cond $X=4.92 $Y=1.62
+ $X2=4.825 $Y2=1.7
r147 44 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=1.62
+ $X2=5.5 $Y2=1.535
r148 44 45 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.415 $Y=1.62
+ $X2=4.92 $Y2=1.62
r149 40 51 2.34704 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=1.865
+ $X2=4.825 $Y2=1.7
r150 40 42 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=4.825 $Y=1.865
+ $X2=4.825 $Y2=2.27
r151 38 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=0.74
+ $X2=5.5 $Y2=0.825
r152 38 39 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.415 $Y=0.74
+ $X2=4.59 $Y2=0.74
r153 34 39 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.415 $Y=0.655
+ $X2=4.59 $Y2=0.74
r154 34 36 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.415 $Y=0.655
+ $X2=4.415 $Y2=0.4
r155 32 59 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.69 $Y2=1.7
r156 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r157 29 51 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.73 $Y=1.7
+ $X2=4.825 $Y2=1.7
r158 29 31 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=4.73 $Y=1.7
+ $X2=3.925 $Y2=1.7
r159 25 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.325
+ $X2=5.97 $Y2=1.16
r160 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.97 $Y=1.325
+ $X2=5.97 $Y2=1.985
r161 22 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=1.16
r162 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=0.56
r163 19 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.55 $Y=0.995
+ $X2=5.55 $Y2=1.16
r164 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.55 $Y=0.995
+ $X2=5.55 $Y2=0.56
r165 15 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.515 $Y=1.325
+ $X2=5.515 $Y2=1.16
r166 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.515 $Y=1.325
+ $X2=5.515 $Y2=1.985
r167 11 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=1.535
+ $X2=3.69 $Y2=1.7
r168 11 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.69 $Y=1.535
+ $X2=3.69 $Y2=0.445
r169 7 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=1.7
r170 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=2.275
r171 2 51 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=1.485 $X2=4.825 $Y2=1.755
r172 2 42 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=1.485 $X2=4.825 $Y2=2.27
r173 1 36 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.295
+ $Y=0.235 $X2=4.42 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%A_560_47# 1 2 9 13 15 16 17 21 26 28 31 34
c86 34 0 1.54454e-19 $X=3.33 $Y=1.025
c87 31 0 1.01992e-19 $X=4.145 $Y=1.16
c88 9 0 6.36774e-20 $X=4.615 $Y=1.985
r89 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=1.16 $X2=4.145 $Y2=1.16
r90 29 34 0.597483 $w=3e-07 $l=3.4187e-07 $layer=LI1_cond $X=3.605 $Y=1.175
+ $X2=3.33 $Y2=1.025
r91 29 31 20.744 $w=2.98e-07 $l=5.4e-07 $layer=LI1_cond $X=3.605 $Y=1.175
+ $X2=4.145 $Y2=1.175
r92 27 34 8.04615 $w=1.7e-07 $l=3.83406e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.33 $Y2=1.025
r93 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=2.255
r94 26 34 8.04615 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.025
+ $X2=3.33 $Y2=1.025
r95 25 26 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=1.025
r96 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r97 21 23 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=2.98 $Y2=0.45
r98 17 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.435 $Y=2.34
+ $X2=3.52 $Y2=2.255
r99 17 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.435 $Y=2.34
+ $X2=2.94 $Y2=2.34
r100 15 32 87.7586 $w=2.7e-07 $l=3.95e-07 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.145 $Y2=1.16
r101 15 16 2.60871 $w=2.7e-07 $l=8.2994e-08 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.622 $Y2=1.162
r102 11 16 32.2453 $w=1.5e-07 $l=1.40943e-07 $layer=POLY_cond $X=4.63 $Y=1.025
+ $X2=4.622 $Y2=1.162
r103 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.63 $Y=1.025
+ $X2=4.63 $Y2=0.56
r104 7 16 32.2453 $w=1.5e-07 $l=1.41457e-07 $layer=POLY_cond $X=4.615 $Y=1.3
+ $X2=4.622 $Y2=1.162
r105 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=4.615 $Y=1.3
+ $X2=4.615 $Y2=1.985
r106 2 19 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=2.94 $Y2=2.34
r107 1 23 182 $w=1.7e-07 $l=2.91419e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.98 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%RESET_B 3 5 7 8 11 12
c40 11 0 1.01992e-19 $X=5.05 $Y=1.16
r41 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.16
+ $X2=5.05 $Y2=1.325
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.16 $X2=5.05 $Y2=1.16
r43 8 12 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.855 $Y=1.16
+ $X2=5.05 $Y2=1.16
r44 5 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=1.16
r45 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.995 $X2=5.05
+ $Y2=0.56
r46 3 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.035 $Y=1.985
+ $X2=5.035 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 43 45
+ 50 55 63 64 68 74 77 84 88
r105 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r106 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r107 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r110 72 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 72 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r112 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r113 69 84 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.46 $Y=2.72
+ $X2=5.275 $Y2=2.72
r114 69 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.46 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 68 87 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.267 $Y2=2.72
r116 68 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r117 67 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 67 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r119 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r120 64 81 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.56 $Y=2.72
+ $X2=4.37 $Y2=2.72
r121 64 66 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.56 $Y=2.72
+ $X2=4.83 $Y2=2.72
r122 63 84 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.09 $Y=2.72
+ $X2=5.275 $Y2=2.72
r123 63 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.09 $Y=2.72
+ $X2=4.83 $Y2=2.72
r124 62 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r127 59 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r128 58 61 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r130 56 77 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r131 56 58 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r132 55 61 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.8 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 54 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 54 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r136 51 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r137 51 53 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r138 50 77 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r139 50 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 45 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r141 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r142 43 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r143 43 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r144 39 87 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.225 $Y=2.635
+ $X2=6.267 $Y2=2.72
r145 39 41 35.4598 $w=2.58e-07 $l=8e-07 $layer=LI1_cond $X=6.225 $Y=2.635
+ $X2=6.225 $Y2=1.835
r146 35 84 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.275 $Y=2.635
+ $X2=5.275 $Y2=2.72
r147 35 37 19.1555 $w=3.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.275 $Y=2.635
+ $X2=5.275 $Y2=2.02
r148 33 81 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.42 $Y=2.34
+ $X2=4.42 $Y2=2.635
r149 27 81 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=4.37 $Y2=2.72
r150 27 55 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=3.8 $Y2=2.72
r151 27 29 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.955 $Y=2.635
+ $X2=3.955 $Y2=2.34
r152 23 77 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r153 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r154 19 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r155 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r156 6 41 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=1.835
r157 5 37 300 $w=1.7e-07 $l=6.11964e-07 $layer=licon1_PDIFF $count=2 $X=5.11
+ $Y=1.485 $X2=5.275 $Y2=2.02
r158 4 33 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.485 $X2=4.405 $Y2=2.34
r159 3 29 600 $w=1.7e-07 $l=3.5373e-07 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=2.065 $X2=3.885 $Y2=2.34
r160 2 25 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r161 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%Q 1 2 8 14 16 17 18 19 20 21 31 37
r48 31 37 0.81742 $w=5.97e-07 $l=4.69042e-08 $layer=LI1_cond $X=6.07 $Y=0.89
+ $X2=6.055 $Y2=0.85
r49 20 37 0.470017 $w=5.97e-07 $l=2.3e-08 $layer=LI1_cond $X=6.055 $Y=0.827
+ $X2=6.055 $Y2=0.85
r50 20 21 5.83351 $w=5.68e-07 $l=2.78e-07 $layer=LI1_cond $X=6.07 $Y=0.912
+ $X2=6.07 $Y2=1.19
r51 20 31 0.461644 $w=5.68e-07 $l=2.2e-08 $layer=LI1_cond $X=6.07 $Y=0.912
+ $X2=6.07 $Y2=0.89
r52 19 29 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=5.79 $Y=2.21 $X2=5.79
+ $Y2=2.3
r53 18 21 4.09185 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.07 $Y=1.385
+ $X2=6.07 $Y2=1.19
r54 16 19 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=5.79 $Y=2.01 $X2=5.79
+ $Y2=2.21
r55 16 17 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.79 $Y=2.01
+ $X2=5.79 $Y2=1.875
r56 12 14 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=5.76 $Y=0.37 $X2=5.84
+ $Y2=0.37
r57 9 18 2.36195 $w=5.94e-07 $l=2.81691e-07 $layer=LI1_cond $X=5.84 $Y=1.5
+ $X2=6.07 $Y2=1.385
r58 9 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.84 $Y=1.5 $X2=5.84
+ $Y2=1.875
r59 8 20 8.23439 $w=5.97e-07 $l=2.44039e-07 $layer=LI1_cond $X=5.84 $Y=0.765
+ $X2=6.055 $Y2=0.827
r60 7 14 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.84 $Y=0.485
+ $X2=5.84 $Y2=0.37
r61 7 8 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.84 $Y=0.485 $X2=5.84
+ $Y2=0.765
r62 2 29 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.59
+ $Y=1.485 $X2=5.74 $Y2=2.3
r63 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.76 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_2%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 56 61 67 70 73 76 80
c105 80 0 2.71124e-20 $X=6.21 $Y=0
c106 30 0 5.5665e-20 $X=5.26 $Y=0.36
c107 22 0 8.7574e-20 $X=2.04 $Y=0.36
r108 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r109 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r110 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r111 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r112 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r113 65 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r114 65 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r115 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r116 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.425 $Y=0 $X2=5.26
+ $Y2=0
r117 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.425 $Y=0
+ $X2=5.75 $Y2=0
r118 61 79 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.267 $Y2=0
r119 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.75
+ $Y2=0
r120 60 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r121 60 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r122 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r123 57 73 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.902
+ $Y2=0
r124 57 59 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.83
+ $Y2=0
r125 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=5.26
+ $Y2=0
r126 56 59 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.095 $Y=0
+ $X2=4.83 $Y2=0
r127 55 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r128 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r129 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r130 52 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r131 51 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r132 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r133 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r134 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r135 48 73 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.902 $Y2=0
r136 48 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.45 $Y2=0
r137 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r138 47 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r139 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r140 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r141 44 46 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r142 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r143 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r144 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r145 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r146 36 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r147 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r148 32 79 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.267 $Y2=0
r149 32 34 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0.38
r150 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.26 $Y=0.085
+ $X2=5.26 $Y2=0
r151 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.26 $Y=0.085
+ $X2=5.26 $Y2=0.36
r152 24 73 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.902 $Y=0.085
+ $X2=3.902 $Y2=0
r153 24 26 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=3.902 $Y=0.085
+ $X2=3.902 $Y2=0.445
r154 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r155 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r156 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r157 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r158 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.38
r159 4 30 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.26 $Y2=0.36
r160 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.235 $X2=3.9 $Y2=0.445
r161 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r162 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


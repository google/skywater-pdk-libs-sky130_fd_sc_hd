* File: sky130_fd_sc_hd__dlrtp_2.spice
* Created: Thu Aug 27 14:17:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlrtp_2.spice.pex"
.subckt sky130_fd_sc_hd__dlrtp_2  VNB VPB GATE D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_GATE_M1020_g N_A_27_47#_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_193_47#_M1012_d N_A_27_47#_M1012_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g N_A_299_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 A_465_47# N_A_299_47#_M1007_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.0567 PD=0.802308 PS=0.69 NRD=32.628 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1017 N_A_560_47#_M1017_d N_A_193_47#_M1017_g A_465_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0603 AS=0.0609231 PD=0.695 PS=0.687692 NRD=0 NRS=38.076 M=1 R=2.4
+ SA=75001.1 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1018 A_657_47# N_A_27_47#_M1018_g N_A_560_47#_M1017_d VNB NSHORT L=0.15 W=0.36
+ AD=0.0609231 AS=0.0603 PD=0.687692 PS=0.695 NRD=38.076 NRS=19.992 M=1 R=2.4
+ SA=75001.6 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1005 N_VGND_M1005_d N_A_711_307#_M1005_g A_657_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 A_940_47# N_A_560_47#_M1019_g N_A_711_307#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=19.38 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_RESET_B_M1015_g A_940_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.099125 AS=0.104 PD=0.955 PS=0.97 NRD=5.532 NRS=19.38 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_Q_M1004_d N_A_711_307#_M1004_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.099125 PD=0.92 PS=0.955 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_Q_M1004_d N_A_711_307#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_GATE_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_D_M1016_g N_A_299_47#_M1016_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1013 A_465_369# N_A_299_47#_M1013_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.115623 AS=0.0864 PD=1.16528 PS=0.91 NRD=38.6711 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_A_560_47#_M1002_d N_A_27_47#_M1002_g A_465_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0758774 PD=0.69 PS=0.764717 NRD=0 NRS=58.9227 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_644_413# N_A_193_47#_M1001_g N_A_560_47#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07035 AS=0.0567 PD=0.755 PS=0.69 NRD=52.7566 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_711_307#_M1011_g A_644_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.07035 PD=1.36 PS=0.755 NRD=0 NRS=52.7566 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_711_307#_M1006_d N_A_560_47#_M1006_g N_VPWR_M1006_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.16 AS=0.27 PD=1.32 PS=2.54 NRD=8.8453 NRS=0.9653 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_RESET_B_M1021_g N_A_711_307#_M1006_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1009 N_Q_M1009_d N_A_711_307#_M1009_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.135 PD=1.305 PS=1.27 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1014 N_Q_M1009_d N_A_711_307#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.26 PD=1.305 PS=2.52 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hd__dlrtp_2.spice.SKY130_FD_SC_HD__DLRTP_2.pxi"
*
.ends
*
*

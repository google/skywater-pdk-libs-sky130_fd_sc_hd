* File: sky130_fd_sc_hd__o311ai_4.spice.SKY130_FD_SC_HD__O311AI_4.pxi
* Created: Thu Aug 27 14:39:41 2020
* 
x_PM_SKY130_FD_SC_HD__O311AI_4%A1 N_A1_M1011_g N_A1_M1001_g N_A1_M1015_g
+ N_A1_M1009_g N_A1_M1024_g N_A1_M1012_g N_A1_M1025_g N_A1_M1027_g A1 A1 A1 A1
+ N_A1_c_157_n PM_SKY130_FD_SC_HD__O311AI_4%A1
x_PM_SKY130_FD_SC_HD__O311AI_4%A2 N_A2_M1020_g N_A2_M1000_g N_A2_M1021_g
+ N_A2_M1003_g N_A2_M1026_g N_A2_M1005_g N_A2_M1035_g N_A2_M1013_g A2 A2 A2 A2
+ N_A2_c_231_n PM_SKY130_FD_SC_HD__O311AI_4%A2
x_PM_SKY130_FD_SC_HD__O311AI_4%A3 N_A3_M1008_g N_A3_M1016_g N_A3_M1006_g
+ N_A3_M1017_g N_A3_M1014_g N_A3_M1031_g N_A3_M1030_g N_A3_M1036_g A3 A3 A3 A3
+ A3 N_A3_c_318_n PM_SKY130_FD_SC_HD__O311AI_4%A3
x_PM_SKY130_FD_SC_HD__O311AI_4%B1 N_B1_M1004_g N_B1_M1018_g N_B1_M1022_g
+ N_B1_M1019_g N_B1_M1033_g N_B1_M1028_g N_B1_M1039_g N_B1_M1032_g B1 B1 B1 B1
+ N_B1_c_408_n PM_SKY130_FD_SC_HD__O311AI_4%B1
x_PM_SKY130_FD_SC_HD__O311AI_4%C1 N_C1_M1007_g N_C1_M1002_g N_C1_M1010_g
+ N_C1_M1029_g N_C1_M1023_g N_C1_M1037_g N_C1_M1034_g N_C1_M1038_g C1 C1 C1
+ N_C1_c_479_n PM_SKY130_FD_SC_HD__O311AI_4%C1
x_PM_SKY130_FD_SC_HD__O311AI_4%A_39_297# N_A_39_297#_M1001_s N_A_39_297#_M1009_s
+ N_A_39_297#_M1027_s N_A_39_297#_M1003_d N_A_39_297#_M1013_d
+ N_A_39_297#_c_537_n N_A_39_297#_c_545_n N_A_39_297#_c_538_n
+ N_A_39_297#_c_575_p N_A_39_297#_c_550_n N_A_39_297#_c_576_p
+ N_A_39_297#_c_556_n N_A_39_297#_c_590_p N_A_39_297#_c_539_n
+ N_A_39_297#_c_540_n N_A_39_297#_c_541_n N_A_39_297#_c_542_n
+ N_A_39_297#_c_543_n PM_SKY130_FD_SC_HD__O311AI_4%A_39_297#
x_PM_SKY130_FD_SC_HD__O311AI_4%VPWR N_VPWR_M1001_d N_VPWR_M1012_d N_VPWR_M1004_s
+ N_VPWR_M1033_s N_VPWR_M1007_d N_VPWR_M1023_d N_VPWR_c_601_n N_VPWR_c_602_n
+ N_VPWR_c_603_n N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n
+ N_VPWR_c_608_n VPWR N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n
+ N_VPWR_c_612_n N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_600_n N_VPWR_c_616_n
+ N_VPWR_c_617_n N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_620_n VPWR
+ PM_SKY130_FD_SC_HD__O311AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O311AI_4%A_461_297# N_A_461_297#_M1000_s
+ N_A_461_297#_M1005_s N_A_461_297#_M1006_s N_A_461_297#_M1030_s
+ N_A_461_297#_c_741_n N_A_461_297#_c_744_n N_A_461_297#_c_746_n
+ N_A_461_297#_c_748_n N_A_461_297#_c_740_n N_A_461_297#_c_755_n
+ N_A_461_297#_c_758_n N_A_461_297#_c_761_n N_A_461_297#_c_752_n
+ N_A_461_297#_c_764_n PM_SKY130_FD_SC_HD__O311AI_4%A_461_297#
x_PM_SKY130_FD_SC_HD__O311AI_4%Y N_Y_M1002_s N_Y_M1037_s N_Y_M1006_d N_Y_M1014_d
+ N_Y_M1036_d N_Y_M1022_d N_Y_M1039_d N_Y_M1010_s N_Y_M1034_s N_Y_c_806_n
+ N_Y_c_817_n N_Y_c_807_n N_Y_c_894_n N_Y_c_823_n N_Y_c_869_n N_Y_c_830_n
+ N_Y_c_873_n N_Y_c_834_n N_Y_c_877_n N_Y_c_841_n N_Y_c_845_n N_Y_c_881_n
+ N_Y_c_851_n N_Y_c_808_n N_Y_c_809_n N_Y_c_810_n N_Y_c_811_n N_Y_c_812_n Y Y Y
+ Y Y N_Y_c_805_n N_Y_c_815_n PM_SKY130_FD_SC_HD__O311AI_4%Y
x_PM_SKY130_FD_SC_HD__O311AI_4%VGND N_VGND_M1011_s N_VGND_M1015_s N_VGND_M1025_s
+ N_VGND_M1021_s N_VGND_M1035_s N_VGND_M1016_s N_VGND_M1031_s N_VGND_c_908_n
+ N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n
+ N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n N_VGND_c_918_n
+ N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n VGND
+ N_VGND_c_923_n N_VGND_c_924_n N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n
+ N_VGND_c_928_n N_VGND_c_929_n VGND PM_SKY130_FD_SC_HD__O311AI_4%VGND
x_PM_SKY130_FD_SC_HD__O311AI_4%A_125_47# N_A_125_47#_M1011_d N_A_125_47#_M1024_d
+ N_A_125_47#_M1020_d N_A_125_47#_M1026_d N_A_125_47#_M1008_d
+ N_A_125_47#_M1017_d N_A_125_47#_M1018_s N_A_125_47#_M1028_s
+ N_A_125_47#_c_1120_n N_A_125_47#_c_1068_n N_A_125_47#_c_1061_n
+ N_A_125_47#_c_1127_n N_A_125_47#_c_1074_n N_A_125_47#_c_1134_n
+ N_A_125_47#_c_1080_n N_A_125_47#_c_1141_n N_A_125_47#_c_1084_n
+ N_A_125_47#_c_1148_n N_A_125_47#_c_1092_n N_A_125_47#_c_1155_n
+ N_A_125_47#_c_1062_n N_A_125_47#_c_1063_n N_A_125_47#_c_1064_n
+ N_A_125_47#_c_1065_n N_A_125_47#_c_1066_n N_A_125_47#_c_1067_n
+ PM_SKY130_FD_SC_HD__O311AI_4%A_125_47#
x_PM_SKY130_FD_SC_HD__O311AI_4%A_1163_47# N_A_1163_47#_M1018_d
+ N_A_1163_47#_M1019_d N_A_1163_47#_M1032_d N_A_1163_47#_M1029_d
+ N_A_1163_47#_M1038_d N_A_1163_47#_c_1167_n N_A_1163_47#_c_1168_n
+ N_A_1163_47#_c_1169_n N_A_1163_47#_c_1198_n
+ PM_SKY130_FD_SC_HD__O311AI_4%A_1163_47#
cc_1 VNB N_A1_M1011_g 0.0234384f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_2 VNB N_A1_M1001_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.985
cc_3 VNB N_A1_M1015_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=0.56
cc_4 VNB N_A1_M1009_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.985
cc_5 VNB N_A1_M1024_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=0.56
cc_6 VNB N_A1_M1012_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.985
cc_7 VNB N_A1_M1025_g 0.0174782f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=0.56
cc_8 VNB N_A1_M1027_g 4.25192e-19 $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.985
cc_9 VNB A1 0.014469f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.105
cc_10 VNB N_A1_c_157_n 0.0734085f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.16
cc_11 VNB N_A2_M1020_g 0.0174782f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_12 VNB N_A2_M1000_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.985
cc_13 VNB N_A2_M1021_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=0.56
cc_14 VNB N_A2_M1003_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.985
cc_15 VNB N_A2_M1026_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=0.56
cc_16 VNB N_A2_M1005_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.985
cc_17 VNB N_A2_M1035_g 0.0176899f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=0.56
cc_18 VNB N_A2_M1013_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.985
cc_19 VNB A2 0.0057236f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.105
cc_20 VNB N_A2_c_231_n 0.0620134f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.16
cc_21 VNB N_A3_M1008_g 0.0176899f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_22 VNB N_A3_M1016_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.985
cc_23 VNB N_A3_M1006_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=0.56
cc_24 VNB N_A3_M1017_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.985
cc_25 VNB N_A3_M1014_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=0.56
cc_26 VNB N_A3_M1031_g 0.0234087f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.985
cc_27 VNB N_A3_M1030_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=0.56
cc_28 VNB N_A3_M1036_g 3.82928e-19 $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.985
cc_29 VNB A3 0.00473476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A3_c_318_n 0.103877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_B1_M1004_g 3.82928e-19 $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_32 VNB N_B1_M1018_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.985
cc_33 VNB N_B1_M1022_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=0.56
cc_34 VNB N_B1_M1019_g 0.017456f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.985
cc_35 VNB N_B1_M1033_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=0.56
cc_36 VNB N_B1_M1028_g 0.017456f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.985
cc_37 VNB N_B1_M1039_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=0.56
cc_38 VNB N_B1_M1032_g 0.0177817f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.985
cc_39 VNB B1 0.00514993f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.105
cc_40 VNB N_B1_c_408_n 0.0651446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_C1_M1007_g 4.25129e-19 $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_42 VNB N_C1_M1002_g 0.0177817f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.985
cc_43 VNB N_C1_M1010_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=0.56
cc_44 VNB N_C1_M1029_g 0.017456f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.985
cc_45 VNB N_C1_M1023_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=0.56
cc_46 VNB N_C1_M1037_g 0.0174509f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.985
cc_47 VNB N_C1_M1034_g 4.54257e-19 $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=0.56
cc_48 VNB N_C1_M1038_g 0.0207559f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.985
cc_49 VNB N_C1_c_479_n 0.069841f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.185
cc_50 VNB N_VPWR_c_600_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB Y 0.0227487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_805_n 0.0112379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_908_n 0.0117482f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.985
cc_54 VNB N_VGND_c_909_n 0.0337587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_910_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_911_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_912_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.105
cc_58 VNB N_VGND_c_913_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_914_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.16
cc_60 VNB N_VGND_c_915_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.16
cc_61 VNB N_VGND_c_916_n 0.00543672f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.16
cc_62 VNB N_VGND_c_917_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=1.595 $Y2=1.16
cc_63 VNB N_VGND_c_918_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.16
cc_64 VNB N_VGND_c_919_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.185
cc_65 VNB N_VGND_c_920_n 0.00462871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_921_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_922_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.185
cc_68 VNB N_VGND_c_923_n 0.0117571f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=1.185
cc_69 VNB N_VGND_c_924_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_925_n 0.0942059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_926_n 0.449402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_927_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_928_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_929_n 0.00545721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_125_47#_c_1061_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.295
cc_76 VNB N_A_125_47#_c_1062_n 0.00705765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_125_47#_c_1063_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.185
cc_78 VNB N_A_125_47#_c_1064_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_125_47#_c_1065_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.185
cc_80 VNB N_A_125_47#_c_1066_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=1.185
cc_81 VNB N_A_125_47#_c_1067_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1163_47#_c_1167_n 0.00313199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1163_47#_c_1168_n 0.00162339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1163_47#_c_1169_n 0.0120148f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.985
cc_85 VPB N_A1_M1001_g 0.0271545f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.985
cc_86 VPB N_A1_M1009_g 0.0192043f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.985
cc_87 VPB N_A1_M1012_g 0.0192043f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.985
cc_88 VPB N_A1_M1027_g 0.0196044f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=1.985
cc_89 VPB A1 0.011511f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.105
cc_90 VPB N_A2_M1000_g 0.019782f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.985
cc_91 VPB N_A2_M1003_g 0.0194315f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.985
cc_92 VPB N_A2_M1005_g 0.0194315f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.985
cc_93 VPB N_A2_M1013_g 0.0273817f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=1.985
cc_94 VPB A2 0.0100369f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.105
cc_95 VPB N_A3_M1006_g 0.0273817f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=0.56
cc_96 VPB N_A3_M1014_g 0.0194315f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=0.56
cc_97 VPB N_A3_M1030_g 0.0194315f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=0.56
cc_98 VPB N_A3_M1036_g 0.0200232f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=1.985
cc_99 VPB A3 0.0189194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_B1_M1004_g 0.019796f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.56
cc_101 VPB N_B1_M1022_g 0.0192043f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=0.56
cc_102 VPB N_B1_M1033_g 0.0192043f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=0.56
cc_103 VPB N_B1_M1039_g 0.0195548f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=0.56
cc_104 VPB B1 0.00973f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.105
cc_105 VPB N_C1_M1007_g 0.0196044f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.56
cc_106 VPB N_C1_M1010_g 0.0192043f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=0.56
cc_107 VPB N_C1_M1023_g 0.0191997f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=0.56
cc_108 VPB N_C1_M1034_g 0.0227748f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=0.56
cc_109 VPB C1 0.00749287f $X=-0.19 $Y=1.305 $X2=1.045 $Y2=1.105
cc_110 VPB N_A_39_297#_c_537_n 0.0312108f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=0.56
cc_111 VPB N_A_39_297#_c_538_n 0.0137466f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.295
cc_112 VPB N_A_39_297#_c_539_n 0.00566527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_39_297#_c_540_n 0.00378316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_39_297#_c_541_n 0.00117749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_39_297#_c_542_n 0.00143675f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.16
cc_116 VPB N_A_39_297#_c_543_n 0.00117596f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.16
cc_117 VPB N_VPWR_c_601_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.295
cc_118 VPB N_VPWR_c_602_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.81 $Y2=1.025
cc_119 VPB N_VPWR_c_603_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.81 $Y2=1.295
cc_120 VPB N_VPWR_c_604_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.125 $Y2=1.105
cc_121 VPB N_VPWR_c_605_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_606_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.16
cc_123 VPB N_VPWR_c_607_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.16
cc_124 VPB N_VPWR_c_608_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.16
cc_125 VPB N_VPWR_c_609_n 0.0170261f $X=-0.19 $Y=1.305 $X2=1.255 $Y2=1.16
cc_126 VPB N_VPWR_c_610_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.595 $Y2=1.16
cc_127 VPB N_VPWR_c_611_n 0.102081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_612_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_613_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_614_n 0.0177474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_600_n 0.0484895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_616_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_617_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_618_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_619_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_620_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_461_297#_c_740_n 0.0109256f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.985
cc_138 VPB N_Y_c_806_n 0.00378316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_Y_c_807_n 0.00364602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_Y_c_808_n 0.00117596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_Y_c_809_n 0.00244254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_Y_c_810_n 0.00117749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_Y_c_811_n 0.00146492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_Y_c_812_n 0.00117749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB Y 0.0100409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB Y 0.0121046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_Y_c_815_n 0.0338711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 N_A1_M1025_g N_A2_M1020_g 0.0233716f $X=1.81 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A1_M1027_g N_A2_M1000_g 0.0233716f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_150 A1 A2 0.0229564f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A1_c_157_n A2 0.00243442f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A1_c_157_n N_A2_c_231_n 0.0233716f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A1_M1001_g N_A_39_297#_c_537_n 0.00791096f $X=0.55 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A1_M1001_g N_A_39_297#_c_545_n 0.0169795f $X=0.55 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A1_M1009_g N_A_39_297#_c_545_n 0.0156665f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_156 A1 N_A_39_297#_c_545_n 0.04366f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A1_c_157_n N_A_39_297#_c_545_n 9.33689e-19 $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_158 A1 N_A_39_297#_c_538_n 0.0274616f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A1_M1012_g N_A_39_297#_c_550_n 0.0156665f $X=1.39 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A1_M1027_g N_A_39_297#_c_550_n 0.0171535f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_161 A1 N_A_39_297#_c_550_n 0.0324797f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A1_c_157_n N_A_39_297#_c_550_n 6.177e-19 $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_163 A1 N_A_39_297#_c_541_n 0.013857f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A1_c_157_n N_A_39_297#_c_541_n 6.77113e-19 $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A1_M1001_g N_VPWR_c_601_n 0.0126048f $X=0.55 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A1_M1009_g N_VPWR_c_601_n 0.0104025f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_M1012_g N_VPWR_c_601_n 6.54417e-19 $X=1.39 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A1_M1009_g N_VPWR_c_602_n 6.54417e-19 $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A1_M1012_g N_VPWR_c_602_n 0.0104025f $X=1.39 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A1_M1027_g N_VPWR_c_602_n 0.0116083f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A1_M1001_g N_VPWR_c_609_n 0.0046653f $X=0.55 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A1_M1009_g N_VPWR_c_610_n 0.0046653f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A1_M1012_g N_VPWR_c_610_n 0.0046653f $X=1.39 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A1_M1027_g N_VPWR_c_611_n 0.0046653f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A1_M1001_g N_VPWR_c_600_n 0.00902958f $X=0.55 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A1_M1009_g N_VPWR_c_600_n 0.00796766f $X=0.97 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A1_M1012_g N_VPWR_c_600_n 0.00796766f $X=1.39 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A1_M1027_g N_VPWR_c_600_n 0.00799591f $X=1.81 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A1_M1011_g N_VGND_c_909_n 0.0122699f $X=0.55 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A1_M1015_g N_VGND_c_909_n 7.34721e-19 $X=0.97 $Y=0.56 $X2=0 $Y2=0
cc_181 A1 N_VGND_c_909_n 0.0327559f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A1_c_157_n N_VGND_c_909_n 0.00132469f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A1_M1011_g N_VGND_c_910_n 5.54209e-19 $X=0.55 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A1_M1015_g N_VGND_c_910_n 0.00685342f $X=0.97 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A1_M1024_g N_VGND_c_910_n 0.00685342f $X=1.39 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A1_M1025_g N_VGND_c_910_n 5.54209e-19 $X=1.81 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A1_M1024_g N_VGND_c_911_n 5.54209e-19 $X=1.39 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A1_M1025_g N_VGND_c_911_n 0.00681952f $X=1.81 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A1_M1011_g N_VGND_c_923_n 0.0046653f $X=0.55 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A1_M1015_g N_VGND_c_923_n 0.00341689f $X=0.97 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A1_M1024_g N_VGND_c_924_n 0.00341689f $X=1.39 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A1_M1025_g N_VGND_c_924_n 0.00341689f $X=1.81 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A1_M1011_g N_VGND_c_926_n 0.00796766f $X=0.55 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A1_M1015_g N_VGND_c_926_n 0.0040262f $X=0.97 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A1_M1024_g N_VGND_c_926_n 0.0040262f $X=1.39 $Y=0.56 $X2=0 $Y2=0
cc_196 N_A1_M1025_g N_VGND_c_926_n 0.0040262f $X=1.81 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A1_M1015_g N_A_125_47#_c_1068_n 0.0122458f $X=0.97 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A1_M1024_g N_A_125_47#_c_1068_n 0.0125517f $X=1.39 $Y=0.56 $X2=0 $Y2=0
cc_199 A1 N_A_125_47#_c_1068_n 0.0408166f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_200 N_A1_c_157_n N_A_125_47#_c_1068_n 0.00202123f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_201 A1 N_A_125_47#_c_1061_n 0.0131017f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A1_c_157_n N_A_125_47#_c_1061_n 0.00208088f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A1_M1025_g N_A_125_47#_c_1074_n 0.0140707f $X=1.81 $Y=0.56 $X2=0 $Y2=0
cc_204 A1 N_A_125_47#_c_1074_n 0.00467597f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_205 A1 N_A_125_47#_c_1063_n 0.0131017f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_206 N_A1_c_157_n N_A_125_47#_c_1063_n 0.00208088f $X=1.81 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A2_M1035_g N_A3_M1008_g 0.0193797f $X=3.49 $Y=0.56 $X2=0 $Y2=0
cc_208 A2 A3 0.0223265f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_209 N_A2_c_231_n A3 0.00100704f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_210 A2 N_A3_c_318_n 8.78793e-19 $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_211 N_A2_c_231_n N_A3_c_318_n 0.0193797f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_M1000_g N_A_39_297#_c_556_n 0.0156313f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A2_M1003_g N_A_39_297#_c_556_n 0.0133553f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_214 A2 N_A_39_297#_c_556_n 0.0423979f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_215 N_A2_c_231_n N_A_39_297#_c_556_n 6.177e-19 $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_M1005_g N_A_39_297#_c_539_n 0.0133553f $X=3.07 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A2_M1013_g N_A_39_297#_c_539_n 0.0145015f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_218 A2 N_A_39_297#_c_539_n 0.0423979f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_219 N_A2_c_231_n N_A_39_297#_c_539_n 6.177e-19 $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_220 A2 N_A_39_297#_c_542_n 0.0133192f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_221 A2 N_A_39_297#_c_543_n 0.0137781f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A2_c_231_n N_A_39_297#_c_543_n 6.69205e-19 $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A2_M1000_g N_VPWR_c_602_n 0.00130728f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A2_M1000_g N_VPWR_c_611_n 0.00539841f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A2_M1003_g N_VPWR_c_611_n 0.00357835f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A2_M1005_g N_VPWR_c_611_n 0.00357835f $X=3.07 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A2_M1013_g N_VPWR_c_611_n 0.00357835f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A2_M1000_g N_VPWR_c_600_n 0.00969144f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A2_M1003_g N_VPWR_c_600_n 0.00522513f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A2_M1005_g N_VPWR_c_600_n 0.00522513f $X=3.07 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A2_M1013_g N_VPWR_c_600_n 0.0066022f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A2_M1000_g N_A_461_297#_c_741_n 0.0045641f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A2_M1003_g N_A_461_297#_c_741_n 0.00581235f $X=2.65 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A2_M1005_g N_A_461_297#_c_741_n 5.92384e-19 $X=3.07 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A2_M1003_g N_A_461_297#_c_744_n 0.00801314f $X=2.65 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A2_M1005_g N_A_461_297#_c_744_n 0.00801314f $X=3.07 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A2_M1000_g N_A_461_297#_c_746_n 0.00202057f $X=2.23 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A2_M1003_g N_A_461_297#_c_746_n 7.04098e-19 $X=2.65 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A2_M1003_g N_A_461_297#_c_748_n 5.92384e-19 $X=2.65 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A2_M1005_g N_A_461_297#_c_748_n 0.00581235f $X=3.07 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A2_M1013_g N_A_461_297#_c_748_n 0.0106522f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A2_M1013_g N_A_461_297#_c_740_n 0.0101161f $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A2_M1005_g N_A_461_297#_c_752_n 7.04098e-19 $X=3.07 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_A2_M1013_g N_A_461_297#_c_752_n 7.04098e-19 $X=3.49 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_A2_M1013_g N_Y_c_807_n 7.60605e-19 $X=3.49 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A2_M1020_g N_VGND_c_911_n 0.00681952f $X=2.23 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A2_M1021_g N_VGND_c_911_n 5.54209e-19 $X=2.65 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A2_M1020_g N_VGND_c_912_n 5.54209e-19 $X=2.23 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A2_M1021_g N_VGND_c_912_n 0.00685342f $X=2.65 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A2_M1026_g N_VGND_c_912_n 0.00685342f $X=3.07 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A2_M1035_g N_VGND_c_912_n 5.54209e-19 $X=3.49 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A2_M1026_g N_VGND_c_913_n 5.5541e-19 $X=3.07 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A2_M1035_g N_VGND_c_913_n 0.00691054f $X=3.49 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A2_M1020_g N_VGND_c_917_n 0.00341689f $X=2.23 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A2_M1021_g N_VGND_c_917_n 0.00341689f $X=2.65 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A2_M1026_g N_VGND_c_919_n 0.00341689f $X=3.07 $Y=0.56 $X2=0 $Y2=0
cc_257 N_A2_M1035_g N_VGND_c_919_n 0.00341689f $X=3.49 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A2_M1020_g N_VGND_c_926_n 0.0040262f $X=2.23 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A2_M1021_g N_VGND_c_926_n 0.0040262f $X=2.65 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A2_M1026_g N_VGND_c_926_n 0.0040262f $X=3.07 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A2_M1035_g N_VGND_c_926_n 0.0040262f $X=3.49 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A2_M1020_g N_A_125_47#_c_1074_n 0.0125517f $X=2.23 $Y=0.56 $X2=0 $Y2=0
cc_263 A2 N_A_125_47#_c_1074_n 0.0268079f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_264 N_A2_M1021_g N_A_125_47#_c_1080_n 0.0126116f $X=2.65 $Y=0.56 $X2=0 $Y2=0
cc_265 N_A2_M1026_g N_A_125_47#_c_1080_n 0.0126116f $X=3.07 $Y=0.56 $X2=0 $Y2=0
cc_266 A2 N_A_125_47#_c_1080_n 0.0408166f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_267 N_A2_c_231_n N_A_125_47#_c_1080_n 0.00202123f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A2_M1035_g N_A_125_47#_c_1084_n 0.0127126f $X=3.49 $Y=0.56 $X2=0 $Y2=0
cc_269 A2 N_A_125_47#_c_1084_n 0.0145686f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_270 A2 N_A_125_47#_c_1064_n 0.0131017f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_271 N_A2_c_231_n N_A_125_47#_c_1064_n 0.00208088f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_272 A2 N_A_125_47#_c_1065_n 0.0131017f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_273 N_A2_c_231_n N_A_125_47#_c_1065_n 0.00208088f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A3_M1036_g N_B1_M1004_g 0.0192069f $X=5.69 $Y=1.985 $X2=0 $Y2=0
cc_275 A3 B1 0.0229595f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_276 N_A3_c_318_n B1 2.61683e-19 $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_277 A3 N_B1_c_408_n 0.00103382f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_278 N_A3_c_318_n N_B1_c_408_n 0.0192069f $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A3_M1006_g N_A_39_297#_c_539_n 7.60605e-19 $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_280 A3 N_A_39_297#_c_539_n 0.0051523f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_281 N_A3_M1036_g N_VPWR_c_603_n 0.00127003f $X=5.69 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A3_M1006_g N_VPWR_c_611_n 0.00357835f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A3_M1014_g N_VPWR_c_611_n 0.00357835f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A3_M1030_g N_VPWR_c_611_n 0.00357835f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A3_M1036_g N_VPWR_c_611_n 0.00539841f $X=5.69 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A3_M1006_g N_VPWR_c_600_n 0.0066022f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A3_M1014_g N_VPWR_c_600_n 0.00522513f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A3_M1030_g N_VPWR_c_600_n 0.00522513f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A3_M1036_g N_VPWR_c_600_n 0.00974189f $X=5.69 $Y=1.985 $X2=0 $Y2=0
cc_290 N_A3_M1006_g N_A_461_297#_c_740_n 0.0101161f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A3_M1006_g N_A_461_297#_c_755_n 0.0106522f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A3_M1014_g N_A_461_297#_c_755_n 0.00581235f $X=4.85 $Y=1.985 $X2=0
+ $Y2=0
cc_293 N_A3_M1030_g N_A_461_297#_c_755_n 5.92384e-19 $X=5.27 $Y=1.985 $X2=0
+ $Y2=0
cc_294 N_A3_M1014_g N_A_461_297#_c_758_n 0.00801314f $X=4.85 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A3_M1030_g N_A_461_297#_c_758_n 0.00871724f $X=5.27 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A3_M1036_g N_A_461_297#_c_758_n 0.00202643f $X=5.69 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_A3_M1014_g N_A_461_297#_c_761_n 5.92384e-19 $X=4.85 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A3_M1030_g N_A_461_297#_c_761_n 0.00581235f $X=5.27 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A3_M1036_g N_A_461_297#_c_761_n 0.00457792f $X=5.69 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A3_M1006_g N_A_461_297#_c_764_n 7.04098e-19 $X=4.43 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A3_M1014_g N_A_461_297#_c_764_n 7.04098e-19 $X=4.85 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A3_M1006_g N_Y_c_817_n 0.0145015f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A3_M1014_g N_Y_c_817_n 0.0133553f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_304 A3 N_Y_c_817_n 0.0423979f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_305 N_A3_c_318_n N_Y_c_817_n 6.08811e-19 $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_306 A3 N_Y_c_807_n 0.0209344f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_307 N_A3_c_318_n N_Y_c_807_n 0.00182127f $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A3_M1030_g N_Y_c_823_n 0.0133553f $X=5.27 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A3_M1036_g N_Y_c_823_n 0.0157258f $X=5.69 $Y=1.985 $X2=0 $Y2=0
cc_310 A3 N_Y_c_823_n 0.0423979f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_311 N_A3_c_318_n N_Y_c_823_n 6.177e-19 $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_312 A3 N_Y_c_808_n 0.0137781f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_313 N_A3_c_318_n N_Y_c_808_n 6.60288e-19 $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_314 A3 N_Y_c_809_n 0.00565044f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_315 N_A3_M1008_g N_VGND_c_913_n 0.00691054f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A3_M1016_g N_VGND_c_913_n 5.5541e-19 $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A3_M1008_g N_VGND_c_914_n 5.54209e-19 $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_318 N_A3_M1016_g N_VGND_c_914_n 0.00685342f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_319 N_A3_M1017_g N_VGND_c_914_n 0.00685342f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_320 N_A3_M1031_g N_VGND_c_914_n 5.54209e-19 $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_321 N_A3_M1017_g N_VGND_c_915_n 0.00341689f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_322 N_A3_M1031_g N_VGND_c_915_n 0.00341689f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_323 N_A3_M1017_g N_VGND_c_916_n 5.5541e-19 $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_324 N_A3_M1031_g N_VGND_c_916_n 0.00799399f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A3_M1008_g N_VGND_c_921_n 0.00341689f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_326 N_A3_M1016_g N_VGND_c_921_n 0.00341689f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_327 N_A3_M1008_g N_VGND_c_926_n 0.0040262f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_328 N_A3_M1016_g N_VGND_c_926_n 0.0040262f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_329 N_A3_M1017_g N_VGND_c_926_n 0.0040262f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_330 N_A3_M1031_g N_VGND_c_926_n 0.0040262f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_331 N_A3_M1008_g N_A_125_47#_c_1084_n 0.0127126f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_332 A3 N_A_125_47#_c_1084_n 0.0145686f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_333 N_A3_M1016_g N_A_125_47#_c_1092_n 0.0126116f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_334 N_A3_M1017_g N_A_125_47#_c_1092_n 0.0126116f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_335 A3 N_A_125_47#_c_1092_n 0.0408166f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_336 N_A3_c_318_n N_A_125_47#_c_1092_n 0.00242163f $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A3_M1031_g N_A_125_47#_c_1062_n 0.0154657f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_338 A3 N_A_125_47#_c_1062_n 0.0572401f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_339 N_A3_c_318_n N_A_125_47#_c_1062_n 0.0131387f $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_340 A3 N_A_125_47#_c_1066_n 0.0131017f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_341 N_A3_c_318_n N_A_125_47#_c_1066_n 0.00208088f $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_342 A3 N_A_125_47#_c_1067_n 0.0131017f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_343 N_A3_c_318_n N_A_125_47#_c_1067_n 0.00248172f $X=5.69 $Y=1.16 $X2=0 $Y2=0
cc_344 N_B1_M1039_g N_C1_M1007_g 0.0280326f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_345 N_B1_M1032_g N_C1_M1002_g 0.0141063f $X=7.43 $Y=0.56 $X2=0 $Y2=0
cc_346 B1 C1 0.0229561f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_347 B1 N_C1_c_479_n 0.00234696f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_348 N_B1_c_408_n N_C1_c_479_n 0.0163259f $X=7.43 $Y=1.16 $X2=0 $Y2=0
cc_349 N_B1_M1004_g N_VPWR_c_603_n 0.0116323f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_350 N_B1_M1022_g N_VPWR_c_603_n 0.0104025f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_351 N_B1_M1033_g N_VPWR_c_603_n 6.54417e-19 $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_352 N_B1_M1022_g N_VPWR_c_604_n 6.54417e-19 $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_353 N_B1_M1033_g N_VPWR_c_604_n 0.0104025f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_354 N_B1_M1039_g N_VPWR_c_604_n 0.0104025f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_355 N_B1_M1039_g N_VPWR_c_605_n 6.54417e-19 $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_356 N_B1_M1004_g N_VPWR_c_611_n 0.0046653f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_357 N_B1_M1022_g N_VPWR_c_612_n 0.0046653f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_358 N_B1_M1033_g N_VPWR_c_612_n 0.0046653f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_359 N_B1_M1039_g N_VPWR_c_613_n 0.0046653f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_360 N_B1_M1004_g N_VPWR_c_600_n 0.00804636f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_361 N_B1_M1022_g N_VPWR_c_600_n 0.00796766f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_362 N_B1_M1033_g N_VPWR_c_600_n 0.00796766f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_363 N_B1_M1039_g N_VPWR_c_600_n 0.00799591f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_364 N_B1_M1004_g N_Y_c_830_n 0.0157258f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_365 N_B1_M1022_g N_Y_c_830_n 0.0156665f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_366 B1 N_Y_c_830_n 0.0403899f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_367 N_B1_c_408_n N_Y_c_830_n 6.13255e-19 $X=7.43 $Y=1.16 $X2=0 $Y2=0
cc_368 N_B1_M1033_g N_Y_c_834_n 0.0156665f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_369 N_B1_M1039_g N_Y_c_834_n 0.0156313f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_370 B1 N_Y_c_834_n 0.0423979f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_371 N_B1_c_408_n N_Y_c_834_n 6.13255e-19 $X=7.43 $Y=1.16 $X2=0 $Y2=0
cc_372 B1 N_Y_c_810_n 0.013857f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_373 N_B1_c_408_n N_Y_c_810_n 6.72654e-19 $X=7.43 $Y=1.16 $X2=0 $Y2=0
cc_374 B1 N_Y_c_811_n 0.0138571f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_375 N_B1_M1018_g N_VGND_c_916_n 0.00229695f $X=6.17 $Y=0.56 $X2=0 $Y2=0
cc_376 N_B1_M1018_g N_VGND_c_925_n 0.00357877f $X=6.17 $Y=0.56 $X2=0 $Y2=0
cc_377 N_B1_M1019_g N_VGND_c_925_n 0.00357877f $X=6.59 $Y=0.56 $X2=0 $Y2=0
cc_378 N_B1_M1028_g N_VGND_c_925_n 0.00357877f $X=7.01 $Y=0.56 $X2=0 $Y2=0
cc_379 N_B1_M1032_g N_VGND_c_925_n 0.00357877f $X=7.43 $Y=0.56 $X2=0 $Y2=0
cc_380 N_B1_M1018_g N_VGND_c_926_n 0.00655123f $X=6.17 $Y=0.56 $X2=0 $Y2=0
cc_381 N_B1_M1019_g N_VGND_c_926_n 0.00522516f $X=6.59 $Y=0.56 $X2=0 $Y2=0
cc_382 N_B1_M1028_g N_VGND_c_926_n 0.00522516f $X=7.01 $Y=0.56 $X2=0 $Y2=0
cc_383 N_B1_M1032_g N_VGND_c_926_n 0.00525237f $X=7.43 $Y=0.56 $X2=0 $Y2=0
cc_384 N_B1_M1018_g N_A_125_47#_c_1062_n 0.0128039f $X=6.17 $Y=0.56 $X2=0 $Y2=0
cc_385 N_B1_M1019_g N_A_125_47#_c_1062_n 0.00994985f $X=6.59 $Y=0.56 $X2=0 $Y2=0
cc_386 N_B1_M1028_g N_A_125_47#_c_1062_n 0.00994985f $X=7.01 $Y=0.56 $X2=0 $Y2=0
cc_387 N_B1_M1032_g N_A_125_47#_c_1062_n 0.00318865f $X=7.43 $Y=0.56 $X2=0 $Y2=0
cc_388 B1 N_A_125_47#_c_1062_n 0.0827969f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_389 N_B1_c_408_n N_A_125_47#_c_1062_n 0.00666428f $X=7.43 $Y=1.16 $X2=0 $Y2=0
cc_390 N_B1_M1018_g N_A_1163_47#_c_1167_n 0.00918728f $X=6.17 $Y=0.56 $X2=0
+ $Y2=0
cc_391 N_B1_M1019_g N_A_1163_47#_c_1167_n 0.00918728f $X=6.59 $Y=0.56 $X2=0
+ $Y2=0
cc_392 N_B1_M1028_g N_A_1163_47#_c_1167_n 0.00918728f $X=7.01 $Y=0.56 $X2=0
+ $Y2=0
cc_393 N_B1_M1032_g N_A_1163_47#_c_1167_n 0.0107429f $X=7.43 $Y=0.56 $X2=0 $Y2=0
cc_394 B1 N_A_1163_47#_c_1167_n 0.00403046f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_395 B1 N_A_1163_47#_c_1168_n 0.0115075f $X=7.525 $Y=1.105 $X2=0 $Y2=0
cc_396 N_C1_M1007_g N_VPWR_c_604_n 6.54417e-19 $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_397 N_C1_M1007_g N_VPWR_c_605_n 0.0104025f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_398 N_C1_M1010_g N_VPWR_c_605_n 0.0104025f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_399 N_C1_M1023_g N_VPWR_c_605_n 6.54417e-19 $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_400 N_C1_M1010_g N_VPWR_c_606_n 6.54417e-19 $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_401 N_C1_M1023_g N_VPWR_c_606_n 0.0104025f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_402 N_C1_M1034_g N_VPWR_c_606_n 0.0123094f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_403 N_C1_M1010_g N_VPWR_c_607_n 0.0046653f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_404 N_C1_M1023_g N_VPWR_c_607_n 0.0046653f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_405 N_C1_M1007_g N_VPWR_c_613_n 0.0046653f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_406 N_C1_M1034_g N_VPWR_c_614_n 0.0046653f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_407 N_C1_M1007_g N_VPWR_c_600_n 0.00799591f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_408 N_C1_M1010_g N_VPWR_c_600_n 0.00796766f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_409 N_C1_M1023_g N_VPWR_c_600_n 0.00796766f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_410 N_C1_M1034_g N_VPWR_c_600_n 0.00905913f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_411 N_C1_M1007_g N_Y_c_841_n 0.0196916f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_412 N_C1_M1010_g N_Y_c_841_n 0.0156665f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_413 C1 N_Y_c_841_n 0.0310415f $X=8.905 $Y=1.105 $X2=0 $Y2=0
cc_414 N_C1_c_479_n N_Y_c_841_n 6.13255e-19 $X=9.11 $Y=1.16 $X2=0 $Y2=0
cc_415 N_C1_M1002_g N_Y_c_845_n 0.00318865f $X=7.85 $Y=0.56 $X2=0 $Y2=0
cc_416 N_C1_M1029_g N_Y_c_845_n 0.00994985f $X=8.27 $Y=0.56 $X2=0 $Y2=0
cc_417 N_C1_M1037_g N_Y_c_845_n 0.00994985f $X=8.69 $Y=0.56 $X2=0 $Y2=0
cc_418 N_C1_M1038_g N_Y_c_845_n 0.0132827f $X=9.11 $Y=0.56 $X2=0 $Y2=0
cc_419 C1 N_Y_c_845_n 0.0745403f $X=8.905 $Y=1.105 $X2=0 $Y2=0
cc_420 N_C1_c_479_n N_Y_c_845_n 0.00666428f $X=9.11 $Y=1.16 $X2=0 $Y2=0
cc_421 N_C1_M1023_g N_Y_c_851_n 0.0156665f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_422 N_C1_M1034_g N_Y_c_851_n 0.0177461f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_423 C1 N_Y_c_851_n 0.0364348f $X=8.905 $Y=1.105 $X2=0 $Y2=0
cc_424 N_C1_c_479_n N_Y_c_851_n 6.13255e-19 $X=9.11 $Y=1.16 $X2=0 $Y2=0
cc_425 C1 N_Y_c_812_n 0.013857f $X=8.905 $Y=1.105 $X2=0 $Y2=0
cc_426 N_C1_c_479_n N_Y_c_812_n 6.72654e-19 $X=9.11 $Y=1.16 $X2=0 $Y2=0
cc_427 N_C1_M1034_g Y 0.00704969f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_428 N_C1_M1038_g Y 0.0143382f $X=9.11 $Y=0.56 $X2=0 $Y2=0
cc_429 C1 Y 0.02153f $X=8.905 $Y=1.105 $X2=0 $Y2=0
cc_430 N_C1_M1002_g N_VGND_c_925_n 0.00357877f $X=7.85 $Y=0.56 $X2=0 $Y2=0
cc_431 N_C1_M1029_g N_VGND_c_925_n 0.00357877f $X=8.27 $Y=0.56 $X2=0 $Y2=0
cc_432 N_C1_M1037_g N_VGND_c_925_n 0.00357877f $X=8.69 $Y=0.56 $X2=0 $Y2=0
cc_433 N_C1_M1038_g N_VGND_c_925_n 0.00357877f $X=9.11 $Y=0.56 $X2=0 $Y2=0
cc_434 N_C1_M1002_g N_VGND_c_926_n 0.00525237f $X=7.85 $Y=0.56 $X2=0 $Y2=0
cc_435 N_C1_M1029_g N_VGND_c_926_n 0.00522516f $X=8.27 $Y=0.56 $X2=0 $Y2=0
cc_436 N_C1_M1037_g N_VGND_c_926_n 0.00522516f $X=8.69 $Y=0.56 $X2=0 $Y2=0
cc_437 N_C1_M1038_g N_VGND_c_926_n 0.00624775f $X=9.11 $Y=0.56 $X2=0 $Y2=0
cc_438 N_C1_M1002_g N_A_1163_47#_c_1169_n 0.0124217f $X=7.85 $Y=0.56 $X2=0 $Y2=0
cc_439 N_C1_M1029_g N_A_1163_47#_c_1169_n 0.00918728f $X=8.27 $Y=0.56 $X2=0
+ $Y2=0
cc_440 N_C1_M1037_g N_A_1163_47#_c_1169_n 0.00918728f $X=8.69 $Y=0.56 $X2=0
+ $Y2=0
cc_441 N_C1_M1038_g N_A_1163_47#_c_1169_n 0.00918728f $X=9.11 $Y=0.56 $X2=0
+ $Y2=0
cc_442 C1 N_A_1163_47#_c_1169_n 7.94104e-19 $X=8.905 $Y=1.105 $X2=0 $Y2=0
cc_443 N_A_39_297#_c_545_n N_VPWR_M1001_d 0.00315342f $X=1.095 $Y=1.605
+ $X2=-0.19 $Y2=1.305
cc_444 N_A_39_297#_c_550_n N_VPWR_M1012_d 0.00315342f $X=1.935 $Y=1.605 $X2=0
+ $Y2=0
cc_445 N_A_39_297#_c_537_n N_VPWR_c_601_n 0.0405143f $X=0.32 $Y=1.815 $X2=0
+ $Y2=0
cc_446 N_A_39_297#_c_545_n N_VPWR_c_601_n 0.017435f $X=1.095 $Y=1.605 $X2=0
+ $Y2=0
cc_447 N_A_39_297#_c_550_n N_VPWR_c_602_n 0.017435f $X=1.935 $Y=1.605 $X2=0
+ $Y2=0
cc_448 N_A_39_297#_c_537_n N_VPWR_c_609_n 0.0225118f $X=0.32 $Y=1.815 $X2=0
+ $Y2=0
cc_449 N_A_39_297#_c_575_p N_VPWR_c_610_n 0.0113958f $X=1.18 $Y=1.815 $X2=0
+ $Y2=0
cc_450 N_A_39_297#_c_576_p N_VPWR_c_611_n 0.0113958f $X=2.02 $Y=1.815 $X2=0
+ $Y2=0
cc_451 N_A_39_297#_M1001_s N_VPWR_c_600_n 0.00472999f $X=0.195 $Y=1.485 $X2=0
+ $Y2=0
cc_452 N_A_39_297#_M1009_s N_VPWR_c_600_n 0.00570907f $X=1.045 $Y=1.485 $X2=0
+ $Y2=0
cc_453 N_A_39_297#_M1027_s N_VPWR_c_600_n 0.00570907f $X=1.885 $Y=1.485 $X2=0
+ $Y2=0
cc_454 N_A_39_297#_M1003_d N_VPWR_c_600_n 0.00216833f $X=2.725 $Y=1.485 $X2=0
+ $Y2=0
cc_455 N_A_39_297#_M1013_d N_VPWR_c_600_n 0.00210147f $X=3.565 $Y=1.485 $X2=0
+ $Y2=0
cc_456 N_A_39_297#_c_537_n N_VPWR_c_600_n 0.0122467f $X=0.32 $Y=1.815 $X2=0
+ $Y2=0
cc_457 N_A_39_297#_c_575_p N_VPWR_c_600_n 0.00646998f $X=1.18 $Y=1.815 $X2=0
+ $Y2=0
cc_458 N_A_39_297#_c_576_p N_VPWR_c_600_n 0.00646998f $X=2.02 $Y=1.815 $X2=0
+ $Y2=0
cc_459 N_A_39_297#_c_556_n N_A_461_297#_M1000_s 0.00315342f $X=2.775 $Y=1.605
+ $X2=-0.19 $Y2=1.305
cc_460 N_A_39_297#_c_539_n N_A_461_297#_M1005_s 0.00315342f $X=3.615 $Y=1.605
+ $X2=0 $Y2=0
cc_461 N_A_39_297#_c_556_n N_A_461_297#_c_741_n 0.0171917f $X=2.775 $Y=1.605
+ $X2=0 $Y2=0
cc_462 N_A_39_297#_M1003_d N_A_461_297#_c_744_n 0.00316374f $X=2.725 $Y=1.485
+ $X2=0 $Y2=0
cc_463 N_A_39_297#_c_556_n N_A_461_297#_c_744_n 0.0030597f $X=2.775 $Y=1.605
+ $X2=0 $Y2=0
cc_464 N_A_39_297#_c_590_p N_A_461_297#_c_744_n 0.0112509f $X=2.86 $Y=1.725
+ $X2=0 $Y2=0
cc_465 N_A_39_297#_c_539_n N_A_461_297#_c_744_n 0.0030597f $X=3.615 $Y=1.605
+ $X2=0 $Y2=0
cc_466 N_A_39_297#_c_539_n N_A_461_297#_c_748_n 0.0171917f $X=3.615 $Y=1.605
+ $X2=0 $Y2=0
cc_467 N_A_39_297#_M1013_d N_A_461_297#_c_740_n 0.00486083f $X=3.565 $Y=1.485
+ $X2=0 $Y2=0
cc_468 N_A_39_297#_c_539_n N_A_461_297#_c_740_n 0.0030597f $X=3.615 $Y=1.605
+ $X2=0 $Y2=0
cc_469 N_A_39_297#_c_540_n N_A_461_297#_c_740_n 0.0175665f $X=3.74 $Y=1.725
+ $X2=0 $Y2=0
cc_470 N_A_39_297#_c_540_n N_Y_c_806_n 0.0287208f $X=3.74 $Y=1.725 $X2=0 $Y2=0
cc_471 N_A_39_297#_c_539_n N_Y_c_807_n 0.0207751f $X=3.615 $Y=1.605 $X2=0 $Y2=0
cc_472 N_A_39_297#_c_550_n N_A_125_47#_c_1074_n 0.00276135f $X=1.935 $Y=1.605
+ $X2=0 $Y2=0
cc_473 N_A_39_297#_c_539_n N_A_125_47#_c_1084_n 0.00576301f $X=3.615 $Y=1.605
+ $X2=0 $Y2=0
cc_474 N_VPWR_c_600_n N_A_461_297#_M1000_s 0.00215201f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_475 N_VPWR_c_600_n N_A_461_297#_M1005_s 0.00215201f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_600_n N_A_461_297#_M1006_s 0.00215201f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_600_n N_A_461_297#_M1030_s 0.00215201f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_611_n N_A_461_297#_c_744_n 0.0286211f $X=6.175 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_600_n N_A_461_297#_c_744_n 0.0178969f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_611_n N_A_461_297#_c_746_n 0.0188514f $X=6.175 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_600_n N_A_461_297#_c_746_n 0.0122326f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_611_n N_A_461_297#_c_740_n 0.0618643f $X=6.175 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_600_n N_A_461_297#_c_740_n 0.0372646f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_611_n N_A_461_297#_c_758_n 0.0474725f $X=6.175 $Y=2.72 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_600_n N_A_461_297#_c_758_n 0.0301295f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_611_n N_A_461_297#_c_752_n 0.0188514f $X=6.175 $Y=2.72 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_600_n N_A_461_297#_c_752_n 0.0122326f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_611_n N_A_461_297#_c_764_n 0.0188514f $X=6.175 $Y=2.72 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_600_n N_A_461_297#_c_764_n 0.0122326f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_600_n N_Y_M1006_d 0.00210147f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_491 N_VPWR_c_600_n N_Y_M1014_d 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_492 N_VPWR_c_600_n N_Y_M1036_d 0.00586967f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_493 N_VPWR_c_600_n N_Y_M1022_d 0.00570907f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_494 N_VPWR_c_600_n N_Y_M1039_d 0.00570907f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_c_600_n N_Y_M1010_s 0.00570907f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_496 N_VPWR_c_600_n N_Y_M1034_s 0.00387172f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_497 N_VPWR_c_611_n N_Y_c_869_n 0.0128022f $X=6.175 $Y=2.72 $X2=0 $Y2=0
cc_498 N_VPWR_c_600_n N_Y_c_869_n 0.00724021f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_499 N_VPWR_M1004_s N_Y_c_830_n 0.00315342f $X=6.205 $Y=1.485 $X2=0 $Y2=0
cc_500 N_VPWR_c_603_n N_Y_c_830_n 0.017435f $X=6.34 $Y=2.02 $X2=0 $Y2=0
cc_501 N_VPWR_c_612_n N_Y_c_873_n 0.0113958f $X=7.015 $Y=2.72 $X2=0 $Y2=0
cc_502 N_VPWR_c_600_n N_Y_c_873_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_503 N_VPWR_M1033_s N_Y_c_834_n 0.00315342f $X=7.045 $Y=1.485 $X2=0 $Y2=0
cc_504 N_VPWR_c_604_n N_Y_c_834_n 0.017435f $X=7.18 $Y=2.02 $X2=0 $Y2=0
cc_505 N_VPWR_c_613_n N_Y_c_877_n 0.0113958f $X=7.855 $Y=2.72 $X2=0 $Y2=0
cc_506 N_VPWR_c_600_n N_Y_c_877_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_507 N_VPWR_M1007_d N_Y_c_841_n 0.00315342f $X=7.885 $Y=1.485 $X2=0 $Y2=0
cc_508 N_VPWR_c_605_n N_Y_c_841_n 0.017435f $X=8.02 $Y=2.02 $X2=0 $Y2=0
cc_509 N_VPWR_c_607_n N_Y_c_881_n 0.0113958f $X=8.695 $Y=2.72 $X2=0 $Y2=0
cc_510 N_VPWR_c_600_n N_Y_c_881_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_511 N_VPWR_M1023_d N_Y_c_851_n 0.00315342f $X=8.725 $Y=1.485 $X2=0 $Y2=0
cc_512 N_VPWR_c_606_n N_Y_c_851_n 0.017435f $X=8.86 $Y=2.02 $X2=0 $Y2=0
cc_513 N_VPWR_c_614_n N_Y_c_815_n 0.0266045f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_514 N_VPWR_c_600_n N_Y_c_815_n 0.0145574f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_515 N_A_461_297#_c_740_n N_Y_M1006_d 0.00486083f $X=4.475 $Y=2.38 $X2=0 $Y2=0
cc_516 N_A_461_297#_c_758_n N_Y_M1014_d 0.00316374f $X=5.315 $Y=2.38 $X2=0 $Y2=0
cc_517 N_A_461_297#_c_740_n N_Y_c_806_n 0.0175665f $X=4.475 $Y=2.38 $X2=0 $Y2=0
cc_518 N_A_461_297#_M1006_s N_Y_c_817_n 0.00315342f $X=4.505 $Y=1.485 $X2=0
+ $Y2=0
cc_519 N_A_461_297#_c_740_n N_Y_c_817_n 0.0030597f $X=4.475 $Y=2.38 $X2=0 $Y2=0
cc_520 N_A_461_297#_c_755_n N_Y_c_817_n 0.0171917f $X=4.64 $Y=2.02 $X2=0 $Y2=0
cc_521 N_A_461_297#_c_758_n N_Y_c_817_n 0.0030597f $X=5.315 $Y=2.38 $X2=0 $Y2=0
cc_522 N_A_461_297#_c_758_n N_Y_c_894_n 0.0112509f $X=5.315 $Y=2.38 $X2=0 $Y2=0
cc_523 N_A_461_297#_M1030_s N_Y_c_823_n 0.00315342f $X=5.345 $Y=1.485 $X2=0
+ $Y2=0
cc_524 N_A_461_297#_c_758_n N_Y_c_823_n 0.0030597f $X=5.315 $Y=2.38 $X2=0 $Y2=0
cc_525 N_A_461_297#_c_761_n N_Y_c_823_n 0.0171917f $X=5.48 $Y=2.02 $X2=0 $Y2=0
cc_526 N_Y_M1002_s N_VGND_c_926_n 0.00216833f $X=7.925 $Y=0.235 $X2=0 $Y2=0
cc_527 N_Y_M1037_s N_VGND_c_926_n 0.00216833f $X=8.765 $Y=0.235 $X2=0 $Y2=0
cc_528 N_Y_c_809_n N_A_125_47#_c_1062_n 0.0037486f $X=5.91 $Y=1.605 $X2=0 $Y2=0
cc_529 N_Y_c_845_n N_A_1163_47#_M1029_d 0.0030829f $X=9.26 $Y=0.77 $X2=0 $Y2=0
cc_530 N_Y_c_845_n N_A_1163_47#_M1038_d 4.94239e-19 $X=9.26 $Y=0.77 $X2=0 $Y2=0
cc_531 N_Y_c_805_n N_A_1163_47#_M1038_d 0.00346845f $X=9.417 $Y=0.885 $X2=0
+ $Y2=0
cc_532 N_Y_M1002_s N_A_1163_47#_c_1169_n 0.0030596f $X=7.925 $Y=0.235 $X2=0
+ $Y2=0
cc_533 N_Y_M1037_s N_A_1163_47#_c_1169_n 0.0030596f $X=8.765 $Y=0.235 $X2=0
+ $Y2=0
cc_534 N_Y_c_845_n N_A_1163_47#_c_1169_n 0.0673613f $X=9.26 $Y=0.77 $X2=0 $Y2=0
cc_535 N_Y_c_805_n N_A_1163_47#_c_1169_n 0.025158f $X=9.417 $Y=0.885 $X2=0 $Y2=0
cc_536 N_VGND_c_926_n N_A_125_47#_M1011_d 0.00412745f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_537 N_VGND_c_926_n N_A_125_47#_M1024_d 0.00254582f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_926_n N_A_125_47#_M1020_d 0.00254582f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_926_n N_A_125_47#_M1026_d 0.00254582f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_926_n N_A_125_47#_M1008_d 0.00254582f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_926_n N_A_125_47#_M1017_d 0.00254582f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_c_926_n N_A_125_47#_M1018_s 0.00216833f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_926_n N_A_125_47#_M1028_s 0.00216833f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_923_n N_A_125_47#_c_1120_n 0.0113346f $X=1.015 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_926_n N_A_125_47#_c_1120_n 0.00645703f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_546 N_VGND_M1015_s N_A_125_47#_c_1068_n 0.00307912f $X=1.045 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_VGND_c_910_n N_A_125_47#_c_1068_n 0.0163853f $X=1.18 $Y=0.36 $X2=0
+ $Y2=0
cc_548 N_VGND_c_923_n N_A_125_47#_c_1068_n 0.00235985f $X=1.015 $Y=0 $X2=0 $Y2=0
cc_549 N_VGND_c_924_n N_A_125_47#_c_1068_n 0.00235985f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_926_n N_A_125_47#_c_1068_n 0.00984999f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_551 N_VGND_c_924_n N_A_125_47#_c_1127_n 0.0113346f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_926_n N_A_125_47#_c_1127_n 0.00645703f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_M1025_s N_A_125_47#_c_1074_n 0.00326179f $X=1.885 $Y=0.235 $X2=0
+ $Y2=0
cc_554 N_VGND_c_911_n N_A_125_47#_c_1074_n 0.0163853f $X=2.02 $Y=0.36 $X2=0
+ $Y2=0
cc_555 N_VGND_c_917_n N_A_125_47#_c_1074_n 0.00235985f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_924_n N_A_125_47#_c_1074_n 0.00235985f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_926_n N_A_125_47#_c_1074_n 0.00984999f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_c_917_n N_A_125_47#_c_1134_n 0.0113346f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_926_n N_A_125_47#_c_1134_n 0.00645703f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_M1021_s N_A_125_47#_c_1080_n 0.00307912f $X=2.725 $Y=0.235 $X2=0
+ $Y2=0
cc_561 N_VGND_c_912_n N_A_125_47#_c_1080_n 0.0163853f $X=2.86 $Y=0.36 $X2=0
+ $Y2=0
cc_562 N_VGND_c_917_n N_A_125_47#_c_1080_n 0.00235985f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_563 N_VGND_c_919_n N_A_125_47#_c_1080_n 0.00235985f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_564 N_VGND_c_926_n N_A_125_47#_c_1080_n 0.00984999f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_565 N_VGND_c_919_n N_A_125_47#_c_1141_n 0.0113346f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_566 N_VGND_c_926_n N_A_125_47#_c_1141_n 0.00645703f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_M1035_s N_A_125_47#_c_1084_n 0.00536163f $X=3.565 $Y=0.235 $X2=0
+ $Y2=0
cc_568 N_VGND_c_913_n N_A_125_47#_c_1084_n 0.0179513f $X=3.72 $Y=0.36 $X2=0
+ $Y2=0
cc_569 N_VGND_c_919_n N_A_125_47#_c_1084_n 0.00235985f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_c_921_n N_A_125_47#_c_1084_n 0.00235985f $X=4.395 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_926_n N_A_125_47#_c_1084_n 0.00993797f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_921_n N_A_125_47#_c_1148_n 0.0113346f $X=4.395 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_926_n N_A_125_47#_c_1148_n 0.00645703f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_M1016_s N_A_125_47#_c_1092_n 0.00307912f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_575 N_VGND_c_914_n N_A_125_47#_c_1092_n 0.0163853f $X=4.56 $Y=0.36 $X2=0
+ $Y2=0
cc_576 N_VGND_c_915_n N_A_125_47#_c_1092_n 0.00235985f $X=5.235 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_c_921_n N_A_125_47#_c_1092_n 0.00235985f $X=4.395 $Y=0 $X2=0 $Y2=0
cc_578 N_VGND_c_926_n N_A_125_47#_c_1092_n 0.00984999f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_579 N_VGND_c_915_n N_A_125_47#_c_1155_n 0.0113346f $X=5.235 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_926_n N_A_125_47#_c_1155_n 0.00645703f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_M1031_s N_A_125_47#_c_1062_n 0.00539394f $X=5.265 $Y=0.235 $X2=0
+ $Y2=0
cc_582 N_VGND_c_915_n N_A_125_47#_c_1062_n 0.00235985f $X=5.235 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_916_n N_A_125_47#_c_1062_n 0.0227163f $X=5.4 $Y=0.36 $X2=0 $Y2=0
cc_584 N_VGND_c_925_n N_A_125_47#_c_1062_n 0.0030357f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_926_n N_A_125_47#_c_1062_n 0.0136387f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_926_n N_A_1163_47#_M1018_d 0.00225742f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_587 N_VGND_c_926_n N_A_1163_47#_M1019_d 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_926_n N_A_1163_47#_M1032_d 0.0021521f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_926_n N_A_1163_47#_M1029_d 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_926_n N_A_1163_47#_M1038_d 0.00225742f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_916_n N_A_1163_47#_c_1167_n 0.0202541f $X=5.4 $Y=0.36 $X2=0
+ $Y2=0
cc_592 N_VGND_c_925_n N_A_1163_47#_c_1167_n 0.102037f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_926_n N_A_1163_47#_c_1167_n 0.0644622f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_925_n N_A_1163_47#_c_1169_n 0.105327f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_926_n N_A_1163_47#_c_1169_n 0.0663367f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_925_n N_A_1163_47#_c_1198_n 0.0114055f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_926_n N_A_1163_47#_c_1198_n 0.00653405f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_598 N_A_125_47#_c_1062_n N_A_1163_47#_M1018_d 0.00736278f $X=7.22 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_599 N_A_125_47#_c_1062_n N_A_1163_47#_M1019_d 0.0030829f $X=7.22 $Y=0.76
+ $X2=0 $Y2=0
cc_600 N_A_125_47#_M1018_s N_A_1163_47#_c_1167_n 0.0030596f $X=6.245 $Y=0.235
+ $X2=0 $Y2=0
cc_601 N_A_125_47#_M1028_s N_A_1163_47#_c_1167_n 0.0030596f $X=7.085 $Y=0.235
+ $X2=0 $Y2=0
cc_602 N_A_125_47#_c_1062_n N_A_1163_47#_c_1167_n 0.0867371f $X=7.22 $Y=0.76
+ $X2=0 $Y2=0

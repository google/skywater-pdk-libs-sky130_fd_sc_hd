# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.740000 1.020000 4.975000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.637500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.635000 4.975000 0.850000 ;
        RECT 3.190000 0.850000 3.570000 1.445000 ;
        RECT 3.190000 1.445000 4.360000 1.615000 ;
        RECT 3.190000 1.615000 3.520000 2.125000 ;
        RECT 4.030000 1.615000 4.360000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.695000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.695000 0.995000 ;
      RECT 0.500000  0.995000 3.020000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.035000  0.255000 1.205000 0.655000 ;
      RECT 1.035000  0.655000 3.020000 0.825000 ;
      RECT 1.075000  1.555000 2.995000 1.725000 ;
      RECT 1.075000  1.725000 1.285000 2.465000 ;
      RECT 1.375000  0.085000 1.705000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.875000  0.255000 2.045000 0.655000 ;
      RECT 1.955000  1.725000 2.125000 2.465000 ;
      RECT 2.215000  0.085000 2.555000 0.485000 ;
      RECT 2.295000  1.895000 2.655000 2.635000 ;
      RECT 2.735000  0.255000 4.975000 0.465000 ;
      RECT 2.735000  0.465000 3.020000 0.655000 ;
      RECT 2.825000  1.725000 2.995000 2.295000 ;
      RECT 2.825000  2.295000 4.975000 2.465000 ;
      RECT 3.690000  1.785000 3.860000 2.295000 ;
      RECT 4.530000  1.445000 4.975000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_4
END LIBRARY

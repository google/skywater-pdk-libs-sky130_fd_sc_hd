* File: sky130_fd_sc_hd__or3_4.spice.SKY130_FD_SC_HD__OR3_4.pxi
* Created: Thu Aug 27 14:43:31 2020
* 
x_PM_SKY130_FD_SC_HD__OR3_4%C N_C_c_78_n N_C_M1012_g N_C_M1008_g C N_C_c_80_n
+ PM_SKY130_FD_SC_HD__OR3_4%C
x_PM_SKY130_FD_SC_HD__OR3_4%B N_B_c_106_n N_B_M1004_g N_B_M1002_g N_B_c_107_n
+ N_B_c_108_n B B PM_SKY130_FD_SC_HD__OR3_4%B
x_PM_SKY130_FD_SC_HD__OR3_4%A N_A_M1007_g N_A_M1000_g A N_A_c_146_n N_A_c_147_n
+ PM_SKY130_FD_SC_HD__OR3_4%A
x_PM_SKY130_FD_SC_HD__OR3_4%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1004_d
+ N_A_27_47#_M1008_s N_A_27_47#_c_185_n N_A_27_47#_M1009_g N_A_27_47#_M1001_g
+ N_A_27_47#_c_186_n N_A_27_47#_M1010_g N_A_27_47#_M1003_g N_A_27_47#_c_187_n
+ N_A_27_47#_M1011_g N_A_27_47#_M1005_g N_A_27_47#_c_188_n N_A_27_47#_M1013_g
+ N_A_27_47#_M1006_g N_A_27_47#_c_189_n N_A_27_47#_c_203_n N_A_27_47#_c_204_n
+ N_A_27_47#_c_190_n N_A_27_47#_c_191_n N_A_27_47#_c_216_n N_A_27_47#_c_217_n
+ N_A_27_47#_c_233_n N_A_27_47#_c_192_n N_A_27_47#_c_237_n N_A_27_47#_c_226_n
+ N_A_27_47#_c_193_n N_A_27_47#_c_194_n N_A_27_47#_c_195_n N_A_27_47#_c_196_n
+ N_A_27_47#_c_197_n N_A_27_47#_c_198_n PM_SKY130_FD_SC_HD__OR3_4%A_27_47#
x_PM_SKY130_FD_SC_HD__OR3_4%VPWR N_VPWR_M1000_d N_VPWR_M1003_s N_VPWR_M1006_s
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n VPWR N_VPWR_c_360_n
+ N_VPWR_c_351_n N_VPWR_c_362_n PM_SKY130_FD_SC_HD__OR3_4%VPWR
x_PM_SKY130_FD_SC_HD__OR3_4%X N_X_M1009_s N_X_M1011_s N_X_M1001_d N_X_M1005_d
+ N_X_c_415_n N_X_c_410_n N_X_c_454_n N_X_c_411_n N_X_c_404_n N_X_c_405_n
+ N_X_c_436_n N_X_c_458_n N_X_c_412_n N_X_c_406_n N_X_c_407_n N_X_c_413_n X
+ N_X_c_409_n PM_SKY130_FD_SC_HD__OR3_4%X
x_PM_SKY130_FD_SC_HD__OR3_4%VGND N_VGND_M1012_d N_VGND_M1007_d N_VGND_M1010_d
+ N_VGND_M1013_d N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n
+ N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n
+ VGND N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n
+ PM_SKY130_FD_SC_HD__OR3_4%VGND
cc_1 VNB N_C_c_78_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB C 0.00896247f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_c_80_n 0.0360339f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B_c_106_n 0.0162239f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_B_c_107_n 0.00449274f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_6 VNB N_B_c_108_n 0.0190353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB A 0.00454089f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_c_146_n 0.0221506f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_9 VNB N_A_c_147_n 0.0199492f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_185_n 0.0190947f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_11 VNB N_A_27_47#_c_186_n 0.0157974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_187_n 0.0157986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_188_n 0.0192362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_189_n 0.0187495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_190_n 0.0035423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_191_n 0.0096461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_192_n 0.00499152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_193_n 0.00291462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_194_n 3.90207e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_195_n 0.0015776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_196_n 0.00311049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_197_n 0.00113699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_198_n 0.0850078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_351_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_404_n 0.00217862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_405_n 0.00222466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_406_n 0.00226423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_407_n 0.00222466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB X 0.0221383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_409_n 0.0100985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_481_n 0.00410729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_482_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_483_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_484_n 0.0171314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_485_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_486_n 0.0176032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_487_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_488_n 0.0169753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_489_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_490_n 0.0116138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_491_n 0.219819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_492_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_493_n 0.019982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VPB N_C_M1008_g 0.0262632f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB C 0.00359492f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_46 VPB N_C_c_80_n 0.00949799f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_47 VPB N_B_M1002_g 0.0182245f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_48 VPB N_B_c_107_n 9.58651e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_B_c_108_n 0.00506541f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB B 0.0019548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_M1000_g 0.0232584f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_52 VPB A 0.00194567f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_53 VPB N_A_c_146_n 0.00451126f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_54 VPB N_A_27_47#_M1001_g 0.0219104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_M1003_g 0.0182177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_M1005_g 0.0182024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_M1006_g 0.0220253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_203_n 0.00759484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_204_n 0.0317434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_194_n 0.00364496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_198_n 0.0202201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_352_n 0.00704479f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_63 VPB N_VPWR_c_353_n 0.00397811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_354_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_355_n 0.0176511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_356_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_357_n 0.0112126f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_358_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_359_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_360_n 0.0363217f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_351_n 0.04719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_362_n 0.0134347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_X_c_410_n 0.00248279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_X_c_411_n 0.00252706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_X_c_412_n 0.0141375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_X_c_413_n 0.00220075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB X 0.00853041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 N_C_c_78_n N_B_c_106_n 0.0258694f $X=0.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_79 N_C_M1008_g N_B_M1002_g 0.0567245f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_80 C N_B_c_107_n 0.0202944f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_81 N_C_c_80_n N_B_c_107_n 0.00190655f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C_c_80_n N_B_c_108_n 0.0216732f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_83 N_C_M1008_g B 0.00636768f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_84 N_C_c_78_n N_A_27_47#_c_189_n 0.00630972f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_85 N_C_M1008_g N_A_27_47#_c_203_n 7.12665e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_86 N_C_M1008_g N_A_27_47#_c_204_n 0.0106949f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_87 C N_A_27_47#_c_204_n 0.0250713f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_88 N_C_c_80_n N_A_27_47#_c_204_n 0.00196424f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_89 N_C_c_78_n N_A_27_47#_c_190_n 0.0123222f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C_c_78_n N_A_27_47#_c_191_n 0.00129702f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_91 C N_A_27_47#_c_191_n 0.0280294f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_92 N_C_c_80_n N_A_27_47#_c_191_n 0.00690502f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_93 N_C_M1008_g N_A_27_47#_c_216_n 0.0100707f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_94 N_C_c_78_n N_A_27_47#_c_217_n 5.22228e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_95 N_C_M1008_g N_VPWR_c_360_n 0.00357835f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_96 N_C_M1008_g N_VPWR_c_351_n 0.00620759f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_97 N_C_c_78_n N_VGND_c_481_n 0.00268723f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_98 N_C_c_78_n N_VGND_c_484_n 0.00423334f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_99 N_C_c_78_n N_VGND_c_491_n 0.00669771f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B_M1002_g N_A_M1000_g 0.0573576f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 B N_A_M1000_g 0.00121961f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_102 N_B_c_107_n A 0.0219556f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_c_108_n A 8.07997e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B_c_107_n N_A_c_146_n 8.42607e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B_c_108_n N_A_c_146_n 0.0220076f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B_c_106_n N_A_c_147_n 0.0124239f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B_c_106_n N_A_27_47#_c_189_n 5.22062e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B_M1002_g N_A_27_47#_c_204_n 0.00115568f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B_c_106_n N_A_27_47#_c_190_n 0.00865686f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B_c_107_n N_A_27_47#_c_190_n 0.0252826f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B_c_108_n N_A_27_47#_c_190_n 0.00148089f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B_M1002_g N_A_27_47#_c_216_n 0.0137123f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_113 B N_A_27_47#_c_216_n 0.0093945f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_114 N_B_c_106_n N_A_27_47#_c_217_n 0.00630972f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_107_n N_A_27_47#_c_226_n 0.00358699f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B_c_108_n N_A_27_47#_c_226_n 5.15355e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B_c_106_n N_A_27_47#_c_196_n 0.00112787f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B_c_107_n N_A_27_47#_c_196_n 0.00987832f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B_c_108_n N_A_27_47#_c_196_n 0.00153559f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_120 B A_109_297# 0.00289592f $X=0.61 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_121 N_B_M1002_g N_VPWR_c_360_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B_M1002_g N_VPWR_c_351_n 0.00532055f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B_c_106_n N_VGND_c_481_n 0.00146339f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_106_n N_VGND_c_491_n 0.00577071f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B_c_106_n N_VGND_c_492_n 0.00423334f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_M1000_g N_A_27_47#_c_216_n 0.00407199f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_c_147_n N_A_27_47#_c_217_n 0.0109565f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_M1000_g N_A_27_47#_c_233_n 0.0179813f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_129 A N_A_27_47#_c_192_n 0.0323643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A_c_146_n N_A_27_47#_c_192_n 0.00345541f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_147_n N_A_27_47#_c_192_n 0.0108831f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_M1000_g N_A_27_47#_c_237_n 0.0127759f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_133 A N_A_27_47#_c_237_n 0.0297381f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_c_146_n N_A_27_47#_c_237_n 0.00301383f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_M1000_g N_A_27_47#_c_226_n 0.00245009f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_136 A N_A_27_47#_c_226_n 0.00274851f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A_c_146_n N_A_27_47#_c_193_n 0.00149709f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_147_n N_A_27_47#_c_193_n 0.00225679f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_A_27_47#_c_194_n 0.00428536f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_140 A N_A_27_47#_c_194_n 0.00655732f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_141 A N_A_27_47#_c_196_n 0.00320352f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_142 N_A_c_147_n N_A_27_47#_c_196_n 0.00112787f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_143 A N_A_27_47#_c_197_n 0.0154158f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A_c_146_n N_A_27_47#_c_197_n 4.82661e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_145 A N_A_27_47#_c_198_n 9.18726e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A_c_146_n N_A_27_47#_c_198_n 0.0101041f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_VPWR_c_352_n 0.0173183f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1000_g N_VPWR_c_360_n 0.00539841f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1000_g N_VPWR_c_351_n 0.0109844f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_c_147_n N_VGND_c_491_n 0.00706711f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_147_n N_VGND_c_492_n 0.00423334f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_147_n N_VGND_c_493_n 0.00336132f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_216_n A_109_297# 0.00341692f $X=1 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_27_47#_c_216_n A_193_297# 0.0015256f $X=1 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_155 N_A_27_47#_c_233_n A_193_297# 8.21952e-19 $X=1.132 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_27_47#_c_226_n A_193_297# 0.0028989f $X=1.265 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A_27_47#_c_237_n N_VPWR_M1000_d 0.0189723f $X=1.87 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_27_47#_c_194_n N_VPWR_M1000_d 2.28327e-19 $X=1.98 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_27_47#_M1001_g N_VPWR_c_352_n 0.00330246f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_237_n N_VPWR_c_352_n 0.0545304f $X=1.87 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_195_n N_VPWR_c_352_n 0.00119333f $X=3.425 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_198_n N_VPWR_c_352_n 0.00155946f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1003_g N_VPWR_c_353_n 0.00163116f $X=2.68 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1005_g N_VPWR_c_353_n 0.00157837f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_27_47#_M1006_g N_VPWR_c_354_n 0.00338128f $X=3.52 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_M1001_g N_VPWR_c_355_n 0.00585385f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_M1003_g N_VPWR_c_355_n 0.00585385f $X=2.68 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_M1005_g N_VPWR_c_358_n 0.00585385f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1006_g N_VPWR_c_358_n 0.00585385f $X=3.52 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_203_n N_VPWR_c_360_n 0.0218588f $X=0.255 $Y=2.295 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_216_n N_VPWR_c_360_n 0.0475457f $X=1 $Y=2.38 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1008_s N_VPWR_c_351_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1001_g N_VPWR_c_351_n 0.0118632f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1003_g N_VPWR_c_351_n 0.0104367f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1005_g N_VPWR_c_351_n 0.0104367f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1006_g N_VPWR_c_351_n 0.011507f $X=3.52 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_203_n N_VPWR_c_351_n 0.0128791f $X=0.255 $Y=2.295 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_216_n N_VPWR_c_351_n 0.0302493f $X=1 $Y=2.38 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_185_n N_X_c_415_n 0.0110125f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_186_n N_X_c_415_n 0.00639222f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_187_n N_X_c_415_n 5.48633e-19 $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_192_n N_X_c_415_n 6.57759e-19 $X=1.87 $Y=0.815 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1001_g N_X_c_410_n 3.12327e-19 $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_194_n N_X_c_410_n 0.00215607f $X=1.98 $Y=1.495 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_195_n N_X_c_410_n 0.0172286f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_198_n N_X_c_410_n 0.00226413f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1003_g N_X_c_411_n 0.0134538f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_27_47#_M1005_g N_X_c_411_n 0.013468f $X=3.1 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_195_n N_X_c_411_n 0.03482f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_198_n N_X_c_411_n 0.00216069f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_186_n N_X_c_404_n 0.00850187f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_187_n N_X_c_404_n 0.00850187f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_195_n N_X_c_404_n 0.0355133f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_198_n N_X_c_404_n 0.00221825f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_185_n N_X_c_405_n 0.00271199f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_186_n N_X_c_405_n 0.00110527f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_192_n N_X_c_405_n 0.0124158f $X=1.87 $Y=0.815 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_195_n N_X_c_405_n 0.0262212f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_198_n N_X_c_405_n 0.00230227f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_186_n N_X_c_436_n 5.48633e-19 $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_187_n N_X_c_436_n 0.00639222f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_188_n N_X_c_436_n 0.0112717f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_27_47#_M1006_g N_X_c_412_n 0.0152886f $X=3.52 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_195_n N_X_c_412_n 0.00916434f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_188_n N_X_c_406_n 0.0102783f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_195_n N_X_c_406_n 0.00809975f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_187_n N_X_c_407_n 0.00110527f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_188_n N_X_c_407_n 0.00110527f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_195_n N_X_c_407_n 0.0262212f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_198_n N_X_c_407_n 0.00230227f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_195_n N_X_c_413_n 0.0172286f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_198_n N_X_c_413_n 0.00226413f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_188_n X 0.00679473f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_195_n X 0.0139618f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_198_n X 0.0094714f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_190_n N_VGND_M1012_d 0.00162089f $X=0.935 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_27_47#_c_192_n N_VGND_M1007_d 0.0115157f $X=1.87 $Y=0.815 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_190_n N_VGND_c_481_n 0.0122559f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_186_n N_VGND_c_482_n 0.00146339f $X=2.68 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_187_n N_VGND_c_482_n 0.00146448f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_188_n N_VGND_c_483_n 0.00316354f $X=3.52 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_189_n N_VGND_c_484_n 0.0216897f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_190_n N_VGND_c_484_n 0.00198695f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_185_n N_VGND_c_486_n 0.00541763f $X=2.26 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_186_n N_VGND_c_486_n 0.0042482f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_187_n N_VGND_c_488_n 0.0042482f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_188_n N_VGND_c_488_n 0.0042482f $X=3.52 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_27_47#_M1012_s N_VGND_c_491_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1004_d N_VGND_c_491_n 0.00215201f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_185_n N_VGND_c_491_n 0.0108255f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_186_n N_VGND_c_491_n 0.00573646f $X=2.68 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_187_n N_VGND_c_491_n 0.00573646f $X=3.1 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_188_n N_VGND_c_491_n 0.00680668f $X=3.52 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_189_n N_VGND_c_491_n 0.0127966f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_190_n N_VGND_c_491_n 0.00835832f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_217_n N_VGND_c_491_n 0.0122069f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_192_n N_VGND_c_491_n 0.00645912f $X=1.87 $Y=0.815 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_190_n N_VGND_c_492_n 0.00198695f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_217_n N_VGND_c_492_n 0.0188551f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_192_n N_VGND_c_492_n 0.00198695f $X=1.87 $Y=0.815 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_185_n N_VGND_c_493_n 0.00336132f $X=2.26 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_192_n N_VGND_c_493_n 0.0523434f $X=1.87 $Y=0.815 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_195_n N_VGND_c_493_n 0.00133125f $X=3.425 $Y=1.16 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_198_n N_VGND_c_493_n 0.00170541f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_245 A_109_297# N_VPWR_c_351_n 0.00216833f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_246 A_193_297# N_VPWR_c_351_n 0.0021681f $X=0.965 $Y=1.485 $X2=0.425
+ $Y2=0.815
cc_247 N_VPWR_c_351_n N_X_M1001_d 0.00284632f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_248 N_VPWR_c_351_n N_X_M1005_d 0.00284632f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_c_355_n N_X_c_454_n 0.0142343f $X=2.765 $Y=2.72 $X2=0 $Y2=0
cc_250 N_VPWR_c_351_n N_X_c_454_n 0.00955092f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_251 N_VPWR_M1003_s N_X_c_411_n 0.00165831f $X=2.755 $Y=1.485 $X2=0 $Y2=0
cc_252 N_VPWR_c_353_n N_X_c_411_n 0.0126919f $X=2.89 $Y=1.96 $X2=0 $Y2=0
cc_253 N_VPWR_c_358_n N_X_c_458_n 0.0142343f $X=3.605 $Y=2.72 $X2=0 $Y2=0
cc_254 N_VPWR_c_351_n N_X_c_458_n 0.00955092f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_255 N_VPWR_M1006_s N_X_c_412_n 0.00812647f $X=3.595 $Y=1.485 $X2=0 $Y2=0
cc_256 N_VPWR_c_354_n N_X_c_412_n 0.0171814f $X=3.73 $Y=1.96 $X2=0 $Y2=0
cc_257 N_X_c_404_n N_VGND_M1010_d 0.00165819f $X=3.145 $Y=0.82 $X2=0 $Y2=0
cc_258 N_X_c_406_n N_VGND_M1013_d 0.00119049f $X=3.765 $Y=0.82 $X2=0 $Y2=0
cc_259 N_X_c_409_n N_VGND_M1013_d 0.00359674f $X=3.91 $Y=0.905 $X2=0 $Y2=0
cc_260 N_X_c_404_n N_VGND_c_482_n 0.0116528f $X=3.145 $Y=0.82 $X2=0 $Y2=0
cc_261 N_X_c_406_n N_VGND_c_483_n 0.00840877f $X=3.765 $Y=0.82 $X2=0 $Y2=0
cc_262 N_X_c_409_n N_VGND_c_483_n 0.00404097f $X=3.91 $Y=0.905 $X2=0 $Y2=0
cc_263 N_X_c_415_n N_VGND_c_486_n 0.017716f $X=2.47 $Y=0.39 $X2=0 $Y2=0
cc_264 N_X_c_404_n N_VGND_c_486_n 0.00193763f $X=3.145 $Y=0.82 $X2=0 $Y2=0
cc_265 N_X_c_404_n N_VGND_c_488_n 0.00193763f $X=3.145 $Y=0.82 $X2=0 $Y2=0
cc_266 N_X_c_436_n N_VGND_c_488_n 0.017716f $X=3.31 $Y=0.39 $X2=0 $Y2=0
cc_267 N_X_c_406_n N_VGND_c_488_n 0.00193763f $X=3.765 $Y=0.82 $X2=0 $Y2=0
cc_268 N_X_c_409_n N_VGND_c_490_n 0.00391203f $X=3.91 $Y=0.905 $X2=0 $Y2=0
cc_269 N_X_M1009_s N_VGND_c_491_n 0.00215535f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_270 N_X_M1011_s N_VGND_c_491_n 0.00215535f $X=3.175 $Y=0.235 $X2=0 $Y2=0
cc_271 N_X_c_415_n N_VGND_c_491_n 0.0121406f $X=2.47 $Y=0.39 $X2=0 $Y2=0
cc_272 N_X_c_404_n N_VGND_c_491_n 0.00827287f $X=3.145 $Y=0.82 $X2=0 $Y2=0
cc_273 N_X_c_436_n N_VGND_c_491_n 0.0121406f $X=3.31 $Y=0.39 $X2=0 $Y2=0
cc_274 N_X_c_406_n N_VGND_c_491_n 0.00426887f $X=3.765 $Y=0.82 $X2=0 $Y2=0
cc_275 N_X_c_409_n N_VGND_c_491_n 0.00696444f $X=3.91 $Y=0.905 $X2=0 $Y2=0

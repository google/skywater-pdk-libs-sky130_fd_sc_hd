* File: sky130_fd_sc_hd__a22o_1.pxi.spice
* Created: Thu Aug 27 14:02:26 2020
* 
x_PM_SKY130_FD_SC_HD__A22O_1%B2 N_B2_M1008_g N_B2_M1004_g B2 N_B2_c_58_n
+ N_B2_c_59_n N_B2_c_60_n PM_SKY130_FD_SC_HD__A22O_1%B2
x_PM_SKY130_FD_SC_HD__A22O_1%B1 N_B1_M1001_g N_B1_M1002_g B1 B1 N_B1_c_86_n
+ N_B1_c_87_n PM_SKY130_FD_SC_HD__A22O_1%B1
x_PM_SKY130_FD_SC_HD__A22O_1%A1 N_A1_c_125_n N_A1_M1006_g N_A1_c_126_n
+ N_A1_M1000_g A1 A1 PM_SKY130_FD_SC_HD__A22O_1%A1
x_PM_SKY130_FD_SC_HD__A22O_1%A2 N_A2_c_162_n N_A2_M1005_g N_A2_c_163_n
+ N_A2_M1007_g A2 N_A2_c_164_n PM_SKY130_FD_SC_HD__A22O_1%A2
x_PM_SKY130_FD_SC_HD__A22O_1%A_27_297# N_A_27_297#_M1001_d N_A_27_297#_M1006_s
+ N_A_27_297#_M1004_s N_A_27_297#_M1002_d N_A_27_297#_M1003_g
+ N_A_27_297#_M1009_g N_A_27_297#_c_208_n N_A_27_297#_c_209_n
+ N_A_27_297#_c_202_n N_A_27_297#_c_210_n N_A_27_297#_c_242_n
+ N_A_27_297#_c_251_n N_A_27_297#_c_243_n N_A_27_297#_c_203_n
+ N_A_27_297#_c_204_n N_A_27_297#_c_205_n N_A_27_297#_c_213_n
+ N_A_27_297#_c_214_n N_A_27_297#_c_215_n N_A_27_297#_c_206_n
+ PM_SKY130_FD_SC_HD__A22O_1%A_27_297#
x_PM_SKY130_FD_SC_HD__A22O_1%A_109_297# N_A_109_297#_M1004_d
+ N_A_109_297#_M1000_d N_A_109_297#_c_311_n N_A_109_297#_c_309_n
+ N_A_109_297#_c_324_p N_A_109_297#_c_310_n
+ PM_SKY130_FD_SC_HD__A22O_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A22O_1%VPWR N_VPWR_M1000_s N_VPWR_M1007_d N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n VPWR N_VPWR_c_339_n N_VPWR_c_340_n
+ N_VPWR_c_335_n N_VPWR_c_342_n N_VPWR_c_343_n PM_SKY130_FD_SC_HD__A22O_1%VPWR
x_PM_SKY130_FD_SC_HD__A22O_1%X N_X_M1003_d N_X_M1009_d N_X_c_382_n X X X
+ PM_SKY130_FD_SC_HD__A22O_1%X
x_PM_SKY130_FD_SC_HD__A22O_1%VGND N_VGND_M1008_s N_VGND_M1005_d N_VGND_c_398_n
+ N_VGND_c_399_n N_VGND_c_400_n VGND N_VGND_c_401_n N_VGND_c_402_n
+ N_VGND_c_403_n N_VGND_c_404_n PM_SKY130_FD_SC_HD__A22O_1%VGND
cc_1 VNB N_B2_c_58_n 0.0271486f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_2 VNB N_B2_c_59_n 0.0144124f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_3 VNB N_B2_c_60_n 0.0202523f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_4 VNB B1 0.00544773f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB B1 0.00543772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_B1_c_86_n 0.023835f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_7 VNB N_B1_c_87_n 0.0190454f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_8 VNB N_A1_c_125_n 0.0199438f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_9 VNB N_A1_c_126_n 0.0296627f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_10 VNB A1 0.00257773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A1 0.00175555f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_A2_c_162_n 0.0155225f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_A2_c_163_n 0.0221813f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_14 VNB N_A2_c_164_n 0.00487814f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_15 VNB N_A_27_297#_c_202_n 0.0121231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_203_n 0.00132262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_204_n 9.16142e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_205_n 0.0316546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_206_n 0.0189156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_335_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_382_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_22 VNB X 0.0303219f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_23 VNB N_VGND_c_398_n 0.0118708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_399_n 0.0280194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_400_n 0.00280379f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_26 VNB N_VGND_c_401_n 0.0434773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_402_n 0.0147189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_403_n 0.182415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_404_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_B2_M1004_g 0.0255531f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_31 VPB N_B2_c_58_n 0.00476222f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_32 VPB N_B1_M1002_g 0.0240877f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB N_B1_c_86_n 0.0048554f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_34 VPB N_A1_c_126_n 0.0347399f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_35 VPB N_A2_c_163_n 0.00427048f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_36 VPB N_A2_M1007_g 0.0198764f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A2_c_164_n 0.00304462f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_38 VPB N_A_27_297#_M1009_g 0.0214778f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.175
cc_39 VPB N_A_27_297#_c_208_n 0.0233212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_297#_c_209_n 0.00948748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_297#_c_210_n 0.0115397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_297#_c_204_n 0.00152104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_297#_c_205_n 0.00884434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_297#_c_213_n 0.00889261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_297#_c_214_n 0.00743097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_297#_c_215_n 0.00519526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_109_297#_c_309_n 0.00355166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_109_297#_c_310_n 0.00459344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_336_n 0.0069237f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_337_n 0.0171091f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_51 VPB N_VPWR_c_338_n 0.00184392f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_52 VPB N_VPWR_c_339_n 0.0405947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_340_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_335_n 0.0461466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_342_n 0.00549283f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_343_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB X 0.0452842f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_58 N_B2_M1004_g N_B1_M1002_g 0.0436496f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_59 N_B2_c_58_n B1 3.38478e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_60 N_B2_c_58_n B1 9.18012e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_61 N_B2_c_59_n B1 0.0162709f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B2_c_58_n N_B1_c_86_n 0.033955f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_63 N_B2_c_59_n N_B1_c_86_n 7.16521e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B2_c_60_n N_B1_c_87_n 0.033955f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_65 N_B2_c_58_n N_A_27_297#_c_209_n 0.00172397f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_66 N_B2_c_59_n N_A_27_297#_c_209_n 0.0206403f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B2_c_60_n N_A_27_297#_c_202_n 6.07844e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_68 N_B2_M1004_g N_A_27_297#_c_213_n 0.00507721f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 N_B2_M1004_g N_A_27_297#_c_214_n 0.0130391f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_70 N_B2_c_58_n N_A_27_297#_c_214_n 0.00117895f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B2_c_59_n N_A_27_297#_c_214_n 0.015462f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B2_M1004_g N_A_27_297#_c_215_n 2.69644e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_73 N_B2_M1004_g N_VPWR_c_339_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_74 N_B2_M1004_g N_VPWR_c_335_n 0.0106826f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_75 N_B2_c_58_n N_VGND_c_399_n 0.00275758f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B2_c_59_n N_VGND_c_399_n 0.0274141f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B2_c_60_n N_VGND_c_399_n 0.0267674f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B2_c_60_n N_VGND_c_403_n 7.20442e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B1_M1002_g N_A1_c_126_n 0.00220187f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_80 B1 N_A1_c_126_n 3.01697e-19 $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_81 B1 N_A1_c_126_n 8.92876e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_82 N_B1_c_86_n N_A1_c_126_n 0.00880991f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_83 B1 A1 0.0238753f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_84 N_B1_c_86_n A1 2.12022e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_85 B1 A1 0.0138885f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B1_c_86_n A1 5.95583e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_87 B1 N_A_27_297#_M1001_d 0.00578233f $X=1.07 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_88 B1 N_A_27_297#_c_202_n 0.0138186f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_89 B1 N_A_27_297#_c_202_n 0.00429942f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B1_c_86_n N_A_27_297#_c_202_n 0.00174563f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B1_c_87_n N_A_27_297#_c_202_n 0.00747225f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B1_M1002_g N_A_27_297#_c_213_n 0.0010873f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 N_B1_M1002_g N_A_27_297#_c_214_n 0.00745625f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_94 B1 N_A_27_297#_c_214_n 0.035387f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B1_c_86_n N_A_27_297#_c_214_n 0.00110462f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B1_M1002_g N_A_27_297#_c_215_n 0.00351756f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B1_c_86_n N_A_27_297#_c_215_n 0.00237455f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_98 N_B1_M1002_g N_A_109_297#_c_311_n 0.00214252f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_99 N_B1_M1002_g N_A_109_297#_c_310_n 0.0128426f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_VPWR_c_336_n 0.00845597f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B1_M1002_g N_VPWR_c_339_n 0.00424683f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_M1002_g N_VPWR_c_335_n 0.00727577f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_103 B1 N_VGND_c_399_n 0.00606901f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_104 N_B1_c_87_n N_VGND_c_399_n 0.00425856f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B1_c_87_n N_VGND_c_401_n 0.0042613f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B1_c_87_n N_VGND_c_403_n 0.0081372f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A1_c_125_n N_A2_c_162_n 0.0267871f $X=1.79 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_108 N_A1_c_125_n N_A2_c_163_n 0.0183693f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A1_c_126_n N_A2_c_163_n 0.00326474f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_110 A1 N_A2_c_163_n 2.5356e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A1_c_126_n N_A2_M1007_g 0.024042f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A1_c_126_n N_A2_c_164_n 0.00319547f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_113 A1 N_A2_c_164_n 0.0017897f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_114 A1 N_A2_c_164_n 0.0169123f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_115 A1 N_A_27_297#_M1006_s 0.00569149f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_116 N_A1_c_125_n N_A_27_297#_c_202_n 0.011544f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A1_c_126_n N_A_27_297#_c_202_n 6.6454e-19 $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_118 A1 N_A_27_297#_c_202_n 0.0107791f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_119 A1 N_A_27_297#_c_202_n 0.00270345f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A1_c_126_n N_A_27_297#_c_210_n 0.0213932f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_121 A1 N_A_27_297#_c_210_n 0.0168877f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A1_c_125_n N_A_27_297#_c_242_n 0.00353591f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A1_c_125_n N_A_27_297#_c_243_n 0.00298703f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A1_c_126_n N_A_27_297#_c_215_n 0.00252921f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_126_n N_A_109_297#_c_309_n 0.0131089f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A1_c_126_n N_VPWR_c_336_n 0.00873033f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A1_c_126_n N_VPWR_c_337_n 0.00311027f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A1_c_126_n N_VPWR_c_335_n 0.00380419f $X=1.82 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A1_c_125_n N_VGND_c_401_n 0.00357877f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A1_c_125_n N_VGND_c_403_n 0.00677073f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_M1007_g N_A_27_297#_M1009_g 0.0249955f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A2_c_162_n N_A_27_297#_c_202_n 0.00249112f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_133 N_A2_c_163_n N_A_27_297#_c_210_n 7.3074e-19 $X=2.29 $Y=1.325 $X2=0 $Y2=0
cc_134 N_A2_M1007_g N_A_27_297#_c_210_n 0.0160837f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A2_c_164_n N_A_27_297#_c_210_n 0.0276239f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A2_c_162_n N_A_27_297#_c_242_n 0.00349096f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_137 N_A2_c_162_n N_A_27_297#_c_251_n 0.0123047f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_138 N_A2_c_163_n N_A_27_297#_c_251_n 0.00207191f $X=2.29 $Y=1.325 $X2=0 $Y2=0
cc_139 N_A2_c_164_n N_A_27_297#_c_251_n 0.0121737f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A2_c_163_n N_A_27_297#_c_243_n 8.52145e-19 $X=2.29 $Y=1.325 $X2=0 $Y2=0
cc_141 N_A2_c_164_n N_A_27_297#_c_243_n 0.00837661f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A2_c_162_n N_A_27_297#_c_203_n 0.00279456f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_143 N_A2_c_162_n N_A_27_297#_c_204_n 0.0016919f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_144 N_A2_c_163_n N_A_27_297#_c_204_n 6.05966e-19 $X=2.29 $Y=1.325 $X2=0 $Y2=0
cc_145 N_A2_M1007_g N_A_27_297#_c_204_n 0.00260422f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A2_c_164_n N_A_27_297#_c_204_n 0.0187519f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_c_163_n N_A_27_297#_c_205_n 0.0210419f $X=2.29 $Y=1.325 $X2=0 $Y2=0
cc_148 N_A2_c_164_n N_A_27_297#_c_205_n 0.001867f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A2_c_162_n N_A_27_297#_c_206_n 0.0219887f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_150 N_A2_M1007_g N_VPWR_c_336_n 5.49415e-19 $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_M1007_g N_VPWR_c_337_n 0.00585385f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A2_M1007_g N_VPWR_c_338_n 0.00437775f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A2_M1007_g N_VPWR_c_335_n 0.0109055f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A2_c_162_n N_VGND_c_400_n 0.00317431f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_155 N_A2_c_162_n N_VGND_c_401_n 0.00422112f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_156 N_A2_c_162_n N_VGND_c_403_n 0.00590531f $X=2.29 $Y=0.96 $X2=0 $Y2=0
cc_157 N_A_27_297#_c_214_n N_A_109_297#_M1004_d 0.00165831f $X=0.935 $Y=1.585
+ $X2=-0.19 $Y2=-0.24
cc_158 N_A_27_297#_c_210_n N_A_109_297#_M1000_d 0.00519899f $X=2.595 $Y=1.6
+ $X2=0 $Y2=0
cc_159 N_A_27_297#_c_214_n N_A_109_297#_c_311_n 0.0124521f $X=0.935 $Y=1.585
+ $X2=0 $Y2=0
cc_160 N_A_27_297#_c_210_n N_A_109_297#_c_309_n 0.0453822f $X=2.595 $Y=1.6 $X2=0
+ $Y2=0
cc_161 N_A_27_297#_M1002_d N_A_109_297#_c_310_n 0.00617549f $X=0.965 $Y=1.485
+ $X2=0 $Y2=0
cc_162 N_A_27_297#_c_210_n N_A_109_297#_c_310_n 0.00707435f $X=2.595 $Y=1.6
+ $X2=0 $Y2=0
cc_163 N_A_27_297#_c_214_n N_A_109_297#_c_310_n 0.00532813f $X=0.935 $Y=1.585
+ $X2=0 $Y2=0
cc_164 N_A_27_297#_c_215_n N_A_109_297#_c_310_n 0.0206661f $X=1.265 $Y=1.585
+ $X2=0 $Y2=0
cc_165 N_A_27_297#_c_210_n N_VPWR_M1000_s 0.00461148f $X=2.595 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_27_297#_c_210_n N_VPWR_M1007_d 0.00851162f $X=2.595 $Y=1.6 $X2=0
+ $Y2=0
cc_167 N_A_27_297#_M1009_g N_VPWR_c_338_n 0.0124779f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_27_297#_c_210_n N_VPWR_c_338_n 0.0155897f $X=2.595 $Y=1.6 $X2=0 $Y2=0
cc_169 N_A_27_297#_c_213_n N_VPWR_c_339_n 0.0212522f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_170 N_A_27_297#_M1009_g N_VPWR_c_340_n 0.0046653f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_27_297#_M1004_s N_VPWR_c_335_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_M1002_d N_VPWR_c_335_n 0.00293129f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_173 N_A_27_297#_M1009_g N_VPWR_c_335_n 0.008846f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_27_297#_c_213_n N_VPWR_c_335_n 0.0125406f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_175 N_A_27_297#_c_205_n N_X_c_382_n 0.00208568f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_27_297#_M1009_g X 0.0103168f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_27_297#_c_210_n X 0.0148838f $X=2.595 $Y=1.6 $X2=0 $Y2=0
cc_178 N_A_27_297#_c_203_n X 0.0194042f $X=2.71 $Y=0.905 $X2=0 $Y2=0
cc_179 N_A_27_297#_c_204_n X 0.0409864f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_205_n X 0.0111991f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_206_n X 0.00817176f $X=2.76 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_251_n N_VGND_M1005_d 0.00493095f $X=2.525 $Y=0.7 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_203_n N_VGND_M1005_d 0.0021798f $X=2.71 $Y=0.905 $X2=0
+ $Y2=0
cc_184 N_A_27_297#_c_202_n N_VGND_c_399_n 0.011553f $X=1.95 $Y=0.36 $X2=0 $Y2=0
cc_185 N_A_27_297#_c_251_n N_VGND_c_400_n 0.00777568f $X=2.525 $Y=0.7 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_c_203_n N_VGND_c_400_n 0.00957953f $X=2.71 $Y=0.905 $X2=0
+ $Y2=0
cc_187 N_A_27_297#_c_206_n N_VGND_c_400_n 0.00808927f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_27_297#_c_202_n N_VGND_c_401_n 0.079152f $X=1.95 $Y=0.36 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_251_n N_VGND_c_401_n 0.00394099f $X=2.525 $Y=0.7 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_c_203_n N_VGND_c_402_n 0.00127967f $X=2.71 $Y=0.905 $X2=0
+ $Y2=0
cc_191 N_A_27_297#_c_206_n N_VGND_c_402_n 0.00380117f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_M1001_d N_VGND_c_403_n 0.00209344f $X=0.925 $Y=0.235 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_M1006_s N_VGND_c_403_n 0.00209344f $X=1.455 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_202_n N_VGND_c_403_n 0.0474779f $X=1.95 $Y=0.36 $X2=0 $Y2=0
cc_195 N_A_27_297#_c_251_n N_VGND_c_403_n 0.00722039f $X=2.525 $Y=0.7 $X2=0
+ $Y2=0
cc_196 N_A_27_297#_c_203_n N_VGND_c_403_n 0.00292689f $X=2.71 $Y=0.905 $X2=0
+ $Y2=0
cc_197 N_A_27_297#_c_206_n N_VGND_c_403_n 0.00599293f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_202_n A_373_47# 0.00588336f $X=1.95 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_199 N_A_27_297#_c_242_n A_373_47# 0.00328891f $X=2.035 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_200 N_A_27_297#_c_251_n A_373_47# 9.949e-19 $X=2.525 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_201 N_A_27_297#_c_243_n A_373_47# 0.00576269f $X=2.12 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_202 N_A_109_297#_c_309_n N_VPWR_M1000_s 0.00471787f $X=2.08 $Y=2.085
+ $X2=-0.19 $Y2=1.305
cc_203 N_A_109_297#_c_309_n N_VPWR_c_336_n 0.022835f $X=2.08 $Y=2.085 $X2=0
+ $Y2=0
cc_204 N_A_109_297#_c_324_p N_VPWR_c_336_n 0.0160476f $X=2.04 $Y=2.3 $X2=0 $Y2=0
cc_205 N_A_109_297#_c_309_n N_VPWR_c_337_n 0.00244585f $X=2.08 $Y=2.085 $X2=0
+ $Y2=0
cc_206 N_A_109_297#_c_324_p N_VPWR_c_337_n 0.015255f $X=2.04 $Y=2.3 $X2=0 $Y2=0
cc_207 N_A_109_297#_c_311_n N_VPWR_c_339_n 0.0040075f $X=0.825 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_109_297#_c_310_n N_VPWR_c_339_n 0.0102405f $X=1.37 $Y=1.98 $X2=0
+ $Y2=0
cc_209 N_A_109_297#_M1004_d N_VPWR_c_335_n 0.00457832f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_210 N_A_109_297#_M1000_d N_VPWR_c_335_n 0.00307681f $X=1.895 $Y=1.485 $X2=0
+ $Y2=0
cc_211 N_A_109_297#_c_311_n N_VPWR_c_335_n 0.0068268f $X=0.825 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_109_297#_c_309_n N_VPWR_c_335_n 0.0059291f $X=2.08 $Y=2.085 $X2=0
+ $Y2=0
cc_213 N_A_109_297#_c_324_p N_VPWR_c_335_n 0.00941222f $X=2.04 $Y=2.3 $X2=0
+ $Y2=0
cc_214 N_A_109_297#_c_310_n N_VPWR_c_335_n 0.0165823f $X=1.37 $Y=1.98 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_335_n N_X_M1009_d 0.00382897f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_c_340_n X 0.018001f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_335_n X 0.00993603f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_218 N_X_c_382_n N_VGND_c_402_n 0.0170867f $X=3.05 $Y=0.42 $X2=0 $Y2=0
cc_219 N_X_M1003_d N_VGND_c_403_n 0.00379446f $X=2.825 $Y=0.235 $X2=0 $Y2=0
cc_220 N_X_c_382_n N_VGND_c_403_n 0.00982816f $X=3.05 $Y=0.42 $X2=0 $Y2=0
cc_221 N_VGND_c_403_n A_109_47# 0.00978874f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_222 N_VGND_c_403_n A_373_47# 0.00312992f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o22a_4.pex.spice
* Created: Thu Aug 27 14:37:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O22A_4%A_96_21# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 50 52 54 55 56 57 61 63 65 66 67 72 83
c153 61 0 6.89549e-20 $X=3.805 $Y=0.73
r154 80 81 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=1.395 $Y2=1.16
r155 72 75 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.145 $Y=1.87
+ $X2=5.145 $Y2=1.96
r156 67 70 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.385 $Y=1.87
+ $X2=3.385 $Y2=1.96
r157 64 67 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.51 $Y=1.87
+ $X2=3.385 $Y2=1.87
r158 63 72 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.02 $Y=1.87
+ $X2=5.145 $Y2=1.87
r159 63 64 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=5.02 $Y=1.87
+ $X2=3.51 $Y2=1.87
r160 59 61 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=2.965 $Y=0.775
+ $X2=3.805 $Y2=0.775
r161 57 66 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.545 $Y=0.775
+ $X2=2.415 $Y2=0.775
r162 57 59 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=2.545 $Y=0.775
+ $X2=2.965 $Y2=0.775
r163 55 67 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.26 $Y=1.87
+ $X2=3.385 $Y2=1.87
r164 55 56 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.26 $Y=1.87
+ $X2=2.23 $Y2=1.87
r165 54 66 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.23 $Y=0.82
+ $X2=2.415 $Y2=0.82
r166 52 65 3.53812 $w=3.1e-07 $l=1.09545e-07 $layer=LI1_cond $X=2.085 $Y=1.075
+ $X2=2.065 $Y2=1.175
r167 51 54 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.085 $Y=0.905
+ $X2=2.23 $Y2=0.82
r168 51 52 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.085 $Y=0.905
+ $X2=2.085 $Y2=1.075
r169 50 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.065 $Y=1.785
+ $X2=2.23 $Y2=1.87
r170 49 65 3.53812 $w=3.1e-07 $l=1e-07 $layer=LI1_cond $X=2.065 $Y=1.275
+ $X2=2.065 $Y2=1.175
r171 49 50 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.065 $Y=1.275
+ $X2=2.065 $Y2=1.785
r172 48 83 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.725 $Y=1.16
+ $X2=1.815 $Y2=1.16
r173 48 81 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.725 $Y=1.16
+ $X2=1.395 $Y2=1.16
r174 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.725
+ $Y=1.16 $X2=1.725 $Y2=1.16
r175 44 80 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.705 $Y=1.16
+ $X2=0.975 $Y2=1.16
r176 44 77 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.705 $Y=1.16
+ $X2=0.555 $Y2=1.16
r177 43 47 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=1.725 $Y2=1.175
r178 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.16 $X2=0.705 $Y2=1.16
r179 41 65 2.95888 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=1.175
+ $X2=2.065 $Y2=1.175
r180 41 47 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=1.9 $Y=1.175
+ $X2=1.725 $Y2=1.175
r181 37 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.16
r182 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.985
r183 34 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r184 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=0.56
r185 30 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.16
r186 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.985
r187 27 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=1.16
r188 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=0.56
r189 23 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.16
r190 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.985
r191 20 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=1.16
r192 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=0.56
r193 16 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.325
+ $X2=0.555 $Y2=1.16
r194 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.555 $Y=1.325
+ $X2=0.555 $Y2=1.985
r195 13 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=1.16
r196 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=0.56
r197 4 75 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.485 $X2=5.145 $Y2=1.96
r198 3 70 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=1.485 $X2=3.385 $Y2=1.96
r199 2 61 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.235 $X2=3.805 $Y2=0.73
r200 1 59 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.235 $X2=2.965 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%B1 1 3 6 8 10 13 15 19 20 22 25 26
c86 26 0 1.81811e-19 $X=2.755 $Y=1.16
r87 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.16 $X2=2.755 $Y2=1.16
r88 22 32 7.60125 $w=5.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.687 $Y=1.19
+ $X2=2.687 $Y2=1.53
r89 22 26 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=2.687 $Y=1.19
+ $X2=2.687 $Y2=1.16
r90 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.015
+ $Y=1.16 $X2=4.015 $Y2=1.16
r91 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.015 $Y=1.445
+ $X2=4.015 $Y2=1.16
r92 16 32 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=2.955 $Y=1.53
+ $X2=2.687 $Y2=1.53
r93 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.85 $Y=1.53
+ $X2=4.015 $Y2=1.445
r94 15 16 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.85 $Y=1.53
+ $X2=2.955 $Y2=1.53
r95 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.16
r96 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.985
r97 8 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=1.16
r98 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=0.56
r99 4 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.325
+ $X2=2.755 $Y2=1.16
r100 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.755 $Y=1.325
+ $X2=2.755 $Y2=1.985
r101 1 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=0.995
+ $X2=2.755 $Y2=1.16
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.755 $Y=0.995
+ $X2=2.755 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%B2 1 3 6 8 10 13 15 22
c41 6 0 1.81811e-19 $X=3.175 $Y=1.985
r42 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.385 $Y=1.16
+ $X2=3.595 $Y2=1.16
r43 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.175 $Y=1.16
+ $X2=3.385 $Y2=1.16
r44 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.16 $X2=3.385 $Y2=1.16
r45 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.325
+ $X2=3.595 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.595 $Y=1.325
+ $X2=3.595 $Y2=1.985
r47 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=0.56
r49 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=1.325
+ $X2=3.175 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.175 $Y=1.325
+ $X2=3.175 $Y2=1.985
r51 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=0.995
+ $X2=3.175 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.175 $Y=0.995
+ $X2=3.175 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%A1 1 3 6 8 10 13 17 18 20 21 23 24 25 29 33
c86 29 0 1.25382e-19 $X=5.775 $Y=1.16
c87 1 0 9.81989e-20 $X=4.515 $Y=0.995
r88 30 33 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=5.775 $Y=1.175
+ $X2=6.21 $Y2=1.175
r89 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.775
+ $Y=1.16 $X2=5.775 $Y2=1.16
r90 25 33 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=6.23 $Y=1.175 $X2=6.21
+ $Y2=1.175
r91 24 30 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=5.735 $Y=1.175
+ $X2=5.775 $Y2=1.175
r92 22 24 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.65 $Y=1.275
+ $X2=5.735 $Y2=1.175
r93 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.65 $Y=1.275
+ $X2=5.65 $Y2=1.445
r94 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.565 $Y=1.53
+ $X2=5.65 $Y2=1.445
r95 20 21 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=5.565 $Y=1.53
+ $X2=4.68 $Y2=1.53
r96 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.515
+ $Y=1.16 $X2=4.515 $Y2=1.16
r97 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.515 $Y=1.445
+ $X2=4.68 $Y2=1.53
r98 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.515 $Y=1.445
+ $X2=4.515 $Y2=1.16
r99 11 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=1.325
+ $X2=5.775 $Y2=1.16
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.775 $Y=1.325
+ $X2=5.775 $Y2=1.985
r101 8 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=0.995
+ $X2=5.775 $Y2=1.16
r102 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.775 $Y=0.995
+ $X2=5.775 $Y2=0.56
r103 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.515 $Y=1.325
+ $X2=4.515 $Y2=1.16
r104 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.515 $Y=1.325
+ $X2=4.515 $Y2=1.985
r105 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.515 $Y=0.995
+ $X2=4.515 $Y2=1.16
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.515 $Y=0.995
+ $X2=4.515 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%A2 1 3 6 8 10 13 15 22
r48 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.145 $Y=1.16
+ $X2=5.355 $Y2=1.16
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=1.16 $X2=5.145 $Y2=1.16
r50 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.935 $Y=1.16
+ $X2=5.145 $Y2=1.16
r51 15 21 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.31 $Y=1.175
+ $X2=5.145 $Y2=1.175
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=1.325
+ $X2=5.355 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.355 $Y=1.325
+ $X2=5.355 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=0.995
+ $X2=5.355 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.355 $Y=0.995
+ $X2=5.355 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.325
+ $X2=4.935 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.935 $Y=1.325
+ $X2=4.935 $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=0.995
+ $X2=4.935 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.935 $Y=0.995
+ $X2=4.935 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%VPWR 1 2 3 4 5 16 18 22 26 30 35 36 37 39 49
+ 62 63 69 74 77 79
r91 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r92 76 77 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.545 $Y=2.465
+ $X2=2.67 $Y2=2.465
r93 72 76 0.263841 $w=6.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.53 $Y=2.465
+ $X2=2.545 $Y2=2.465
r94 72 74 18.8554 $w=6.78e-07 $l=6.3e-07 $layer=LI1_cond $X=2.53 $Y=2.465
+ $X2=1.9 $Y2=2.465
r95 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r96 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r97 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r98 60 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r99 60 80 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=2.72
+ $X2=4.265 $Y2=2.72
r102 57 59 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=4.43 $Y=2.72
+ $X2=5.75 $Y2=2.72
r103 56 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r104 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r105 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 53 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 52 55 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r108 52 77 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.67 $Y2=2.72
r109 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r110 49 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=2.72
+ $X2=4.265 $Y2=2.72
r111 49 55 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.1 $Y=2.72
+ $X2=3.91 $Y2=2.72
r112 48 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r113 48 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r114 47 74 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.9 $Y2=2.72
r115 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 45 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.31 $Y=2.72
+ $X2=1.185 $Y2=2.72
r117 45 47 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.31 $Y=2.72 $X2=1.61
+ $Y2=2.72
r118 43 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r119 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 40 66 3.90382 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=0.235 $Y2=2.72
r121 40 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 39 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.06 $Y=2.72
+ $X2=1.185 $Y2=2.72
r123 39 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 37 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 37 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 35 59 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.75 $Y2=2.72
r127 35 36 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=6.007 $Y2=2.72
r128 34 62 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.11 $Y=2.72 $X2=6.21
+ $Y2=2.72
r129 34 36 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=6.11 $Y=2.72
+ $X2=6.007 $Y2=2.72
r130 30 33 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.007 $Y=1.62
+ $X2=6.007 $Y2=2.3
r131 28 36 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.007 $Y=2.635
+ $X2=6.007 $Y2=2.72
r132 28 33 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=6.007 $Y=2.635
+ $X2=6.007 $Y2=2.3
r133 24 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=2.635
+ $X2=4.265 $Y2=2.72
r134 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.265 $Y=2.635
+ $X2=4.265 $Y2=2.3
r135 20 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=2.72
r136 20 22 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=1.99
r137 16 66 3.23934 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.235 $Y2=2.72
r138 16 18 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.345 $Y2=1.99
r139 5 33 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=1.485 $X2=5.99 $Y2=2.3
r140 5 30 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=1.485 $X2=5.99 $Y2=1.62
r141 4 26 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=1.485 $X2=4.225 $Y2=2.3
r142 3 76 300 $w=1.7e-07 $l=1.09455e-06 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=1.485 $X2=2.545 $Y2=2.3
r143 2 22 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.485 $X2=1.185 $Y2=1.99
r144 1 18 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=1.485 $X2=0.345 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43 44
+ 45
r73 42 45 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.227 $Y=1.445
+ $X2=0.227 $Y2=1.19
r74 41 45 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=0.227 $Y=0.905
+ $X2=0.227 $Y2=1.19
r75 37 39 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=1.62
+ $X2=1.605 $Y2=2.3
r76 35 37 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=1.615
+ $X2=1.605 $Y2=1.62
r77 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.605 $Y=0.725
+ $X2=1.605 $Y2=0.39
r78 30 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=0.815
+ $X2=0.765 $Y2=0.815
r79 29 31 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.44 $Y=0.815
+ $X2=1.605 $Y2=0.725
r80 29 30 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.44 $Y=0.815
+ $X2=0.93 $Y2=0.815
r81 28 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.89 $Y=1.53
+ $X2=0.765 $Y2=1.53
r82 27 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.48 $Y=1.53
+ $X2=1.605 $Y2=1.615
r83 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.48 $Y=1.53 $X2=0.89
+ $Y2=1.53
r84 23 25 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.765 $Y=1.62
+ $X2=0.765 $Y2=2.3
r85 21 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.615
+ $X2=0.765 $Y2=1.53
r86 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.765 $Y=1.615
+ $X2=0.765 $Y2=1.62
r87 17 43 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.765 $Y=0.725
+ $X2=0.765 $Y2=0.815
r88 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.765 $Y=0.725
+ $X2=0.765 $Y2=0.39
r89 16 42 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.37 $Y=1.53
+ $X2=0.227 $Y2=1.445
r90 15 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.64 $Y=1.53
+ $X2=0.765 $Y2=1.53
r91 15 16 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.64 $Y=1.53 $X2=0.37
+ $Y2=1.53
r92 14 41 7.27854 $w=1.8e-07 $l=1.82535e-07 $layer=LI1_cond $X=0.37 $Y=0.815
+ $X2=0.227 $Y2=0.905
r93 13 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=0.815
+ $X2=0.765 $Y2=0.815
r94 13 14 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.6 $Y=0.815
+ $X2=0.37 $Y2=0.815
r95 4 39 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.485 $X2=1.605 $Y2=2.3
r96 4 37 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.485 $X2=1.605 $Y2=1.62
r97 3 25 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.485 $X2=0.765 $Y2=2.3
r98 3 23 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.485 $X2=0.765 $Y2=1.62
r99 2 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.47
+ $Y=0.235 $X2=1.605 $Y2=0.39
r100 1 19 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.235 $X2=0.765 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%A_566_297# 1 2 7 10 15
r21 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.805 $Y=2.3 $X2=3.805
+ $Y2=2.38
r22 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.965 $Y=2.3 $X2=2.965
+ $Y2=2.38
r23 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=2.38
+ $X2=2.965 $Y2=2.38
r24 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.68 $Y=2.38
+ $X2=3.805 $Y2=2.38
r25 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.68 $Y=2.38 $X2=3.09
+ $Y2=2.38
r26 2 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.485 $X2=3.805 $Y2=2.3
r27 1 10 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.485 $X2=2.965 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%A_918_297# 1 2 7 11 14
c17 11 0 1.25382e-19 $X=5.565 $Y=1.96
r18 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.725 $Y=2.3 $X2=4.725
+ $Y2=2.38
r19 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.565 $Y=2.295
+ $X2=5.565 $Y2=1.96
r20 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=2.38
+ $X2=4.725 $Y2=2.38
r21 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.44 $Y=2.38
+ $X2=5.565 $Y2=2.295
r22 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.44 $Y=2.38 $X2=4.85
+ $Y2=2.38
r23 2 11 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.43
+ $Y=1.485 $X2=5.565 $Y2=1.96
r24 1 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=1.485 $X2=4.725 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%VGND 1 2 3 4 5 18 20 21 24 28 32 36 39 40 42
+ 43 44 46 59 60 68 71
r100 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r101 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r102 63 66 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.345 $Y2=0
r103 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r104 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r105 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r106 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r107 54 72 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=2.07
+ $Y2=0
r108 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r109 51 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.025
+ $Y2=0
r110 51 53 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=2.11 $Y=0 $X2=4.37
+ $Y2=0
r111 50 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r112 50 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r113 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r114 47 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.185
+ $Y2=0
r115 47 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.61
+ $Y2=0
r116 46 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.025
+ $Y2=0
r117 46 49 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.61
+ $Y2=0
r118 44 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r119 44 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 42 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.48 $Y=0 $X2=5.29
+ $Y2=0
r121 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0 $X2=5.565
+ $Y2=0
r122 41 59 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.65 $Y=0 $X2=6.21
+ $Y2=0
r123 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=0 $X2=5.565
+ $Y2=0
r124 39 53 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.37
+ $Y2=0
r125 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.725
+ $Y2=0
r126 38 56 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.81 $Y=0 $X2=5.29
+ $Y2=0
r127 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=0 $X2=4.725
+ $Y2=0
r128 34 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.085
+ $X2=5.565 $Y2=0
r129 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.565 $Y=0.085
+ $X2=5.565 $Y2=0.39
r130 30 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=0.085
+ $X2=4.725 $Y2=0
r131 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.725 $Y=0.085
+ $X2=4.725 $Y2=0.39
r132 26 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r133 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.39
r134 22 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r135 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.39
r136 21 66 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.345
+ $Y2=0
r137 20 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0 $X2=1.185
+ $Y2=0
r138 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=0.43
+ $Y2=0
r139 16 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0
r140 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.39
r141 5 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.235 $X2=5.565 $Y2=0.39
r142 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.59
+ $Y=0.235 $X2=4.725 $Y2=0.39
r143 3 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.235 $X2=2.025 $Y2=0.39
r144 2 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.235 $X2=1.185 $Y2=0.39
r145 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.345 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_4%A_484_47# 1 2 3 4 5 16 22 25 26 27 30 32 36
+ 40
c75 40 0 2.9244e-20 $X=5.145 $Y=0.815
r76 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.985 $Y=0.725
+ $X2=5.985 $Y2=0.39
r77 33 40 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=5.31 $Y=0.815
+ $X2=5.145 $Y2=0.815
r78 32 34 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.82 $Y=0.815
+ $X2=5.985 $Y2=0.725
r79 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.82 $Y=0.815
+ $X2=5.31 $Y2=0.815
r80 28 40 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.145 $Y=0.725
+ $X2=5.145 $Y2=0.815
r81 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.145 $Y=0.725
+ $X2=5.145 $Y2=0.39
r82 26 40 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.98 $Y=0.82
+ $X2=5.145 $Y2=0.815
r83 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.98 $Y=0.82
+ $X2=4.47 $Y2=0.82
r84 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.305 $Y=0.735
+ $X2=4.47 $Y2=0.82
r85 23 25 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.305 $Y=0.735
+ $X2=4.305 $Y2=0.73
r86 22 39 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.305 $Y=0.475
+ $X2=4.305 $Y2=0.365
r87 22 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=0.475
+ $X2=4.305 $Y2=0.73
r88 18 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=2.545 $Y=0.365
+ $X2=3.385 $Y2=0.365
r89 16 39 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0.365
+ $X2=4.305 $Y2=0.365
r90 16 21 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=4.14 $Y=0.365
+ $X2=3.385 $Y2=0.365
r91 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.85
+ $Y=0.235 $X2=5.985 $Y2=0.39
r92 4 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.01
+ $Y=0.235 $X2=5.145 $Y2=0.39
r93 3 39 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.235 $X2=4.27 $Y2=0.39
r94 3 25 182 $w=1.7e-07 $l=5.78035e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.235 $X2=4.27 $Y2=0.73
r95 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.235 $X2=3.385 $Y2=0.39
r96 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.235 $X2=2.545 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__o32ai_4.spice.SKY130_FD_SC_HD__O32AI_4.pxi
* Created: Thu Aug 27 14:41:33 2020
* 
x_PM_SKY130_FD_SC_HD__O32AI_4%B2 N_B2_M1013_g N_B2_M1004_g N_B2_M1022_g
+ N_B2_M1006_g N_B2_M1023_g N_B2_M1025_g N_B2_M1035_g N_B2_M1034_g B2 B2 B2
+ N_B2_c_129_n N_B2_c_130_n PM_SKY130_FD_SC_HD__O32AI_4%B2
x_PM_SKY130_FD_SC_HD__O32AI_4%B1 N_B1_M1024_g N_B1_M1008_g N_B1_M1031_g
+ N_B1_M1011_g N_B1_M1036_g N_B1_M1012_g N_B1_M1038_g N_B1_M1029_g B1 B1 B1
+ N_B1_c_199_n PM_SKY130_FD_SC_HD__O32AI_4%B1
x_PM_SKY130_FD_SC_HD__O32AI_4%A3 N_A3_M1002_g N_A3_M1003_g N_A3_M1000_g
+ N_A3_M1027_g N_A3_M1007_g N_A3_M1014_g N_A3_M1037_g N_A3_M1030_g A3 A3 A3 A3
+ N_A3_c_264_n PM_SKY130_FD_SC_HD__O32AI_4%A3
x_PM_SKY130_FD_SC_HD__O32AI_4%A2 N_A2_M1009_g N_A2_M1015_g N_A2_M1016_g
+ N_A2_M1021_g N_A2_M1019_g N_A2_M1033_g N_A2_M1028_g N_A2_M1039_g A2 A2 A2
+ N_A2_c_349_n PM_SKY130_FD_SC_HD__O32AI_4%A2
x_PM_SKY130_FD_SC_HD__O32AI_4%A1 N_A1_M1010_g N_A1_M1001_g N_A1_M1017_g
+ N_A1_M1005_g N_A1_M1018_g N_A1_M1026_g N_A1_c_424_n N_A1_c_425_n N_A1_M1020_g
+ N_A1_M1032_g A1 A1 A1 A1 N_A1_c_428_n A1 PM_SKY130_FD_SC_HD__O32AI_4%A1
x_PM_SKY130_FD_SC_HD__O32AI_4%A_27_297# N_A_27_297#_M1004_s N_A_27_297#_M1006_s
+ N_A_27_297#_M1034_s N_A_27_297#_M1011_d N_A_27_297#_M1029_d
+ N_A_27_297#_c_502_n N_A_27_297#_c_503_n N_A_27_297#_c_508_n
+ N_A_27_297#_c_521_p N_A_27_297#_c_510_n N_A_27_297#_c_534_p
+ N_A_27_297#_c_513_n N_A_27_297#_c_512_n N_A_27_297#_c_546_p
+ N_A_27_297#_c_515_n N_A_27_297#_c_504_n N_A_27_297#_c_505_n
+ N_A_27_297#_c_544_p N_A_27_297#_c_529_p PM_SKY130_FD_SC_HD__O32AI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__O32AI_4%Y N_Y_M1013_s N_Y_M1023_s N_Y_M1024_s N_Y_M1036_s
+ N_Y_M1004_d N_Y_M1025_d N_Y_M1000_s N_Y_M1014_s N_Y_c_567_n N_Y_c_578_n
+ N_Y_c_568_n N_Y_c_569_n N_Y_c_571_n N_Y_c_584_n N_Y_c_613_n N_Y_c_587_n
+ N_Y_c_666_p N_Y_c_617_n N_Y_c_622_n Y PM_SKY130_FD_SC_HD__O32AI_4%Y
x_PM_SKY130_FD_SC_HD__O32AI_4%VPWR N_VPWR_M1008_s N_VPWR_M1012_s N_VPWR_M1001_d
+ N_VPWR_M1005_d N_VPWR_M1032_d N_VPWR_c_684_n N_VPWR_c_685_n N_VPWR_c_686_n
+ N_VPWR_c_687_n N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_690_n N_VPWR_c_691_n
+ N_VPWR_c_692_n N_VPWR_c_693_n N_VPWR_c_694_n N_VPWR_c_695_n N_VPWR_c_696_n
+ N_VPWR_c_697_n VPWR N_VPWR_c_698_n N_VPWR_c_683_n
+ PM_SKY130_FD_SC_HD__O32AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O32AI_4%A_806_297# N_A_806_297#_M1000_d
+ N_A_806_297#_M1007_d N_A_806_297#_M1030_d N_A_806_297#_M1021_d
+ N_A_806_297#_M1039_d N_A_806_297#_c_827_n N_A_806_297#_c_828_n
+ N_A_806_297#_c_831_n N_A_806_297#_c_849_n N_A_806_297#_c_833_n
+ N_A_806_297#_c_835_n N_A_806_297#_c_882_p N_A_806_297#_c_837_n
+ N_A_806_297#_c_829_n N_A_806_297#_c_830_n N_A_806_297#_c_872_n
+ N_A_806_297#_c_874_n N_A_806_297#_c_876_n
+ PM_SKY130_FD_SC_HD__O32AI_4%A_806_297#
x_PM_SKY130_FD_SC_HD__O32AI_4%A_1224_297# N_A_1224_297#_M1015_s
+ N_A_1224_297#_M1033_s N_A_1224_297#_M1001_s N_A_1224_297#_M1026_s
+ N_A_1224_297#_c_891_n N_A_1224_297#_c_889_n N_A_1224_297#_c_907_n
+ N_A_1224_297#_c_910_n N_A_1224_297#_c_914_n N_A_1224_297#_c_918_n
+ N_A_1224_297#_c_890_n N_A_1224_297#_c_901_n N_A_1224_297#_c_921_n
+ PM_SKY130_FD_SC_HD__O32AI_4%A_1224_297#
x_PM_SKY130_FD_SC_HD__O32AI_4%A_27_47# N_A_27_47#_M1013_d N_A_27_47#_M1022_d
+ N_A_27_47#_M1035_d N_A_27_47#_M1031_d N_A_27_47#_M1038_d N_A_27_47#_M1003_s
+ N_A_27_47#_M1037_s N_A_27_47#_M1016_s N_A_27_47#_M1028_s N_A_27_47#_M1017_s
+ N_A_27_47#_M1020_s N_A_27_47#_c_952_n N_A_27_47#_c_953_n N_A_27_47#_c_970_n
+ N_A_27_47#_c_980_n N_A_27_47#_c_954_n N_A_27_47#_c_955_n N_A_27_47#_c_988_n
+ N_A_27_47#_c_956_n N_A_27_47#_c_1007_n N_A_27_47#_c_957_n N_A_27_47#_c_1027_n
+ N_A_27_47#_c_958_n N_A_27_47#_c_959_n N_A_27_47#_c_960_n N_A_27_47#_c_961_n
+ N_A_27_47#_c_962_n N_A_27_47#_c_963_n N_A_27_47#_c_964_n N_A_27_47#_c_965_n
+ N_A_27_47#_c_966_n PM_SKY130_FD_SC_HD__O32AI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O32AI_4%VGND N_VGND_M1002_d N_VGND_M1027_d N_VGND_M1009_d
+ N_VGND_M1019_d N_VGND_M1010_d N_VGND_M1018_d N_VGND_c_1118_n N_VGND_c_1119_n
+ N_VGND_c_1120_n N_VGND_c_1121_n N_VGND_c_1122_n N_VGND_c_1123_n
+ N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n
+ N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n VGND N_VGND_c_1131_n
+ N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n
+ N_VGND_c_1136_n N_VGND_c_1137_n PM_SKY130_FD_SC_HD__O32AI_4%VGND
cc_1 VNB N_B2_M1013_g 0.0229701f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_B2_M1022_g 0.0168049f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_B2_M1023_g 0.0167831f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_4 VNB N_B2_M1035_g 0.0171462f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_5 VNB N_B2_c_129_n 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.16
cc_6 VNB N_B2_c_130_n 0.0818978f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_7 VNB N_B1_M1024_g 0.0171464f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_8 VNB N_B1_M1031_g 0.0167833f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_9 VNB N_B1_M1036_g 0.0168049f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_10 VNB N_B1_M1038_g 0.0171822f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_11 VNB B1 0.00242518f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_12 VNB N_B1_c_199_n 0.0597713f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_13 VNB N_A3_M1002_g 0.0170334f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_14 VNB N_A3_M1003_g 0.0168007f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_A3_M1027_g 0.0183205f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_16 VNB N_A3_M1037_g 0.0213409f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_17 VNB A3 0.00140887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A3_c_264_n 0.0889036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_M1009_g 0.0198211f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_A2_M1016_g 0.0168007f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_21 VNB N_A2_M1019_g 0.0168007f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_22 VNB N_A2_M1028_g 0.023095f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_23 VNB N_A2_c_349_n 0.0713692f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_24 VNB N_A1_M1010_g 0.023095f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_25 VNB N_A1_M1017_g 0.0168007f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_26 VNB N_A1_M1018_g 0.0177544f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_27 VNB N_A1_c_424_n 0.0154558f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.015
cc_28 VNB N_A1_c_425_n 0.0506654f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_29 VNB N_A1_M1020_g 0.0240303f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.305
cc_30 VNB A1 0.0110416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A1_c_428_n 0.0264065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_567_n 0.00727592f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.015
cc_33 VNB N_Y_c_568_n 0.00727175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_569_n 0.007346f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_35 VNB N_VPWR_c_683_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_952_n 0.00922242f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_37 VNB N_A_27_47#_c_953_n 0.0184482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_954_n 0.00368718f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.16
cc_39 VNB N_A_27_47#_c_955_n 0.00218177f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.16
cc_40 VNB N_A_27_47#_c_956_n 0.00218177f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.175
cc_41 VNB N_A_27_47#_c_957_n 0.00421299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_958_n 0.0129648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_959_n 0.0206947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_27_47#_c_960_n 0.00222843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_27_47#_c_961_n 0.00314926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_27_47#_c_962_n 0.0145559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_27_47#_c_963_n 0.00222843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_27_47#_c_964_n 0.00218177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_27_47#_c_965_n 0.011017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_27_47#_c_966_n 0.00222843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1118_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.305
cc_52 VNB N_VGND_c_1119_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_53 VNB N_VGND_c_1120_n 0.00499469f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_54 VNB N_VGND_c_1121_n 0.00415222f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_55 VNB N_VGND_c_1122_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_56 VNB N_VGND_c_1123_n 0.00415222f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_57 VNB N_VGND_c_1124_n 0.00463836f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_58 VNB N_VGND_c_1125_n 0.0918935f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_59 VNB N_VGND_c_1126_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.16
cc_60 VNB N_VGND_c_1127_n 0.0294016f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.16
cc_61 VNB N_VGND_c_1128_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_62 VNB N_VGND_c_1129_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_63 VNB N_VGND_c_1130_n 0.00496831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1131_n 0.0248982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1132_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1133_n 0.0184038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1134_n 0.467574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1135_n 0.00631235f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1136_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1137_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VPB N_B2_M1004_g 0.0275854f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_72 VPB N_B2_M1006_g 0.0195069f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_73 VPB N_B2_M1025_g 0.0194992f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_74 VPB N_B2_M1034_g 0.0199889f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_75 VPB N_B2_c_130_n 0.0147273f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_76 VPB N_B1_M1008_g 0.0197621f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_77 VPB N_B1_M1011_g 0.0192722f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_78 VPB N_B1_M1012_g 0.0192797f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_79 VPB N_B1_M1029_g 0.0273582f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_80 VPB N_B1_c_199_n 0.00651607f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_81 VPB N_A3_M1000_g 0.0275854f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_82 VPB N_A3_M1007_g 0.0195069f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_83 VPB N_A3_M1014_g 0.0195069f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_84 VPB N_A3_M1030_g 0.0198722f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_85 VPB N_A3_c_264_n 0.0202847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A2_M1015_g 0.0198722f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_87 VPB N_A2_M1021_g 0.0195069f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_88 VPB N_A2_M1033_g 0.0195069f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_89 VPB N_A2_M1039_g 0.0275854f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_90 VPB N_A2_c_349_n 0.00651342f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_91 VPB N_A1_M1001_g 0.0275854f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_92 VPB N_A1_M1005_g 0.0195069f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_93 VPB N_A1_M1026_g 0.0206539f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_94 VPB N_A1_c_424_n 0.00446199f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.015
cc_95 VPB N_A1_c_425_n 0.00434272f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_96 VPB N_A1_M1032_g 0.0277543f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_97 VPB N_A1_c_428_n 0.00494437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_27_297#_c_502_n 0.00922995f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_297#_c_503_n 0.0291185f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_100 VPB N_A_27_297#_c_504_n 0.00184354f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_101 VPB N_A_27_297#_c_505_n 0.0043399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_Y_c_568_n 0.00333735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_Y_c_571_n 0.0108306f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_104 VPB N_VPWR_c_684_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_105 VPB N_VPWR_c_685_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_106 VPB N_VPWR_c_686_n 0.0108453f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_107 VPB N_VPWR_c_687_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_108 VPB N_VPWR_c_688_n 0.011345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_689_n 0.0454352f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_110 VPB N_VPWR_c_690_n 0.0519394f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_111 VPB N_VPWR_c_691_n 0.00436611f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_112 VPB N_VPWR_c_692_n 0.0113044f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_693_n 0.00436611f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_114 VPB N_VPWR_c_694_n 0.103099f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_115 VPB N_VPWR_c_695_n 0.00477947f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_116 VPB N_VPWR_c_696_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_117 VPB N_VPWR_c_697_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_118 VPB N_VPWR_c_698_n 0.0169988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_683_n 0.0610369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_806_297#_c_827_n 0.00217929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_806_297#_c_828_n 0.00399114f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_122 VPB N_A_806_297#_c_829_n 0.00217929f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_123 VPB N_A_806_297#_c_830_n 0.00408452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_1224_297#_c_889_n 0.0132401f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_125 N_B2_M1035_g N_B1_M1024_g 0.0252948f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_126 N_B2_M1034_g N_B1_M1008_g 0.0252948f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B2_c_130_n N_B1_c_199_n 0.0252948f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B2_c_129_n N_A_27_297#_c_503_n 0.0151342f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B2_c_130_n N_A_27_297#_c_503_n 0.00534919f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B2_M1004_g N_A_27_297#_c_508_n 0.0124471f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B2_M1006_g N_A_27_297#_c_508_n 0.0102593f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B2_M1025_g N_A_27_297#_c_510_n 0.0102319f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_133 N_B2_M1034_g N_A_27_297#_c_510_n 0.0110304f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_134 N_B2_M1034_g N_A_27_297#_c_512_n 0.0012299f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B2_M1013_g N_Y_c_567_n 0.00378792f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_136 N_B2_M1022_g N_Y_c_567_n 0.0108206f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_137 N_B2_M1023_g N_Y_c_567_n 0.0108206f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_138 N_B2_M1035_g N_Y_c_567_n 0.0123906f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_139 N_B2_c_129_n N_Y_c_567_n 0.0859305f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B2_c_130_n N_Y_c_567_n 0.00639054f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B2_M1006_g N_Y_c_578_n 0.00891221f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B2_M1025_g N_Y_c_578_n 0.00891221f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B2_c_129_n N_Y_c_578_n 0.0412785f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B2_c_130_n N_Y_c_578_n 0.00197018f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B2_M1035_g N_Y_c_568_n 0.0112495f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_146 N_B2_c_129_n N_Y_c_568_n 0.0158866f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B2_M1025_g N_Y_c_584_n 0.0010018f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B2_M1034_g N_Y_c_584_n 0.0109782f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B2_c_130_n N_Y_c_584_n 0.00197018f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_150 N_B2_M1004_g N_Y_c_587_n 0.00734464f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B2_M1006_g N_Y_c_587_n 0.00687399f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B2_M1025_g N_Y_c_587_n 5.07492e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B2_c_129_n N_Y_c_587_n 0.0169697f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B2_c_130_n N_Y_c_587_n 0.00205111f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B2_M1006_g Y 5.08048e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B2_M1025_g Y 0.00604703f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B2_M1034_g Y 0.00697479f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_158 N_B2_M1034_g N_VPWR_c_684_n 0.00122467f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B2_M1004_g N_VPWR_c_690_n 0.00357877f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B2_M1006_g N_VPWR_c_690_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B2_M1025_g N_VPWR_c_690_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_162 N_B2_M1034_g N_VPWR_c_690_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_163 N_B2_M1004_g N_VPWR_c_683_n 0.00617937f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_B2_M1006_g N_VPWR_c_683_n 0.00522516f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B2_M1025_g N_VPWR_c_683_n 0.00522516f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_166 N_B2_M1034_g N_VPWR_c_683_n 0.0053303f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_167 N_B2_M1013_g N_A_27_47#_c_953_n 4.62114e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_168 N_B2_c_129_n N_A_27_47#_c_953_n 0.0190063f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B2_c_130_n N_A_27_47#_c_953_n 0.00569691f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B2_M1013_g N_A_27_47#_c_970_n 0.0103559f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_171 N_B2_M1022_g N_A_27_47#_c_970_n 0.00878931f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_172 N_B2_M1023_g N_A_27_47#_c_970_n 0.00878931f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_173 N_B2_M1035_g N_A_27_47#_c_970_n 0.00878931f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_174 N_B2_c_129_n N_A_27_47#_c_970_n 0.00349599f $X=1.52 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B2_M1013_g N_VGND_c_1125_n 0.00357877f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_176 N_B2_M1022_g N_VGND_c_1125_n 0.00357877f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_177 N_B2_M1023_g N_VGND_c_1125_n 0.00357877f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_178 N_B2_M1035_g N_VGND_c_1125_n 0.00357877f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_179 N_B2_M1013_g N_VGND_c_1134_n 0.00617937f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_180 N_B2_M1022_g N_VGND_c_1134_n 0.00522516f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_181 N_B2_M1023_g N_VGND_c_1134_n 0.00522516f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_182 N_B2_M1035_g N_VGND_c_1134_n 0.00528897f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_183 N_B1_M1038_g N_A3_M1002_g 0.0144883f $X=3.425 $Y=0.56 $X2=0 $Y2=0
cc_184 B1 A3 0.0140536f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_185 N_B1_c_199_n A3 2.32892e-19 $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_186 B1 N_A3_c_264_n 8.49417e-19 $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_187 N_B1_c_199_n N_A3_c_264_n 0.0144883f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B1_M1008_g N_A_27_297#_c_513_n 0.0110101f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B1_M1011_g N_A_27_297#_c_513_n 0.00967544f $X=2.585 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_B1_M1012_g N_A_27_297#_c_515_n 0.00971959f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_B1_M1029_g N_A_27_297#_c_515_n 0.00971959f $X=3.425 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_B1_M1024_g N_Y_c_568_n 0.01117f $X=2.165 $Y=0.56 $X2=0 $Y2=0
cc_193 B1 N_Y_c_568_n 0.0158867f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_194 N_B1_M1024_g N_Y_c_569_n 0.012328f $X=2.165 $Y=0.56 $X2=0 $Y2=0
cc_195 N_B1_M1031_g N_Y_c_569_n 0.0108206f $X=2.585 $Y=0.56 $X2=0 $Y2=0
cc_196 N_B1_M1036_g N_Y_c_569_n 0.0108206f $X=3.005 $Y=0.56 $X2=0 $Y2=0
cc_197 N_B1_M1038_g N_Y_c_569_n 0.0036445f $X=3.425 $Y=0.56 $X2=0 $Y2=0
cc_198 B1 N_Y_c_569_n 0.0862841f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_199 N_B1_c_199_n N_Y_c_569_n 0.00639054f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B1_M1008_g N_Y_c_571_n 0.01195f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B1_M1011_g N_Y_c_571_n 0.0106666f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B1_M1012_g N_Y_c_571_n 0.0106666f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_M1029_g N_Y_c_571_n 0.0127696f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_204 B1 N_Y_c_571_n 0.0653269f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_205 N_B1_c_199_n N_Y_c_571_n 0.00591053f $X=3.425 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B1_M1008_g Y 9.76831e-19 $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1008_g N_VPWR_c_684_n 0.0086771f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_M1011_g N_VPWR_c_684_n 0.00775986f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1012_g N_VPWR_c_684_n 6.13129e-19 $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1011_g N_VPWR_c_685_n 6.13129e-19 $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1012_g N_VPWR_c_685_n 0.00775986f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1029_g N_VPWR_c_685_n 0.00922945f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1008_g N_VPWR_c_690_n 0.00348405f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1011_g N_VPWR_c_692_n 0.00348405f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1012_g N_VPWR_c_692_n 0.00348405f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_M1029_g N_VPWR_c_694_n 0.00348405f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B1_M1008_g N_VPWR_c_683_n 0.00421182f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_M1011_g N_VPWR_c_683_n 0.00414556f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B1_M1012_g N_VPWR_c_683_n 0.00414556f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B1_M1029_g N_VPWR_c_683_n 0.00552264f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B1_M1024_g N_A_27_47#_c_970_n 0.00878931f $X=2.165 $Y=0.56 $X2=0 $Y2=0
cc_222 N_B1_M1031_g N_A_27_47#_c_970_n 0.00878931f $X=2.585 $Y=0.56 $X2=0 $Y2=0
cc_223 N_B1_M1036_g N_A_27_47#_c_970_n 0.00878931f $X=3.005 $Y=0.56 $X2=0 $Y2=0
cc_224 N_B1_M1038_g N_A_27_47#_c_970_n 0.0103559f $X=3.425 $Y=0.56 $X2=0 $Y2=0
cc_225 B1 N_A_27_47#_c_970_n 0.0035277f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_226 N_B1_M1024_g N_VGND_c_1125_n 0.00357877f $X=2.165 $Y=0.56 $X2=0 $Y2=0
cc_227 N_B1_M1031_g N_VGND_c_1125_n 0.00357877f $X=2.585 $Y=0.56 $X2=0 $Y2=0
cc_228 N_B1_M1036_g N_VGND_c_1125_n 0.00357877f $X=3.005 $Y=0.56 $X2=0 $Y2=0
cc_229 N_B1_M1038_g N_VGND_c_1125_n 0.00357877f $X=3.425 $Y=0.56 $X2=0 $Y2=0
cc_230 N_B1_M1024_g N_VGND_c_1134_n 0.00528897f $X=2.165 $Y=0.56 $X2=0 $Y2=0
cc_231 N_B1_M1031_g N_VGND_c_1134_n 0.00522516f $X=2.585 $Y=0.56 $X2=0 $Y2=0
cc_232 N_B1_M1036_g N_VGND_c_1134_n 0.00522516f $X=3.005 $Y=0.56 $X2=0 $Y2=0
cc_233 N_B1_M1038_g N_VGND_c_1134_n 0.00525237f $X=3.425 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A3_M1037_g N_A2_M1009_g 0.00519413f $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_235 N_A3_M1030_g N_A2_M1015_g 0.0234554f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A3_c_264_n A2 0.00115296f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_237 A3 N_A2_c_349_n 8.14015e-19 $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_238 N_A3_c_264_n N_A2_c_349_n 0.0234554f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A3_M1000_g N_Y_c_571_n 0.0110152f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_240 A3 N_Y_c_571_n 0.0356382f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_241 N_A3_c_264_n N_Y_c_571_n 0.0131362f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A3_M1007_g N_Y_c_613_n 0.00891221f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A3_M1014_g N_Y_c_613_n 0.00891221f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_244 A3 N_Y_c_613_n 0.025666f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_245 N_A3_c_264_n N_Y_c_613_n 0.00197018f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A3_M1000_g N_Y_c_617_n 0.0114674f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A3_M1007_g N_Y_c_617_n 0.00687399f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A3_M1014_g N_Y_c_617_n 5.07492e-19 $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_249 A3 N_Y_c_617_n 0.0169697f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_250 N_A3_c_264_n N_Y_c_617_n 0.00245031f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A3_M1007_g N_Y_c_622_n 5.07492e-19 $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A3_M1014_g N_Y_c_622_n 0.00687399f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A3_M1030_g N_Y_c_622_n 0.00958948f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_254 A3 N_Y_c_622_n 0.0062218f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_255 N_A3_c_264_n N_Y_c_622_n 0.00243034f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A3_M1000_g N_VPWR_c_694_n 0.00357877f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A3_M1007_g N_VPWR_c_694_n 0.00357877f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A3_M1014_g N_VPWR_c_694_n 0.00357877f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A3_M1030_g N_VPWR_c_694_n 0.00357877f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A3_M1000_g N_VPWR_c_683_n 0.00655123f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A3_M1007_g N_VPWR_c_683_n 0.00522516f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A3_M1014_g N_VPWR_c_683_n 0.00522516f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A3_M1030_g N_VPWR_c_683_n 0.00525237f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A3_M1000_g N_A_806_297#_c_831_n 0.0102593f $X=4.365 $Y=1.985 $X2=0
+ $Y2=0
cc_265 N_A3_M1007_g N_A_806_297#_c_831_n 0.0102593f $X=4.785 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_A3_M1014_g N_A_806_297#_c_833_n 0.0102593f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_A3_M1030_g N_A_806_297#_c_833_n 0.0124471f $X=5.625 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A3_M1030_g N_A_1224_297#_c_890_n 0.00100442f $X=5.625 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A3_M1002_g N_A_27_47#_c_980_n 0.00244813f $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_270 N_A3_M1002_g N_A_27_47#_c_954_n 0.00517044f $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_271 N_A3_M1003_g N_A_27_47#_c_954_n 5.17008e-19 $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_272 A3 N_A_27_47#_c_954_n 0.00230247f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_273 N_A3_M1002_g N_A_27_47#_c_955_n 0.00850187f $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A3_M1003_g N_A_27_47#_c_955_n 0.00845772f $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_275 A3 N_A_27_47#_c_955_n 0.0359511f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_276 N_A3_c_264_n N_A_27_47#_c_955_n 0.00210947f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A3_M1002_g N_A_27_47#_c_988_n 5.77985e-19 $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A3_M1003_g N_A_27_47#_c_988_n 0.00655349f $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A3_M1027_g N_A_27_47#_c_988_n 0.00724486f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A3_M1037_g N_A_27_47#_c_988_n 6.55335e-19 $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A3_M1003_g N_A_27_47#_c_960_n 0.00110555f $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A3_M1027_g N_A_27_47#_c_960_n 0.00110555f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_283 A3 N_A_27_47#_c_960_n 0.0265407f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_284 N_A3_c_264_n N_A_27_47#_c_960_n 0.00262649f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A3_M1027_g N_A_27_47#_c_961_n 0.00932519f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A3_M1037_g N_A_27_47#_c_961_n 0.00932519f $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_287 A3 N_A_27_47#_c_961_n 0.0530561f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_288 N_A3_c_264_n N_A_27_47#_c_961_n 0.00663278f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A3_M1027_g N_A_27_47#_c_962_n 6.53424e-19 $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A3_M1037_g N_A_27_47#_c_962_n 0.00855266f $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A3_c_264_n N_A_27_47#_c_962_n 0.0139698f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A3_M1002_g N_VGND_c_1118_n 0.00268723f $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A3_M1003_g N_VGND_c_1118_n 0.00146448f $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A3_M1003_g N_VGND_c_1119_n 0.00424416f $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_295 N_A3_M1027_g N_VGND_c_1119_n 0.00424416f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_296 N_A3_M1027_g N_VGND_c_1120_n 0.00367224f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A3_M1037_g N_VGND_c_1120_n 0.00499979f $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A3_M1002_g N_VGND_c_1125_n 0.00422898f $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A3_M1037_g N_VGND_c_1131_n 0.0042294f $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_300 N_A3_M1002_g N_VGND_c_1134_n 0.00577235f $X=3.845 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A3_M1003_g N_VGND_c_1134_n 0.00573607f $X=4.265 $Y=0.56 $X2=0 $Y2=0
cc_302 N_A3_M1027_g N_VGND_c_1134_n 0.00616144f $X=4.685 $Y=0.56 $X2=0 $Y2=0
cc_303 N_A3_M1037_g N_VGND_c_1134_n 0.00685106f $X=5.265 $Y=0.56 $X2=0 $Y2=0
cc_304 N_A2_M1015_g N_Y_c_622_n 0.00100442f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A2_M1039_g N_VPWR_c_686_n 0.00229957f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A2_M1015_g N_VPWR_c_694_n 0.00357877f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A2_M1021_g N_VPWR_c_694_n 0.00357877f $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A2_M1033_g N_VPWR_c_694_n 0.00357877f $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A2_M1039_g N_VPWR_c_694_n 0.00357877f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A2_M1015_g N_VPWR_c_683_n 0.00525237f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A2_M1021_g N_VPWR_c_683_n 0.00522516f $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A2_M1033_g N_VPWR_c_683_n 0.00522516f $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A2_M1039_g N_VPWR_c_683_n 0.00655123f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A2_M1015_g N_A_806_297#_c_835_n 0.0124471f $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A2_M1021_g N_A_806_297#_c_835_n 0.0102593f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A2_M1033_g N_A_806_297#_c_837_n 0.0102593f $X=6.885 $Y=1.985 $X2=0
+ $Y2=0
cc_317 N_A2_M1039_g N_A_806_297#_c_837_n 0.0102593f $X=7.305 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A2_M1021_g N_A_1224_297#_c_891_n 0.00891221f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_319 N_A2_M1033_g N_A_1224_297#_c_891_n 0.00891221f $X=6.885 $Y=1.985 $X2=0
+ $Y2=0
cc_320 A2 N_A_1224_297#_c_891_n 0.025666f $X=7.05 $Y=1.105 $X2=0 $Y2=0
cc_321 N_A2_c_349_n N_A_1224_297#_c_891_n 0.00197018f $X=7.305 $Y=1.16 $X2=0
+ $Y2=0
cc_322 N_A2_M1039_g N_A_1224_297#_c_889_n 0.0123686f $X=7.305 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A2_M1015_g N_A_1224_297#_c_890_n 0.00937398f $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A2_M1021_g N_A_1224_297#_c_890_n 0.00687399f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A2_M1033_g N_A_1224_297#_c_890_n 5.07492e-19 $X=6.885 $Y=1.985 $X2=0
+ $Y2=0
cc_326 A2 N_A_1224_297#_c_890_n 0.0169697f $X=7.05 $Y=1.105 $X2=0 $Y2=0
cc_327 N_A2_c_349_n N_A_1224_297#_c_890_n 0.00205111f $X=7.305 $Y=1.16 $X2=0
+ $Y2=0
cc_328 N_A2_M1021_g N_A_1224_297#_c_901_n 5.07492e-19 $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A2_M1033_g N_A_1224_297#_c_901_n 0.00687399f $X=6.885 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_A2_M1039_g N_A_1224_297#_c_901_n 0.0114674f $X=7.305 $Y=1.985 $X2=0
+ $Y2=0
cc_331 A2 N_A_1224_297#_c_901_n 0.0169697f $X=7.05 $Y=1.105 $X2=0 $Y2=0
cc_332 N_A2_c_349_n N_A_1224_297#_c_901_n 0.00205111f $X=7.305 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_A2_M1009_g N_A_27_47#_c_956_n 0.012933f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_334 N_A2_M1016_g N_A_27_47#_c_956_n 0.00850187f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_335 A2 N_A_27_47#_c_956_n 0.0298075f $X=7.05 $Y=1.105 $X2=0 $Y2=0
cc_336 N_A2_c_349_n N_A_27_47#_c_956_n 0.00210947f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A2_M1009_g N_A_27_47#_c_1007_n 5.82624e-19 $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_338 N_A2_M1016_g N_A_27_47#_c_1007_n 0.00660544f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A2_M1019_g N_A_27_47#_c_1007_n 0.00654251f $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A2_M1028_g N_A_27_47#_c_1007_n 5.77739e-19 $X=7.305 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A2_M1009_g N_A_27_47#_c_962_n 0.00697849f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A2_M1016_g N_A_27_47#_c_962_n 5.64169e-19 $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_343 N_A2_M1016_g N_A_27_47#_c_963_n 0.00110555f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A2_M1019_g N_A_27_47#_c_963_n 0.00110555f $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_345 A2 N_A_27_47#_c_963_n 0.0265407f $X=7.05 $Y=1.105 $X2=0 $Y2=0
cc_346 N_A2_c_349_n N_A_27_47#_c_963_n 0.00219112f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A2_M1019_g N_A_27_47#_c_964_n 0.00850187f $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A2_M1028_g N_A_27_47#_c_964_n 0.00969146f $X=7.305 $Y=0.56 $X2=0 $Y2=0
cc_349 A2 N_A_27_47#_c_964_n 0.0298075f $X=7.05 $Y=1.105 $X2=0 $Y2=0
cc_350 N_A2_c_349_n N_A_27_47#_c_964_n 0.00210947f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A2_M1019_g N_A_27_47#_c_965_n 5.74673e-19 $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_352 N_A2_M1028_g N_A_27_47#_c_965_n 0.00835358f $X=7.305 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A2_M1009_g N_VGND_c_1121_n 0.00268723f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A2_M1016_g N_VGND_c_1121_n 0.00146448f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A2_M1019_g N_VGND_c_1122_n 0.00146448f $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A2_M1028_g N_VGND_c_1122_n 0.00268723f $X=7.305 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A2_M1028_g N_VGND_c_1127_n 0.0042294f $X=7.305 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A2_M1009_g N_VGND_c_1131_n 0.00433784f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A2_M1016_g N_VGND_c_1132_n 0.00424416f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A2_M1019_g N_VGND_c_1132_n 0.00424416f $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A2_M1009_g N_VGND_c_1134_n 0.00654026f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A2_M1016_g N_VGND_c_1134_n 0.00573607f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A2_M1019_g N_VGND_c_1134_n 0.00573607f $X=6.885 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A2_M1028_g N_VGND_c_1134_n 0.00707125f $X=7.305 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A1_M1001_g N_VPWR_c_686_n 0.00321269f $X=8.245 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A1_M1005_g N_VPWR_c_687_n 0.00146448f $X=8.665 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A1_M1026_g N_VPWR_c_687_n 0.00146448f $X=9.085 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A1_M1026_g N_VPWR_c_689_n 4.74261e-19 $X=9.085 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A1_M1032_g N_VPWR_c_689_n 0.018019f $X=9.6 $Y=1.985 $X2=0 $Y2=0
cc_370 A1 N_VPWR_c_689_n 0.0248908f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_371 N_A1_c_428_n N_VPWR_c_689_n 0.00449407f $X=9.715 $Y=1.16 $X2=0 $Y2=0
cc_372 N_A1_M1001_g N_VPWR_c_696_n 0.00541359f $X=8.245 $Y=1.985 $X2=0 $Y2=0
cc_373 N_A1_M1005_g N_VPWR_c_696_n 0.00541359f $X=8.665 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A1_M1026_g N_VPWR_c_698_n 0.00541359f $X=9.085 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A1_M1032_g N_VPWR_c_698_n 0.00407992f $X=9.6 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A1_M1001_g N_VPWR_c_683_n 0.0108276f $X=8.245 $Y=1.985 $X2=0 $Y2=0
cc_377 N_A1_M1005_g N_VPWR_c_683_n 0.00950154f $X=8.665 $Y=1.985 $X2=0 $Y2=0
cc_378 N_A1_M1026_g N_VPWR_c_683_n 0.00973281f $X=9.085 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A1_M1032_g N_VPWR_c_683_n 0.00728641f $X=9.6 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A1_M1001_g N_A_1224_297#_c_889_n 0.0144124f $X=8.245 $Y=1.985 $X2=0
+ $Y2=0
cc_381 N_A1_M1001_g N_A_1224_297#_c_907_n 0.0145598f $X=8.245 $Y=1.985 $X2=0
+ $Y2=0
cc_382 N_A1_M1005_g N_A_1224_297#_c_907_n 0.00975139f $X=8.665 $Y=1.985 $X2=0
+ $Y2=0
cc_383 N_A1_M1026_g N_A_1224_297#_c_907_n 6.1949e-19 $X=9.085 $Y=1.985 $X2=0
+ $Y2=0
cc_384 N_A1_M1005_g N_A_1224_297#_c_910_n 0.0109561f $X=8.665 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_A1_M1026_g N_A_1224_297#_c_910_n 0.0109561f $X=9.085 $Y=1.985 $X2=0
+ $Y2=0
cc_386 N_A1_c_425_n N_A_1224_297#_c_910_n 0.00197018f $X=9.16 $Y=1.16 $X2=0
+ $Y2=0
cc_387 A1 N_A_1224_297#_c_910_n 0.025666f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_388 N_A1_M1026_g N_A_1224_297#_c_914_n 9.46316e-19 $X=9.085 $Y=1.985 $X2=0
+ $Y2=0
cc_389 N_A1_c_424_n N_A_1224_297#_c_914_n 0.00424668f $X=9.525 $Y=1.16 $X2=0
+ $Y2=0
cc_390 N_A1_M1032_g N_A_1224_297#_c_914_n 0.00152598f $X=9.6 $Y=1.985 $X2=0
+ $Y2=0
cc_391 A1 N_A_1224_297#_c_914_n 0.0193333f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_392 N_A1_M1005_g N_A_1224_297#_c_918_n 6.1949e-19 $X=8.665 $Y=1.985 $X2=0
+ $Y2=0
cc_393 N_A1_M1026_g N_A_1224_297#_c_918_n 0.00975139f $X=9.085 $Y=1.985 $X2=0
+ $Y2=0
cc_394 N_A1_M1032_g N_A_1224_297#_c_918_n 0.00668144f $X=9.6 $Y=1.985 $X2=0
+ $Y2=0
cc_395 N_A1_M1001_g N_A_1224_297#_c_921_n 9.46316e-19 $X=8.245 $Y=1.985 $X2=0
+ $Y2=0
cc_396 N_A1_M1005_g N_A_1224_297#_c_921_n 9.46316e-19 $X=8.665 $Y=1.985 $X2=0
+ $Y2=0
cc_397 N_A1_c_425_n N_A_1224_297#_c_921_n 0.00206595f $X=9.16 $Y=1.16 $X2=0
+ $Y2=0
cc_398 A1 N_A_1224_297#_c_921_n 0.0171311f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_399 N_A1_M1010_g N_A_27_47#_c_957_n 0.0158613f $X=8.245 $Y=0.56 $X2=0 $Y2=0
cc_400 N_A1_M1017_g N_A_27_47#_c_957_n 0.00850187f $X=8.665 $Y=0.56 $X2=0 $Y2=0
cc_401 N_A1_c_425_n N_A_27_47#_c_957_n 0.00210947f $X=9.16 $Y=1.16 $X2=0 $Y2=0
cc_402 A1 N_A_27_47#_c_957_n 0.0298075f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_403 N_A1_M1010_g N_A_27_47#_c_1027_n 6.15105e-19 $X=8.245 $Y=0.56 $X2=0 $Y2=0
cc_404 N_A1_M1017_g N_A_27_47#_c_1027_n 0.00699928f $X=8.665 $Y=0.56 $X2=0 $Y2=0
cc_405 N_A1_M1018_g N_A_27_47#_c_1027_n 0.00698027f $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_406 N_A1_M1020_g N_A_27_47#_c_1027_n 5.84711e-19 $X=9.6 $Y=0.56 $X2=0 $Y2=0
cc_407 N_A1_M1018_g N_A_27_47#_c_958_n 0.00903265f $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_408 N_A1_c_424_n N_A_27_47#_c_958_n 0.00433613f $X=9.525 $Y=1.16 $X2=0 $Y2=0
cc_409 N_A1_M1020_g N_A_27_47#_c_958_n 0.0103171f $X=9.6 $Y=0.56 $X2=0 $Y2=0
cc_410 A1 N_A_27_47#_c_958_n 0.0749003f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_411 N_A1_c_428_n N_A_27_47#_c_958_n 0.00499088f $X=9.715 $Y=1.16 $X2=0 $Y2=0
cc_412 N_A1_M1018_g N_A_27_47#_c_959_n 5.85693e-19 $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A1_M1020_g N_A_27_47#_c_959_n 0.00701441f $X=9.6 $Y=0.56 $X2=0 $Y2=0
cc_414 N_A1_M1010_g N_A_27_47#_c_965_n 0.0121897f $X=8.245 $Y=0.56 $X2=0 $Y2=0
cc_415 N_A1_M1017_g N_A_27_47#_c_966_n 0.00110555f $X=8.665 $Y=0.56 $X2=0 $Y2=0
cc_416 N_A1_M1018_g N_A_27_47#_c_966_n 0.00110555f $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_417 N_A1_c_425_n N_A_27_47#_c_966_n 0.00219112f $X=9.16 $Y=1.16 $X2=0 $Y2=0
cc_418 A1 N_A_27_47#_c_966_n 0.0265407f $X=9.83 $Y=1.105 $X2=0 $Y2=0
cc_419 N_A1_M1010_g N_VGND_c_1123_n 0.00268723f $X=8.245 $Y=0.56 $X2=0 $Y2=0
cc_420 N_A1_M1017_g N_VGND_c_1123_n 0.00146448f $X=8.665 $Y=0.56 $X2=0 $Y2=0
cc_421 N_A1_M1018_g N_VGND_c_1124_n 0.00165665f $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_422 N_A1_M1020_g N_VGND_c_1124_n 0.002917f $X=9.6 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A1_M1010_g N_VGND_c_1127_n 0.00439206f $X=8.245 $Y=0.56 $X2=0 $Y2=0
cc_424 N_A1_M1017_g N_VGND_c_1129_n 0.00424416f $X=8.665 $Y=0.56 $X2=0 $Y2=0
cc_425 N_A1_M1018_g N_VGND_c_1129_n 0.00424416f $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_426 N_A1_M1020_g N_VGND_c_1133_n 0.00424416f $X=9.6 $Y=0.56 $X2=0 $Y2=0
cc_427 N_A1_M1010_g N_VGND_c_1134_n 0.00733298f $X=8.245 $Y=0.56 $X2=0 $Y2=0
cc_428 N_A1_M1017_g N_VGND_c_1134_n 0.00573607f $X=8.665 $Y=0.56 $X2=0 $Y2=0
cc_429 N_A1_M1018_g N_VGND_c_1134_n 0.00596734f $X=9.085 $Y=0.56 $X2=0 $Y2=0
cc_430 N_A1_M1020_g N_VGND_c_1134_n 0.00697875f $X=9.6 $Y=0.56 $X2=0 $Y2=0
cc_431 N_A_27_297#_c_508_n N_Y_M1004_d 0.0031439f $X=1.015 $Y=2.36 $X2=0 $Y2=0
cc_432 N_A_27_297#_c_510_n N_Y_M1025_d 0.0031439f $X=1.87 $Y=2.36 $X2=0 $Y2=0
cc_433 N_A_27_297#_M1006_s N_Y_c_578_n 0.00328413f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_434 N_A_27_297#_c_508_n N_Y_c_578_n 0.0029342f $X=1.015 $Y=2.36 $X2=0 $Y2=0
cc_435 N_A_27_297#_c_521_p N_Y_c_578_n 0.0126131f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_436 N_A_27_297#_c_510_n N_Y_c_578_n 0.00577832f $X=1.87 $Y=2.36 $X2=0 $Y2=0
cc_437 N_A_27_297#_M1034_s N_Y_c_568_n 5.05631e-19 $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_438 N_A_27_297#_M1011_d N_Y_c_571_n 0.00328413f $X=2.66 $Y=1.485 $X2=0 $Y2=0
cc_439 N_A_27_297#_M1029_d N_Y_c_571_n 0.00690355f $X=3.5 $Y=1.485 $X2=0 $Y2=0
cc_440 N_A_27_297#_c_513_n N_Y_c_571_n 0.031631f $X=2.71 $Y=1.92 $X2=0 $Y2=0
cc_441 N_A_27_297#_c_515_n N_Y_c_571_n 0.0315971f $X=3.55 $Y=1.92 $X2=0 $Y2=0
cc_442 N_A_27_297#_c_504_n N_Y_c_571_n 0.0197708f $X=3.675 $Y=2.005 $X2=0 $Y2=0
cc_443 N_A_27_297#_c_529_p N_Y_c_571_n 0.012546f $X=2.795 $Y=1.92 $X2=0 $Y2=0
cc_444 N_A_27_297#_M1034_s N_Y_c_584_n 0.0023962f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_445 N_A_27_297#_c_512_n N_Y_c_584_n 0.013179f $X=2.04 $Y=1.92 $X2=0 $Y2=0
cc_446 N_A_27_297#_c_508_n N_Y_c_587_n 0.0161525f $X=1.015 $Y=2.36 $X2=0 $Y2=0
cc_447 N_A_27_297#_c_510_n Y 0.0168004f $X=1.87 $Y=2.36 $X2=0 $Y2=0
cc_448 N_A_27_297#_c_534_p Y 0.00589108f $X=1.955 $Y=2.17 $X2=0 $Y2=0
cc_449 N_A_27_297#_c_512_n Y 0.0140822f $X=2.04 $Y=1.92 $X2=0 $Y2=0
cc_450 N_A_27_297#_c_513_n N_VPWR_M1008_s 0.00317944f $X=2.71 $Y=1.92 $X2=-0.19
+ $Y2=1.305
cc_451 N_A_27_297#_c_515_n N_VPWR_M1012_s 0.00317944f $X=3.55 $Y=1.92 $X2=0
+ $Y2=0
cc_452 N_A_27_297#_c_513_n N_VPWR_c_684_n 0.0163351f $X=2.71 $Y=1.92 $X2=0 $Y2=0
cc_453 N_A_27_297#_c_515_n N_VPWR_c_685_n 0.0163351f $X=3.55 $Y=1.92 $X2=0 $Y2=0
cc_454 N_A_27_297#_c_502_n N_VPWR_c_690_n 0.0177497f $X=0.217 $Y=2.255 $X2=0
+ $Y2=0
cc_455 N_A_27_297#_c_508_n N_VPWR_c_690_n 0.0362386f $X=1.015 $Y=2.36 $X2=0
+ $Y2=0
cc_456 N_A_27_297#_c_510_n N_VPWR_c_690_n 0.0486447f $X=1.87 $Y=2.36 $X2=0 $Y2=0
cc_457 N_A_27_297#_c_513_n N_VPWR_c_690_n 0.0020257f $X=2.71 $Y=1.92 $X2=0 $Y2=0
cc_458 N_A_27_297#_c_544_p N_VPWR_c_690_n 0.0114055f $X=1.1 $Y=2.34 $X2=0 $Y2=0
cc_459 N_A_27_297#_c_513_n N_VPWR_c_692_n 0.0020257f $X=2.71 $Y=1.92 $X2=0 $Y2=0
cc_460 N_A_27_297#_c_546_p N_VPWR_c_692_n 0.0089773f $X=2.795 $Y=2.26 $X2=0
+ $Y2=0
cc_461 N_A_27_297#_c_515_n N_VPWR_c_692_n 0.0020257f $X=3.55 $Y=1.92 $X2=0 $Y2=0
cc_462 N_A_27_297#_c_515_n N_VPWR_c_694_n 0.0020257f $X=3.55 $Y=1.92 $X2=0 $Y2=0
cc_463 N_A_27_297#_c_505_n N_VPWR_c_694_n 0.0171883f $X=3.635 $Y=2.26 $X2=0
+ $Y2=0
cc_464 N_A_27_297#_M1004_s N_VPWR_c_683_n 0.00209324f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_465 N_A_27_297#_M1006_s N_VPWR_c_683_n 0.0021521f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_466 N_A_27_297#_M1034_s N_VPWR_c_683_n 0.00252971f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_A_27_297#_M1011_d N_VPWR_c_683_n 0.00264883f $X=2.66 $Y=1.485 $X2=0
+ $Y2=0
cc_468 N_A_27_297#_M1029_d N_VPWR_c_683_n 0.00233432f $X=3.5 $Y=1.485 $X2=0
+ $Y2=0
cc_469 N_A_27_297#_c_502_n N_VPWR_c_683_n 0.00981527f $X=0.217 $Y=2.255 $X2=0
+ $Y2=0
cc_470 N_A_27_297#_c_508_n N_VPWR_c_683_n 0.023553f $X=1.015 $Y=2.36 $X2=0 $Y2=0
cc_471 N_A_27_297#_c_510_n N_VPWR_c_683_n 0.0307184f $X=1.87 $Y=2.36 $X2=0 $Y2=0
cc_472 N_A_27_297#_c_513_n N_VPWR_c_683_n 0.00913773f $X=2.71 $Y=1.92 $X2=0
+ $Y2=0
cc_473 N_A_27_297#_c_546_p N_VPWR_c_683_n 0.00631544f $X=2.795 $Y=2.26 $X2=0
+ $Y2=0
cc_474 N_A_27_297#_c_515_n N_VPWR_c_683_n 0.00913773f $X=3.55 $Y=1.92 $X2=0
+ $Y2=0
cc_475 N_A_27_297#_c_505_n N_VPWR_c_683_n 0.00953181f $X=3.635 $Y=2.26 $X2=0
+ $Y2=0
cc_476 N_A_27_297#_c_544_p N_VPWR_c_683_n 0.00653405f $X=1.1 $Y=2.34 $X2=0 $Y2=0
cc_477 N_A_27_297#_c_505_n N_A_806_297#_c_827_n 0.0168365f $X=3.635 $Y=2.26
+ $X2=0 $Y2=0
cc_478 N_A_27_297#_c_504_n N_A_806_297#_c_828_n 0.0136295f $X=3.675 $Y=2.005
+ $X2=0 $Y2=0
cc_479 N_A_27_297#_c_505_n N_A_806_297#_c_828_n 0.0183843f $X=3.635 $Y=2.26
+ $X2=0 $Y2=0
cc_480 N_A_27_297#_c_503_n N_A_27_47#_c_953_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0
+ $Y2=0
cc_481 N_Y_c_571_n N_VPWR_M1008_s 0.00328818f $X=4.41 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_482 N_Y_c_571_n N_VPWR_M1012_s 0.00328818f $X=4.41 $Y=1.58 $X2=0 $Y2=0
cc_483 N_Y_M1004_d N_VPWR_c_683_n 0.00216833f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_484 N_Y_M1025_d N_VPWR_c_683_n 0.00216833f $X=1.385 $Y=1.485 $X2=0 $Y2=0
cc_485 N_Y_M1000_s N_VPWR_c_683_n 0.00216833f $X=4.44 $Y=1.485 $X2=0 $Y2=0
cc_486 N_Y_M1014_s N_VPWR_c_683_n 0.00216833f $X=5.28 $Y=1.485 $X2=0 $Y2=0
cc_487 N_Y_c_571_n N_A_806_297#_M1000_d 0.00479405f $X=4.41 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_488 N_Y_c_613_n N_A_806_297#_M1007_d 0.00328413f $X=5.25 $Y=1.58 $X2=0 $Y2=0
cc_489 N_Y_c_571_n N_A_806_297#_c_828_n 0.0196863f $X=4.41 $Y=1.58 $X2=0 $Y2=0
cc_490 N_Y_M1000_s N_A_806_297#_c_831_n 0.0031439f $X=4.44 $Y=1.485 $X2=0 $Y2=0
cc_491 N_Y_c_571_n N_A_806_297#_c_831_n 0.0029342f $X=4.41 $Y=1.58 $X2=0 $Y2=0
cc_492 N_Y_c_613_n N_A_806_297#_c_831_n 0.0029342f $X=5.25 $Y=1.58 $X2=0 $Y2=0
cc_493 N_Y_c_617_n N_A_806_297#_c_831_n 0.0161525f $X=4.575 $Y=1.66 $X2=0 $Y2=0
cc_494 N_Y_c_613_n N_A_806_297#_c_849_n 0.0126131f $X=5.25 $Y=1.58 $X2=0 $Y2=0
cc_495 N_Y_M1014_s N_A_806_297#_c_833_n 0.0031439f $X=5.28 $Y=1.485 $X2=0 $Y2=0
cc_496 N_Y_c_613_n N_A_806_297#_c_833_n 0.0029342f $X=5.25 $Y=1.58 $X2=0 $Y2=0
cc_497 N_Y_c_622_n N_A_806_297#_c_833_n 0.0161525f $X=5.415 $Y=1.66 $X2=0 $Y2=0
cc_498 N_Y_c_622_n N_A_1224_297#_c_890_n 0.011001f $X=5.415 $Y=1.66 $X2=0 $Y2=0
cc_499 N_Y_c_567_n N_A_27_47#_M1022_d 0.00169911f $X=1.855 $Y=0.78 $X2=0 $Y2=0
cc_500 N_Y_c_666_p N_A_27_47#_M1035_d 0.00191657f $X=1.945 $Y=0.78 $X2=0 $Y2=0
cc_501 N_Y_c_569_n N_A_27_47#_M1031_d 0.00169911f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_502 N_Y_c_567_n N_A_27_47#_c_953_n 0.01117f $X=1.855 $Y=0.78 $X2=0 $Y2=0
cc_503 N_Y_M1013_s N_A_27_47#_c_970_n 0.00312712f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_504 N_Y_M1023_s N_A_27_47#_c_970_n 0.00312712f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_505 N_Y_M1024_s N_A_27_47#_c_970_n 0.00312712f $X=2.24 $Y=0.235 $X2=0 $Y2=0
cc_506 N_Y_M1036_s N_A_27_47#_c_970_n 0.00312712f $X=3.08 $Y=0.235 $X2=0 $Y2=0
cc_507 N_Y_c_567_n N_A_27_47#_c_970_n 0.0597391f $X=1.855 $Y=0.78 $X2=0 $Y2=0
cc_508 N_Y_c_569_n N_A_27_47#_c_970_n 0.0597391f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_509 N_Y_c_666_p N_A_27_47#_c_970_n 0.0121347f $X=1.945 $Y=0.78 $X2=0 $Y2=0
cc_510 N_Y_c_569_n N_A_27_47#_c_954_n 0.00799569f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_511 N_Y_c_571_n N_A_27_47#_c_954_n 0.00735546f $X=4.41 $Y=1.58 $X2=0 $Y2=0
cc_512 N_Y_c_622_n N_A_27_47#_c_962_n 0.00620948f $X=5.415 $Y=1.66 $X2=0 $Y2=0
cc_513 N_Y_M1013_s N_VGND_c_1134_n 0.00216833f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_514 N_Y_M1023_s N_VGND_c_1134_n 0.00216833f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_515 N_Y_M1024_s N_VGND_c_1134_n 0.00216833f $X=2.24 $Y=0.235 $X2=0 $Y2=0
cc_516 N_Y_M1036_s N_VGND_c_1134_n 0.00216833f $X=3.08 $Y=0.235 $X2=0 $Y2=0
cc_517 N_VPWR_c_683_n N_A_806_297#_M1000_d 0.00209324f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_518 N_VPWR_c_683_n N_A_806_297#_M1007_d 0.0021521f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_683_n N_A_806_297#_M1030_d 0.0021521f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_683_n N_A_806_297#_M1021_d 0.0021521f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_683_n N_A_806_297#_M1039_d 0.00209324f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_694_n N_A_806_297#_c_827_n 0.0172955f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_683_n N_A_806_297#_c_827_n 0.00960883f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_694_n N_A_806_297#_c_831_n 0.0362386f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_683_n N_A_806_297#_c_831_n 0.023553f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_526 N_VPWR_c_694_n N_A_806_297#_c_833_n 0.0362386f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_683_n N_A_806_297#_c_833_n 0.023553f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_528 N_VPWR_c_694_n N_A_806_297#_c_835_n 0.0362386f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_683_n N_A_806_297#_c_835_n 0.023553f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_530 N_VPWR_c_694_n N_A_806_297#_c_837_n 0.0362386f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_683_n N_A_806_297#_c_837_n 0.023553f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_c_686_n N_A_806_297#_c_829_n 0.0168365f $X=8.035 $Y=2 $X2=0 $Y2=0
cc_533 N_VPWR_c_694_n N_A_806_297#_c_829_n 0.0172955f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_683_n N_A_806_297#_c_829_n 0.00960883f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_686_n N_A_806_297#_c_830_n 0.0309727f $X=8.035 $Y=2 $X2=0 $Y2=0
cc_536 N_VPWR_c_694_n N_A_806_297#_c_872_n 0.0114055f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_683_n N_A_806_297#_c_872_n 0.00653405f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_694_n N_A_806_297#_c_874_n 0.0114055f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_683_n N_A_806_297#_c_874_n 0.00653405f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_694_n N_A_806_297#_c_876_n 0.0114055f $X=7.87 $Y=2.72 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_683_n N_A_806_297#_c_876_n 0.00653405f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_683_n N_A_1224_297#_M1015_s 0.00216833f $X=9.89 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_543 N_VPWR_c_683_n N_A_1224_297#_M1033_s 0.00216833f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_683_n N_A_1224_297#_M1001_s 0.00215201f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_683_n N_A_1224_297#_M1026_s 0.00521412f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_546 N_VPWR_M1001_d N_A_1224_297#_c_889_n 0.00690717f $X=7.91 $Y=1.485 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_686_n N_A_1224_297#_c_889_n 0.0198097f $X=8.035 $Y=2 $X2=0 $Y2=0
cc_548 N_VPWR_c_696_n N_A_1224_297#_c_907_n 0.0189039f $X=8.79 $Y=2.72 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_683_n N_A_1224_297#_c_907_n 0.0122217f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_550 N_VPWR_M1005_d N_A_1224_297#_c_910_n 0.00328413f $X=8.74 $Y=1.485 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_687_n N_A_1224_297#_c_910_n 0.0126919f $X=8.875 $Y=2 $X2=0 $Y2=0
cc_552 N_VPWR_c_689_n N_A_1224_297#_c_914_n 0.0142425f $X=9.81 $Y=1.66 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_689_n N_A_1224_297#_c_918_n 0.063015f $X=9.81 $Y=1.66 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_698_n N_A_1224_297#_c_918_n 0.0209845f $X=9.63 $Y=2.72 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_683_n N_A_1224_297#_c_918_n 0.0124268f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_556 N_A_806_297#_c_835_n N_A_1224_297#_M1015_s 0.0031439f $X=6.59 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_557 N_A_806_297#_c_837_n N_A_1224_297#_M1033_s 0.0031439f $X=7.43 $Y=2.36
+ $X2=0 $Y2=0
cc_558 N_A_806_297#_M1021_d N_A_1224_297#_c_891_n 0.00328413f $X=6.54 $Y=1.485
+ $X2=0 $Y2=0
cc_559 N_A_806_297#_c_835_n N_A_1224_297#_c_891_n 0.0029342f $X=6.59 $Y=2.36
+ $X2=0 $Y2=0
cc_560 N_A_806_297#_c_882_p N_A_1224_297#_c_891_n 0.0126131f $X=6.675 $Y=2 $X2=0
+ $Y2=0
cc_561 N_A_806_297#_c_837_n N_A_1224_297#_c_891_n 0.0029342f $X=7.43 $Y=2.36
+ $X2=0 $Y2=0
cc_562 N_A_806_297#_M1039_d N_A_1224_297#_c_889_n 0.00690717f $X=7.38 $Y=1.485
+ $X2=0 $Y2=0
cc_563 N_A_806_297#_c_837_n N_A_1224_297#_c_889_n 0.0029342f $X=7.43 $Y=2.36
+ $X2=0 $Y2=0
cc_564 N_A_806_297#_c_830_n N_A_1224_297#_c_889_n 0.0196863f $X=7.515 $Y=2 $X2=0
+ $Y2=0
cc_565 N_A_806_297#_c_835_n N_A_1224_297#_c_890_n 0.0161525f $X=6.59 $Y=2.36
+ $X2=0 $Y2=0
cc_566 N_A_806_297#_c_837_n N_A_1224_297#_c_901_n 0.0161525f $X=7.43 $Y=2.36
+ $X2=0 $Y2=0
cc_567 N_A_1224_297#_c_889_n N_A_27_47#_c_964_n 0.0308414f $X=8.29 $Y=1.58 $X2=0
+ $Y2=0
cc_568 N_A_27_47#_c_955_n N_VGND_M1002_d 0.00169589f $X=4.31 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_569 N_A_27_47#_c_961_n N_VGND_M1027_d 0.00401257f $X=5.31 $Y=0.58 $X2=0 $Y2=0
cc_570 N_A_27_47#_c_956_n N_VGND_M1009_d 0.00169589f $X=6.51 $Y=0.82 $X2=0 $Y2=0
cc_571 N_A_27_47#_c_964_n N_VGND_M1019_d 0.00169589f $X=7.35 $Y=0.58 $X2=0 $Y2=0
cc_572 N_A_27_47#_c_957_n N_VGND_M1010_d 0.00169589f $X=8.71 $Y=0.82 $X2=0 $Y2=0
cc_573 N_A_27_47#_c_958_n N_VGND_M1018_d 0.00276988f $X=9.645 $Y=0.82 $X2=0
+ $Y2=0
cc_574 N_A_27_47#_c_955_n N_VGND_c_1118_n 0.0111177f $X=4.31 $Y=0.82 $X2=0 $Y2=0
cc_575 N_A_27_47#_c_955_n N_VGND_c_1119_n 0.00193763f $X=4.31 $Y=0.82 $X2=0
+ $Y2=0
cc_576 N_A_27_47#_c_988_n N_VGND_c_1119_n 0.0188551f $X=4.475 $Y=0.38 $X2=0
+ $Y2=0
cc_577 N_A_27_47#_c_961_n N_VGND_c_1119_n 0.00193763f $X=5.31 $Y=0.58 $X2=0
+ $Y2=0
cc_578 N_A_27_47#_c_961_n N_VGND_c_1120_n 0.0225205f $X=5.31 $Y=0.58 $X2=0 $Y2=0
cc_579 N_A_27_47#_c_956_n N_VGND_c_1121_n 0.0111177f $X=6.51 $Y=0.82 $X2=0 $Y2=0
cc_580 N_A_27_47#_c_964_n N_VGND_c_1122_n 0.0111177f $X=7.35 $Y=0.58 $X2=0 $Y2=0
cc_581 N_A_27_47#_c_957_n N_VGND_c_1123_n 0.0111177f $X=8.71 $Y=0.82 $X2=0 $Y2=0
cc_582 N_A_27_47#_c_958_n N_VGND_c_1124_n 0.0178881f $X=9.645 $Y=0.82 $X2=0
+ $Y2=0
cc_583 N_A_27_47#_c_952_n N_VGND_c_1125_n 0.0176918f $X=0.217 $Y=0.465 $X2=0
+ $Y2=0
cc_584 N_A_27_47#_c_970_n N_VGND_c_1125_n 0.177492f $X=3.55 $Y=0.36 $X2=0 $Y2=0
cc_585 N_A_27_47#_c_980_n N_VGND_c_1125_n 0.0152108f $X=3.675 $Y=0.465 $X2=0
+ $Y2=0
cc_586 N_A_27_47#_c_955_n N_VGND_c_1125_n 0.00193763f $X=4.31 $Y=0.82 $X2=0
+ $Y2=0
cc_587 N_A_27_47#_c_957_n N_VGND_c_1127_n 0.0037967f $X=8.71 $Y=0.82 $X2=0 $Y2=0
cc_588 N_A_27_47#_c_964_n N_VGND_c_1127_n 0.00193763f $X=7.35 $Y=0.58 $X2=0
+ $Y2=0
cc_589 N_A_27_47#_c_965_n N_VGND_c_1127_n 0.0459879f $X=8.04 $Y=0.58 $X2=0 $Y2=0
cc_590 N_A_27_47#_c_957_n N_VGND_c_1129_n 0.00193763f $X=8.71 $Y=0.82 $X2=0
+ $Y2=0
cc_591 N_A_27_47#_c_1027_n N_VGND_c_1129_n 0.0188551f $X=8.875 $Y=0.38 $X2=0
+ $Y2=0
cc_592 N_A_27_47#_c_958_n N_VGND_c_1129_n 0.00193763f $X=9.645 $Y=0.82 $X2=0
+ $Y2=0
cc_593 N_A_27_47#_c_956_n N_VGND_c_1131_n 0.00219975f $X=6.51 $Y=0.82 $X2=0
+ $Y2=0
cc_594 N_A_27_47#_c_961_n N_VGND_c_1131_n 0.00193763f $X=5.31 $Y=0.58 $X2=0
+ $Y2=0
cc_595 N_A_27_47#_c_962_n N_VGND_c_1131_n 0.0425836f $X=5.98 $Y=0.58 $X2=0 $Y2=0
cc_596 N_A_27_47#_c_956_n N_VGND_c_1132_n 0.00193763f $X=6.51 $Y=0.82 $X2=0
+ $Y2=0
cc_597 N_A_27_47#_c_1007_n N_VGND_c_1132_n 0.0188551f $X=6.675 $Y=0.38 $X2=0
+ $Y2=0
cc_598 N_A_27_47#_c_964_n N_VGND_c_1132_n 0.00193763f $X=7.35 $Y=0.58 $X2=0
+ $Y2=0
cc_599 N_A_27_47#_c_958_n N_VGND_c_1133_n 0.00197543f $X=9.645 $Y=0.82 $X2=0
+ $Y2=0
cc_600 N_A_27_47#_c_959_n N_VGND_c_1133_n 0.0252622f $X=9.81 $Y=0.38 $X2=0 $Y2=0
cc_601 N_A_27_47#_M1013_d N_VGND_c_1134_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_27_47#_M1022_d N_VGND_c_1134_n 0.00215227f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_603 N_A_27_47#_M1035_d N_VGND_c_1134_n 0.00227273f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_604 N_A_27_47#_M1031_d N_VGND_c_1134_n 0.00215227f $X=2.66 $Y=0.235 $X2=0
+ $Y2=0
cc_605 N_A_27_47#_M1038_d N_VGND_c_1134_n 0.00215206f $X=3.5 $Y=0.235 $X2=0
+ $Y2=0
cc_606 N_A_27_47#_M1003_s N_VGND_c_1134_n 0.00215201f $X=4.34 $Y=0.235 $X2=0
+ $Y2=0
cc_607 N_A_27_47#_M1037_s N_VGND_c_1134_n 0.00508876f $X=5.34 $Y=0.235 $X2=0
+ $Y2=0
cc_608 N_A_27_47#_M1016_s N_VGND_c_1134_n 0.00215201f $X=6.54 $Y=0.235 $X2=0
+ $Y2=0
cc_609 N_A_27_47#_M1028_s N_VGND_c_1134_n 0.00707417f $X=7.38 $Y=0.235 $X2=0
+ $Y2=0
cc_610 N_A_27_47#_M1017_s N_VGND_c_1134_n 0.00215201f $X=8.74 $Y=0.235 $X2=0
+ $Y2=0
cc_611 N_A_27_47#_M1020_s N_VGND_c_1134_n 0.00209319f $X=9.675 $Y=0.235 $X2=0
+ $Y2=0
cc_612 N_A_27_47#_c_952_n N_VGND_c_1134_n 0.00980895f $X=0.217 $Y=0.465 $X2=0
+ $Y2=0
cc_613 N_A_27_47#_c_970_n N_VGND_c_1134_n 0.11388f $X=3.55 $Y=0.36 $X2=0 $Y2=0
cc_614 N_A_27_47#_c_980_n N_VGND_c_1134_n 0.00940698f $X=3.675 $Y=0.465 $X2=0
+ $Y2=0
cc_615 N_A_27_47#_c_955_n N_VGND_c_1134_n 0.00828806f $X=4.31 $Y=0.82 $X2=0
+ $Y2=0
cc_616 N_A_27_47#_c_988_n N_VGND_c_1134_n 0.0122069f $X=4.475 $Y=0.38 $X2=0
+ $Y2=0
cc_617 N_A_27_47#_c_956_n N_VGND_c_1134_n 0.00871293f $X=6.51 $Y=0.82 $X2=0
+ $Y2=0
cc_618 N_A_27_47#_c_1007_n N_VGND_c_1134_n 0.0122069f $X=6.675 $Y=0.38 $X2=0
+ $Y2=0
cc_619 N_A_27_47#_c_957_n N_VGND_c_1134_n 0.012333f $X=8.71 $Y=0.82 $X2=0 $Y2=0
cc_620 N_A_27_47#_c_1027_n N_VGND_c_1134_n 0.0122069f $X=8.875 $Y=0.38 $X2=0
+ $Y2=0
cc_621 N_A_27_47#_c_958_n N_VGND_c_1134_n 0.00877231f $X=9.645 $Y=0.82 $X2=0
+ $Y2=0
cc_622 N_A_27_47#_c_959_n N_VGND_c_1134_n 0.0147199f $X=9.81 $Y=0.38 $X2=0 $Y2=0
cc_623 N_A_27_47#_c_961_n N_VGND_c_1134_n 0.00899121f $X=5.31 $Y=0.58 $X2=0
+ $Y2=0
cc_624 N_A_27_47#_c_962_n N_VGND_c_1134_n 0.0254304f $X=5.98 $Y=0.58 $X2=0 $Y2=0
cc_625 N_A_27_47#_c_964_n N_VGND_c_1134_n 0.00828806f $X=7.35 $Y=0.58 $X2=0
+ $Y2=0
cc_626 N_A_27_47#_c_965_n N_VGND_c_1134_n 0.0263174f $X=8.04 $Y=0.58 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__and3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
M1000 VPWR a_215_311# X VPB phighvt w=1e+06u l=150000u
+  ad=7.741e+11p pd=7.93e+06u as=2.7e+11p ps=2.54e+06u
M1001 X a_215_311# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_301_53# a_109_53# a_215_311# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u
M1003 a_373_53# B a_301_53# VNB nshort w=420000u l=150000u
+  ad=1.071e+11p pd=1.35e+06u as=0p ps=0u
M1004 VGND C a_373_53# VNB nshort w=420000u l=150000u
+  ad=5.325e+11p pd=5.37e+06u as=0p ps=0u
M1005 a_109_53# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1006 a_109_53# A_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 a_215_311# B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.5795e+11p pd=2.99e+06u as=0p ps=0u
M1008 VPWR C a_215_311# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_215_311# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1010 VPWR a_109_53# a_215_311# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_215_311# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__macro_sparecell.spice.pex
* Created: Thu Aug 27 14:27:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_1/A 1 2 3 10
+ 12 15 17 19 22 24 25 28 30 34 41 44 47 49 50 56 57 63
c117 47 0 1.29151e-19 $X=1.15 $Y=1.19
c118 41 0 1.19433e-19 $X=2.14 $Y=1.62
r119 61 63 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.9 $Y=1.16
+ $X2=1.11 $Y2=1.16
r120 59 61 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.48 $Y=1.16
+ $X2=0.9 $Y2=1.16
r121 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.655 $Y=1.19
+ $X2=1.655 $Y2=1.19
r122 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.315 $Y=1.19
+ $X2=1.17 $Y2=1.19
r123 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.51 $Y=1.19
+ $X2=1.655 $Y2=1.19
r124 49 50 0.241336 $w=1.4e-07 $l=1.95e-07 $layer=MET1_cond $X=1.51 $Y=1.19
+ $X2=1.315 $Y2=1.19
r125 47 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.16 $X2=1.11 $Y2=1.16
r126 47 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.17 $Y=1.19
+ $X2=1.17 $Y2=1.19
r127 38 57 13.6685 $w=2.13e-07 $l=2.55e-07 $layer=LI1_cond $X=1.652 $Y=1.445
+ $X2=1.652 $Y2=1.19
r128 37 41 25.5633 $w=2.18e-07 $l=4.88e-07 $layer=LI1_cond $X=1.652 $Y=1.555
+ $X2=2.14 $Y2=1.555
r129 37 38 0.884026 $w=2.15e-07 $l=1.1e-07 $layer=LI1_cond $X=1.652 $Y=1.555
+ $X2=1.652 $Y2=1.445
r130 36 57 15.2766 $w=2.13e-07 $l=2.85e-07 $layer=LI1_cond $X=1.652 $Y=0.905
+ $X2=1.652 $Y2=1.19
r131 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.98 $Y=0.725
+ $X2=2.98 $Y2=0.39
r132 31 44 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.815
+ $X2=2.14 $Y2=0.815
r133 30 32 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.815 $Y=0.815
+ $X2=2.98 $Y2=0.725
r134 30 31 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.815 $Y=0.815
+ $X2=2.305 $Y2=0.815
r135 26 44 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.14 $Y=0.725
+ $X2=2.14 $Y2=0.815
r136 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=0.725
+ $X2=2.14 $Y2=0.39
r137 25 36 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=1.76 $Y=0.82
+ $X2=1.652 $Y2=0.905
r138 24 44 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=2.14 $Y2=0.815
r139 24 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.975 $Y=0.82
+ $X2=1.76 $Y2=0.82
r140 20 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=1.325
+ $X2=0.9 $Y2=1.16
r141 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.9 $Y=1.325
+ $X2=0.9 $Y2=1.985
r142 17 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.9 $Y2=1.16
r143 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.9 $Y2=0.56
r144 13 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r145 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.985
r146 10 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r147 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=0.56
r148 3 41 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.005
+ $Y=1.485 $X2=2.14 $Y2=1.62
r149 2 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.845
+ $Y=0.235 $X2=2.98 $Y2=0.39
r150 1 28 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__NOR2_2_1/B 1 2 3 10
+ 12 15 17 19 22 24 26 29 31 33 36 40 42 46 48 50 52 55 65 67 69 74 75 76 77 86
+ 94 101 111 112
c157 69 0 1.4808e-19 $X=3.905 $Y=0.835
c158 40 0 9.09144e-20 $X=4.46 $Y=0.74
c159 29 0 1.19433e-19 $X=2.77 $Y=1.985
r160 99 101 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.035 $Y=1.16
+ $X2=3.19 $Y2=1.16
r161 96 99 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=2.77 $Y=1.16
+ $X2=3.035 $Y2=1.16
r162 92 94 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.14 $Y=1.16
+ $X2=2.35 $Y2=1.16
r163 89 92 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.93 $Y=1.16
+ $X2=2.14 $Y2=1.16
r164 77 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.19 $Y=1.19
+ $X2=3.045 $Y2=1.19
r165 76 86 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.76 $Y=1.19
+ $X2=3.905 $Y2=1.19
r166 76 77 0.705444 $w=1.4e-07 $l=5.7e-07 $layer=MET1_cond $X=3.76 $Y=1.19
+ $X2=3.19 $Y2=1.19
r167 75 79 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.33 $Y=1.19
+ $X2=2.185 $Y2=1.19
r168 74 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.9 $Y=1.19
+ $X2=3.045 $Y2=1.19
r169 74 75 0.705444 $w=1.4e-07 $l=5.7e-07 $layer=MET1_cond $X=2.9 $Y=1.19
+ $X2=2.33 $Y2=1.19
r170 72 112 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=1.58
+ $X2=3.905 $Y2=1.495
r171 72 112 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.905 $Y=1.47
+ $X2=3.905 $Y2=1.495
r172 71 72 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=3.905 $Y=1.19
+ $X2=3.905 $Y2=1.47
r173 71 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.905 $Y=1.19
+ $X2=3.905 $Y2=1.19
r174 69 111 3.22874 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=0.78
+ $X2=3.905 $Y2=0.905
r175 69 71 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.905 $Y=0.92
+ $X2=3.905 $Y2=1.19
r176 69 111 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.905 $Y=0.92
+ $X2=3.905 $Y2=0.905
r177 67 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=1.16 $X2=3.035 $Y2=1.16
r178 67 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.045 $Y=1.19
+ $X2=3.045 $Y2=1.19
r179 65 92 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r180 65 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.185 $Y=1.19
+ $X2=2.185 $Y2=1.19
r181 50 57 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=1.665 $X2=5.3
+ $Y2=1.58
r182 50 52 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.3 $Y=1.665
+ $X2=5.3 $Y2=2.34
r183 49 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=1.58
+ $X2=4.46 $Y2=1.58
r184 48 57 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=1.58
+ $X2=5.3 $Y2=1.58
r185 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.135 $Y=1.58
+ $X2=4.625 $Y2=1.58
r186 44 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=1.665
+ $X2=4.46 $Y2=1.58
r187 44 46 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.46 $Y=1.665
+ $X2=4.46 $Y2=2.34
r188 43 72 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.045 $Y=1.58
+ $X2=3.905 $Y2=1.58
r189 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=1.58
+ $X2=4.46 $Y2=1.58
r190 42 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.295 $Y=1.58
+ $X2=4.045 $Y2=1.58
r191 38 69 3.61619 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=4.045 $Y=0.78
+ $X2=3.905 $Y2=0.78
r192 38 40 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=4.045 $Y=0.78
+ $X2=4.46 $Y2=0.78
r193 34 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.325
+ $X2=3.19 $Y2=1.16
r194 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.19 $Y=1.325
+ $X2=3.19 $Y2=1.985
r195 31 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=0.995
+ $X2=3.19 $Y2=1.16
r196 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.19 $Y=0.995
+ $X2=3.19 $Y2=0.56
r197 27 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.325
+ $X2=2.77 $Y2=1.16
r198 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.77 $Y=1.325
+ $X2=2.77 $Y2=1.985
r199 24 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=0.995
+ $X2=2.77 $Y2=1.16
r200 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.77 $Y=0.995
+ $X2=2.77 $Y2=0.56
r201 20 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.325
+ $X2=2.35 $Y2=1.16
r202 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.35 $Y=1.325
+ $X2=2.35 $Y2=1.985
r203 17 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.16
r204 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r205 13 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=1.325
+ $X2=1.93 $Y2=1.16
r206 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.93 $Y=1.325
+ $X2=1.93 $Y2=1.985
r207 10 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.16
r208 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r209 3 57 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=1.66
r210 3 52 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2.34
r211 2 55 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=1.66
r212 2 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2.34
r213 1 40 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%LO 1 3 6 8 10 13 15 17 20 22 24 27
+ 29 31 34 36 38 41 43 45 48 50 52 55 67 69 72 75 76 77 78 79 80 81 82 94 97 99
+ 101 109 116 123 129 130 142
c232 75 0 1.95213e-19 $X=5.645 $Y=1.19
c233 43 0 5.77853e-20 $X=8.67 $Y=0.995
c234 36 0 9.09144e-20 $X=8.25 $Y=0.995
c235 15 0 9.09144e-20 $X=5.09 $Y=0.995
c236 8 0 5.77853e-20 $X=4.67 $Y=0.995
r237 128 130 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.88 $Y=1.16
+ $X2=9.09 $Y2=1.16
r238 128 129 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.88
+ $Y=1.16 $X2=8.88 $Y2=1.16
r239 125 128 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.67 $Y=1.16
+ $X2=8.88 $Y2=1.16
r240 121 123 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.04 $Y=1.16
+ $X2=8.25 $Y2=1.16
r241 118 121 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.83 $Y=1.16
+ $X2=8.04 $Y2=1.16
r242 114 116 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.3 $Y=1.16
+ $X2=5.51 $Y2=1.16
r243 111 114 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.3 $Y2=1.16
r244 107 109 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.46 $Y=1.16
+ $X2=4.67 $Y2=1.16
r245 107 108 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r246 104 107 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.46 $Y2=1.16
r247 101 102 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.92
+ $Y=1.995 $X2=6.92 $Y2=1.995
r248 99 101 88.0569 $w=4.8e-07 $l=7.9e-07 $layer=POLY_cond $X=7.015 $Y=1.205
+ $X2=7.015 $Y2=1.995
r249 97 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.85 $Y=1.19
+ $X2=6.85 $Y2=1.19
r250 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.71 $Y=1.19
+ $X2=7.71 $Y2=1.19
r251 82 91 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.855 $Y=1.19
+ $X2=7.71 $Y2=1.19
r252 81 94 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.425 $Y=1.19
+ $X2=8.57 $Y2=1.19
r253 81 82 0.705444 $w=1.4e-07 $l=5.7e-07 $layer=MET1_cond $X=8.425 $Y=1.19
+ $X2=7.855 $Y2=1.19
r254 80 97 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.995 $Y=1.19
+ $X2=6.85 $Y2=1.19
r255 79 91 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.565 $Y=1.19
+ $X2=7.71 $Y2=1.19
r256 79 80 0.705444 $w=1.4e-07 $l=5.7e-07 $layer=MET1_cond $X=7.565 $Y=1.19
+ $X2=6.995 $Y2=1.19
r257 78 88 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.935 $Y=1.19
+ $X2=5.79 $Y2=1.19
r258 77 97 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.705 $Y=1.19
+ $X2=6.85 $Y2=1.19
r259 77 78 0.952968 $w=1.4e-07 $l=7.7e-07 $layer=MET1_cond $X=6.705 $Y=1.19
+ $X2=5.935 $Y2=1.19
r260 76 84 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.005 $Y=1.19
+ $X2=4.86 $Y2=1.19
r261 75 88 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.645 $Y=1.19
+ $X2=5.79 $Y2=1.19
r262 75 76 0.792078 $w=1.4e-07 $l=6.4e-07 $layer=MET1_cond $X=5.645 $Y=1.19
+ $X2=5.005 $Y2=1.19
r263 73 129 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=8.515 $Y=1.2
+ $X2=8.88 $Y2=1.2
r264 73 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.57 $Y=1.19
+ $X2=8.57 $Y2=1.19
r265 72 92 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=8.04 $Y=1.2
+ $X2=7.71 $Y2=1.2
r266 72 121 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.04
+ $Y=1.16 $X2=8.04 $Y2=1.16
r267 70 102 10.6957 $w=5.18e-07 $l=4.65e-07 $layer=LI1_cond $X=7.015 $Y=1.53
+ $X2=7.015 $Y2=1.995
r268 70 142 7.82051 $w=5.18e-07 $l=3.4e-07 $layer=LI1_cond $X=7.015 $Y=1.53
+ $X2=7.015 $Y2=1.19
r269 69 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.79 $Y=1.19
+ $X2=5.79 $Y2=1.19
r270 68 69 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=5.285 $Y=1.2
+ $X2=5.745 $Y2=1.2
r271 68 114 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.3
+ $Y=1.16 $X2=5.3 $Y2=1.16
r272 67 108 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=4.825 $Y=1.2
+ $X2=4.46 $Y2=1.2
r273 67 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.86 $Y=1.19
+ $X2=4.86 $Y2=1.19
r274 53 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.09 $Y=1.325
+ $X2=9.09 $Y2=1.16
r275 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.09 $Y=1.325
+ $X2=9.09 $Y2=1.985
r276 50 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.09 $Y=0.995
+ $X2=9.09 $Y2=1.16
r277 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.09 $Y=0.995
+ $X2=9.09 $Y2=0.56
r278 46 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.325
+ $X2=8.67 $Y2=1.16
r279 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.67 $Y=1.325
+ $X2=8.67 $Y2=1.985
r280 43 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=0.995
+ $X2=8.67 $Y2=1.16
r281 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.67 $Y=0.995
+ $X2=8.67 $Y2=0.56
r282 39 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.25 $Y=1.325
+ $X2=8.25 $Y2=1.16
r283 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.25 $Y=1.325
+ $X2=8.25 $Y2=1.985
r284 36 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.25 $Y=0.995
+ $X2=8.25 $Y2=1.16
r285 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.25 $Y=0.995
+ $X2=8.25 $Y2=0.56
r286 32 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.83 $Y=1.325
+ $X2=7.83 $Y2=1.16
r287 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.83 $Y=1.325
+ $X2=7.83 $Y2=1.985
r288 29 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.83 $Y=0.995
+ $X2=7.83 $Y2=1.16
r289 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.83 $Y=0.995
+ $X2=7.83 $Y2=0.56
r290 25 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=1.325
+ $X2=5.51 $Y2=1.16
r291 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.51 $Y=1.325
+ $X2=5.51 $Y2=1.985
r292 22 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=0.995
+ $X2=5.51 $Y2=1.16
r293 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.51 $Y=0.995
+ $X2=5.51 $Y2=0.56
r294 18 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.325
+ $X2=5.09 $Y2=1.16
r295 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.09 $Y=1.325
+ $X2=5.09 $Y2=1.985
r296 15 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=0.995
+ $X2=5.09 $Y2=1.16
r297 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.09 $Y=0.995
+ $X2=5.09 $Y2=0.56
r298 11 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=1.325
+ $X2=4.67 $Y2=1.16
r299 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.67 $Y=1.325
+ $X2=4.67 $Y2=1.985
r300 8 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=0.995
+ $X2=4.67 $Y2=1.16
r301 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.67 $Y=0.995
+ $X2=4.67 $Y2=0.56
r302 4 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.325
+ $X2=4.25 $Y2=1.16
r303 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.25 $Y=1.325
+ $X2=4.25 $Y2=1.985
r304 1 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=1.16
r305 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37
+ 39 45 51 53 57 59 63 67 73 74 78 84 88 92 96 100 102 107 108 110 111 113 114
+ 115 131 134 139 147 156 167 171 179 188 191 194 197 200 203 206 209 213
c198 67 0 6.22404e-20 $X=5.72 $Y=1.66
c199 9 0 1.4808e-19 $X=9.165 $Y=1.485
c200 4 0 1.4808e-19 $X=3.915 $Y=1.485
r201 212 213 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r202 206 207 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r203 197 198 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r204 195 198 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r205 194 195 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r206 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r207 183 213 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r208 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r209 180 209 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.315 $Y=2.72
+ $X2=12.2 $Y2=2.72
r210 180 182 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.315 $Y=2.72
+ $X2=12.65 $Y2=2.72
r211 179 212 3.66464 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=12.985 $Y=2.72
+ $X2=13.162 $Y2=2.72
r212 179 182 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.985 $Y=2.72
+ $X2=12.65 $Y2=2.72
r213 177 178 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r214 175 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r215 175 207 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r216 174 177 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r217 174 175 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r218 172 206 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=2.72
+ $X2=10.36 $Y2=2.72
r219 172 174 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.525 $Y=2.72
+ $X2=10.81 $Y2=2.72
r220 171 209 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.085 $Y=2.72
+ $X2=12.2 $Y2=2.72
r221 171 177 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.085 $Y=2.72
+ $X2=11.73 $Y2=2.72
r222 167 206 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.195 $Y=2.72
+ $X2=10.36 $Y2=2.72
r223 167 169 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.195 $Y=2.72
+ $X2=9.89 $Y2=2.72
r224 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r225 163 166 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r226 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r227 160 203 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=7.575 $Y2=2.72
r228 160 162 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=8.05 $Y2=2.72
r229 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r230 156 203 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.445 $Y=2.72
+ $X2=7.575 $Y2=2.72
r231 156 158 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.445 $Y=2.72
+ $X2=7.13 $Y2=2.72
r232 152 200 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.895 $Y=2.72
+ $X2=5.765 $Y2=2.72
r233 152 154 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.895 $Y=2.72
+ $X2=6.21 $Y2=2.72
r234 151 198 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r235 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r236 148 197 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=4.88 $Y2=2.72
r237 148 150 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=5.29 $Y2=2.72
r238 147 200 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.765 $Y2=2.72
r239 147 150 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.29 $Y2=2.72
r240 146 192 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r241 145 146 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r242 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r243 142 145 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r244 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r245 140 188 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.14 $Y2=2.72
r246 140 142 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.61 $Y2=2.72
r247 139 191 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.98 $Y2=2.72
r248 139 145 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.53 $Y2=2.72
r249 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r250 135 185 3.6634 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.177 $Y2=2.72
r251 135 137 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.69 $Y2=2.72
r252 134 188 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=1.14 $Y2=2.72
r253 134 137 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=0.69 $Y2=2.72
r254 130 183 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=12.65 $Y2=2.72
r255 130 178 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r256 130 209 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r257 129 207 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r258 129 166 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=8.97 $Y2=2.72
r259 129 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r260 128 163 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r261 128 159 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r262 128 203 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r263 127 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r264 127 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r265 126 127 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=5.745 $Y=2.72
+ $X2=6.21 $Y2=2.72
r266 126 151 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=5.745 $Y=2.72
+ $X2=5.29 $Y2=2.72
r267 126 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r268 125 195 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=3.445 $Y=2.72
+ $X2=3.91 $Y2=2.72
r269 125 192 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=3.445 $Y=2.72
+ $X2=2.99 $Y2=2.72
r270 124 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r271 124 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r272 124 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r273 115 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r274 115 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r275 113 165 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.215 $Y=2.72
+ $X2=8.97 $Y2=2.72
r276 113 114 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.215 $Y=2.72
+ $X2=9.342 $Y2=2.72
r277 112 169 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.47 $Y=2.72
+ $X2=9.89 $Y2=2.72
r278 112 114 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.47 $Y=2.72
+ $X2=9.342 $Y2=2.72
r279 110 162 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.375 $Y=2.72
+ $X2=8.05 $Y2=2.72
r280 110 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.375 $Y=2.72
+ $X2=8.46 $Y2=2.72
r281 109 165 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.545 $Y=2.72
+ $X2=8.97 $Y2=2.72
r282 109 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=2.72
+ $X2=8.46 $Y2=2.72
r283 107 154 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.255 $Y=2.72
+ $X2=6.21 $Y2=2.72
r284 107 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=2.72
+ $X2=6.42 $Y2=2.72
r285 106 158 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=7.13 $Y2=2.72
r286 106 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=2.72
+ $X2=6.42 $Y2=2.72
r287 102 105 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=13.09 $Y=1.66
+ $X2=13.09 $Y2=2.34
r288 100 212 3.25055 $w=2.1e-07 $l=1.15521e-07 $layer=LI1_cond $X=13.09 $Y=2.635
+ $X2=13.162 $Y2=2.72
r289 100 105 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=13.09 $Y=2.635
+ $X2=13.09 $Y2=2.34
r290 96 99 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=12.2 $Y=1.66
+ $X2=12.2 $Y2=2.34
r291 94 209 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=2.635
+ $X2=12.2 $Y2=2.72
r292 94 99 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.2 $Y=2.635
+ $X2=12.2 $Y2=2.34
r293 90 206 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=2.635
+ $X2=10.36 $Y2=2.72
r294 90 92 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=10.36 $Y=2.635
+ $X2=10.36 $Y2=2
r295 86 114 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.342 $Y=2.635
+ $X2=9.342 $Y2=2.72
r296 86 88 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=9.342 $Y=2.635
+ $X2=9.342 $Y2=2
r297 82 111 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=2.635
+ $X2=8.46 $Y2=2.72
r298 82 84 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.46 $Y=2.635
+ $X2=8.46 $Y2=2
r299 78 81 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=7.575 $Y=1.66
+ $X2=7.575 $Y2=2.34
r300 76 203 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=2.635
+ $X2=7.575 $Y2=2.72
r301 76 81 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=7.575 $Y=2.635
+ $X2=7.575 $Y2=2.34
r302 74 131 88.0569 $w=4.8e-07 $l=7.9e-07 $layer=POLY_cond $X=6.325 $Y=1.995
+ $X2=6.325 $Y2=1.205
r303 73 74 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.42
+ $Y=1.995 $X2=6.42 $Y2=1.995
r304 71 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r305 71 73 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=1.995
r306 67 70 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=5.765 $Y=1.66
+ $X2=5.765 $Y2=2.34
r307 65 200 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.765 $Y=2.635
+ $X2=5.765 $Y2=2.72
r308 65 70 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.765 $Y=2.635
+ $X2=5.765 $Y2=2.34
r309 61 197 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2.72
r310 61 63 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2
r311 60 194 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.125 $Y=2.72
+ $X2=3.997 $Y2=2.72
r312 59 197 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.88 $Y2=2.72
r313 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.125 $Y2=2.72
r314 55 194 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.997 $Y=2.635
+ $X2=3.997 $Y2=2.72
r315 55 57 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=3.997 $Y=2.635
+ $X2=3.997 $Y2=2
r316 54 191 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=2.72
+ $X2=2.98 $Y2=2.72
r317 53 194 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.87 $Y=2.72
+ $X2=3.997 $Y2=2.72
r318 53 54 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.87 $Y=2.72
+ $X2=3.145 $Y2=2.72
r319 49 191 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.635
+ $X2=2.98 $Y2=2.72
r320 49 51 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.98 $Y=2.635
+ $X2=2.98 $Y2=2
r321 45 48 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.14 $Y=1.66
+ $X2=1.14 $Y2=2.34
r322 43 188 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.72
r323 43 48 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.34
r324 39 42 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.25 $Y=1.66
+ $X2=0.25 $Y2=2.34
r325 37 185 3.25179 $w=2.1e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.25 $Y=2.635
+ $X2=0.177 $Y2=2.72
r326 37 42 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.25 $Y=2.635
+ $X2=0.25 $Y2=2.34
r327 12 105 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.935
+ $Y=1.485 $X2=13.07 $Y2=2.34
r328 12 102 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=12.935
+ $Y=1.485 $X2=13.07 $Y2=1.66
r329 11 99 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=12.105
+ $Y=1.485 $X2=12.23 $Y2=2.34
r330 11 96 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=12.105
+ $Y=1.485 $X2=12.23 $Y2=1.66
r331 10 92 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=10.225
+ $Y=1.485 $X2=10.36 $Y2=2
r332 9 88 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.165
+ $Y=1.485 $X2=9.3 $Y2=2
r333 8 84 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=1.485 $X2=8.46 $Y2=2
r334 7 81 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=7.495
+ $Y=1.485 $X2=7.62 $Y2=2.34
r335 7 78 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=7.495
+ $Y=1.485 $X2=7.62 $Y2=1.66
r336 6 70 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=2.34
r337 6 67 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=1.66
r338 5 63 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2
r339 4 57 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=3.915
+ $Y=1.485 $X2=4.04 $Y2=2
r340 3 51 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=1.485 $X2=2.98 $Y2=2
r341 2 48 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.485 $X2=1.11 $Y2=2.34
r342 2 45 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.485 $X2=1.11 $Y2=1.66
r343 1 42 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.34
r344 1 39 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37
+ 39 43 45 49 51 55 59 63 67 68 72 76 80 84 86 90 92 94 97 98 100 101 102 118
+ 121 126 131 143 147 156 160 169 172 175 178 181 184 187 190 193 197
r214 196 197 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r215 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r216 184 185 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r217 181 182 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r218 175 176 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r219 173 176 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r220 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r221 164 197 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r222 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r223 161 193 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.315 $Y=0
+ $X2=12.2 $Y2=0
r224 161 163 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.315 $Y=0
+ $X2=12.65 $Y2=0
r225 160 196 3.66464 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=12.985 $Y=0
+ $X2=13.162 $Y2=0
r226 160 163 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.985 $Y=0
+ $X2=12.65 $Y2=0
r227 159 191 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r228 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r229 156 190 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.535 $Y=0
+ $X2=11.68 $Y2=0
r230 156 158 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.535 $Y=0
+ $X2=11.27 $Y2=0
r231 155 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r232 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r233 152 187 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.025 $Y=0
+ $X2=9.887 $Y2=0
r234 152 154 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.025 $Y=0
+ $X2=10.35 $Y2=0
r235 151 185 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.05 $Y2=0
r236 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r237 148 184 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.125 $Y=0
+ $X2=8.04 $Y2=0
r238 148 150 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=8.125 $Y=0
+ $X2=9.43 $Y2=0
r239 147 187 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=9.75 $Y=0
+ $X2=9.887 $Y2=0
r240 147 150 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.75 $Y=0 $X2=9.43
+ $Y2=0
r241 143 184 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=0
+ $X2=8.04 $Y2=0
r242 143 145 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.955 $Y=0
+ $X2=7.59 $Y2=0
r243 141 142 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r244 138 141 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r245 136 181 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.3
+ $Y2=0
r246 136 138 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.385 $Y=0
+ $X2=5.75 $Y2=0
r247 135 182 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r248 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r249 132 178 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.59 $Y=0
+ $X2=3.452 $Y2=0
r250 132 134 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.91
+ $Y2=0
r251 131 181 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.3
+ $Y2=0
r252 131 134 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=3.91 $Y2=0
r253 130 176 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.53 $Y2=0
r254 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r255 127 175 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=2.56 $Y2=0
r256 127 129 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=2.99 $Y2=0
r257 126 178 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.452 $Y2=0
r258 126 129 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=2.99 $Y2=0
r259 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r260 122 166 3.6634 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0
+ $X2=0.177 $Y2=0
r261 122 124 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0
+ $X2=0.69 $Y2=0
r262 121 169 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.025 $Y=0
+ $X2=1.14 $Y2=0
r263 121 124 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=0
+ $X2=0.69 $Y2=0
r264 117 164 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=12.65 $Y2=0
r265 117 191 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r266 117 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r267 116 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r268 116 151 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=9.43 $Y2=0
r269 116 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r270 115 185 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r271 115 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=6.67 $Y2=0
r272 115 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r273 114 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r274 113 114 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=5.745 $Y=0
+ $X2=6.21 $Y2=0
r275 113 182 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=5.745 $Y=0
+ $X2=5.29 $Y2=0
r276 113 138 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r277 112 135 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=3.445 $Y=0
+ $X2=3.91 $Y2=0
r278 112 130 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=3.445 $Y=0
+ $X2=2.99 $Y2=0
r279 112 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r280 111 173 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r281 111 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r282 111 169 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r283 102 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r284 102 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r285 100 154 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.695 $Y=0
+ $X2=10.35 $Y2=0
r286 100 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.695 $Y=0
+ $X2=10.78 $Y2=0
r287 99 158 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=10.865 $Y=0
+ $X2=11.27 $Y2=0
r288 99 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.865 $Y=0
+ $X2=10.78 $Y2=0
r289 97 141 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.67 $Y2=0
r290 97 98 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.925
+ $Y2=0
r291 96 145 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.095 $Y=0
+ $X2=7.59 $Y2=0
r292 96 98 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=6.925
+ $Y2=0
r293 92 196 3.25055 $w=2.1e-07 $l=1.15521e-07 $layer=LI1_cond $X=13.09 $Y=0.085
+ $X2=13.162 $Y2=0
r294 92 94 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=13.09 $Y=0.085
+ $X2=13.09 $Y2=0.38
r295 88 193 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0
r296 88 90 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0.38
r297 87 190 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=11.68 $Y2=0
r298 86 193 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.085 $Y=0
+ $X2=12.2 $Y2=0
r299 86 87 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.085 $Y=0
+ $X2=11.825 $Y2=0
r300 82 190 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0
r301 82 84 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0.39
r302 78 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.78 $Y=0.085
+ $X2=10.78 $Y2=0
r303 78 80 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.78 $Y=0.085
+ $X2=10.78 $Y2=0.39
r304 74 187 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.887 $Y=0.085
+ $X2=9.887 $Y2=0
r305 74 76 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=9.887 $Y=0.085
+ $X2=9.887 $Y2=0.39
r306 70 184 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=0.085
+ $X2=8.04 $Y2=0
r307 70 72 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.04 $Y=0.085
+ $X2=8.04 $Y2=0.38
r308 68 118 93.6302 $w=4.8e-07 $l=8.4e-07 $layer=POLY_cond $X=7.015 $Y=0.32
+ $X2=7.015 $Y2=1.16
r309 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.92
+ $Y=0.32 $X2=6.92 $Y2=0.32
r310 65 98 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=0.085
+ $X2=6.925 $Y2=0
r311 65 67 7.96542 $w=3.38e-07 $l=2.35e-07 $layer=LI1_cond $X=6.925 $Y=0.085
+ $X2=6.925 $Y2=0.32
r312 61 181 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0
r313 61 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0.38
r314 57 178 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.452 $Y=0.085
+ $X2=3.452 $Y2=0
r315 57 59 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=3.452 $Y=0.085
+ $X2=3.452 $Y2=0.39
r316 53 175 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r317 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.39
r318 52 172 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=1.66 $Y2=0
r319 51 175 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.56
+ $Y2=0
r320 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=1.805 $Y2=0
r321 47 172 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0
r322 47 49 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0.39
r323 46 169 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.255 $Y=0
+ $X2=1.14 $Y2=0
r324 45 172 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=1.66 $Y2=0
r325 45 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=1.255 $Y2=0
r326 41 169 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r327 41 43 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.38
r328 37 166 3.25179 $w=2.1e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.25 $Y=0.085
+ $X2=0.177 $Y2=0
r329 37 39 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.25 $Y=0.085
+ $X2=0.25 $Y2=0.38
r330 12 94 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.935
+ $Y=0.235 $X2=13.07 $Y2=0.38
r331 11 90 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=12.105
+ $Y=0.235 $X2=12.23 $Y2=0.38
r332 10 84 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=11.485
+ $Y=0.235 $X2=11.62 $Y2=0.39
r333 9 80 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.645
+ $Y=0.235 $X2=10.78 $Y2=0.39
r334 8 76 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=9.795
+ $Y=0.235 $X2=9.94 $Y2=0.39
r335 7 72 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.905
+ $Y=0.235 $X2=8.04 $Y2=0.38
r336 6 63 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.165
+ $Y=0.235 $X2=5.3 $Y2=0.38
r337 5 59 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.265
+ $Y=0.235 $X2=3.4 $Y2=0.39
r338 4 55 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.56 $Y2=0.39
r339 3 49 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.39
r340 2 43 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.235 $X2=1.11 $Y2=0.38
r341 1 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__NOR2_2_0/A 1 2 3 10
+ 12 15 17 19 22 24 26 29 31 33 36 38 40 42 44 50 52 57 65 71 73 74 75 76 77 86
+ 94 101 103 104
c161 75 0 7.35574e-20 $X=9.575 $Y=1.19
c162 65 0 1.4808e-19 $X=9.435 $Y=0.835
c163 44 0 9.09144e-20 $X=9.295 $Y=0.78
c164 22 0 1.19433e-19 $X=10.57 $Y=1.985
r165 99 101 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=11.2 $Y=1.16
+ $X2=11.41 $Y2=1.16
r166 96 99 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=10.99 $Y=1.16
+ $X2=11.2 $Y2=1.16
r167 92 94 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=10.305 $Y=1.16
+ $X2=10.57 $Y2=1.16
r168 89 92 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=10.15 $Y=1.16
+ $X2=10.305 $Y2=1.16
r169 77 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.435 $Y=1.19
+ $X2=10.29 $Y2=1.19
r170 76 86 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.005 $Y=1.19
+ $X2=11.15 $Y2=1.19
r171 76 77 0.705444 $w=1.4e-07 $l=5.7e-07 $layer=MET1_cond $X=11.005 $Y=1.19
+ $X2=10.435 $Y2=1.19
r172 75 79 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.575 $Y=1.19
+ $X2=9.43 $Y2=1.19
r173 74 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.145 $Y=1.19
+ $X2=10.29 $Y2=1.19
r174 74 75 0.705444 $w=1.4e-07 $l=5.7e-07 $layer=MET1_cond $X=10.145 $Y=1.19
+ $X2=9.575 $Y2=1.19
r175 73 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.2
+ $Y=1.16 $X2=11.2 $Y2=1.16
r176 73 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.15 $Y=1.19
+ $X2=11.15 $Y2=1.19
r177 71 92 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.305
+ $Y=1.16 $X2=10.305 $Y2=1.16
r178 71 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.29 $Y=1.19
+ $X2=10.29 $Y2=1.19
r179 68 104 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.435 $Y=1.58
+ $X2=9.435 $Y2=1.495
r180 68 104 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=9.435 $Y=1.47
+ $X2=9.435 $Y2=1.495
r181 67 68 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=9.435 $Y=1.19
+ $X2=9.435 $Y2=1.47
r182 67 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=1.19
+ $X2=9.43 $Y2=1.19
r183 65 103 3.22874 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=9.435 $Y=0.78
+ $X2=9.435 $Y2=0.905
r184 65 67 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=9.435 $Y=0.92
+ $X2=9.435 $Y2=1.19
r185 65 103 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=9.435 $Y=0.92
+ $X2=9.435 $Y2=0.905
r186 53 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.58
+ $X2=8.88 $Y2=1.58
r187 52 68 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.295 $Y=1.58
+ $X2=9.435 $Y2=1.58
r188 52 53 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=9.295 $Y=1.58
+ $X2=9.045 $Y2=1.58
r189 48 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.58
r190 48 50 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=2.34
r191 44 65 3.61619 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=9.295 $Y=0.78
+ $X2=9.435 $Y2=0.78
r192 44 46 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=9.295 $Y=0.78
+ $X2=8.88 $Y2=0.78
r193 43 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=1.58
+ $X2=8.04 $Y2=1.58
r194 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.715 $Y=1.58
+ $X2=8.88 $Y2=1.58
r195 42 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.715 $Y=1.58
+ $X2=8.205 $Y2=1.58
r196 38 55 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=1.665
+ $X2=8.04 $Y2=1.58
r197 38 40 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.04 $Y=1.665
+ $X2=8.04 $Y2=2.34
r198 34 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.41 $Y=1.325
+ $X2=11.41 $Y2=1.16
r199 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.41 $Y=1.325
+ $X2=11.41 $Y2=1.985
r200 31 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.41 $Y=0.995
+ $X2=11.41 $Y2=1.16
r201 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.41 $Y=0.995
+ $X2=11.41 $Y2=0.56
r202 27 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.99 $Y=1.325
+ $X2=10.99 $Y2=1.16
r203 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.99 $Y=1.325
+ $X2=10.99 $Y2=1.985
r204 24 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.99 $Y=0.995
+ $X2=10.99 $Y2=1.16
r205 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.99 $Y=0.995
+ $X2=10.99 $Y2=0.56
r206 20 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.57 $Y=1.325
+ $X2=10.57 $Y2=1.16
r207 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.57 $Y=1.325
+ $X2=10.57 $Y2=1.985
r208 17 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.57 $Y=0.995
+ $X2=10.57 $Y2=1.16
r209 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.57 $Y=0.995
+ $X2=10.57 $Y2=0.56
r210 13 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.15 $Y=1.325
+ $X2=10.15 $Y2=1.16
r211 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.15 $Y=1.325
+ $X2=10.15 $Y2=1.985
r212 10 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.15 $Y=0.995
+ $X2=10.15 $Y2=1.16
r213 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.15 $Y=0.995
+ $X2=10.15 $Y2=0.56
r214 3 57 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.485 $X2=8.88 $Y2=1.66
r215 3 50 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.485 $X2=8.88 $Y2=2.34
r216 2 55 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.905
+ $Y=1.485 $X2=8.04 $Y2=1.66
r217 2 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.905
+ $Y=1.485 $X2=8.04 $Y2=2.34
r218 1 46 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=8.745
+ $Y=0.235 $X2=8.88 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_0/A 1 2 3 10
+ 12 15 17 19 22 26 28 29 32 34 36 38 41 48 49 50 53 56 64
c120 48 0 1.29151e-19 $X=12.19 $Y=1.19
c121 41 0 1.19433e-19 $X=11.687 $Y=1.555
r122 63 64 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.44 $Y=1.16
+ $X2=12.86 $Y2=1.16
r123 60 63 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=12.23 $Y=1.16
+ $X2=12.44 $Y2=1.16
r124 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.69 $Y=1.19
+ $X2=11.69 $Y2=1.19
r125 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.835 $Y=1.19
+ $X2=11.69 $Y2=1.19
r126 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.03 $Y=1.19
+ $X2=12.175 $Y2=1.19
r127 49 50 0.241336 $w=1.4e-07 $l=1.95e-07 $layer=MET1_cond $X=12.03 $Y=1.19
+ $X2=11.835 $Y2=1.19
r128 48 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.23
+ $Y=1.16 $X2=12.23 $Y2=1.16
r129 48 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.175 $Y=1.19
+ $X2=12.175 $Y2=1.19
r130 44 53 15.2766 $w=2.13e-07 $l=2.85e-07 $layer=LI1_cond $X=11.687 $Y=0.905
+ $X2=11.687 $Y2=1.19
r131 42 53 13.6685 $w=2.13e-07 $l=2.55e-07 $layer=LI1_cond $X=11.687 $Y=1.445
+ $X2=11.687 $Y2=1.19
r132 41 42 0.884026 $w=2.15e-07 $l=1.1e-07 $layer=LI1_cond $X=11.687 $Y=1.555
+ $X2=11.687 $Y2=1.445
r133 38 41 25.5109 $w=2.18e-07 $l=4.87e-07 $layer=LI1_cond $X=11.2 $Y=1.555
+ $X2=11.687 $Y2=1.555
r134 35 36 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=11.365 $Y=0.82
+ $X2=11.2 $Y2=0.815
r135 34 44 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=11.58 $Y=0.82
+ $X2=11.687 $Y2=0.905
r136 34 35 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.58 $Y=0.82
+ $X2=11.365 $Y2=0.82
r137 30 36 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=11.2 $Y=0.725
+ $X2=11.2 $Y2=0.815
r138 30 32 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.2 $Y=0.725
+ $X2=11.2 $Y2=0.39
r139 28 36 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=11.035 $Y=0.815
+ $X2=11.2 $Y2=0.815
r140 28 29 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=11.035 $Y=0.815
+ $X2=10.525 $Y2=0.815
r141 24 29 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=10.36 $Y=0.725
+ $X2=10.525 $Y2=0.815
r142 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.36 $Y=0.725
+ $X2=10.36 $Y2=0.39
r143 20 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.86 $Y=1.325
+ $X2=12.86 $Y2=1.16
r144 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.86 $Y=1.325
+ $X2=12.86 $Y2=1.985
r145 17 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.86 $Y=0.995
+ $X2=12.86 $Y2=1.16
r146 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.86 $Y=0.995
+ $X2=12.86 $Y2=0.56
r147 13 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.44 $Y=1.325
+ $X2=12.44 $Y2=1.16
r148 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.44 $Y=1.325
+ $X2=12.44 $Y2=1.985
r149 10 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.44 $Y=0.995
+ $X2=12.44 $Y2=1.16
r150 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.44 $Y=0.995
+ $X2=12.44 $Y2=0.56
r151 3 38 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=11.065
+ $Y=1.485 $X2=11.2 $Y2=1.62
r152 2 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=11.065
+ $Y=0.235 $X2=11.2 $Y2=0.39
r153 1 26 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.225
+ $Y=0.235 $X2=10.36 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_1/Y 1 2 9 13
+ 20 22 23
r26 23 38 2.97463 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=0.69 $Y=1.55
+ $X2=0.69 $Y2=1.485
r27 23 38 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=0.65 $Y=1.465
+ $X2=0.65 $Y2=1.485
r28 22 23 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.65 $Y=1.19
+ $X2=0.65 $Y2=1.465
r29 20 36 2.80002 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.69 $Y=0.825 $X2=0.69
+ $Y2=0.885
r30 20 22 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.65 $Y=0.91
+ $X2=0.65 $Y2=1.19
r31 20 36 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.65 $Y=0.91
+ $X2=0.65 $Y2=0.885
r32 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.66
+ $X2=0.69 $Y2=2.34
r33 11 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=1.65 $X2=0.69
+ $Y2=1.55
r34 11 13 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.69 $Y=1.65 $X2=0.69
+ $Y2=1.66
r35 7 20 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.69 $Y=0.72
+ $X2=0.69 $Y2=0.825
r36 7 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.69 $Y=0.72 $X2=0.69
+ $Y2=0.38
r37 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.485 $X2=0.69 $Y2=2.34
r38 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.485 $X2=0.69 $Y2=1.66
r39 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#
+ 1 2 3 12 14 15 16 17 18 20 22
r48 20 29 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=3.452 $Y=1.665
+ $X2=3.452 $Y2=1.56
r49 20 22 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=3.452 $Y=1.665
+ $X2=3.452 $Y2=2.3
r50 19 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=1.56
+ $X2=2.56 $Y2=1.56
r51 18 29 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=3.315 $Y=1.56
+ $X2=3.452 $Y2=1.56
r52 18 19 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=3.315 $Y=1.56
+ $X2=2.645 $Y2=1.56
r53 17 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=2.295
+ $X2=2.56 $Y2=2.38
r54 16 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.56 $Y=1.665
+ $X2=2.56 $Y2=1.56
r55 16 17 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.56 $Y=1.665
+ $X2=2.56 $Y2=2.295
r56 14 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=2.38
+ $X2=2.56 $Y2=2.38
r57 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=2.38
+ $X2=1.805 $Y2=2.38
r58 10 15 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.655 $Y=2.295
+ $X2=1.805 $Y2=2.38
r59 10 12 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=1.655 $Y=2.295
+ $X2=1.655 $Y2=2
r60 3 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.485 $X2=3.4 $Y2=1.62
r61 3 22 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.485 $X2=3.4 $Y2=2.3
r62 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.485 $X2=2.56 $Y2=2.3
r63 2 25 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.485 $X2=2.56 $Y2=1.62
r64 1 12 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#
+ 1 2 3 10 12 14 16 17 18 22
r48 20 22 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=11.685 $Y=2.295
+ $X2=11.685 $Y2=2
r49 19 29 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.865 $Y=2.38
+ $X2=10.78 $Y2=2.38
r50 18 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=11.535 $Y=2.38
+ $X2=11.685 $Y2=2.295
r51 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.535 $Y=2.38
+ $X2=10.865 $Y2=2.38
r52 17 29 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.78 $Y=2.295
+ $X2=10.78 $Y2=2.38
r53 16 27 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=10.78 $Y=1.665
+ $X2=10.78 $Y2=1.56
r54 16 17 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.78 $Y=1.665
+ $X2=10.78 $Y2=2.295
r55 15 25 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=10.025 $Y=1.56
+ $X2=9.887 $Y2=1.56
r56 14 27 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=10.695 $Y=1.56
+ $X2=10.78 $Y2=1.56
r57 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=10.695 $Y=1.56
+ $X2=10.025 $Y2=1.56
r58 10 25 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=9.887 $Y=1.665
+ $X2=9.887 $Y2=1.56
r59 10 12 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=9.887 $Y=1.665
+ $X2=9.887 $Y2=2.3
r60 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=11.485
+ $Y=1.485 $X2=11.62 $Y2=2
r61 2 29 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=10.645
+ $Y=1.485 $X2=10.78 $Y2=2.3
r62 2 27 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=10.645
+ $Y=1.485 $X2=10.78 $Y2=1.62
r63 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.795
+ $Y=1.485 $X2=9.94 $Y2=1.62
r64 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.795
+ $Y=1.485 $X2=9.94 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%SKY130_FD_SC_HD__INV_2_0/Y 1 2 9 13
+ 20 22 23
r26 23 38 2.97463 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=12.65 $Y=1.55
+ $X2=12.65 $Y2=1.485
r27 23 38 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=12.69 $Y=1.465
+ $X2=12.69 $Y2=1.485
r28 22 23 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=12.69 $Y=1.19
+ $X2=12.69 $Y2=1.465
r29 20 36 2.80002 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=12.65 $Y=0.825
+ $X2=12.65 $Y2=0.885
r30 20 22 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=12.69 $Y=0.91
+ $X2=12.69 $Y2=1.19
r31 20 36 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=12.69 $Y=0.91
+ $X2=12.69 $Y2=0.885
r32 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=12.65 $Y=1.66
+ $X2=12.65 $Y2=2.34
r33 11 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=12.65 $Y=1.65
+ $X2=12.65 $Y2=1.55
r34 11 13 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=12.65 $Y=1.65
+ $X2=12.65 $Y2=1.66
r35 7 20 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=12.65 $Y=0.72
+ $X2=12.65 $Y2=0.825
r36 7 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=12.65 $Y=0.72
+ $X2=12.65 $Y2=0.38
r37 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.515
+ $Y=1.485 $X2=12.65 $Y2=2.34
r38 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=12.515
+ $Y=1.485 $X2=12.65 $Y2=1.66
r39 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.515
+ $Y=0.235 $X2=12.65 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#
+ 1 2 3 10 12 13 14 18 23
c49 23 0 5.77853e-20 $X=4.205 $Y=0.37
r50 21 23 8.37661 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=0.37
+ $X2=4.205 $Y2=0.37
r51 16 18 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=5.725 $Y=0.715
+ $X2=5.725 $Y2=0.38
r52 15 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.045 $Y=0.8
+ $X2=4.92 $Y2=0.8
r53 14 16 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=5.555 $Y=0.8
+ $X2=5.725 $Y2=0.715
r54 14 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.555 $Y=0.8
+ $X2=5.045 $Y2=0.8
r55 13 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=0.715
+ $X2=4.92 $Y2=0.8
r56 12 25 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.92 $Y=0.465
+ $X2=4.92 $Y2=0.36
r57 12 13 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.92 $Y=0.465
+ $X2=4.92 $Y2=0.715
r58 10 25 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.795 $Y=0.36
+ $X2=4.92 $Y2=0.36
r59 10 23 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.795 $Y=0.36
+ $X2=4.205 $Y2=0.36
r60 3 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.38
r61 2 27 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.72
r62 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.38
r63 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.235 $X2=4.04 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MACRO_SPARECELL%XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#
+ 1 2 3 12 14 15 16 17 25 26
c55 25 0 5.77853e-20 $X=9.3 $Y=0.38
r56 25 26 8.37661 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.3 $Y=0.37
+ $X2=9.135 $Y2=0.37
r57 19 21 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=0.36
+ $X2=8.42 $Y2=0.36
r58 19 26 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=8.545 $Y=0.36
+ $X2=9.135 $Y2=0.36
r59 17 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.715
+ $X2=8.42 $Y2=0.8
r60 16 21 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=8.42 $Y=0.465
+ $X2=8.42 $Y2=0.36
r61 16 17 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=8.42 $Y=0.465
+ $X2=8.42 $Y2=0.715
r62 14 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=0.8
+ $X2=8.42 $Y2=0.8
r63 14 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.295 $Y=0.8
+ $X2=7.785 $Y2=0.8
r64 10 15 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=7.615 $Y=0.715
+ $X2=7.785 $Y2=0.8
r65 10 12 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=7.615 $Y=0.715
+ $X2=7.615 $Y2=0.38
r66 3 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=9.165
+ $Y=0.235 $X2=9.3 $Y2=0.38
r67 2 23 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.235 $X2=8.46 $Y2=0.72
r68 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.235 $X2=8.46 $Y2=0.38
r69 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=7.495
+ $Y=0.235 $X2=7.62 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a21bo_2.pex.spice
* Created: Thu Aug 27 14:00:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BO_2%A_79_21# 1 2 9 13 17 21 24 25 26 29 32 33 35
+ 36 37 38 44 46 47 50 55
c103 29 0 2.81618e-19 $X=0.735 $Y=1.16
c104 21 0 9.19488e-20 $X=0.9 $Y=1.985
r105 52 55 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.43 $Y=0.73
+ $X2=2.575 $Y2=0.73
r106 48 50 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.14 $Y=1.59
+ $X2=2.43 $Y2=1.59
r107 46 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=1.505
+ $X2=2.43 $Y2=1.59
r108 45 52 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.43 $Y=0.825 $X2=2.43
+ $Y2=0.73
r109 45 46 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.43 $Y=0.825
+ $X2=2.43 $Y2=1.505
r110 42 47 5.16603 $w=2.1e-07 $l=1.2339e-07 $layer=LI1_cond $X=2.14 $Y=1.895
+ $X2=2.1 $Y2=2
r111 42 44 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.14 $Y=1.895
+ $X2=2.14 $Y2=1.77
r112 41 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.675
+ $X2=2.14 $Y2=1.59
r113 41 44 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.14 $Y=1.675
+ $X2=2.14 $Y2=1.77
r114 38 47 5.16603 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=2.1 $Y=2.105
+ $X2=2.1 $Y2=2
r115 38 40 0.244 $w=2.5e-07 $l=5e-09 $layer=LI1_cond $X=2.1 $Y=2.105 $X2=2.1
+ $Y2=2.11
r116 36 47 1.34256 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.975 $Y=2 $X2=2.1
+ $Y2=2
r117 36 37 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.975 $Y=2
+ $X2=1.285 $Y2=2
r118 35 37 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.2 $Y=1.895
+ $X2=1.285 $Y2=2
r119 34 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.895
r120 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=1.2 $Y2=1.665
r121 32 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=0.9 $Y2=1.58
r122 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.735
+ $Y=1.16 $X2=0.735 $Y2=1.16
r123 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.735 $Y=1.495
+ $X2=0.9 $Y2=1.58
r124 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.735 $Y=1.495
+ $X2=0.735 $Y2=1.16
r125 25 30 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.825 $Y=1.16
+ $X2=0.735 $Y2=1.16
r126 25 26 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.825 $Y=1.16
+ $X2=0.9 $Y2=1.16
r127 23 30 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.735 $Y2=1.16
r128 23 24 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.47 $Y2=1.16
r129 19 26 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.9 $Y=1.295
+ $X2=0.9 $Y2=1.16
r130 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.9 $Y=1.295
+ $X2=0.9 $Y2=1.985
r131 15 26 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.9 $Y=1.025
+ $X2=0.9 $Y2=1.16
r132 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.9 $Y=1.025
+ $X2=0.9 $Y2=0.56
r133 11 24 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r134 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.985
r135 7 24 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r136 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
r137 2 44 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.14 $Y2=1.77
r138 2 40 600 $w=1.7e-07 $l=6.84653e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.14 $Y2=2.11
r139 1 55 182 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.575 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%B1_N 3 6 8 11 13
c36 13 0 2.03766e-19 $X=1.44 $Y=0.995
c37 11 0 1.99872e-19 $X=1.44 $Y=1.16
c38 6 0 1.34885e-19 $X=1.41 $Y=1.695
r39 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.16
+ $X2=1.44 $Y2=1.325
r40 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.16
+ $X2=1.44 $Y2=0.995
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.44
+ $Y=1.16 $X2=1.44 $Y2=1.16
r42 8 12 11.3257 $w=3.07e-07 $l=2.85e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.44 $Y2=1.16
r43 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.41 $Y=1.695
+ $X2=1.41 $Y2=1.325
r44 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.41 $Y=0.675
+ $X2=1.41 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%A_297_93# 1 2 7 9 12 15 17 21 26 31
c56 26 0 9.19488e-20 $X=1.78 $Y=1.64
c57 7 0 8.15699e-20 $X=2.35 $Y=0.99
r58 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.16 $X2=2.09 $Y2=1.16
r59 28 31 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.78 $Y=1.16 $X2=2.09
+ $Y2=1.16
r60 24 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.62 $Y=1.64
+ $X2=1.78 $Y2=1.64
r61 19 21 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.62 $Y=0.74
+ $X2=1.78 $Y2=0.74
r62 17 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=1.555
+ $X2=1.78 $Y2=1.64
r63 16 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.16
r64 16 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.555
r65 15 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0.995
+ $X2=1.78 $Y2=1.16
r66 14 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.825
+ $X2=1.78 $Y2=0.74
r67 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.78 $Y=0.825
+ $X2=1.78 $Y2=0.995
r68 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.35 $Y=1.325
+ $X2=2.35 $Y2=1.985
r69 7 10 21.5811 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.35 $Y=1.157
+ $X2=2.35 $Y2=1.325
r70 7 32 44.7854 $w=3.35e-07 $l=2.6e-07 $layer=POLY_cond $X=2.35 $Y=1.157
+ $X2=2.09 $Y2=1.157
r71 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.35 $Y=0.99 $X2=2.35
+ $Y2=0.56
r72 2 24 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.64
r73 1 19 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.465 $X2=1.62 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%A1 3 7 8 11 12 13
c38 11 0 1.34089e-19 $X=2.77 $Y=1.16
r39 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.16
+ $X2=2.77 $Y2=0.995
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.16 $X2=2.77 $Y2=1.16
r41 8 12 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.892 $Y=1.53
+ $X2=2.892 $Y2=1.16
r42 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.83 $Y=0.56 $X2=2.83
+ $Y2=0.995
r43 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.325
+ $X2=2.77 $Y2=1.16
r44 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.77 $Y=1.325 $X2=2.77
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%A2 3 6 8 11 13 18
r26 12 18 2.21853 $w=6.18e-07 $l=1.15e-07 $layer=LI1_cond $X=3.355 $Y=1.305
+ $X2=3.47 $Y2=1.305
r27 11 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.302 $Y=1.16
+ $X2=3.302 $Y2=1.325
r28 11 13 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.302 $Y=1.16
+ $X2=3.302 $Y2=0.995
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.355
+ $Y=1.16 $X2=3.355 $Y2=1.16
r30 8 18 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=3.475 $Y=1.305
+ $X2=3.47 $Y2=1.305
r31 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.19 $Y=1.985
+ $X2=3.19 $Y2=1.325
r32 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.19 $Y=0.56 $X2=3.19
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%VPWR 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r64 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r68 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 35 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=2.72
+ $X2=1.205 $Y2=2.72
r73 32 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.37 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 31 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 28 44 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r77 28 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=2.72
+ $X2=1.205 $Y2=2.72
r79 27 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.04 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 25 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r82 23 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.895 $Y=2.72
+ $X2=2.53 $Y2=2.72
r83 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=2.72
+ $X2=2.98 $Y2=2.72
r84 22 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.065 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=2.72
+ $X2=2.98 $Y2=2.72
r86 18 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.635
+ $X2=2.98 $Y2=2.72
r87 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.98 $Y=2.635
+ $X2=2.98 $Y2=2.36
r88 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=2.635
+ $X2=1.205 $Y2=2.72
r89 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.205 $Y=2.635
+ $X2=1.205 $Y2=2.36
r90 10 44 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r91 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r92 3 20 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.485 $X2=2.98 $Y2=2.36
r93 2 16 600 $w=1.7e-07 $l=9.83298e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.485 $X2=1.205 $Y2=2.36
r94 1 12 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%X 1 2 7 9 11 13 15 24 27
c38 15 0 2.40354e-20 $X=0.685 $Y=2.26
c39 13 0 1.10849e-19 $X=0.722 $Y=2.005
c40 9 0 1.22196e-19 $X=0.685 $Y=0.715
c41 2 0 2.14206e-20 $X=0.545 $Y=1.485
r42 24 27 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.92
+ $X2=0.265 $Y2=1.835
r43 24 27 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=1.81
+ $X2=0.265 $Y2=1.835
r44 18 24 46.3483 $w=2.28e-07 $l=9.25e-07 $layer=LI1_cond $X=0.265 $Y=0.885
+ $X2=0.265 $Y2=1.81
r45 13 23 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.722 $Y=2.005
+ $X2=0.722 $Y2=1.92
r46 13 15 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.722 $Y=2.005
+ $X2=0.722 $Y2=2.26
r47 9 18 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.685 $Y=0.8
+ $X2=0.265 $Y2=0.8
r48 9 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.685 $Y=0.715
+ $X2=0.685 $Y2=0.4
r49 8 24 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.38 $Y=1.92
+ $X2=0.265 $Y2=1.92
r50 7 23 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.595 $Y=1.92
+ $X2=0.722 $Y2=1.92
r51 7 8 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.595 $Y=1.92
+ $X2=0.38 $Y2=1.92
r52 2 23 600 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.685 $Y2=1.92
r53 2 15 600 $w=1.7e-07 $l=8.42096e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.685 $Y2=2.26
r54 1 11 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.685 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%A_485_297# 1 2 9 14 16
c28 9 0 1.34089e-19 $X=3.235 $Y=1.93
r29 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.93
+ $X2=2.56 $Y2=1.93
r30 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=1.93 $X2=3.4
+ $Y2=1.93
r31 9 10 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.235 $Y=1.93
+ $X2=2.725 $Y2=1.93
r32 2 16 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=1.485 $X2=3.4 $Y2=2
r33 1 14 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.425
+ $Y=1.485 $X2=2.56 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_2%VGND 1 2 3 4 13 15 19 23 25 27 30 31 32 38
+ 42 51 55
r53 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r55 46 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r56 46 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r57 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 43 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.14
+ $Y2=0
r59 43 45 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.99
+ $Y2=0
r60 42 54 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.457
+ $Y2=0
r61 42 45 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=2.99
+ $Y2=0
r62 41 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r63 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r64 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.14
+ $Y2=0
r65 38 40 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.61
+ $Y2=0
r66 37 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r67 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r68 34 48 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r69 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r70 32 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r71 32 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r72 30 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.69
+ $Y2=0
r73 30 31 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.12
+ $Y2=0
r74 29 40 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.61
+ $Y2=0
r75 29 31 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.12
+ $Y2=0
r76 25 54 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.4 $Y=0.085
+ $X2=3.457 $Y2=0
r77 25 27 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.4 $Y=0.085
+ $X2=3.4 $Y2=0.74
r78 21 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r79 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.38
r80 17 31 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085 $X2=1.12
+ $Y2=0
r81 17 19 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r82 13 48 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r83 13 15 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.38
r84 4 27 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.235 $X2=3.4 $Y2=0.74
r85 3 23 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.235 $X2=2.14 $Y2=0.38
r86 2 19 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.235 $X2=1.115 $Y2=0.36
r87 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


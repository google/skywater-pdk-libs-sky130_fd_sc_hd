* File: sky130_fd_sc_hd__sdfxtp_4.spice.pex
* Created: Thu Aug 27 14:47:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%CLK 1 2 3 5 6 8 11 13
c42 1 0 2.71124e-20 $X=0.31 $Y=1.325
r43 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.475 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=2.135
r47 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r50 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_27_47# 1 2 9 13 17 19 20 25 29 31 35 39
+ 43 44 45 49 50 52 55 56 57 58 59 60 69 75 78 79 80 82 86
c246 86 0 1.77381e-19 $X=6.7 $Y=1.41
c247 52 0 8.70797e-20 $X=0.76 $Y=1.235
c248 50 0 1.81794e-19 $X=0.73 $Y=1.795
c249 45 0 3.29888e-20 $X=0.615 $Y=1.88
c250 29 0 4.21632e-20 $X=6.705 $Y=2.275
c251 19 0 1.57835e-19 $X=5.015 $Y=1.32
r252 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.41
+ $X2=6.7 $Y2=1.575
r253 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=1.41 $X2=6.7 $Y2=1.41
r254 82 85 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.7 $Y=1.32 $X2=6.7
+ $Y2=1.41
r255 78 81 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=1.74
+ $X2=5.15 $Y2=1.905
r256 78 80 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=1.74
+ $X2=5.15 $Y2=1.575
r257 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.15
+ $Y=1.74 $X2=5.15 $Y2=1.74
r258 74 75 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=0.89 $Y=1.235
+ $X2=0.895 $Y2=1.235
r259 70 86 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.71 $Y=1.87
+ $X2=6.71 $Y2=1.41
r260 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=1.87
+ $X2=6.71 $Y2=1.87
r261 66 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.3 $Y=1.87 $X2=5.3
+ $Y2=1.87
r262 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.7 $Y=1.87 $X2=0.7
+ $Y2=1.87
r263 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.445 $Y=1.87
+ $X2=5.3 $Y2=1.87
r264 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.565 $Y=1.87
+ $X2=6.71 $Y2=1.87
r265 59 60 1.38614 $w=1.4e-07 $l=1.12e-06 $layer=MET1_cond $X=6.565 $Y=1.87
+ $X2=5.445 $Y2=1.87
r266 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.845 $Y=1.87
+ $X2=0.7 $Y2=1.87
r267 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.155 $Y=1.87
+ $X2=5.3 $Y2=1.87
r268 57 58 5.33415 $w=1.4e-07 $l=4.31e-06 $layer=MET1_cond $X=5.155 $Y=1.87
+ $X2=0.845 $Y2=1.87
r269 53 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r270 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r271 50 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r272 50 52 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r273 49 56 6.0623 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=0.97
r274 49 52 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=1.235
r275 47 56 9.38461 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=0.805
+ $X2=0.712 $Y2=0.97
r276 46 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r277 45 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r278 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.35 $Y2=1.88
r279 43 47 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.712 $Y2=0.805
r280 43 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r281 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r282 37 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r283 33 35 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.35 $Y=1.245
+ $X2=7.35 $Y2=0.415
r284 32 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.835 $Y=1.32
+ $X2=6.7 $Y2=1.32
r285 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.275 $Y=1.32
+ $X2=7.35 $Y2=1.245
r286 31 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.275 $Y=1.32
+ $X2=6.835 $Y2=1.32
r287 29 87 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.705 $Y=2.275
+ $X2=6.705 $Y2=1.575
r288 25 81 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.09 $Y=2.275
+ $X2=5.09 $Y2=1.905
r289 21 80 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.09 $Y=1.395
+ $X2=5.09 $Y2=1.575
r290 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.015 $Y=1.32
+ $X2=5.09 $Y2=1.395
r291 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=5.015 $Y=1.32
+ $X2=4.705 $Y2=1.32
r292 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.63 $Y=1.245
+ $X2=4.705 $Y2=1.32
r293 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.63 $Y=1.245
+ $X2=4.63 $Y2=0.415
r294 11 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=1.235
r295 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=2.135
r296 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r297 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r298 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r299 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%SCE 3 7 11 15 19 20 22 23 24 28 29 32 33
c110 24 0 1.66251e-19 $X=3.085 $Y=0.7
c111 22 0 1.76484e-19 $X=2.475 $Y=0.7
r112 35 36 3.41038 $w=2.12e-07 $l=1.5e-08 $layer=POLY_cond $X=1.835 $Y=1.52
+ $X2=1.85 $Y2=1.52
r113 31 33 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.51
r114 31 32 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.7
r115 29 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=0.95
+ $X2=3.17 $Y2=0.785
r116 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=0.95 $X2=3.17 $Y2=0.95
r117 26 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0.785
+ $X2=3.17 $Y2=0.95
r118 25 32 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.65 $Y=0.7
+ $X2=2.562 $Y2=0.7
r119 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=0.7
+ $X2=3.17 $Y2=0.785
r120 24 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.085 $Y=0.7
+ $X2=2.65 $Y2=0.7
r121 22 32 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=2.562 $Y2=0.7
r122 22 23 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=1.95 $Y2=0.7
r123 20 38 88.6698 $w=2.12e-07 $l=3.9e-07 $layer=POLY_cond $X=1.865 $Y=1.52
+ $X2=2.255 $Y2=1.52
r124 20 36 3.41038 $w=2.12e-07 $l=1.5e-08 $layer=POLY_cond $X=1.865 $Y=1.52
+ $X2=1.85 $Y2=1.52
r125 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=1.52 $X2=1.865 $Y2=1.52
r126 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=0.785
+ $X2=1.95 $Y2=0.7
r127 17 19 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.865 $Y=0.785
+ $X2=1.865 $Y2=1.52
r128 15 40 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.23 $Y=0.445
+ $X2=3.23 $Y2=0.785
r129 9 38 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.255 $Y=1.655
+ $X2=2.255 $Y2=1.52
r130 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.255 $Y=1.655
+ $X2=2.255 $Y2=2.165
r131 5 36 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.85 $Y=1.385
+ $X2=1.85 $Y2=1.52
r132 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.85 $Y=1.385 $X2=1.85
+ $Y2=0.445
r133 1 35 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.835 $Y=1.655
+ $X2=1.835 $Y2=1.52
r134 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.835 $Y=1.655
+ $X2=1.835 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_299_47# 1 2 9 13 16 19 21 24 25 28 32 34
+ 38 39 41 43 44
c126 43 0 1.84493e-19 $X=3.19 $Y=1.52
c127 39 0 1.12087e-19 $X=2.3 $Y=1.04
c128 24 0 1.60762e-19 $X=2.205 $Y=1.86
c129 9 0 1.20015e-19 $X=2.36 $Y=0.445
r130 44 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.52
+ $X2=3.19 $Y2=1.685
r131 43 46 9.59627 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.177 $Y=1.52
+ $X2=3.177 $Y2=1.685
r132 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.52 $X2=3.19 $Y2=1.52
r133 39 48 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.3 $Y=1.04
+ $X2=2.3 $Y2=0.905
r134 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.04 $X2=2.3 $Y2=1.04
r135 35 38 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.205 $Y=1.04
+ $X2=2.3 $Y2=1.04
r136 29 32 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.52 $Y=0.36
+ $X2=1.64 $Y2=0.36
r137 28 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.165 $Y=1.86
+ $X2=3.165 $Y2=1.685
r138 26 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=1.967
+ $X2=2.205 $Y2=1.967
r139 25 28 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.08 $Y=1.967
+ $X2=3.165 $Y2=1.86
r140 25 26 42.3456 $w=2.13e-07 $l=7.9e-07 $layer=LI1_cond $X=3.08 $Y=1.967
+ $X2=2.29 $Y2=1.967
r141 24 41 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.205 $Y=1.86
+ $X2=2.205 $Y2=1.967
r142 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=1.125
+ $X2=2.205 $Y2=1.04
r143 23 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.205 $Y=1.125
+ $X2=2.205 $Y2=1.86
r144 22 34 1.46632 $w=2.15e-07 $l=1.38e-07 $layer=LI1_cond $X=1.71 $Y=1.967
+ $X2=1.572 $Y2=1.967
r145 21 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=1.967
+ $X2=2.205 $Y2=1.967
r146 21 22 21.9768 $w=2.13e-07 $l=4.1e-07 $layer=LI1_cond $X=2.12 $Y=1.967
+ $X2=1.71 $Y2=1.967
r147 17 34 5.02022 $w=2.22e-07 $l=1.08e-07 $layer=LI1_cond $X=1.572 $Y=2.075
+ $X2=1.572 $Y2=1.967
r148 17 19 4.1907 $w=2.73e-07 $l=1e-07 $layer=LI1_cond $X=1.572 $Y=2.075
+ $X2=1.572 $Y2=2.175
r149 16 34 5.02022 $w=2.22e-07 $l=1.30434e-07 $layer=LI1_cond $X=1.52 $Y=1.86
+ $X2=1.572 $Y2=1.967
r150 15 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.445
+ $X2=1.52 $Y2=0.36
r151 15 16 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.52 $Y=0.445
+ $X2=1.52 $Y2=1.86
r152 13 52 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.145 $Y=2.165
+ $X2=3.145 $Y2=1.685
r153 9 48 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.36 $Y=0.445
+ $X2=2.36 $Y2=0.905
r154 2 19 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.845 $X2=1.625 $Y2=2.175
r155 1 32 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.64 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%D 3 7 9 12 19
c49 19 0 2.8857e-19 $X=2.64 $Y=1.53
r50 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.52
+ $X2=2.71 $Y2=1.685
r51 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.52
+ $X2=2.71 $Y2=1.355
r52 12 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.52 $X2=2.71 $Y2=1.52
r53 9 19 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=1.52 $X2=2.64
+ $Y2=1.52
r54 7 14 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.75 $Y=0.445
+ $X2=2.75 $Y2=1.355
r55 3 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.725 $Y=2.165
+ $X2=2.725 $Y2=1.685
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%SCD 3 7 9 12
c48 7 0 1.84493e-19 $X=3.61 $Y=2.165
c49 3 0 1.66251e-19 $X=3.61 $Y=0.445
r50 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.355
+ $X2=3.67 $Y2=1.52
r51 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.355
+ $X2=3.67 $Y2=1.19
r52 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.67
+ $Y=1.355 $X2=3.67 $Y2=1.355
r53 9 13 4.62998 $w=6.18e-07 $l=2.4e-07 $layer=LI1_cond $X=3.91 $Y=1.345
+ $X2=3.67 $Y2=1.345
r54 7 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.61 $Y=2.165
+ $X2=3.61 $Y2=1.52
r55 3 14 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.61 $Y=0.445
+ $X2=3.61 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_193_47# 1 2 9 13 14 16 19 23 24 27 30 33
+ 37 38 40 41 42 43 46 52 59 60 61 66
c214 66 0 1.77381e-19 $X=6.93 $Y=0.87
c215 42 0 1.57835e-19 $X=6.565 $Y=0.85
r216 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=0.87 $X2=6.93 $Y2=0.87
r217 63 66 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.835 $Y=0.87
+ $X2=6.93 $Y2=0.87
r218 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=0.87
+ $X2=5.05 $Y2=0.705
r219 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=0.87 $X2=5.05 $Y2=0.87
r220 53 67 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.71 $Y=0.87
+ $X2=6.93 $Y2=0.87
r221 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=0.85
+ $X2=6.71 $Y2=0.85
r222 50 60 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.84 $Y=0.87
+ $X2=5.05 $Y2=0.87
r223 50 80 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=0.87
+ $X2=4.675 $Y2=0.87
r224 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.84 $Y=0.85
+ $X2=4.84 $Y2=0.85
r225 46 75 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.132 $Y=0.85
+ $X2=1.132 $Y2=1.96
r226 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=0.85
+ $X2=1.14 $Y2=0.85
r227 43 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.985 $Y=0.85
+ $X2=4.84 $Y2=0.85
r228 42 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.565 $Y=0.85
+ $X2=6.71 $Y2=0.85
r229 42 43 1.95544 $w=1.4e-07 $l=1.58e-06 $layer=MET1_cond $X=6.565 $Y=0.85
+ $X2=4.985 $Y2=0.85
r230 41 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.285 $Y=0.85
+ $X2=1.14 $Y2=0.85
r231 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.695 $Y=0.85
+ $X2=4.84 $Y2=0.85
r232 40 41 4.22029 $w=1.4e-07 $l=3.41e-06 $layer=MET1_cond $X=4.695 $Y=0.85
+ $X2=1.285 $Y2=0.85
r233 38 69 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=7.21 $Y=1.74
+ $X2=7.125 $Y2=1.74
r234 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=1.74 $X2=7.21 $Y2=1.74
r235 34 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.07 $Y=1.74
+ $X2=7.21 $Y2=1.74
r236 33 67 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.975 $Y=0.87
+ $X2=6.93 $Y2=0.87
r237 32 46 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=1.132 $Y=0.715
+ $X2=1.132 $Y2=0.85
r238 30 32 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.13 $Y=0.51
+ $X2=1.13 $Y2=0.715
r239 27 34 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.07 $Y=1.575
+ $X2=7.07 $Y2=1.74
r240 26 33 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.07 $Y=1.035
+ $X2=6.975 $Y2=0.87
r241 26 27 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.07 $Y=1.035
+ $X2=7.07 $Y2=1.575
r242 24 57 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.64 $Y=1.74
+ $X2=4.64 $Y2=1.875
r243 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=1.74 $X2=4.64 $Y2=1.74
r244 21 80 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=1.035
+ $X2=4.675 $Y2=0.87
r245 21 23 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.675 $Y=1.035
+ $X2=4.675 $Y2=1.74
r246 17 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.125 $Y=1.875
+ $X2=7.125 $Y2=1.74
r247 17 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.125 $Y=1.875
+ $X2=7.125 $Y2=2.275
r248 14 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.835 $Y=0.705
+ $X2=6.835 $Y2=0.87
r249 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.835 $Y=0.705
+ $X2=6.835 $Y2=0.415
r250 13 61 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.11 $Y=0.415
+ $X2=5.11 $Y2=0.705
r251 9 57 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.625 $Y=2.275
+ $X2=4.625 $Y2=1.875
r252 2 75 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.815 $X2=1.105 $Y2=1.96
r253 1 30 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_1099_183# 1 2 9 13 15 18 21 23 29 30 32
+ 33 36
r95 35 36 5.54023 $w=2.61e-07 $l=3e-08 $layer=POLY_cond $X=5.57 $Y=0.93 $X2=5.6
+ $Y2=0.93
r96 32 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.4 $Y=2.3 $X2=6.4
+ $Y2=2.135
r97 27 36 24.0077 $w=2.61e-07 $l=1.3e-07 $layer=POLY_cond $X=5.73 $Y=0.93
+ $X2=5.6 $Y2=0.93
r98 26 29 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=0.93
+ $X2=5.815 $Y2=0.93
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=0.93 $X2=5.73 $Y2=0.93
r100 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.445 $Y=0.45
+ $X2=6.57 $Y2=0.45
r101 19 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.36 $Y=1.065
+ $X2=6.36 $Y2=0.915
r102 19 33 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.36 $Y=1.065
+ $X2=6.36 $Y2=2.135
r103 18 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.36 $Y=0.765
+ $X2=6.36 $Y2=0.915
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.36 $Y=0.535
+ $X2=6.445 $Y2=0.45
r105 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.36 $Y=0.535
+ $X2=6.36 $Y2=0.765
r106 15 30 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=0.915
+ $X2=6.36 $Y2=0.915
r107 15 29 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.275 $Y=0.915
+ $X2=5.815 $Y2=0.915
r108 11 36 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.6 $Y=0.795
+ $X2=5.6 $Y2=0.93
r109 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.6 $Y=0.795
+ $X2=5.6 $Y2=0.445
r110 7 35 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.57 $Y=1.065
+ $X2=5.57 $Y2=0.93
r111 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.57 $Y=1.065
+ $X2=5.57 $Y2=2.275
r112 2 32 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.735 $X2=6.44 $Y2=2.3
r113 1 23 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.405
+ $Y=0.235 $X2=6.57 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_940_413# 1 2 8 11 13 15 18 20 21 22 26 31
+ 33 35
c109 31 0 1.42307e-19 $X=5.39 $Y=1.315
r110 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.02
+ $Y=1.41 $X2=6.02 $Y2=1.41
r111 35 37 17.1405 $w=2.42e-07 $l=3.4e-07 $layer=LI1_cond $X=5.68 $Y=1.41
+ $X2=6.02 $Y2=1.41
r112 32 35 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=1.575
+ $X2=5.68 $Y2=1.41
r113 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.68 $Y=1.575
+ $X2=5.68 $Y2=2.19
r114 31 35 14.6198 $w=2.42e-07 $l=2.9e-07 $layer=LI1_cond $X=5.39 $Y=1.41
+ $X2=5.68 $Y2=1.41
r115 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.39 $Y=0.535
+ $X2=5.39 $Y2=1.315
r116 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.305 $Y=0.45
+ $X2=5.39 $Y2=0.535
r117 26 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.305 $Y=0.45
+ $X2=4.9 $Y2=0.45
r118 22 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.595 $Y=2.275
+ $X2=5.68 $Y2=2.19
r119 22 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.595 $Y=2.275
+ $X2=4.86 $Y2=2.275
r120 20 38 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.155 $Y=1.41
+ $X2=6.02 $Y2=1.41
r121 20 21 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.155 $Y=1.41
+ $X2=6.23 $Y2=1.41
r122 16 18 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.23 $Y=1.025
+ $X2=6.33 $Y2=1.025
r123 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.33 $Y=0.95
+ $X2=6.33 $Y2=1.025
r124 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.33 $Y=0.95
+ $X2=6.33 $Y2=0.555
r125 9 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.23 $Y=1.545
+ $X2=6.23 $Y2=1.41
r126 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.23 $Y=1.545
+ $X2=6.23 $Y2=2.11
r127 8 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.23 $Y=1.275
+ $X2=6.23 $Y2=1.41
r128 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.23 $Y=1.1 $X2=6.23
+ $Y2=1.025
r129 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.23 $Y=1.1 $X2=6.23
+ $Y2=1.275
r130 2 24 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=4.7
+ $Y=2.065 $X2=4.86 $Y2=2.275
r131 1 28 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=4.705
+ $Y=0.235 $X2=4.9 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_1527_315# 1 2 9 13 15 17 20 22 24 27 29
+ 31 34 36 38 41 43 46 50 53 55 61 65 68 69 81
r145 78 79 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.66 $Y=1.16
+ $X2=10.09 $Y2=1.16
r146 70 72 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.71 $Y=1.74
+ $X2=7.825 $Y2=1.74
r147 65 67 16.9646 $w=3.58e-07 $l=4.4e-07 $layer=LI1_cond $X=8.57 $Y=0.385
+ $X2=8.57 $Y2=0.825
r148 62 81 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=10.32 $Y=1.16
+ $X2=10.51 $Y2=1.16
r149 62 79 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=10.32 $Y=1.16
+ $X2=10.09 $Y2=1.16
r150 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.32
+ $Y=1.16 $X2=10.32 $Y2=1.16
r151 59 78 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=9.3 $Y=1.16
+ $X2=9.66 $Y2=1.16
r152 59 75 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=9.3 $Y=1.16 $X2=9.24
+ $Y2=1.16
r153 58 61 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=9.3 $Y=1.2
+ $X2=10.32 $Y2=1.2
r154 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.3
+ $Y=1.16 $X2=9.3 $Y2=1.16
r155 56 69 0.237926 $w=2.5e-07 $l=9.3e-08 $layer=LI1_cond $X=8.755 $Y=1.2
+ $X2=8.662 $Y2=1.2
r156 56 58 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=8.755 $Y=1.2
+ $X2=9.3 $Y2=1.2
r157 55 68 6.7841 $w=2.35e-07 $l=1.88348e-07 $layer=LI1_cond $X=8.662 $Y=1.575
+ $X2=8.612 $Y2=1.74
r158 54 69 6.65529 $w=1.82e-07 $l=1.25e-07 $layer=LI1_cond $X=8.662 $Y=1.325
+ $X2=8.662 $Y2=1.2
r159 54 55 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=8.662 $Y=1.325
+ $X2=8.662 $Y2=1.575
r160 53 69 6.65529 $w=1.82e-07 $l=1.25996e-07 $layer=LI1_cond $X=8.66 $Y=1.075
+ $X2=8.662 $Y2=1.2
r161 53 67 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=8.66 $Y=1.075
+ $X2=8.66 $Y2=0.825
r162 48 68 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=8.612 $Y=1.905
+ $X2=8.612 $Y2=1.74
r163 48 50 1.81965 $w=2.83e-07 $l=4.5e-08 $layer=LI1_cond $X=8.612 $Y=1.905
+ $X2=8.612 $Y2=1.95
r164 46 72 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.89 $Y=1.74
+ $X2=7.825 $Y2=1.74
r165 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.74 $X2=7.89 $Y2=1.74
r166 43 68 0.153733 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=8.47 $Y=1.74
+ $X2=8.612 $Y2=1.74
r167 43 45 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=8.47 $Y=1.74
+ $X2=7.89 $Y2=1.74
r168 39 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.51 $Y=1.325
+ $X2=10.51 $Y2=1.16
r169 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.51 $Y=1.325
+ $X2=10.51 $Y2=1.985
r170 36 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.51 $Y=0.995
+ $X2=10.51 $Y2=1.16
r171 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.51 $Y=0.995
+ $X2=10.51 $Y2=0.56
r172 32 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.09 $Y=1.325
+ $X2=10.09 $Y2=1.16
r173 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.09 $Y=1.325
+ $X2=10.09 $Y2=1.985
r174 29 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.09 $Y=0.995
+ $X2=10.09 $Y2=1.16
r175 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.09 $Y=0.995
+ $X2=10.09 $Y2=0.56
r176 25 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.66 $Y=1.325
+ $X2=9.66 $Y2=1.16
r177 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.66 $Y=1.325
+ $X2=9.66 $Y2=1.985
r178 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.66 $Y=0.995
+ $X2=9.66 $Y2=1.16
r179 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.66 $Y=0.995
+ $X2=9.66 $Y2=0.56
r180 18 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=1.325
+ $X2=9.24 $Y2=1.16
r181 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.24 $Y=1.325
+ $X2=9.24 $Y2=1.985
r182 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=0.995
+ $X2=9.24 $Y2=1.16
r183 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.24 $Y=0.995
+ $X2=9.24 $Y2=0.56
r184 11 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.825 $Y=1.575
+ $X2=7.825 $Y2=1.74
r185 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.825 $Y=1.575
+ $X2=7.825 $Y2=0.445
r186 7 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.71 $Y=1.905
+ $X2=7.71 $Y2=1.74
r187 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.71 $Y=1.905
+ $X2=7.71 $Y2=2.275
r188 2 50 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=8.43
+ $Y=1.485 $X2=8.555 $Y2=1.95
r189 1 65 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=8.43
+ $Y=0.235 $X2=8.555 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_1356_413# 1 2 7 9 12 14 15 16 20 27 30 33
+ 34
c91 27 0 4.21632e-20 $X=7.55 $Y=2.165
c92 7 0 1.60992e-19 $X=8.765 $Y=0.995
r93 33 35 11.5578 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=7.485 $Y=1.16
+ $X2=7.485 $Y2=1.405
r94 33 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=1.16
+ $X2=7.485 $Y2=0.995
r95 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.315
+ $Y=1.16 $X2=8.315 $Y2=1.16
r96 28 33 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.635 $Y=1.16
+ $X2=7.485 $Y2=1.16
r97 28 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.635 $Y=1.16
+ $X2=8.315 $Y2=1.16
r98 27 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.55 $Y=2.165
+ $X2=7.55 $Y2=1.405
r99 24 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.42 $Y=0.535
+ $X2=7.42 $Y2=0.995
r100 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.335 $Y=0.45
+ $X2=7.42 $Y2=0.535
r101 20 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.335 $Y=0.45
+ $X2=7.13 $Y2=0.45
r102 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.465 $Y=2.25
+ $X2=7.55 $Y2=2.165
r103 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.465 $Y=2.25
+ $X2=6.915 $Y2=2.25
r104 14 31 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=8.69 $Y=1.16
+ $X2=8.315 $Y2=1.16
r105 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.69 $Y=1.16
+ $X2=8.765 $Y2=1.16
r106 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=1.325
+ $X2=8.765 $Y2=1.16
r107 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.765 $Y=1.325
+ $X2=8.765 $Y2=1.985
r108 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=0.995
+ $X2=8.765 $Y2=1.16
r109 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.765 $Y=0.995
+ $X2=8.765 $Y2=0.56
r110 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=6.78
+ $Y=2.065 $X2=6.915 $Y2=2.25
r111 1 22 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=6.91
+ $Y=0.235 $X2=7.13 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 45 49
+ 53 55 57 60 61 63 64 65 67 72 77 89 100 105 108 111 114 117 121
c179 121 0 1.81794e-19 $X=10.81 $Y=2.72
c180 2 0 1.60762e-19 $X=1.91 $Y=1.845
c181 1 0 3.29888e-20 $X=0.55 $Y=1.815
r182 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r183 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r184 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r185 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r186 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r187 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r188 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r189 103 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r190 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r191 100 120 3.40825 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=10.635 $Y=2.72
+ $X2=10.837 $Y2=2.72
r192 100 102 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.635 $Y=2.72
+ $X2=10.35 $Y2=2.72
r193 99 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r194 99 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r195 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r196 96 117 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.105 $Y=2.72
+ $X2=9.015 $Y2=2.72
r197 96 98 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.105 $Y=2.72
+ $X2=9.43 $Y2=2.72
r198 95 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r199 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r200 92 95 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r201 91 94 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r202 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r203 89 114 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.815 $Y=2.72
+ $X2=7.967 $Y2=2.72
r204 89 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.815 $Y=2.72
+ $X2=7.59 $Y2=2.72
r205 88 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r206 88 112 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r207 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r208 85 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=2.72
+ $X2=3.845 $Y2=2.72
r209 85 87 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=3.93 $Y=2.72
+ $X2=5.75 $Y2=2.72
r210 84 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r211 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r212 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r213 81 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r214 80 83 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r215 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r216 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.045 $Y2=2.72
r217 78 80 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.53 $Y2=2.72
r218 77 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=2.72
+ $X2=3.845 $Y2=2.72
r219 77 83 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=2.72
+ $X2=3.45 $Y2=2.72
r220 76 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r221 76 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r222 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r223 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=0.685 $Y2=2.72
r224 73 75 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r225 72 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=2.045 $Y2=2.72
r226 72 75 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=1.61 $Y2=2.72
r227 67 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.685 $Y2=2.72
r228 67 69 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r229 65 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r230 65 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r231 63 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=9.43 $Y2=2.72
r232 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=9.88 $Y2=2.72
r233 62 102 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.965 $Y=2.72
+ $X2=10.35 $Y2=2.72
r234 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.965 $Y=2.72
+ $X2=9.88 $Y2=2.72
r235 60 87 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.935 $Y=2.72
+ $X2=5.75 $Y2=2.72
r236 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.935 $Y=2.72
+ $X2=6.02 $Y2=2.72
r237 59 91 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.105 $Y=2.72
+ $X2=6.21 $Y2=2.72
r238 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.105 $Y=2.72
+ $X2=6.02 $Y2=2.72
r239 55 120 3.40825 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=10.72 $Y=2.635
+ $X2=10.837 $Y2=2.72
r240 55 57 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=10.72 $Y=2.635
+ $X2=10.72 $Y2=2.01
r241 51 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.88 $Y=2.635
+ $X2=9.88 $Y2=2.72
r242 51 53 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=9.88 $Y=2.635
+ $X2=9.88 $Y2=2.01
r243 47 117 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.015 $Y=2.635
+ $X2=9.015 $Y2=2.72
r244 47 49 52.0657 $w=1.78e-07 $l=8.45e-07 $layer=LI1_cond $X=9.015 $Y=2.635
+ $X2=9.015 $Y2=1.79
r245 46 114 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.12 $Y=2.72
+ $X2=7.967 $Y2=2.72
r246 45 117 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.925 $Y=2.72
+ $X2=9.015 $Y2=2.72
r247 45 46 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.925 $Y=2.72
+ $X2=8.12 $Y2=2.72
r248 41 114 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.967 $Y=2.635
+ $X2=7.967 $Y2=2.72
r249 41 43 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=7.967 $Y=2.635
+ $X2=7.967 $Y2=2.3
r250 37 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=2.635
+ $X2=6.02 $Y2=2.72
r251 37 39 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.02 $Y=2.635
+ $X2=6.02 $Y2=2
r252 33 111 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.72
r253 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.33
r254 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.72
r255 29 31 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.33
r256 25 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.72
r257 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.22
r258 8 57 300 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_PDIFF $count=2 $X=10.585
+ $Y=1.485 $X2=10.72 $Y2=2.01
r259 7 53 300 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_PDIFF $count=2 $X=9.735
+ $Y=1.485 $X2=9.88 $Y2=2.01
r260 6 49 300 $w=1.7e-07 $l=3.80624e-07 $layer=licon1_PDIFF $count=2 $X=8.84
+ $Y=1.485 $X2=9.01 $Y2=1.79
r261 5 43 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=7.785
+ $Y=2.065 $X2=8.03 $Y2=2.3
r262 4 39 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=5.645
+ $Y=2.065 $X2=6.02 $Y2=2
r263 3 35 600 $w=1.7e-07 $l=5.59308e-07 $layer=licon1_PDIFF $count=1 $X=3.685
+ $Y=1.845 $X2=3.845 $Y2=2.33
r264 2 31 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.845 $X2=2.045 $Y2=2.33
r265 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.815 $X2=0.685 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%A_560_369# 1 2 3 4 13 17 22 24 25 26 27 28
+ 30 32 36 38 39
c112 17 0 1.20015e-19 $X=3.425 $Y=0.36
r113 39 41 21.3062 $w=2.09e-07 $l=3.65e-07 $layer=LI1_cond $X=4.332 $Y=1.91
+ $X2=4.332 $Y2=2.275
r114 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.3 $Y=0.45 $X2=4.4
+ $Y2=0.45
r115 32 39 5.42244 $w=2.09e-07 $l=9.97246e-08 $layer=LI1_cond $X=4.3 $Y=1.825
+ $X2=4.332 $Y2=1.91
r116 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.865 $X2=4.3
+ $Y2=0.78
r117 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.3 $Y=0.865 $X2=4.3
+ $Y2=1.825
r118 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.695 $X2=4.3
+ $Y2=0.78
r119 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0.535
+ $X2=4.3 $Y2=0.45
r120 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.3 $Y=0.535
+ $X2=4.3 $Y2=0.695
r121 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.78
+ $X2=4.3 $Y2=0.78
r122 27 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.215 $Y=0.78
+ $X2=3.595 $Y2=0.78
r123 25 39 1.94907 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.215 $Y=1.91
+ $X2=4.332 $Y2=1.91
r124 25 26 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.215 $Y=1.91
+ $X2=3.59 $Y2=1.91
r125 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.51 $Y=0.695
+ $X2=3.595 $Y2=0.78
r126 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.51 $Y=0.445
+ $X2=3.51 $Y2=0.695
r127 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=1.995
+ $X2=3.59 $Y2=1.91
r128 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.505 $Y=1.995
+ $X2=3.505 $Y2=2.245
r129 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=0.36
+ $X2=3.51 $Y2=0.445
r130 17 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.425 $Y=0.36
+ $X2=3.015 $Y2=0.36
r131 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=2.33
+ $X2=3.505 $Y2=2.245
r132 13 15 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.42 $Y=2.33
+ $X2=2.935 $Y2=2.33
r133 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=2.065 $X2=4.365 $Y2=2.275
r134 3 15 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.845 $X2=2.935 $Y2=2.33
r135 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.275
+ $Y=0.235 $X2=4.4 $Y2=0.45
r136 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=3.015 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 31 33 35 39
+ 41 44
c87 15 0 1.60992e-19 $X=9.45 $Y=0.395
r88 43 44 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=10.805 $Y=1.505
+ $X2=10.805 $Y2=1.19
r89 42 44 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=10.805 $Y=0.905
+ $X2=10.805 $Y2=1.19
r90 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=1.59
+ $X2=10.3 $Y2=1.59
r91 35 43 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.655 $Y=1.59
+ $X2=10.805 $Y2=1.505
r92 35 36 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.655 $Y=1.59
+ $X2=10.465 $Y2=1.59
r93 34 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=0.82
+ $X2=10.3 $Y2=0.82
r94 33 42 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.655 $Y=0.82
+ $X2=10.805 $Y2=0.905
r95 33 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.655 $Y=0.82
+ $X2=10.465 $Y2=0.82
r96 29 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=1.675
+ $X2=10.3 $Y2=1.59
r97 29 31 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=10.3 $Y=1.675
+ $X2=10.3 $Y2=2.31
r98 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=0.735
+ $X2=10.3 $Y2=0.82
r99 25 27 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.3 $Y=0.735
+ $X2=10.3 $Y2=0.395
r100 24 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.615 $Y=1.59
+ $X2=9.45 $Y2=1.59
r101 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.135 $Y=1.59
+ $X2=10.3 $Y2=1.59
r102 23 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=10.135 $Y=1.59
+ $X2=9.615 $Y2=1.59
r103 21 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.135 $Y=0.82
+ $X2=10.3 $Y2=0.82
r104 21 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=10.135 $Y=0.82
+ $X2=9.615 $Y2=0.82
r105 17 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.45 $Y=1.675
+ $X2=9.45 $Y2=1.59
r106 17 19 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=9.45 $Y=1.675
+ $X2=9.45 $Y2=2.31
r107 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.45 $Y=0.735
+ $X2=9.615 $Y2=0.82
r108 13 15 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=9.45 $Y=0.735
+ $X2=9.45 $Y2=0.395
r109 4 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.165
+ $Y=1.485 $X2=10.3 $Y2=1.63
r110 4 31 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=10.165
+ $Y=1.485 $X2=10.3 $Y2=2.31
r111 3 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.315
+ $Y=1.485 $X2=9.45 $Y2=1.63
r112 3 19 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.315
+ $Y=1.485 $X2=9.45 $Y2=2.31
r113 2 27 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=10.165
+ $Y=0.235 $X2=10.3 $Y2=0.395
r114 1 15 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=9.315
+ $Y=0.235 $X2=9.45 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 37 41 45 47
+ 51 55 57 59 62 63 64 66 71 76 84 96 101 104 107 110 113 116 120
c183 120 0 2.71124e-20 $X=10.81 $Y=0
r184 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r185 116 117 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r186 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r187 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r188 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r189 108 111 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r190 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r191 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r192 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r193 99 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r194 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r195 96 119 3.40825 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.837 $Y2=0
r196 96 98 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.635 $Y=0
+ $X2=10.35 $Y2=0
r197 95 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r198 95 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r199 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r200 92 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.095 $Y=0 $X2=9.01
+ $Y2=0
r201 92 94 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=9.43 $Y2=0
r202 91 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r203 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r204 88 91 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r205 88 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r206 87 90 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=7.59
+ $Y2=0
r207 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r208 85 110 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=5.91 $Y2=0
r209 85 87 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.21 $Y2=0
r210 84 113 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.75 $Y=0
+ $X2=7.935 $Y2=0
r211 84 90 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.75 $Y=0 $X2=7.59
+ $Y2=0
r212 83 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r213 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r214 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r215 80 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r216 79 82 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r217 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r218 77 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.14 $Y2=0
r219 77 79 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r220 76 107 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.865
+ $Y2=0
r221 76 82 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.765 $Y=0
+ $X2=3.45 $Y2=0
r222 75 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r223 75 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r224 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r225 72 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r226 72 74 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r227 71 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=2.14 $Y2=0
r228 71 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r229 66 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r230 66 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r231 64 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r232 64 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r233 62 94 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.795 $Y=0
+ $X2=9.43 $Y2=0
r234 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=0 $X2=9.88
+ $Y2=0
r235 61 98 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.965 $Y=0
+ $X2=10.35 $Y2=0
r236 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.965 $Y=0 $X2=9.88
+ $Y2=0
r237 57 119 3.40825 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=10.72 $Y=0.085
+ $X2=10.837 $Y2=0
r238 57 59 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.72 $Y=0.085
+ $X2=10.72 $Y2=0.395
r239 53 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.88 $Y=0.085
+ $X2=9.88 $Y2=0
r240 53 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.88 $Y=0.085
+ $X2=9.88 $Y2=0.395
r241 49 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0
r242 49 51 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0.53
r243 48 113 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.12 $Y=0
+ $X2=7.935 $Y2=0
r244 47 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.925 $Y=0 $X2=9.01
+ $Y2=0
r245 47 48 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.925 $Y=0
+ $X2=8.12 $Y2=0
r246 43 113 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=0.085
+ $X2=7.935 $Y2=0
r247 43 45 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.935 $Y=0.085
+ $X2=7.935 $Y2=0.45
r248 39 110 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=0.085
+ $X2=5.91 $Y2=0
r249 39 41 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.91 $Y=0.085
+ $X2=5.91 $Y2=0.42
r250 38 107 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.865
+ $Y2=0
r251 37 110 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.725 $Y=0
+ $X2=5.91 $Y2=0
r252 37 38 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=5.725 $Y=0
+ $X2=3.965 $Y2=0
r253 33 107 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0
r254 33 35 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0.36
r255 29 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r256 29 31 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.36
r257 25 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r258 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r259 8 59 182 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=1 $X=10.585
+ $Y=0.235 $X2=10.72 $Y2=0.395
r260 7 55 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=9.735
+ $Y=0.235 $X2=9.88 $Y2=0.395
r261 6 51 182 $w=1.7e-07 $l=3.70371e-07 $layer=licon1_NDIFF $count=1 $X=8.84
+ $Y=0.235 $X2=9.01 $Y2=0.53
r262 5 45 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=7.9
+ $Y=0.235 $X2=8.035 $Y2=0.45
r263 4 41 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=5.675
+ $Y=0.235 $X2=5.98 $Y2=0.42
r264 3 35 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.235 $X2=3.85 $Y2=0.36
r265 2 31 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.14 $Y2=0.36
r266 1 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlxbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.955000 1.810000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215000 0.415000 5.465000 0.660000 ;
        RECT 5.215000 0.660000 5.500000 0.825000 ;
        RECT 5.215000 1.495000 5.500000 1.710000 ;
        RECT 5.215000 1.710000 5.465000 2.455000 ;
        RECT 5.330000 0.825000 5.500000 0.995000 ;
        RECT 5.330000 0.995000 5.905000 1.325000 ;
        RECT 5.330000 1.325000 5.500000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.050000 0.255000 7.305000 0.825000 ;
        RECT 7.050000 1.445000 7.305000 2.465000 ;
        RECT 7.095000 0.825000 7.305000 1.055000 ;
        RECT 7.095000 1.055000 7.735000 1.325000 ;
        RECT 7.095000 1.325000 7.305000 1.445000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.895000  0.085000 2.225000 0.445000 ;
        RECT 3.760000  0.085000 4.090000 0.825000 ;
        RECT 4.760000  0.085000 5.045000 0.825000 ;
        RECT 5.635000  0.085000 5.905000 0.545000 ;
        RECT 6.585000  0.085000 6.880000 0.545000 ;
        RECT 7.475000  0.085000 7.735000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.975000 1.835000 2.290000 2.635000 ;
        RECT 3.840000 2.135000 4.140000 2.635000 ;
        RECT 4.760000 1.495000 5.045000 2.635000 ;
        RECT 5.635000 1.835000 5.905000 2.635000 ;
        RECT 6.585000 1.835000 6.880000 2.635000 ;
        RECT 7.475000 1.495000 7.735000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.780000 0.805000 ;
      RECT 0.175000 1.795000 0.780000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.780000 1.070000 ;
      RECT 0.610000 1.070000 0.840000 1.400000 ;
      RECT 0.610000 1.400000 0.780000 1.795000 ;
      RECT 1.015000 0.345000 1.185000 1.685000 ;
      RECT 1.015000 1.685000 1.240000 2.465000 ;
      RECT 1.475000 1.495000 2.160000 1.665000 ;
      RECT 1.475000 1.665000 1.805000 2.415000 ;
      RECT 1.555000 0.345000 1.725000 0.615000 ;
      RECT 1.555000 0.615000 2.160000 0.765000 ;
      RECT 1.555000 0.765000 2.360000 0.785000 ;
      RECT 1.990000 0.785000 2.360000 1.095000 ;
      RECT 1.990000 1.095000 2.160000 1.495000 ;
      RECT 2.490000 1.355000 2.775000 2.005000 ;
      RECT 2.735000 0.705000 3.115000 1.035000 ;
      RECT 2.860000 0.365000 3.520000 0.535000 ;
      RECT 2.920000 2.255000 3.670000 2.425000 ;
      RECT 2.945000 1.035000 3.115000 1.415000 ;
      RECT 2.945000 1.415000 3.285000 1.995000 ;
      RECT 3.350000 0.535000 3.520000 0.995000 ;
      RECT 3.350000 0.995000 4.220000 1.165000 ;
      RECT 3.500000 1.165000 4.220000 1.325000 ;
      RECT 3.500000 1.325000 3.670000 2.255000 ;
      RECT 3.860000 1.535000 4.580000 1.865000 ;
      RECT 4.360000 0.415000 4.580000 0.825000 ;
      RECT 4.360000 1.865000 4.580000 2.435000 ;
      RECT 4.410000 0.825000 4.580000 0.995000 ;
      RECT 4.410000 0.995000 5.160000 1.325000 ;
      RECT 4.410000 1.325000 4.580000 1.535000 ;
      RECT 6.075000 0.255000 6.405000 0.995000 ;
      RECT 6.075000 0.995000 6.925000 1.325000 ;
      RECT 6.075000 1.325000 6.405000 2.465000 ;
    LAYER mcon ;
      RECT 0.610000 1.445000 0.780000 1.615000 ;
      RECT 1.070000 1.785000 1.240000 1.955000 ;
      RECT 2.490000 1.785000 2.660000 1.955000 ;
      RECT 2.950000 1.445000 3.120000 1.615000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.720000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.430000 1.755000 2.720000 1.800000 ;
      RECT 2.430000 1.940000 2.720000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxbn_2
END LIBRARY

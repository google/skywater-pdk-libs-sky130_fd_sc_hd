# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__xor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505000 1.075000 7.915000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685000 0.995000 6.855000 1.445000 ;
        RECT 6.685000 1.445000 7.265000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.995000 2.495000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.590000 0.925000 ;
        RECT 0.085000 0.925000 0.400000 1.440000 ;
        RECT 0.085000 1.440000 0.610000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.740000 0.085000 ;
        RECT 0.760000  0.085000 1.010000 0.525000 ;
        RECT 3.930000  0.085000 4.100000 0.865000 ;
        RECT 7.935000  0.085000 8.105000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.740000 2.805000 ;
        RECT 0.780000 2.215000 1.115000 2.635000 ;
        RECT 3.685000 2.235000 4.015000 2.635000 ;
        RECT 7.855000 2.275000 8.190000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.750000 0.995000 0.950000 1.325000 ;
      RECT 0.780000 0.695000 1.350000 0.865000 ;
      RECT 0.780000 0.865000 0.950000 0.995000 ;
      RECT 0.780000 1.325000 0.950000 1.875000 ;
      RECT 0.780000 1.875000 1.470000 2.045000 ;
      RECT 1.180000 0.255000 2.740000 0.425000 ;
      RECT 1.180000 0.425000 1.350000 0.695000 ;
      RECT 1.185000 1.535000 2.835000 1.705000 ;
      RECT 1.300000 2.045000 1.470000 2.235000 ;
      RECT 1.300000 2.235000 2.895000 2.405000 ;
      RECT 1.520000 0.595000 1.690000 1.535000 ;
      RECT 1.870000 1.895000 3.175000 2.065000 ;
      RECT 1.970000 0.655000 3.080000 0.825000 ;
      RECT 2.390000 0.425000 2.740000 0.455000 ;
      RECT 2.665000 0.995000 2.940000 1.325000 ;
      RECT 2.665000 1.325000 2.835000 1.535000 ;
      RECT 2.910000 0.255000 3.760000 0.425000 ;
      RECT 2.910000 0.425000 3.080000 0.655000 ;
      RECT 3.005000 1.525000 3.535000 1.695000 ;
      RECT 3.005000 1.695000 3.175000 1.895000 ;
      RECT 3.110000 2.235000 3.515000 2.405000 ;
      RECT 3.250000 0.595000 3.420000 1.375000 ;
      RECT 3.250000 1.375000 3.535000 1.525000 ;
      RECT 3.345000 1.895000 4.520000 2.065000 ;
      RECT 3.345000 2.065000 3.515000 2.235000 ;
      RECT 3.590000 0.425000 3.760000 1.035000 ;
      RECT 3.590000 1.035000 3.875000 1.205000 ;
      RECT 3.705000 1.205000 3.875000 1.895000 ;
      RECT 4.105000 1.445000 4.520000 1.715000 ;
      RECT 4.280000 0.415000 4.520000 1.445000 ;
      RECT 4.350000 2.065000 4.520000 2.275000 ;
      RECT 4.350000 2.275000 7.445000 2.445000 ;
      RECT 4.695000 0.265000 5.110000 0.485000 ;
      RECT 4.695000 0.485000 4.915000 0.595000 ;
      RECT 4.695000 0.595000 4.865000 2.105000 ;
      RECT 5.035000 0.720000 5.450000 0.825000 ;
      RECT 5.035000 0.825000 5.255000 0.890000 ;
      RECT 5.035000 0.890000 5.205000 2.275000 ;
      RECT 5.085000 0.655000 5.450000 0.720000 ;
      RECT 5.280000 0.320000 5.450000 0.655000 ;
      RECT 5.395000 1.445000 6.175000 1.615000 ;
      RECT 5.395000 1.615000 5.810000 2.045000 ;
      RECT 5.410000 0.995000 5.835000 1.270000 ;
      RECT 5.620000 0.630000 5.835000 0.995000 ;
      RECT 6.005000 0.255000 7.150000 0.425000 ;
      RECT 6.005000 0.425000 6.175000 1.445000 ;
      RECT 6.345000 0.595000 6.515000 1.935000 ;
      RECT 6.345000 1.935000 8.655000 2.105000 ;
      RECT 6.685000 0.425000 7.150000 0.465000 ;
      RECT 7.025000 0.730000 7.230000 0.945000 ;
      RECT 7.025000 0.945000 7.335000 1.275000 ;
      RECT 7.435000 1.495000 8.255000 1.705000 ;
      RECT 7.475000 0.295000 7.765000 0.735000 ;
      RECT 7.475000 0.735000 8.255000 0.750000 ;
      RECT 7.515000 0.750000 8.255000 0.905000 ;
      RECT 8.085000 0.905000 8.255000 0.995000 ;
      RECT 8.085000 0.995000 8.315000 1.325000 ;
      RECT 8.085000 1.325000 8.255000 1.495000 ;
      RECT 8.170000 1.875000 8.655000 1.935000 ;
      RECT 8.355000 0.255000 8.655000 0.585000 ;
      RECT 8.360000 2.105000 8.655000 2.465000 ;
      RECT 8.485000 0.585000 8.655000 1.875000 ;
    LAYER mcon ;
      RECT 3.365000 1.445000 3.535000 1.615000 ;
      RECT 4.285000 0.765000 4.455000 0.935000 ;
      RECT 4.745000 0.425000 4.915000 0.595000 ;
      RECT 5.665000 0.765000 5.835000 0.935000 ;
      RECT 5.665000 1.445000 5.835000 1.615000 ;
      RECT 7.045000 0.765000 7.215000 0.935000 ;
      RECT 7.505000 0.425000 7.675000 0.595000 ;
    LAYER met1 ;
      RECT 3.305000 1.415000 3.595000 1.460000 ;
      RECT 3.305000 1.460000 5.895000 1.600000 ;
      RECT 3.305000 1.600000 3.595000 1.645000 ;
      RECT 4.225000 0.735000 4.515000 0.780000 ;
      RECT 4.225000 0.780000 7.275000 0.920000 ;
      RECT 4.225000 0.920000 4.515000 0.965000 ;
      RECT 4.685000 0.395000 4.975000 0.440000 ;
      RECT 4.685000 0.440000 7.735000 0.580000 ;
      RECT 4.685000 0.580000 4.975000 0.625000 ;
      RECT 5.605000 0.735000 5.895000 0.780000 ;
      RECT 5.605000 0.920000 5.895000 0.965000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.985000 0.735000 7.275000 0.780000 ;
      RECT 6.985000 0.920000 7.275000 0.965000 ;
      RECT 7.445000 0.395000 7.735000 0.440000 ;
      RECT 7.445000 0.580000 7.735000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_1
END LIBRARY

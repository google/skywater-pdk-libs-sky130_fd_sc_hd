* File: sky130_fd_sc_hd__nand3_2.spice
* Created: Tue Sep  1 19:16:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand3_2.pex.spice"
.subckt sky130_fd_sc_hd__nand3_2  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_47#_M1003_d N_A_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1011 N_A_27_47#_M1011_d N_A_M1011_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1011_d N_B_M1007_g N_A_277_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_27_47#_M1008_d N_B_M1008_g N_A_277_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g N_A_277_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_C_M1005_g N_A_277_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1010 N_Y_M1000_d N_B_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75000.2 A=0.15
+ P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_C_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.31
+ AS=0.135 PD=2.62 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__nand3_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a221oi_1.pex.spice
* Created: Tue Sep  1 18:52:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A221OI_1%C1 1 3 6 8 14
c27 8 0 1.69525e-19 $X=0.23 $Y=1.19
r28 11 14 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.25 $Y=1.16
+ $X2=0.47 $Y2=1.16
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r30 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r31 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r32 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r33 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%B2 3 7 8 11 12 13
c29 11 0 1.69525e-19 $X=0.89 $Y=1.16
c30 3 0 1.18612e-19 $X=0.89 $Y=1.985
r31 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r33 8 12 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=0.7 $Y=1.18 $X2=0.89
+ $Y2=1.18
r34 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.56
+ $X2=0.945 $Y2=0.995
r35 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r36 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%B1 3 6 8 9 13 15
r42 14 17 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.18
+ $X2=1.555 $Y2=1.18
r43 13 16 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.382 $Y=1.16
+ $X2=1.382 $Y2=1.325
r44 13 15 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.382 $Y=1.16
+ $X2=1.382 $Y2=0.995
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.16 $X2=1.39 $Y2=1.16
r46 9 17 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=1.61 $Y=1.18
+ $X2=1.555 $Y2=1.18
r47 8 17 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=1.555 $Y=0.85
+ $X2=1.555 $Y2=1.075
r48 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=1.325
r49 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.56 $X2=1.31
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%A1 3 6 8 9 13 15
c39 8 0 7.4301e-20 $X=2.07 $Y=0.85
r40 13 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.15 $Y2=1.325
r41 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.15 $Y2=0.995
r42 9 22 3.5937 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=1.16 $X2=2.11
+ $Y2=1.075
r43 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.16 $X2=2.11 $Y2=1.16
r44 8 22 10.1686 $w=2.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.072 $Y=0.85
+ $X2=2.072 $Y2=1.075
r45 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.985
+ $X2=2.25 $Y2=1.325
r46 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.25 $Y=0.56 $X2=2.25
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%A2 3 6 8 11 12 13
c32 11 0 7.4301e-20 $X=2.67 $Y=1.16
c33 6 0 1.46456e-19 $X=2.705 $Y=1.985
r34 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.67 $Y2=1.325
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.67 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.16 $X2=2.67 $Y2=1.16
r37 8 12 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.555 $Y=1.16
+ $X2=2.67 $Y2=1.16
r38 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.705 $Y=1.985
+ $X2=2.705 $Y2=1.325
r39 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.705 $Y=0.56
+ $X2=2.705 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%Y 1 2 3 4 15 19 21 22 24 27 28 33 37 38 39
+ 40 41 42 43 49 50 52
c101 52 0 1.83134e-19 $X=3.015 $Y=0.85
c102 40 0 2.94484e-19 $X=2.3 $Y=1.56
r103 49 52 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=3.03 $Y=0.825
+ $X2=3.03 $Y2=0.85
r104 43 50 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=1.58
+ $X2=3.03 $Y2=1.495
r105 43 50 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=3.03 $Y=1.47
+ $X2=3.03 $Y2=1.495
r106 42 43 14.7879 $w=2.08e-07 $l=2.8e-07 $layer=LI1_cond $X=3.03 $Y=1.19
+ $X2=3.03 $Y2=1.47
r107 41 49 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=0.74
+ $X2=3.03 $Y2=0.825
r108 41 42 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=3.03 $Y=0.88
+ $X2=3.03 $Y2=1.19
r109 41 52 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=3.03 $Y=0.88 $X2=3.03
+ $Y2=0.85
r110 39 40 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.15 $Y=1.56
+ $X2=2.3 $Y2=1.56
r111 37 41 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.925 $Y=0.74
+ $X2=3.03 $Y2=0.74
r112 37 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.925 $Y=0.74
+ $X2=2.58 $Y2=0.74
r113 36 38 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.48 $Y=0.655
+ $X2=2.58 $Y2=0.74
r114 35 36 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.48 $Y=0.505
+ $X2=2.48 $Y2=0.655
r115 33 43 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=3.03 $Y2=1.58
r116 33 40 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=2.3 $Y2=1.58
r117 30 32 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=1.52 $Y=0.38
+ $X2=2.04 $Y2=0.38
r118 28 30 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=1.235 $Y=0.38
+ $X2=1.52 $Y2=0.38
r119 27 35 6.92652 $w=2.5e-07 $l=1.67705e-07 $layer=LI1_cond $X=2.38 $Y=0.38
+ $X2=2.48 $Y2=0.505
r120 27 32 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.38 $Y=0.38
+ $X2=2.04 $Y2=0.38
r121 25 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.15 $Y=0.505
+ $X2=1.235 $Y2=0.38
r122 25 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.15 $Y=0.505
+ $X2=1.15 $Y2=0.735
r123 24 39 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=0.345 $Y=1.54
+ $X2=2.15 $Y2=1.54
r124 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=0.82
+ $X2=1.15 $Y2=0.735
r125 21 22 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.065 $Y=0.82
+ $X2=0.345 $Y2=0.82
r126 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.345 $Y2=1.54
r127 17 19 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.65
r128 13 22 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.345 $Y2=0.82
r129 13 15 11.0909 $w=1.73e-07 $l=1.75e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.56
r130 4 19 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r131 3 32 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.04 $Y2=0.42
r132 2 30 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.42
r133 1 15 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%A_109_297# 1 2 9 12 14 15
c22 14 0 1.18612e-19 $X=1.52 $Y=2.34
r23 14 15 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=2.36
+ $X2=1.355 $Y2=2.36
r24 12 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.765 $Y=2.38
+ $X2=1.355 $Y2=2.38
r25 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.64 $Y=2.295
+ $X2=0.765 $Y2=2.38
r26 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.64 $Y=2.295
+ $X2=0.64 $Y2=1.96
r27 2 14 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r28 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%A_193_297# 1 2 7 9 11 13 18 19
r28 16 18 5.59382 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.1 $Y=1.96 $X2=1.24
+ $Y2=1.96
r29 11 21 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.5 $Y=2.045 $X2=2.5
+ $Y2=1.94
r30 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.5 $Y=2.045
+ $X2=2.5 $Y2=2.3
r31 9 21 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.375 $Y=1.94 $X2=2.5
+ $Y2=1.94
r32 9 19 18.4848 $w=2.08e-07 $l=3.5e-07 $layer=LI1_cond $X=2.375 $Y=1.94
+ $X2=2.025 $Y2=1.94
r33 7 19 6.09095 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.9 $Y=1.92
+ $X2=2.025 $Y2=1.92
r34 7 18 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=1.9 $Y=1.92 $X2=1.24
+ $Y2=1.92
r35 2 21 600 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.95
r36 2 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.3
r37 1 16 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%VPWR 1 2 9 11 13 15 17 25 31 35
c48 2 0 1.83134e-19 $X=2.78 $Y=1.485
r49 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.04 $Y2=2.72
r55 26 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 25 34 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=3.007 $Y2=2.72
r57 25 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 24 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 19 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=2.04 $Y2=2.72
r62 17 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 15 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 15 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 11 34 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=3.007 $Y2=2.72
r66 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=2.96 $Y2=1.96
r67 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635 $X2=2.04
+ $Y2=2.72
r68 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=2.635 $X2=2.04
+ $Y2=2.3
r69 2 13 300 $w=1.7e-07 $l=5.57786e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=1.485 $X2=2.96 $Y2=1.96
r70 1 9 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.485 $X2=2.04 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_1%VGND 1 2 9 11 13 15 17 22 31 35
r46 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r47 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r49 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r51 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r52 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r55 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r56 22 34 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.985
+ $Y2=0
r57 22 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.53
+ $Y2=0
r58 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r59 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r60 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 11 34 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.985 $Y2=0
r63 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.4
r64 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r65 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.44
r66 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.235 $X2=2.915 $Y2=0.4
r67 1 9 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.44
.ends


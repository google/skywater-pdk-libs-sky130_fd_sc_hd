* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4.spice.SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4.pxi
* Created: Thu Aug 27 14:26:26 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VGND N_VGND_M1014_s
+ N_VGND_M1003_s N_VGND_M1004_s N_VGND_M1010_s N_VGND_M1005_s N_VGND_M1020_s
+ N_VGND_M1012_s N_VGND_M1007_s N_VGND_M1018_s N_VGND_M1014_b N_VGND_c_30_p
+ N_VGND_c_9_p N_VGND_c_31_p N_VGND_c_13_p N_VGND_c_55_p N_VGND_c_25_p
+ N_VGND_c_49_p N_VGND_c_125_p N_VGND_c_141_p N_VGND_c_32_p N_VGND_c_10_p
+ N_VGND_c_40_p N_VGND_c_50_p N_VGND_c_126_p N_VGND_c_135_p VGND VGND
+ N_VGND_c_21_p N_VGND_c_104_p N_VGND_c_33_p N_VGND_c_11_p
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPB N_VPB_X22_noxref_D1
+ N_VPB_M1021_b N_VPB_c_249_p N_VPB_c_166_n VPB N_VPB_c_167_n N_VPB_c_168_n VPB
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPB
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPWRIN N_VPWRIN_M1013_s
+ N_VPWRIN_M1013_b N_VPWRIN_c_281_p N_VPWRIN_c_260_n N_VPWRIN_c_273_p
+ N_VPWRIN_c_255_n N_VPWRIN_c_256_n N_VPWRIN_c_271_p N_VPWRIN_c_257_n VPWRIN
+ N_VPWRIN_c_258_n PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPWRIN
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_505_297#
+ N_A_505_297#_M1014_d N_A_505_297#_M1013_d N_A_505_297#_c_319_n
+ N_A_505_297#_M1003_g N_A_505_297#_c_323_n N_A_505_297#_M1010_g
+ N_A_505_297#_c_327_n N_A_505_297#_c_329_n N_A_505_297#_c_330_n
+ N_A_505_297#_M1019_g N_A_505_297#_c_334_n N_A_505_297#_c_335_n
+ N_A_505_297#_M1020_g N_A_505_297#_c_339_n N_A_505_297#_c_340_n
+ N_A_505_297#_c_345_n N_A_505_297#_c_356_n N_A_505_297#_c_346_n
+ N_A_505_297#_c_347_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_505_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_714_47#
+ N_A_714_47#_M1004_d N_A_714_47#_M1009_d N_A_714_47#_M1000_s
+ N_A_714_47#_c_427_n N_A_714_47#_c_405_n N_A_714_47#_M1021_g
+ N_A_714_47#_c_406_n N_A_714_47#_c_408_n N_A_714_47#_c_409_n
+ N_A_714_47#_c_410_n N_A_714_47#_c_411_n N_A_714_47#_c_412_n
+ N_A_714_47#_c_413_n N_A_714_47#_c_418_n N_A_714_47#_c_434_n
+ N_A_714_47#_c_424_n N_A_714_47#_c_426_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_714_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A N_A_M1013_g N_A_c_507_n
+ N_A_M1014_g N_A_c_512_n N_A_M1004_g N_A_c_518_n N_A_c_519_n N_A_M1005_g
+ N_A_c_526_n N_A_M1009_g N_A_c_532_n N_A_M1012_g N_A_c_538_n N_A_c_539_n
+ N_A_c_540_n A N_A_c_541_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_620_911#
+ N_A_620_911#_M1003_d N_A_620_911#_M1019_d N_A_620_911#_M1021_s
+ N_A_620_911#_c_601_n N_A_620_911#_c_579_n N_A_620_911#_c_580_n
+ N_A_620_911#_M1000_g N_A_620_911#_c_607_n N_A_620_911#_c_608_n
+ N_A_620_911#_M1011_g N_A_620_911#_M1001_g N_A_620_911#_c_612_n
+ N_A_620_911#_c_613_n N_A_620_911#_c_614_n N_A_620_911#_c_585_n
+ N_A_620_911#_c_589_n N_A_620_911#_c_616_n N_A_620_911#_c_591_n
+ N_A_620_911#_c_617_n N_A_620_911#_c_595_n N_A_620_911#_c_596_n
+ N_A_620_911#_c_597_n N_A_620_911#_c_598_n N_A_620_911#_c_623_n
+ N_A_620_911#_c_599_n N_A_620_911#_c_600_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_620_911#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_1032_911#
+ N_A_1032_911#_M1011_d N_A_1032_911#_M1001_d N_A_1032_911#_M1006_g
+ N_A_1032_911#_c_734_n N_A_1032_911#_M1002_g N_A_1032_911#_c_710_n
+ N_A_1032_911#_M1007_g N_A_1032_911#_M1008_g N_A_1032_911#_c_737_n
+ N_A_1032_911#_c_739_n N_A_1032_911#_M1017_g N_A_1032_911#_M1015_g
+ N_A_1032_911#_c_742_n N_A_1032_911#_c_719_n N_A_1032_911#_M1018_g
+ N_A_1032_911#_M1016_g N_A_1032_911#_c_726_n N_A_1032_911#_c_747_n
+ N_A_1032_911#_c_748_n N_A_1032_911#_c_749_n N_A_1032_911#_c_727_n
+ N_A_1032_911#_c_728_n N_A_1032_911#_c_732_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%A_1032_911#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPWR N_VPWR_M1000_d
+ N_VPWR_M1021_d N_VPWR_M1008_s N_VPWR_M1016_s N_VPWR_c_809_n N_VPWR_c_810_n
+ N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n
+ N_VPWR_c_817_n N_VPWR_c_818_n VPWR N_VPWR_c_806_n N_VPWR_c_821_n
+ N_VPWR_c_807_n VPWR PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%X N_X_M1006_d N_X_M1017_d
+ N_X_M1002_d N_X_M1015_d N_X_c_916_n N_X_c_919_n N_X_c_927_n N_X_c_920_n
+ N_X_c_940_n X X N_X_c_924_n X
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4%X
cc_1 N_VGND_M1014_b N_VPB_c_166_n 0.0790644f $X=-0.19 $Y=-0.24 $X2=6.93 $Y2=3.57
cc_2 N_VGND_M1014_b N_VPB_c_167_n 0.0100791f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=3.29
cc_3 N_VGND_M1014_b N_VPB_c_168_n 0.00990609f $X=-0.19 $Y=-0.24 $X2=7.13
+ $Y2=3.29
cc_4 N_VGND_M1014_b N_VPWRIN_c_255_n 0.00447854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 N_VGND_M1014_b N_VPWRIN_c_256_n 0.0244366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 N_VGND_M1014_b N_VPWRIN_c_257_n 0.0306316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 N_VGND_M1014_b N_VPWRIN_c_258_n 0.0344347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 N_VGND_M1014_b N_A_505_297#_c_319_n 0.0179052f $X=-0.19 $Y=-0.24 $X2=-0.19
+ $Y2=1.305
cc_9 N_VGND_c_9_p N_A_505_297#_c_319_n 0.00414737f $X=2.81 $Y=4.7 $X2=-0.19
+ $Y2=1.305
cc_10 N_VGND_c_10_p N_A_505_297#_c_319_n 0.0054895f $X=3.575 $Y=5.44 $X2=-0.19
+ $Y2=1.305
cc_11 N_VGND_c_11_p N_A_505_297#_c_319_n 0.0110264f $X=7.13 $Y=5.44 $X2=-0.19
+ $Y2=1.305
cc_12 N_VGND_M1014_b N_A_505_297#_c_323_n 0.0140848f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_13 N_VGND_c_13_p N_A_505_297#_c_323_n 0.00179869f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_14 N_VGND_c_10_p N_A_505_297#_c_323_n 0.0054895f $X=3.575 $Y=5.44 $X2=0 $Y2=0
cc_15 N_VGND_c_11_p N_A_505_297#_c_323_n 0.00972667f $X=7.13 $Y=5.44 $X2=0 $Y2=0
cc_16 N_VGND_M1014_b N_A_505_297#_c_327_n 0.0130779f $X=-0.19 $Y=-0.24 $X2=0.225
+ $Y2=3.57
cc_17 N_VGND_c_13_p N_A_505_297#_c_327_n 0.00240634f $X=3.67 $Y=4.735 $X2=0.225
+ $Y2=3.57
cc_18 N_VGND_M1014_b N_A_505_297#_c_329_n 0.0294363f $X=-0.19 $Y=-0.24 $X2=0.225
+ $Y2=3.57
cc_19 N_VGND_M1014_b N_A_505_297#_c_330_n 0.0140848f $X=-0.19 $Y=-0.24 $X2=6.93
+ $Y2=3.57
cc_20 N_VGND_c_13_p N_A_505_297#_c_330_n 0.00304527f $X=3.67 $Y=4.735 $X2=6.93
+ $Y2=3.57
cc_21 N_VGND_c_21_p N_A_505_297#_c_330_n 0.0054895f $X=4.445 $Y=5.44 $X2=6.93
+ $Y2=3.57
cc_22 N_VGND_c_11_p N_A_505_297#_c_330_n 0.00972667f $X=7.13 $Y=5.44 $X2=6.93
+ $Y2=3.57
cc_23 N_VGND_M1014_b N_A_505_297#_c_334_n 0.0195784f $X=-0.19 $Y=-0.24 $X2=7.075
+ $Y2=3.57
cc_24 N_VGND_M1014_b N_A_505_297#_c_335_n 0.0162763f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_25 N_VGND_c_25_p N_A_505_297#_c_335_n 0.00390324f $X=4.87 $Y=4.735 $X2=0
+ $Y2=0
cc_26 N_VGND_c_21_p N_A_505_297#_c_335_n 0.0054895f $X=4.445 $Y=5.44 $X2=0 $Y2=0
cc_27 N_VGND_c_11_p N_A_505_297#_c_335_n 0.0103929f $X=7.13 $Y=5.44 $X2=0 $Y2=0
cc_28 N_VGND_M1014_b N_A_505_297#_c_339_n 0.00569361f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_29 N_VGND_M1014_b N_A_505_297#_c_340_n 0.00997858f $X=-0.19 $Y=-0.24
+ $X2=0.557 $Y2=3.57
cc_30 N_VGND_c_30_p N_A_505_297#_c_340_n 0.0068636f $X=2.245 $Y=0.62 $X2=0.557
+ $Y2=3.57
cc_31 N_VGND_c_31_p N_A_505_297#_c_340_n 0.0271827f $X=3.28 $Y=0.42 $X2=0.557
+ $Y2=3.57
cc_32 N_VGND_c_32_p N_A_505_297#_c_340_n 0.00966373f $X=3.115 $Y=0 $X2=0.557
+ $Y2=3.57
cc_33 N_VGND_c_33_p N_A_505_297#_c_340_n 0.00857725f $X=7.13 $Y=0 $X2=0.557
+ $Y2=3.57
cc_34 N_VGND_M1014_b N_A_505_297#_c_345_n 0.016089f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_35 N_VGND_M1014_b N_A_505_297#_c_346_n 0.034685f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_36 N_VGND_M1014_b N_A_505_297#_c_347_n 0.0845171f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_37 N_VGND_c_33_p N_A_714_47#_M1004_d 0.00397884f $X=7.13 $Y=0 $X2=0.145
+ $Y2=3.04
cc_38 N_VGND_c_33_p N_A_714_47#_M1009_d 0.00400851f $X=7.13 $Y=0 $X2=7.045
+ $Y2=3.04
cc_39 N_VGND_M1014_b N_A_714_47#_c_405_n 0.0129761f $X=-0.19 $Y=-0.24 $X2=0.37
+ $Y2=3.57
cc_40 N_VGND_c_40_p N_A_714_47#_c_406_n 0.0121541f $X=3.975 $Y=0 $X2=0.49
+ $Y2=3.5
cc_41 N_VGND_c_33_p N_A_714_47#_c_406_n 0.00717399f $X=7.13 $Y=0 $X2=0.49
+ $Y2=3.5
cc_42 N_VGND_M1014_b N_A_714_47#_c_408_n 0.0175549f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.29
cc_43 N_VGND_M1014_b N_A_714_47#_c_409_n 0.00209323f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_44 N_VGND_M1014_b N_A_714_47#_c_410_n 0.00298088f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.57
cc_45 N_VGND_M1014_b N_A_714_47#_c_411_n 0.0397033f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_46 N_VGND_M1014_b N_A_714_47#_c_412_n 0.0516547f $X=-0.19 $Y=-0.24 $X2=7.13
+ $Y2=3.57
cc_47 N_VGND_M1005_s N_A_714_47#_c_413_n 3.36085e-19 $X=4 $Y=0.235 $X2=0 $Y2=0
cc_48 N_VGND_M1014_b N_A_714_47#_c_413_n 0.00893993f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_49 N_VGND_c_49_p N_A_714_47#_c_413_n 0.00706177f $X=5 $Y=0.42 $X2=0 $Y2=0
cc_50 N_VGND_c_50_p N_A_714_47#_c_413_n 0.00202943f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_51 N_VGND_c_33_p N_A_714_47#_c_413_n 0.00389716f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_52 N_VGND_M1005_s N_A_714_47#_c_418_n 0.00139685f $X=4 $Y=0.235 $X2=0.557
+ $Y2=3.57
cc_53 N_VGND_M1014_b N_A_714_47#_c_418_n 0.00805719f $X=-0.19 $Y=-0.24 $X2=0.557
+ $Y2=3.57
cc_54 N_VGND_c_31_p N_A_714_47#_c_418_n 0.00702407f $X=3.28 $Y=0.42 $X2=0.557
+ $Y2=3.57
cc_55 N_VGND_c_55_p N_A_714_47#_c_418_n 0.0168391f $X=4.14 $Y=0.42 $X2=0.557
+ $Y2=3.57
cc_56 N_VGND_c_40_p N_A_714_47#_c_418_n 0.00204475f $X=3.975 $Y=0 $X2=0.557
+ $Y2=3.57
cc_57 N_VGND_c_33_p N_A_714_47#_c_418_n 0.00522015f $X=7.13 $Y=0 $X2=0.557
+ $Y2=3.57
cc_58 N_VGND_c_50_p N_A_714_47#_c_424_n 0.0124538f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_59 N_VGND_c_33_p N_A_714_47#_c_424_n 0.00724021f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_60 N_VGND_M1014_b N_A_714_47#_c_426_n 0.00576889f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_61 N_VGND_M1014_b N_A_M1013_g 0.00675179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 N_VGND_M1014_b N_A_c_507_n 0.0408343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 N_VGND_c_30_p N_A_c_507_n 0.0135915f $X=2.245 $Y=0.62 $X2=0 $Y2=0
cc_64 N_VGND_c_31_p N_A_c_507_n 0.00625119f $X=3.28 $Y=0.42 $X2=0 $Y2=0
cc_65 N_VGND_c_32_p N_A_c_507_n 0.00585385f $X=3.115 $Y=0 $X2=0 $Y2=0
cc_66 N_VGND_c_33_p N_A_c_507_n 0.0134051f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_67 N_VGND_M1014_b N_A_c_512_n 0.0352506f $X=-0.19 $Y=-0.24 $X2=4.25 $Y2=1.305
cc_68 N_VGND_M1014_b N_A_M1004_g 0.0240979f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=3.57
cc_69 N_VGND_c_31_p N_A_M1004_g 0.0129916f $X=3.28 $Y=0.42 $X2=0.225 $Y2=3.57
cc_70 N_VGND_c_55_p N_A_M1004_g 5.31107e-19 $X=4.14 $Y=0.42 $X2=0.225 $Y2=3.57
cc_71 N_VGND_c_40_p N_A_M1004_g 0.00486043f $X=3.975 $Y=0 $X2=0.225 $Y2=3.57
cc_72 N_VGND_c_33_p N_A_M1004_g 0.00822531f $X=7.13 $Y=0 $X2=0.225 $Y2=3.57
cc_73 N_VGND_M1014_b N_A_c_518_n 0.0168496f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=3.57
cc_74 N_VGND_M1014_b N_A_c_519_n 0.0656946f $X=-0.19 $Y=-0.24 $X2=6.93 $Y2=3.57
cc_75 N_VGND_c_31_p N_A_c_519_n 0.00306309f $X=3.28 $Y=0.42 $X2=6.93 $Y2=3.57
cc_76 N_VGND_M1014_b N_A_M1005_g 0.0189456f $X=-0.19 $Y=-0.24 $X2=7.075 $Y2=3.57
cc_77 N_VGND_c_31_p N_A_M1005_g 6.36276e-19 $X=3.28 $Y=0.42 $X2=7.075 $Y2=3.57
cc_78 N_VGND_c_55_p N_A_M1005_g 0.00741971f $X=4.14 $Y=0.42 $X2=7.075 $Y2=3.57
cc_79 N_VGND_c_40_p N_A_M1005_g 0.00364644f $X=3.975 $Y=0 $X2=7.075 $Y2=3.57
cc_80 N_VGND_c_33_p N_A_M1005_g 0.00430798f $X=7.13 $Y=0 $X2=7.075 $Y2=3.57
cc_81 N_VGND_M1014_b N_A_c_526_n 0.0149976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 N_VGND_M1014_b N_A_M1009_g 0.018948f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=3.57
cc_83 N_VGND_c_55_p N_A_M1009_g 0.00741971f $X=4.14 $Y=0.42 $X2=0.23 $Y2=3.57
cc_84 N_VGND_c_49_p N_A_M1009_g 6.33842e-19 $X=5 $Y=0.42 $X2=0.23 $Y2=3.57
cc_85 N_VGND_c_50_p N_A_M1009_g 0.00364644f $X=4.835 $Y=0 $X2=0.23 $Y2=3.57
cc_86 N_VGND_c_33_p N_A_M1009_g 0.00430798f $X=7.13 $Y=0 $X2=0.23 $Y2=3.57
cc_87 N_VGND_M1014_b N_A_c_532_n 0.0255444f $X=-0.19 $Y=-0.24 $X2=7.13 $Y2=3.29
cc_88 N_VGND_M1014_b N_A_M1012_g 0.0204702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 N_VGND_c_55_p N_A_M1012_g 5.31107e-19 $X=4.14 $Y=0.42 $X2=0 $Y2=0
cc_90 N_VGND_c_49_p N_A_M1012_g 0.0112243f $X=5 $Y=0.42 $X2=0 $Y2=0
cc_91 N_VGND_c_50_p N_A_M1012_g 0.00486043f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_92 N_VGND_c_33_p N_A_M1012_g 0.00822531f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_93 N_VGND_M1014_b N_A_c_538_n 0.017446f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=3.57
cc_94 N_VGND_M1014_b N_A_c_539_n 0.00933068f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=3.57
cc_95 N_VGND_M1014_b N_A_c_540_n 0.0106787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 N_VGND_M1014_b N_A_c_541_n 0.0169952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 N_VGND_c_31_p N_A_c_541_n 0.0150235f $X=3.28 $Y=0.42 $X2=0 $Y2=0
cc_98 N_VGND_c_11_p N_A_620_911#_M1003_d 0.00223231f $X=7.13 $Y=5.44 $X2=0.145
+ $Y2=3.04
cc_99 N_VGND_c_11_p N_A_620_911#_M1019_d 0.00223231f $X=7.13 $Y=5.44 $X2=7.045
+ $Y2=3.04
cc_100 N_VGND_M1014_b N_A_620_911#_c_579_n 0.0127228f $X=-0.19 $Y=-0.24 $X2=0.37
+ $Y2=3.57
cc_101 N_VGND_c_25_p N_A_620_911#_c_580_n 0.0183082f $X=4.87 $Y=4.735 $X2=0.225
+ $Y2=3.57
cc_102 N_VGND_M1014_b N_A_620_911#_M1011_g 0.0484682f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.57
cc_103 N_VGND_c_25_p N_A_620_911#_M1011_g 0.00390249f $X=4.87 $Y=4.735 $X2=0.23
+ $Y2=3.57
cc_104 N_VGND_c_104_p N_A_620_911#_M1011_g 0.00548296f $X=6.985 $Y=5.44 $X2=0.23
+ $Y2=3.57
cc_105 N_VGND_c_11_p N_A_620_911#_M1011_g 0.0116568f $X=7.13 $Y=5.44 $X2=0.23
+ $Y2=3.57
cc_106 N_VGND_c_9_p N_A_620_911#_c_585_n 0.0267051f $X=2.81 $Y=4.7 $X2=0 $Y2=0
cc_107 N_VGND_c_13_p N_A_620_911#_c_585_n 0.0266323f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_108 N_VGND_c_10_p N_A_620_911#_c_585_n 0.0189253f $X=3.575 $Y=5.44 $X2=0
+ $Y2=0
cc_109 N_VGND_c_11_p N_A_620_911#_c_585_n 0.0122674f $X=7.13 $Y=5.44 $X2=0 $Y2=0
cc_110 N_VGND_M1014_b N_A_620_911#_c_589_n 0.0128475f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_111 N_VGND_c_13_p N_A_620_911#_c_589_n 0.0146667f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_112 N_VGND_c_13_p N_A_620_911#_c_591_n 0.0266323f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_113 N_VGND_c_25_p N_A_620_911#_c_591_n 0.025678f $X=4.87 $Y=4.735 $X2=0 $Y2=0
cc_114 N_VGND_c_21_p N_A_620_911#_c_591_n 0.0189253f $X=4.445 $Y=5.44 $X2=0
+ $Y2=0
cc_115 N_VGND_c_11_p N_A_620_911#_c_591_n 0.0122674f $X=7.13 $Y=5.44 $X2=0 $Y2=0
cc_116 N_VGND_M1014_b N_A_620_911#_c_595_n 0.0561622f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_117 N_VGND_M1014_b N_A_620_911#_c_596_n 0.0016479f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_118 N_VGND_M1014_b N_A_620_911#_c_597_n 7.55444e-19 $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_119 N_VGND_M1014_b N_A_620_911#_c_598_n 9.83343e-19 $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_120 N_VGND_M1014_b N_A_620_911#_c_599_n 0.00835191f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_121 N_VGND_M1014_b N_A_620_911#_c_600_n 0.0133087f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_122 N_VGND_c_11_p N_A_1032_911#_M1011_d 0.00214546f $X=7.13 $Y=5.44 $X2=0.145
+ $Y2=3.04
cc_123 N_VGND_M1014_b N_A_1032_911#_M1006_g 0.0226878f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_124 N_VGND_c_49_p N_A_1032_911#_M1006_g 0.00189452f $X=5 $Y=0.42 $X2=0 $Y2=0
cc_125 N_VGND_c_125_p N_A_1032_911#_M1006_g 5.88421e-19 $X=5.99 $Y=0.42 $X2=0
+ $Y2=0
cc_126 N_VGND_c_126_p N_A_1032_911#_M1006_g 0.00585385f $X=5.825 $Y=0 $X2=0
+ $Y2=0
cc_127 N_VGND_c_33_p N_A_1032_911#_M1006_g 0.010837f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_128 N_VGND_M1014_b N_A_1032_911#_c_710_n 0.0140243f $X=-0.19 $Y=-0.24
+ $X2=0.225 $Y2=3.57
cc_129 N_VGND_M1014_b N_A_1032_911#_M1007_g 0.0216078f $X=-0.19 $Y=-0.24
+ $X2=7.075 $Y2=3.57
cc_130 N_VGND_c_125_p N_A_1032_911#_M1007_g 0.0110235f $X=5.99 $Y=0.42 $X2=7.075
+ $Y2=3.57
cc_131 N_VGND_c_126_p N_A_1032_911#_M1007_g 0.00486043f $X=5.825 $Y=0 $X2=7.075
+ $Y2=3.57
cc_132 N_VGND_c_33_p N_A_1032_911#_M1007_g 0.00852643f $X=7.13 $Y=0 $X2=7.075
+ $Y2=3.57
cc_133 N_VGND_M1014_b N_A_1032_911#_M1017_g 0.0205125f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_134 N_VGND_c_125_p N_A_1032_911#_M1017_g 0.010662f $X=5.99 $Y=0.42 $X2=0
+ $Y2=0
cc_135 N_VGND_c_135_p N_A_1032_911#_M1017_g 0.00486043f $X=6.755 $Y=0 $X2=0
+ $Y2=0
cc_136 N_VGND_c_33_p N_A_1032_911#_M1017_g 0.00822531f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_137 N_VGND_M1014_b N_A_1032_911#_c_719_n 0.0411217f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_138 N_VGND_c_125_p N_A_1032_911#_c_719_n 0.00223674f $X=5.99 $Y=0.42 $X2=0
+ $Y2=0
cc_139 N_VGND_M1014_b N_A_1032_911#_M1018_g 0.0282249f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_140 N_VGND_c_125_p N_A_1032_911#_M1018_g 6.48459e-19 $X=5.99 $Y=0.42 $X2=0
+ $Y2=0
cc_141 N_VGND_c_141_p N_A_1032_911#_M1018_g 0.00407687f $X=6.85 $Y=0.42 $X2=0
+ $Y2=0
cc_142 N_VGND_c_135_p N_A_1032_911#_M1018_g 0.00585385f $X=6.755 $Y=0 $X2=0
+ $Y2=0
cc_143 N_VGND_c_33_p N_A_1032_911#_M1018_g 0.011676f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_144 N_VGND_M1014_b N_A_1032_911#_c_726_n 0.0111194f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_145 N_VGND_M1014_b N_A_1032_911#_c_727_n 0.00998896f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_146 N_VGND_M1014_b N_A_1032_911#_c_728_n 0.0492761f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_147 N_VGND_c_25_p N_A_1032_911#_c_728_n 0.0259447f $X=4.87 $Y=4.735 $X2=0
+ $Y2=0
cc_148 N_VGND_c_104_p N_A_1032_911#_c_728_n 0.0239189f $X=6.985 $Y=5.44 $X2=0
+ $Y2=0
cc_149 N_VGND_c_11_p N_A_1032_911#_c_728_n 0.0195213f $X=7.13 $Y=5.44 $X2=0
+ $Y2=0
cc_150 N_VGND_M1014_b N_A_1032_911#_c_732_n 0.0384737f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_151 N_VGND_M1014_b N_VPWR_c_806_n 0.0363208f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 N_VGND_M1014_b N_VPWR_c_807_n 0.0368329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 N_VGND_c_33_p N_X_M1006_d 0.00542784f $X=7.13 $Y=0 $X2=0.145 $Y2=3.04
cc_154 N_VGND_c_33_p N_X_M1017_d 0.00431525f $X=7.13 $Y=0 $X2=7.045 $Y2=3.04
cc_155 N_VGND_c_125_p N_X_c_916_n 0.0406307f $X=5.99 $Y=0.42 $X2=6.93 $Y2=3.57
cc_156 N_VGND_c_126_p N_X_c_916_n 0.0191787f $X=5.825 $Y=0 $X2=6.93 $Y2=3.57
cc_157 N_VGND_c_33_p N_X_c_916_n 0.0114765f $X=7.13 $Y=0 $X2=6.93 $Y2=3.57
cc_158 N_VGND_c_125_p N_X_c_919_n 0.0165907f $X=5.99 $Y=0.42 $X2=7.075 $Y2=3.57
cc_159 N_VGND_M1014_b N_X_c_920_n 0.00373262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_160 N_VGND_c_141_p N_X_c_920_n 0.00274856f $X=6.85 $Y=0.42 $X2=0 $Y2=0
cc_161 N_VGND_c_135_p N_X_c_920_n 0.0135183f $X=6.755 $Y=0 $X2=0 $Y2=0
cc_162 N_VGND_c_33_p N_X_c_920_n 0.00839034f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_163 N_VGND_M1014_b N_X_c_924_n 0.00503584f $X=-0.19 $Y=-0.24 $X2=0.56
+ $Y2=3.57
cc_164 N_VGND_c_49_p N_X_c_924_n 0.001162f $X=5 $Y=0.42 $X2=0.56 $Y2=3.57
cc_165 N_VGND_c_125_p N_X_c_924_n 0.00106574f $X=5.99 $Y=0.42 $X2=0.56 $Y2=3.57
cc_166 N_VPB_c_166_n N_VPWRIN_M1013_b 0.0152996f $X=6.93 $Y=3.57 $X2=4.86
+ $Y2=0.235
cc_167 N_VPB_c_166_n N_VPWRIN_c_260_n 0.0727088f $X=6.93 $Y=3.57 $X2=0 $Y2=0
cc_168 N_VPB_M1021_b N_VPWRIN_c_256_n 0.0251748f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_169 N_VPB_X22_noxref_D1 N_VPWRIN_c_257_n 0.0309709f $X=-0.19 $Y=1.305 $X2=0
+ $Y2=0
cc_170 N_VPB_c_166_n N_A_505_297#_c_346_n 0.0247683f $X=6.93 $Y=3.57 $X2=0 $Y2=0
cc_171 N_VPB_c_166_n N_A_505_297#_c_347_n 6.63876e-19 $X=6.93 $Y=3.57 $X2=-0.19
+ $Y2=-0.24
cc_172 N_VPB_M1021_b N_A_714_47#_c_427_n 0.0256732f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_173 N_VPB_M1021_b N_A_714_47#_c_405_n 5.34541e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_174 N_VPB_M1021_b N_A_714_47#_M1021_g 0.0198732f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_175 N_VPB_M1021_b N_A_714_47#_c_409_n 0.0045246f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_176 N_VPB_c_166_n N_A_714_47#_c_409_n 0.0451176f $X=6.93 $Y=3.57 $X2=0 $Y2=0
cc_177 N_VPB_c_166_n N_A_714_47#_c_410_n 0.010882f $X=6.93 $Y=3.57 $X2=0 $Y2=0
cc_178 N_VPB_M1021_b N_A_714_47#_c_412_n 0.0149067f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_179 N_VPB_M1021_b N_A_714_47#_c_434_n 0.00449536f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_180 N_VPB_M1021_b N_A_620_911#_c_601_n 0.0169344f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_181 N_VPB_M1021_b N_A_620_911#_c_579_n 5.21411e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_182 N_VPB_M1021_b N_A_620_911#_c_580_n 0.0246766f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_183 N_VPB_c_166_n N_A_620_911#_c_580_n 5.78421e-19 $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_184 N_VPB_M1021_b N_A_620_911#_M1000_g 0.00259316f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_185 N_VPB_c_166_n N_A_620_911#_M1000_g 0.00720206f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_186 N_VPB_M1021_b N_A_620_911#_c_607_n 0.0249303f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_187 N_VPB_M1021_b N_A_620_911#_c_608_n 0.0094712f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_188 N_VPB_M1021_b N_A_620_911#_M1011_g 0.00114838f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_189 N_VPB_M1021_b N_A_620_911#_M1001_g 0.0064606f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_190 N_VPB_c_166_n N_A_620_911#_M1001_g 0.00821798f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_191 N_VPB_M1021_b N_A_620_911#_c_612_n 0.00400906f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_192 N_VPB_M1021_b N_A_620_911#_c_613_n 0.00698872f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_193 N_VPB_M1021_b N_A_620_911#_c_614_n 0.0141637f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_194 N_VPB_c_166_n N_A_620_911#_c_589_n 0.0118014f $X=6.93 $Y=3.57 $X2=-0.19
+ $Y2=-0.24
cc_195 N_VPB_c_166_n N_A_620_911#_c_616_n 0.00154646f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_196 N_VPB_c_166_n N_A_620_911#_c_617_n 7.52174e-19 $X=6.93 $Y=3.57 $X2=0.23
+ $Y2=4.8
cc_197 N_VPB_M1021_b N_A_620_911#_c_595_n 0.0188917f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_198 N_VPB_c_166_n N_A_620_911#_c_595_n 0.00519139f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_199 N_VPB_c_166_n N_A_620_911#_c_596_n 0.00368761f $X=6.93 $Y=3.57 $X2=2.185
+ $Y2=0.62
cc_200 N_VPB_M1021_b N_A_620_911#_c_597_n 0.00337762f $X=4.25 $Y=1.305 $X2=2.775
+ $Y2=5.355
cc_201 N_VPB_c_166_n N_A_620_911#_c_597_n 8.12088e-19 $X=6.93 $Y=3.57 $X2=2.775
+ $Y2=5.355
cc_202 N_VPB_M1021_b N_A_620_911#_c_623_n 0.00324872f $X=4.25 $Y=1.305 $X2=3.28
+ $Y2=0.085
cc_203 N_VPB_c_166_n N_A_620_911#_c_599_n 0.00167232f $X=6.93 $Y=3.57 $X2=3.28
+ $Y2=0.42
cc_204 N_VPB_M1021_b N_A_620_911#_c_600_n 6.57859e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_205 N_VPB_c_166_n N_A_1032_911#_M1001_d 0.00329366f $X=6.93 $Y=3.57 $X2=2.685
+ $Y2=4.555
cc_206 N_VPB_M1021_b N_A_1032_911#_c_734_n 0.0147881f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_207 N_VPB_M1021_b N_A_1032_911#_c_710_n 0.00953288f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_208 N_VPB_M1021_b N_A_1032_911#_M1008_g 0.0277715f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_209 N_VPB_M1021_b N_A_1032_911#_c_737_n 0.063957f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_210 N_VPB_c_166_n N_A_1032_911#_c_737_n 0.00877695f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_211 N_VPB_M1021_b N_A_1032_911#_c_739_n 0.0172775f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_212 N_VPB_c_166_n N_A_1032_911#_c_739_n 0.0145367f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_213 N_VPB_M1021_b N_A_1032_911#_M1015_g 0.0202696f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_214 N_VPB_M1021_b N_A_1032_911#_c_742_n 0.0299183f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_215 N_VPB_M1021_b N_A_1032_911#_c_719_n 0.0223728f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_216 N_VPB_M1021_b N_A_1032_911#_M1016_g 0.035372f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_217 N_VPB_c_168_n N_A_1032_911#_M1016_g 0.00604195f $X=7.13 $Y=3.29 $X2=0
+ $Y2=0
cc_218 N_VPB_M1021_b N_A_1032_911#_c_726_n 0.00747506f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_219 N_VPB_M1021_b N_A_1032_911#_c_747_n 0.00596971f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_220 N_VPB_M1021_b N_A_1032_911#_c_748_n 0.00843141f $X=4.25 $Y=1.305
+ $X2=2.185 $Y2=0.085
cc_221 N_VPB_M1021_b N_A_1032_911#_c_749_n 0.00808952f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_222 N_VPB_c_166_n N_A_1032_911#_c_749_n 0.0241804f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_223 N_VPB_M1021_b N_A_1032_911#_c_727_n 8.50392e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_224 N_VPB_c_166_n N_A_1032_911#_c_727_n 0.00972995f $X=6.93 $Y=3.57 $X2=0
+ $Y2=0
cc_225 N_VPB_M1021_b N_A_1032_911#_c_728_n 0.00293548f $X=4.25 $Y=1.305 $X2=3.28
+ $Y2=0.42
cc_226 N_VPB_c_166_n N_A_1032_911#_c_728_n 0.00771994f $X=6.93 $Y=3.57 $X2=3.28
+ $Y2=0.42
cc_227 N_VPB_M1021_b N_A_1032_911#_c_732_n 0.0209772f $X=4.25 $Y=1.305 $X2=3.67
+ $Y2=4.735
cc_228 N_VPB_c_166_n N_A_1032_911#_c_732_n 0.00445361f $X=6.93 $Y=3.57 $X2=3.67
+ $Y2=4.735
cc_229 N_VPB_c_166_n N_VPWR_M1000_d 0.00370825f $X=6.93 $Y=3.57 $X2=2.12
+ $Y2=0.41
cc_230 N_VPB_M1021_b N_VPWR_c_809_n 0.00429074f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_231 N_VPB_M1021_b N_VPWR_c_810_n 0.00447924f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_232 N_VPB_c_166_n N_VPWR_c_810_n 0.0205244f $X=6.93 $Y=3.57 $X2=0 $Y2=0
cc_233 N_VPB_M1021_b N_VPWR_c_812_n 0.00379002f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_234 N_VPB_M1021_b N_VPWR_c_813_n 0.00404706f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_235 N_VPB_M1021_b N_VPWR_c_814_n 0.00101664f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_236 N_VPB_M1021_b N_VPWR_c_815_n 0.0107502f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_237 N_VPB_M1021_b N_VPWR_c_816_n 0.0021751f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_238 N_VPB_M1021_b N_VPWR_c_817_n 0.00753446f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_239 N_VPB_M1021_b N_VPWR_c_818_n 0.00258752f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_240 N_VPB_X22_noxref_D1 N_VPWR_c_806_n 0.0202024f $X=-0.19 $Y=1.305 $X2=0
+ $Y2=0
cc_241 N_VPB_c_167_n N_VPWR_c_806_n 0.0194225f $X=0.23 $Y=3.29 $X2=0 $Y2=0
cc_242 N_VPB_M1021_b N_VPWR_c_821_n 0.0130106f $X=4.25 $Y=1.305 $X2=2.245
+ $Y2=0.62
cc_243 N_VPB_c_168_n N_VPWR_c_821_n 0.0194225f $X=7.13 $Y=3.29 $X2=2.245
+ $Y2=0.62
cc_244 N_VPB_X22_noxref_D1 N_VPWR_c_807_n 0.0368104f $X=-0.19 $Y=1.305 $X2=0
+ $Y2=0
cc_245 N_VPB_M1021_b N_VPWR_c_807_n 0.0461017f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_246 N_VPB_c_249_p N_VPWR_c_807_n 0.0152864f $X=0.37 $Y=3.57 $X2=0 $Y2=0
cc_247 N_VPB_c_166_n N_VPWR_c_807_n 0.338819f $X=6.93 $Y=3.57 $X2=0 $Y2=0
cc_248 N_VPB_c_167_n N_VPWR_c_807_n 0.00501853f $X=0.23 $Y=3.29 $X2=0 $Y2=0
cc_249 N_VPB_c_168_n N_VPWR_c_807_n 0.00506082f $X=7.13 $Y=3.29 $X2=0 $Y2=0
cc_250 N_VPB_M1021_b N_X_c_927_n 0.00374381f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_251 N_VPB_M1021_b X 0.00132567f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_252 N_VPWRIN_c_256_n N_A_505_297#_M1013_d 0.00144688f $X=2.225 $Y=2.2
+ $X2=2.685 $Y2=4.555
cc_253 N_VPWRIN_M1013_b N_A_505_297#_c_340_n 0.0037173f $X=1.92 $Y=1.305 $X2=0
+ $Y2=0
cc_254 N_VPWRIN_c_256_n N_A_505_297#_c_340_n 3.15819e-19 $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_255 N_VPWRIN_M1013_b N_A_505_297#_c_345_n 0.00974718f $X=1.92 $Y=1.305 $X2=0
+ $Y2=0
cc_256 N_VPWRIN_c_260_n N_A_505_297#_c_345_n 3.29394e-19 $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_257 N_VPWRIN_c_256_n N_A_505_297#_c_345_n 0.0372262f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_258 N_VPWRIN_c_260_n N_A_505_297#_c_356_n 0.00924483f $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_259 N_VPWRIN_c_256_n N_A_505_297#_c_356_n 0.0204768f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_260 N_VPWRIN_c_271_p N_A_505_297#_c_356_n 0.0100174f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_261 N_VPWRIN_c_260_n N_A_505_297#_c_346_n 0.0654251f $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_262 N_VPWRIN_c_273_p N_A_505_297#_c_346_n 0.00525651f $X=2.435 $Y=2.66 $X2=0
+ $Y2=0
cc_263 N_VPWRIN_c_260_n N_A_505_297#_c_347_n 0.00169032f $X=2.645 $Y=3.49
+ $X2=-0.19 $Y2=-0.24
cc_264 N_VPWRIN_c_256_n N_A_714_47#_c_427_n 5.4797e-19 $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_265 N_VPWRIN_c_256_n N_A_714_47#_M1021_g 0.00777495f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_266 N_VPWRIN_c_256_n N_A_714_47#_c_411_n 0.0182669f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_267 N_VPWRIN_c_256_n N_A_714_47#_c_412_n 0.0104851f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_268 N_VPWRIN_c_256_n N_A_714_47#_c_426_n 0.00926075f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_269 N_VPWRIN_M1013_b N_A_M1013_g 0.0304234f $X=1.92 $Y=1.305 $X2=3.135
+ $Y2=0.235
cc_270 N_VPWRIN_c_281_p N_A_M1013_g 0.00523247f $X=2.225 $Y=1.79 $X2=3.135
+ $Y2=0.235
cc_271 N_VPWRIN_c_260_n N_A_M1013_g 0.0055008f $X=2.645 $Y=3.49 $X2=3.135
+ $Y2=0.235
cc_272 N_VPWRIN_c_273_p N_A_M1013_g 0.00938999f $X=2.435 $Y=2.66 $X2=3.135
+ $Y2=0.235
cc_273 N_VPWRIN_c_256_n N_A_M1013_g 0.00645994f $X=2.225 $Y=2.2 $X2=3.135
+ $Y2=0.235
cc_274 N_VPWRIN_c_271_p N_A_M1013_g 0.00218038f $X=2.225 $Y=2.2 $X2=3.135
+ $Y2=0.235
cc_275 N_VPWRIN_M1013_b N_A_c_519_n 0.00316885f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_276 N_VPWRIN_M1013_b N_A_c_541_n 0.00111856f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_277 N_VPWRIN_c_256_n N_A_c_541_n 0.00229296f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_278 N_VPWRIN_c_256_n N_A_620_911#_M1021_s 0.00479759f $X=2.225 $Y=2.2
+ $X2=3.135 $Y2=0.235
cc_279 N_VPWRIN_c_256_n N_A_620_911#_c_597_n 0.0011695f $X=2.225 $Y=2.2
+ $X2=2.775 $Y2=5.355
cc_280 N_VPWRIN_c_256_n N_A_620_911#_c_623_n 0.0174341f $X=2.225 $Y=2.2 $X2=3.28
+ $Y2=0.085
cc_281 N_VPWRIN_c_256_n N_A_1032_911#_c_734_n 0.00737951f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_282 N_VPWRIN_c_256_n N_A_1032_911#_M1008_g 0.00870505f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_283 N_VPWRIN_c_256_n N_A_1032_911#_M1015_g 0.00715996f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_284 N_VPWRIN_c_256_n N_A_1032_911#_M1016_g 0.00712859f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_285 N_VPWRIN_c_256_n N_VPWR_M1021_d 0.00413567f $X=2.225 $Y=2.2 $X2=2.685
+ $Y2=4.555
cc_286 N_VPWRIN_c_256_n N_VPWR_M1008_s 0.00463513f $X=2.225 $Y=2.2 $X2=3.135
+ $Y2=0.235
cc_287 N_VPWRIN_c_256_n N_VPWR_M1016_s 0.00454198f $X=2.225 $Y=2.2 $X2=3.53
+ $Y2=4.555
cc_288 N_VPWRIN_c_256_n N_VPWR_c_809_n 0.0221365f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_289 N_VPWRIN_c_256_n N_VPWR_c_812_n 0.0172645f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_290 N_VPWRIN_c_256_n N_VPWR_c_813_n 0.0200894f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_291 N_VPWRIN_c_256_n N_VPWR_c_815_n 0.00466952f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_292 N_VPWRIN_c_256_n N_VPWR_c_817_n 0.00411278f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_293 N_VPWRIN_c_273_p N_VPWR_c_806_n 0.0123972f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_294 N_VPWRIN_c_255_n N_VPWR_c_806_n 5.76636e-19 $X=1.475 $Y=2.2 $X2=0 $Y2=0
cc_295 N_VPWRIN_c_257_n N_VPWR_c_806_n 0.00675753f $X=1.36 $Y=2.2 $X2=0 $Y2=0
cc_296 N_VPWRIN_c_258_n N_VPWR_c_806_n 0.01865f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_297 N_VPWRIN_c_256_n N_VPWR_c_821_n 0.00185735f $X=2.225 $Y=2.2 $X2=2.245
+ $Y2=0.62
cc_298 N_VPWRIN_M1013_b N_VPWR_c_807_n 0.00623335f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_299 N_VPWRIN_c_260_n N_VPWR_c_807_n 0.0659883f $X=2.645 $Y=3.49 $X2=0 $Y2=0
cc_300 N_VPWRIN_c_273_p N_VPWR_c_807_n 0.02138f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_301 N_VPWRIN_c_255_n N_VPWR_c_807_n 0.0948062f $X=1.475 $Y=2.2 $X2=0 $Y2=0
cc_302 N_VPWRIN_c_256_n N_VPWR_c_807_n 0.418194f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_303 N_VPWRIN_c_257_n N_VPWR_c_807_n 0.116739f $X=1.36 $Y=2.2 $X2=0 $Y2=0
cc_304 N_VPWRIN_c_258_n N_VPWR_c_807_n 0.00970859f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_305 N_VPWRIN_c_256_n N_X_M1002_d 0.0041104f $X=2.225 $Y=2.2 $X2=3.135
+ $Y2=0.235
cc_306 N_VPWRIN_c_256_n N_X_c_927_n 0.0245217f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_307 N_VPWRIN_c_256_n X 0.0251052f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_308 N_A_505_297#_c_346_n N_A_714_47#_c_408_n 0.0441264f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_309 N_A_505_297#_c_334_n N_A_714_47#_c_409_n 6.95188e-19 $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_310 N_A_505_297#_c_339_n N_A_714_47#_c_409_n 3.7852e-19 $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_311 N_A_505_297#_c_346_n N_A_714_47#_c_410_n 0.00788518f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_312 N_A_505_297#_c_345_n N_A_714_47#_c_411_n 0.0048486f $X=3.06 $Y=2.25 $X2=0
+ $Y2=0
cc_313 N_A_505_297#_c_346_n N_A_714_47#_c_411_n 9.66994e-19 $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_314 N_A_505_297#_c_345_n N_A_714_47#_c_412_n 0.00327676f $X=3.06 $Y=2.25
+ $X2=0 $Y2=0
cc_315 N_A_505_297#_c_346_n N_A_714_47#_c_412_n 0.00125462f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_316 N_A_505_297#_c_346_n N_A_714_47#_c_426_n 0.0084582f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_317 N_A_505_297#_c_340_n N_A_M1013_g 0.0110528f $X=2.675 $Y=0.62 $X2=3.135
+ $Y2=0.235
cc_318 N_A_505_297#_c_346_n N_A_M1013_g 0.0027023f $X=3.225 $Y=3.84 $X2=3.135
+ $Y2=0.235
cc_319 N_A_505_297#_c_340_n N_A_c_507_n 0.010267f $X=2.675 $Y=0.62 $X2=4
+ $Y2=0.235
cc_320 N_A_505_297#_c_340_n N_A_c_512_n 0.0218308f $X=2.675 $Y=0.62 $X2=5.85
+ $Y2=0.235
cc_321 N_A_505_297#_c_340_n N_A_M1004_g 0.00480585f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_322 N_A_505_297#_c_340_n N_A_c_519_n 0.00146935f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_323 N_A_505_297#_c_340_n N_A_c_541_n 0.0360803f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_324 N_A_505_297#_c_345_n N_A_c_541_n 0.00941491f $X=3.06 $Y=2.25 $X2=0 $Y2=0
cc_325 N_A_505_297#_c_334_n N_A_620_911#_c_580_n 0.0155516f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_326 N_A_505_297#_c_334_n N_A_620_911#_M1011_g 0.00777355f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_327 N_A_505_297#_c_319_n N_A_620_911#_c_585_n 0.00968676f $X=3.025 $Y=4.48
+ $X2=0 $Y2=0
cc_328 N_A_505_297#_c_323_n N_A_620_911#_c_585_n 0.00843936f $X=3.455 $Y=4.48
+ $X2=0 $Y2=0
cc_329 N_A_505_297#_c_329_n N_A_620_911#_c_585_n 0.0169132f $X=3.53 $Y=4.405
+ $X2=0 $Y2=0
cc_330 N_A_505_297#_c_330_n N_A_620_911#_c_585_n 2.89638e-19 $X=3.885 $Y=4.48
+ $X2=0 $Y2=0
cc_331 N_A_505_297#_c_329_n N_A_620_911#_c_589_n 0.021891f $X=3.53 $Y=4.405
+ $X2=-0.19 $Y2=-0.24
cc_332 N_A_505_297#_c_347_n N_A_620_911#_c_589_n 0.00420454f $X=3.225 $Y=3.84
+ $X2=-0.19 $Y2=-0.24
cc_333 N_A_505_297#_c_346_n N_A_620_911#_c_616_n 0.0218015f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_334 N_A_505_297#_c_347_n N_A_620_911#_c_616_n 0.0175078f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_335 N_A_505_297#_c_323_n N_A_620_911#_c_591_n 2.89638e-19 $X=3.455 $Y=4.48
+ $X2=0 $Y2=0
cc_336 N_A_505_297#_c_330_n N_A_620_911#_c_591_n 0.00843936f $X=3.885 $Y=4.48
+ $X2=0 $Y2=0
cc_337 N_A_505_297#_c_334_n N_A_620_911#_c_591_n 0.0149859f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_338 N_A_505_297#_c_335_n N_A_620_911#_c_591_n 0.00985995f $X=4.315 $Y=4.48
+ $X2=0 $Y2=0
cc_339 N_A_505_297#_c_339_n N_A_620_911#_c_591_n 0.00418634f $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_340 N_A_505_297#_c_346_n N_A_620_911#_c_595_n 0.00421035f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_341 N_A_505_297#_c_347_n N_A_620_911#_c_595_n 0.0112331f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_342 N_A_505_297#_c_346_n N_A_620_911#_c_596_n 0.00372705f $X=3.225 $Y=3.84
+ $X2=2.185 $Y2=0.62
cc_343 N_A_505_297#_c_347_n N_A_620_911#_c_596_n 0.0022314f $X=3.225 $Y=3.84
+ $X2=2.185 $Y2=0.62
cc_344 N_A_505_297#_c_339_n N_A_620_911#_c_600_n 0.0155516f $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_345 N_A_505_297#_M1013_d N_VPWR_c_807_n 0.00146082f $X=2.525 $Y=1.485 $X2=0
+ $Y2=0
cc_346 N_A_505_297#_c_345_n N_VPWR_c_807_n 0.00782153f $X=3.06 $Y=2.25 $X2=0
+ $Y2=0
cc_347 N_A_505_297#_c_356_n N_VPWR_c_807_n 0.00276885f $X=2.8 $Y=2.25 $X2=0
+ $Y2=0
cc_348 N_A_505_297#_c_346_n N_VPWR_c_807_n 0.0490709f $X=3.225 $Y=3.84 $X2=0
+ $Y2=0
cc_349 N_A_714_47#_c_418_n N_A_M1004_g 0.00265062f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_350 N_A_714_47#_c_418_n N_A_c_518_n 0.00391065f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_351 N_A_714_47#_c_411_n N_A_M1005_g 0.00224176f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_352 N_A_714_47#_c_418_n N_A_M1005_g 0.0169165f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_353 N_A_714_47#_c_411_n N_A_c_526_n 0.0205035f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_354 N_A_714_47#_c_418_n N_A_c_526_n 6.96042e-19 $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_355 N_A_714_47#_c_411_n N_A_M1009_g 0.00205104f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_356 N_A_714_47#_c_413_n N_A_M1009_g 0.0169165f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_357 N_A_714_47#_M1021_g N_A_c_532_n 0.0124308f $X=4.78 $Y=1.955 $X2=0 $Y2=0
cc_358 N_A_714_47#_c_413_n N_A_c_532_n 0.00296321f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_359 N_A_714_47#_c_413_n N_A_M1012_g 0.00146631f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_360 N_A_714_47#_c_412_n N_A_c_539_n 0.0062571f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_361 N_A_714_47#_c_427_n N_A_620_911#_c_601_n 0.0315412f $X=4.705 $Y=2.58
+ $X2=0 $Y2=0
cc_362 N_A_714_47#_c_409_n N_A_620_911#_c_601_n 4.83528e-19 $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_363 N_A_714_47#_c_434_n N_A_620_911#_c_601_n 0.00503951f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_364 N_A_714_47#_c_405_n N_A_620_911#_c_579_n 0.0315412f $X=4.27 $Y=2.58 $X2=0
+ $Y2=0
cc_365 N_A_714_47#_c_408_n N_A_620_911#_c_579_n 0.0158995f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_366 N_A_714_47#_c_426_n N_A_620_911#_c_579_n 9.48385e-19 $X=4.105 $Y=2.49
+ $X2=0 $Y2=0
cc_367 N_A_714_47#_c_409_n N_A_620_911#_c_580_n 0.00905183f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_368 N_A_714_47#_c_409_n N_A_620_911#_M1000_g 0.00273734f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_369 N_A_714_47#_c_434_n N_A_620_911#_M1000_g 0.00383717f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_370 N_A_714_47#_c_409_n N_A_620_911#_c_589_n 0.00177263f $X=4.39 $Y=3.555
+ $X2=-0.19 $Y2=-0.24
cc_371 N_A_714_47#_c_410_n N_A_620_911#_c_589_n 0.0036785f $X=3.85 $Y=3.555
+ $X2=-0.19 $Y2=-0.24
cc_372 N_A_714_47#_c_408_n N_A_620_911#_c_617_n 0.0272967f $X=3.765 $Y=3.47
+ $X2=0.23 $Y2=4.8
cc_373 N_A_714_47#_c_409_n N_A_620_911#_c_617_n 0.0109877f $X=4.39 $Y=3.555
+ $X2=0.23 $Y2=4.8
cc_374 N_A_714_47#_c_434_n N_A_620_911#_c_617_n 0.014378f $X=4.555 $Y=3.235
+ $X2=0.23 $Y2=4.8
cc_375 N_A_714_47#_c_409_n N_A_620_911#_c_595_n 0.0241447f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_376 N_A_714_47#_c_434_n N_A_620_911#_c_595_n 0.00429612f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_377 N_A_714_47#_c_409_n N_A_620_911#_c_596_n 0.0112348f $X=4.39 $Y=3.555
+ $X2=2.185 $Y2=0.62
cc_378 N_A_714_47#_c_405_n N_A_620_911#_c_597_n 0.00516777f $X=4.27 $Y=2.58
+ $X2=2.775 $Y2=5.355
cc_379 N_A_714_47#_c_409_n N_A_620_911#_c_597_n 0.00294758f $X=4.39 $Y=3.555
+ $X2=2.775 $Y2=5.355
cc_380 N_A_714_47#_c_434_n N_A_620_911#_c_597_n 0.0174384f $X=4.555 $Y=3.235
+ $X2=2.775 $Y2=5.355
cc_381 N_A_714_47#_c_405_n N_A_620_911#_c_598_n 9.46557e-19 $X=4.27 $Y=2.58
+ $X2=2.775 $Y2=4.7
cc_382 N_A_714_47#_c_408_n N_A_620_911#_c_598_n 0.0121174f $X=3.765 $Y=3.47
+ $X2=2.775 $Y2=4.7
cc_383 N_A_714_47#_c_426_n N_A_620_911#_c_598_n 0.0118139f $X=4.105 $Y=2.49
+ $X2=2.775 $Y2=4.7
cc_384 N_A_714_47#_c_427_n N_A_620_911#_c_623_n 0.0110028f $X=4.705 $Y=2.58
+ $X2=3.28 $Y2=0.085
cc_385 N_A_714_47#_M1021_g N_A_620_911#_c_623_n 0.0043455f $X=4.78 $Y=1.955
+ $X2=3.28 $Y2=0.085
cc_386 N_A_714_47#_c_408_n N_A_620_911#_c_623_n 0.00251195f $X=3.765 $Y=3.47
+ $X2=3.28 $Y2=0.085
cc_387 N_A_714_47#_c_411_n N_A_620_911#_c_623_n 0.0372645f $X=4.105 $Y=2.07
+ $X2=3.28 $Y2=0.085
cc_388 N_A_714_47#_c_412_n N_A_620_911#_c_623_n 0.00490309f $X=4.105 $Y=2.07
+ $X2=3.28 $Y2=0.085
cc_389 N_A_714_47#_c_413_n N_A_620_911#_c_623_n 0.00567249f $X=4.475 $Y=0.855
+ $X2=3.28 $Y2=0.085
cc_390 N_A_714_47#_c_426_n N_A_620_911#_c_623_n 0.00754333f $X=4.105 $Y=2.49
+ $X2=3.28 $Y2=0.085
cc_391 N_A_714_47#_c_409_n N_A_620_911#_c_599_n 0.00345728f $X=4.39 $Y=3.555
+ $X2=3.28 $Y2=0.42
cc_392 N_A_714_47#_M1021_g N_A_1032_911#_c_734_n 0.0177359f $X=4.78 $Y=1.955
+ $X2=0 $Y2=0
cc_393 N_A_714_47#_M1021_g N_VPWR_c_809_n 0.00295399f $X=4.78 $Y=1.955 $X2=0
+ $Y2=0
cc_394 N_A_714_47#_c_409_n N_VPWR_c_810_n 0.0121345f $X=4.39 $Y=3.555 $X2=0
+ $Y2=0
cc_395 N_A_714_47#_c_434_n N_VPWR_c_810_n 0.0145663f $X=4.555 $Y=3.235 $X2=0
+ $Y2=0
cc_396 N_A_714_47#_c_427_n N_VPWR_c_807_n 0.00492007f $X=4.705 $Y=2.58 $X2=0
+ $Y2=0
cc_397 N_A_714_47#_c_405_n N_VPWR_c_807_n 0.00298594f $X=4.27 $Y=2.58 $X2=0
+ $Y2=0
cc_398 N_A_714_47#_M1021_g N_VPWR_c_807_n 0.00197299f $X=4.78 $Y=1.955 $X2=0
+ $Y2=0
cc_399 N_A_714_47#_c_408_n N_VPWR_c_807_n 0.0244983f $X=3.765 $Y=3.47 $X2=0
+ $Y2=0
cc_400 N_A_714_47#_c_409_n N_VPWR_c_807_n 0.0055128f $X=4.39 $Y=3.555 $X2=0
+ $Y2=0
cc_401 N_A_714_47#_c_411_n N_VPWR_c_807_n 2.07821e-19 $X=4.105 $Y=2.07 $X2=0
+ $Y2=0
cc_402 N_A_714_47#_c_412_n N_VPWR_c_807_n 0.00102999f $X=4.105 $Y=2.07 $X2=0
+ $Y2=0
cc_403 N_A_714_47#_c_434_n N_VPWR_c_807_n 0.00647659f $X=4.555 $Y=3.235 $X2=0
+ $Y2=0
cc_404 N_A_714_47#_c_426_n N_VPWR_c_807_n 0.0186535f $X=4.105 $Y=2.49 $X2=0
+ $Y2=0
cc_405 N_A_714_47#_c_413_n N_X_c_924_n 0.00263398f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_406 N_A_c_532_n N_A_620_911#_c_623_n 0.0037239f $X=4.71 $Y=1.145 $X2=3.28
+ $Y2=0.085
cc_407 N_A_M1012_g N_A_1032_911#_M1006_g 0.00987876f $X=4.785 $Y=0.56 $X2=6.71
+ $Y2=0.235
cc_408 N_A_c_532_n N_A_1032_911#_c_726_n 0.00987876f $X=4.71 $Y=1.145 $X2=0
+ $Y2=0
cc_409 N_A_M1013_g N_VPWR_c_807_n 0.00543198f $X=2.45 $Y=1.985 $X2=0 $Y2=0
cc_410 N_A_c_532_n N_X_c_924_n 7.02896e-19 $X=4.71 $Y=1.145 $X2=0 $Y2=0
cc_411 N_A_620_911#_c_607_n N_A_1032_911#_c_734_n 0.00897291f $X=5.16 $Y=2.94
+ $X2=0 $Y2=0
cc_412 N_A_620_911#_c_607_n N_A_1032_911#_M1008_g 0.00864604f $X=5.16 $Y=2.94
+ $X2=0 $Y2=0
cc_413 N_A_620_911#_c_614_n N_A_1032_911#_c_737_n 0.00864604f $X=5.235 $Y=4.045
+ $X2=0 $Y2=0
cc_414 N_A_620_911#_M1001_g N_A_1032_911#_c_747_n 0.00864604f $X=5.235 $Y=3.485
+ $X2=0 $Y2=0
cc_415 N_A_620_911#_M1001_g N_A_1032_911#_c_749_n 0.00786959f $X=5.235 $Y=3.485
+ $X2=0 $Y2=0
cc_416 N_A_620_911#_M1011_g N_A_1032_911#_c_728_n 0.0254294f $X=5.085 $Y=4.88
+ $X2=3.28 $Y2=0.42
cc_417 N_A_620_911#_c_614_n N_A_1032_911#_c_728_n 0.00641748f $X=5.235 $Y=4.045
+ $X2=3.28 $Y2=0.42
cc_418 N_A_620_911#_M1011_g N_A_1032_911#_c_732_n 0.00384336f $X=5.085 $Y=4.88
+ $X2=3.67 $Y2=4.735
cc_419 N_A_620_911#_c_623_n N_VPWR_c_809_n 0.035645f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_420 N_A_620_911#_c_607_n N_VPWR_c_810_n 0.0189101f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_421 N_A_620_911#_c_608_n N_VPWR_c_810_n 0.00521099f $X=5.01 $Y=4.045 $X2=0
+ $Y2=0
cc_422 N_A_620_911#_c_597_n N_VPWR_c_810_n 0.00509169f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_423 N_A_620_911#_c_597_n N_VPWR_c_814_n 0.00305029f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_424 N_A_620_911#_c_623_n N_VPWR_c_814_n 0.00537241f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_425 N_A_620_911#_c_607_n N_VPWR_c_815_n 0.004734f $X=5.16 $Y=2.94 $X2=0 $Y2=0
cc_426 N_A_620_911#_c_601_n N_VPWR_c_807_n 0.00365797f $X=4.705 $Y=2.94 $X2=0
+ $Y2=0
cc_427 N_A_620_911#_c_579_n N_VPWR_c_807_n 0.00398455f $X=4.27 $Y=2.94 $X2=0
+ $Y2=0
cc_428 N_A_620_911#_c_607_n N_VPWR_c_807_n 0.00671142f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_429 N_A_620_911#_c_612_n N_VPWR_c_807_n 0.00339161f $X=4.78 $Y=2.94 $X2=0
+ $Y2=0
cc_430 N_A_620_911#_c_617_n N_VPWR_c_807_n 0.00622378f $X=4.105 $Y=3.135 $X2=0
+ $Y2=0
cc_431 N_A_620_911#_c_597_n N_VPWR_c_807_n 0.0219288f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_432 N_A_620_911#_c_598_n N_VPWR_c_807_n 0.00663704f $X=4.19 $Y=2.83 $X2=0
+ $Y2=0
cc_433 N_A_620_911#_c_623_n N_VPWR_c_807_n 0.0165665f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_434 N_A_1032_911#_c_734_n N_VPWR_c_809_n 0.00897993f $X=5.255 $Y=1.41 $X2=0
+ $Y2=0
cc_435 N_A_1032_911#_M1008_g N_VPWR_c_810_n 0.00163667f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_436 N_A_1032_911#_c_747_n N_VPWR_c_810_n 8.67432e-19 $X=5.775 $Y=3.065 $X2=0
+ $Y2=0
cc_437 N_A_1032_911#_c_749_n N_VPWR_c_810_n 0.00470553f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_438 N_A_1032_911#_M1008_g N_VPWR_c_812_n 0.00377671f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_439 N_A_1032_911#_M1015_g N_VPWR_c_812_n 0.00372221f $X=6.205 $Y=1.985 $X2=0
+ $Y2=0
cc_440 N_A_1032_911#_c_719_n N_VPWR_c_812_n 0.00228736f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_441 N_A_1032_911#_M1016_g N_VPWR_c_813_n 0.00741785f $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_442 N_A_1032_911#_c_734_n N_VPWR_c_815_n 0.00545125f $X=5.255 $Y=1.41 $X2=0
+ $Y2=0
cc_443 N_A_1032_911#_M1008_g N_VPWR_c_815_n 0.0154662f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_1032_911#_c_749_n N_VPWR_c_815_n 0.00839873f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_445 N_A_1032_911#_c_739_n N_VPWR_c_816_n 0.00325633f $X=6.13 $Y=3.065 $X2=0
+ $Y2=0
cc_446 N_A_1032_911#_M1015_g N_VPWR_c_817_n 0.0132738f $X=6.205 $Y=1.985 $X2=0
+ $Y2=0
cc_447 N_A_1032_911#_c_742_n N_VPWR_c_817_n 0.00299145f $X=6.56 $Y=3.065 $X2=0
+ $Y2=0
cc_448 N_A_1032_911#_M1016_g N_VPWR_c_817_n 0.0152247f $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_449 N_A_1032_911#_c_734_n N_VPWR_c_807_n 0.00412295f $X=5.255 $Y=1.41 $X2=0
+ $Y2=0
cc_450 N_A_1032_911#_M1008_g N_VPWR_c_807_n 0.00920492f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_451 N_A_1032_911#_c_739_n N_VPWR_c_807_n 0.00181102f $X=6.13 $Y=3.065 $X2=0
+ $Y2=0
cc_452 N_A_1032_911#_M1015_g N_VPWR_c_807_n 0.00691128f $X=6.205 $Y=1.985 $X2=0
+ $Y2=0
cc_453 N_A_1032_911#_c_742_n N_VPWR_c_807_n 0.00181102f $X=6.56 $Y=3.065 $X2=0
+ $Y2=0
cc_454 N_A_1032_911#_M1016_g N_VPWR_c_807_n 0.00988127f $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_1032_911#_c_749_n N_VPWR_c_807_n 0.00327036f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_456 N_A_1032_911#_M1007_g N_X_c_916_n 0.00498668f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_457 N_A_1032_911#_c_710_n N_X_c_919_n 0.00792257f $X=5.7 $Y=1.247 $X2=0 $Y2=0
cc_458 N_A_1032_911#_c_719_n N_X_c_919_n 0.0552661f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_459 N_A_1032_911#_M1016_g N_X_c_927_n 7.94882e-19 $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_460 N_A_1032_911#_M1017_g N_X_c_920_n 0.00496787f $X=6.205 $Y=0.56 $X2=0
+ $Y2=0
cc_461 N_A_1032_911#_M1018_g N_X_c_920_n 0.00458369f $X=6.635 $Y=0.56 $X2=0
+ $Y2=0
cc_462 N_A_1032_911#_c_719_n N_X_c_940_n 0.0308881f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_463 N_A_1032_911#_M1006_g N_X_c_924_n 0.00446469f $X=5.255 $Y=0.56 $X2=0
+ $Y2=0
cc_464 N_A_1032_911#_c_710_n N_X_c_924_n 0.0290305f $X=5.7 $Y=1.247 $X2=0 $Y2=0
cc_465 N_A_1032_911#_M1007_g N_X_c_924_n 0.00667268f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_466 N_A_1032_911#_c_734_n X 0.00308224f $X=5.255 $Y=1.41 $X2=0 $Y2=0
cc_467 N_A_1032_911#_M1008_g X 0.0103699f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_468 N_VPWR_c_807_n N_X_M1002_d 0.00216609f $X=7.13 $Y=2.72 $X2=3.135
+ $Y2=0.235
cc_469 N_VPWR_c_807_n N_X_M1015_d 0.00133453f $X=7.13 $Y=2.72 $X2=3.53 $Y2=4.555
cc_470 N_VPWR_c_812_n N_X_c_919_n 0.0121443f $X=5.99 $Y=1.79 $X2=0 $Y2=0
cc_471 N_VPWR_c_812_n N_X_c_927_n 0.0273305f $X=5.99 $Y=1.79 $X2=0 $Y2=0
cc_472 N_VPWR_c_813_n N_X_c_927_n 0.00424153f $X=6.85 $Y=1.79 $X2=0 $Y2=0
cc_473 N_VPWR_c_817_n N_X_c_927_n 0.00966848f $X=6.755 $Y=2.72 $X2=0 $Y2=0
cc_474 N_VPWR_c_807_n N_X_c_927_n 0.00302523f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_475 N_VPWR_c_809_n X 0.0230063f $X=5.005 $Y=1.79 $X2=0 $Y2=0
cc_476 N_VPWR_c_812_n X 0.021786f $X=5.99 $Y=1.79 $X2=0 $Y2=0
cc_477 N_VPWR_c_815_n X 0.0113333f $X=5.905 $Y=2.72 $X2=0 $Y2=0
cc_478 N_VPWR_c_807_n X 0.00302523f $X=7.13 $Y=2.72 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a311oi_2.spice
* Created: Thu Aug 27 14:04:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a311oi_2.spice.pex"
.subckt sky130_fd_sc_hd__a311oi_2  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1009 N_A_27_47#_M1009_d N_A3_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1019 N_A_27_47#_M1019_d N_A3_M1019_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1015 N_A_27_47#_M1019_d N_A2_M1015_g N_A_277_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_27_47#_M1016_d N_A2_M1016_g N_A_277_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1010_d N_A1_M1010_g N_A_277_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1012_d N_A1_M1012_g N_A_277_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.0975 AS=0.08775 PD=0.95 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_B1_M1007_g N_Y_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.0975 PD=0.92 PS=0.95 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75001.1
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1007_d N_B1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.17 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1011_s N_C1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.17 PS=0.92 NRD=45.228 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_C1_M1013_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A3_M1006_g N_A_109_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A3_M1017_g N_A_109_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1002 N_A_109_297#_M1002_d N_A2_M1002_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1018 N_A_109_297#_M1002_d N_A2_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.145 PD=1.28 PS=1.29 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1018_s N_A1_M1000_g N_A_109_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.135 PD=1.29 PS=1.27 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_109_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_641_297#_M1001_d N_B1_M1001_g N_A_109_297#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1005 N_A_641_297#_M1005_d N_B1_M1005_g N_A_109_297#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=1.52 PS=1.27 NRD=19.7 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g N_A_641_297#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=1.52 NRD=0 NRS=27.5603 M=1 R=6.66667 SA=75001.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1014 N_Y_M1004_d N_C1_M1014_g N_A_641_297#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__a311oi_2.spice.SKY130_FD_SC_HD__A311OI_2.pxi"
*
.ends
*
*

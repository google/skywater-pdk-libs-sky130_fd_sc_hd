* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4.pxi.spice
* Created: Tue Sep  1 19:13:28 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%LOWLVPWR N_LOWLVPWR_M1013_s
+ N_LOWLVPWR_M1013_b N_LOWLVPWR_c_122_p N_LOWLVPWR_c_108_p N_LOWLVPWR_c_114_p
+ N_LOWLVPWR_c_98_n N_LOWLVPWR_c_99_n N_LOWLVPWR_c_112_p N_LOWLVPWR_c_100_n
+ LOWLVPWR N_LOWLVPWR_c_101_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%LOWLVPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_505_297# N_A_505_297#_M1014_d
+ N_A_505_297#_M1013_d N_A_505_297#_c_211_n N_A_505_297#_M1003_g
+ N_A_505_297#_c_212_n N_A_505_297#_M1010_g N_A_505_297#_c_213_n
+ N_A_505_297#_c_214_n N_A_505_297#_c_215_n N_A_505_297#_M1019_g
+ N_A_505_297#_c_216_n N_A_505_297#_c_217_n N_A_505_297#_M1020_g
+ N_A_505_297#_c_218_n N_A_505_297#_c_219_n N_A_505_297#_c_220_n
+ N_A_505_297#_c_229_n N_A_505_297#_c_221_n N_A_505_297#_c_222_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_505_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_714_47# N_A_714_47#_M1004_d
+ N_A_714_47#_M1009_d N_A_714_47#_M1000_s N_A_714_47#_c_302_n
+ N_A_714_47#_c_293_n N_A_714_47#_M1021_g N_A_714_47#_c_383_p
+ N_A_714_47#_c_294_n N_A_714_47#_c_295_n N_A_714_47#_c_296_n
+ N_A_714_47#_c_297_n N_A_714_47#_c_298_n N_A_714_47#_c_299_n
+ N_A_714_47#_c_300_n N_A_714_47#_c_312_n N_A_714_47#_c_386_p
+ N_A_714_47#_c_301_n PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_714_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A N_A_M1013_g N_A_c_394_n
+ N_A_M1014_g N_A_c_395_n N_A_M1004_g N_A_c_397_n N_A_c_398_n N_A_M1005_g
+ N_A_c_400_n N_A_M1009_g N_A_c_402_n N_A_M1012_g N_A_c_404_n N_A_c_405_n
+ N_A_c_406_n A N_A_c_407_n PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_620_911# N_A_620_911#_M1003_d
+ N_A_620_911#_M1019_d N_A_620_911#_M1021_s N_A_620_911#_c_476_n
+ N_A_620_911#_c_464_n N_A_620_911#_c_478_n N_A_620_911#_M1000_g
+ N_A_620_911#_c_480_n N_A_620_911#_c_481_n N_A_620_911#_M1011_g
+ N_A_620_911#_M1001_g N_A_620_911#_c_484_n N_A_620_911#_c_485_n
+ N_A_620_911#_c_486_n N_A_620_911#_c_493_n N_A_620_911#_c_466_n
+ N_A_620_911#_c_499_n N_A_620_911#_c_501_n N_A_620_911#_c_522_n
+ N_A_620_911#_c_467_n N_A_620_911#_c_468_n N_A_620_911#_c_469_n
+ N_A_620_911#_c_470_n N_A_620_911#_c_475_n N_A_620_911#_c_471_n
+ N_A_620_911#_c_472_n PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_620_911#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_1032_911#
+ N_A_1032_911#_M1011_d N_A_1032_911#_M1001_d N_A_1032_911#_M1006_g
+ N_A_1032_911#_c_591_n N_A_1032_911#_M1002_g N_A_1032_911#_c_582_n
+ N_A_1032_911#_M1007_g N_A_1032_911#_M1008_g N_A_1032_911#_c_598_n
+ N_A_1032_911#_c_599_n N_A_1032_911#_M1017_g N_A_1032_911#_M1015_g
+ N_A_1032_911#_c_601_n N_A_1032_911#_c_585_n N_A_1032_911#_M1018_g
+ N_A_1032_911#_M1016_g N_A_1032_911#_c_587_n N_A_1032_911#_c_605_n
+ N_A_1032_911#_c_606_n N_A_1032_911#_c_607_n N_A_1032_911#_c_588_n
+ N_A_1032_911#_c_589_n N_A_1032_911#_c_590_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%A_1032_911#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%VPWR N_VPWR_M1000_d
+ N_VPWR_M1021_d N_VPWR_M1008_s N_VPWR_M1016_s N_VPWR_c_682_n N_VPWR_c_700_n
+ N_VPWR_c_683_n N_VPWR_c_684_n N_VPWR_c_703_n N_VPWR_c_685_n N_VPWR_c_705_n
+ N_VPWR_c_686_n N_VPWR_c_707_n VPWR N_VPWR_c_675_n N_VPWR_c_691_n
+ N_VPWR_c_676_n VPWR PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%X N_X_M1006_d N_X_M1017_d
+ N_X_M1002_d N_X_M1015_d N_X_c_783_n N_X_c_784_n N_X_c_777_n N_X_c_774_n
+ N_X_c_789_n X X N_X_c_775_n X PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%X
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%VGND N_VGND_M1014_s
+ N_VGND_M1003_s N_VGND_M1004_s N_VGND_M1010_s N_VGND_M1005_s N_VGND_M1020_s
+ N_VGND_M1012_s N_VGND_M1007_s N_VGND_M1018_s N_VGND_c_817_n N_VGND_c_818_n
+ N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n
+ N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n
+ N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n
+ N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n
+ N_VGND_c_839_n VGND VGND N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n
+ N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4%VGND
cc_1 VNB N_LOWLVPWR_c_98_n 0.00447854f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=2.2
cc_2 VNB N_LOWLVPWR_c_99_n 0.0244366f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.2
cc_3 VNB N_LOWLVPWR_c_100_n 0.0306316f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=2.2
cc_4 VNB N_LOWLVPWR_c_101_n 0.0344347f $X=-0.19 $Y=-0.24 $X2=2.06 $Y2=2.2
cc_5 VNB N_A_505_297#_c_211_n 0.0179052f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.305
cc_6 VNB N_A_505_297#_c_212_n 0.0140848f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.79
cc_7 VNB N_A_505_297#_c_213_n 0.0130779f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.335
cc_8 VNB N_A_505_297#_c_214_n 0.0294363f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.66
cc_9 VNB N_A_505_297#_c_215_n 0.0140848f $X=-0.19 $Y=-0.24 $X2=2.435 $Y2=3.49
cc_10 VNB N_A_505_297#_c_216_n 0.0195784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_505_297#_c_217_n 0.0162763f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=2.2
cc_12 VNB N_A_505_297#_c_218_n 0.00569361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_505_297#_c_219_n 0.00997858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_505_297#_c_220_n 0.016089f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=2.2
cc_15 VNB N_A_505_297#_c_221_n 0.0360066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_505_297#_c_222_n 0.0848642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_714_47#_c_293_n 0.0129761f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.79
cc_18 VNB N_A_714_47#_c_294_n 0.0175549f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=2.2
cc_19 VNB N_A_714_47#_c_295_n 0.00241554f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=2.2
cc_20 VNB N_A_714_47#_c_296_n 0.00454289f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.2
cc_21 VNB N_A_714_47#_c_297_n 0.0397033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_714_47#_c_298_n 0.0516547f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=2.21
cc_23 VNB N_A_714_47#_c_299_n 0.00893993f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=2.2
cc_24 VNB N_A_714_47#_c_300_n 0.00805719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_714_47#_c_301_n 0.00576889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_M1013_g 0.00675179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_c_394_n 0.0408343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_c_395_n 0.0352506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_M1004_g 0.0240979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_c_397_n 0.0168496f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.66
cc_31 VNB N_A_c_398_n 0.0656946f $X=-0.19 $Y=-0.24 $X2=2.435 $Y2=3.49
cc_32 VNB N_A_M1005_g 0.0189456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_c_400_n 0.0149976f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=2.2
cc_34 VNB N_A_M1009_g 0.018948f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.2
cc_35 VNB N_A_c_402_n 0.0255444f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.2
cc_36 VNB N_A_M1012_g 0.0204702f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=2.2
cc_37 VNB N_A_c_404_n 0.017446f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=2.14
cc_38 VNB N_A_c_405_n 0.00933068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_c_406_n 0.0106787f $X=-0.19 $Y=-0.24 $X2=2.06 $Y2=2.2
cc_40 VNB N_A_c_407_n 0.0169952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_620_911#_c_464_n 0.0127228f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.79
cc_42 VNB N_A_620_911#_M1011_g 0.0484682f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.2
cc_43 VNB N_A_620_911#_c_466_n 0.0181882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_620_911#_c_467_n 0.0561622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_620_911#_c_468_n 0.0016479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_620_911#_c_469_n 7.55444e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_620_911#_c_470_n 9.83343e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_620_911#_c_471_n 0.00843783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_620_911#_c_472_n 0.0133087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1032_911#_M1006_g 0.0226878f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.065
cc_51 VNB N_A_1032_911#_c_582_n 0.0140243f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.66
cc_52 VNB N_A_1032_911#_M1007_g 0.0216078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1032_911#_M1017_g 0.0205125f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=2.2
cc_54 VNB N_A_1032_911#_c_585_n 0.0411217f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=2.21
cc_55 VNB N_A_1032_911#_M1018_g 0.0282249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1032_911#_c_587_n 0.0111194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1032_911#_c_588_n 0.00998896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1032_911#_c_589_n 0.0492761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1032_911#_c_590_n 0.0384737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VPWR_c_675_n 0.0363208f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VPWR_c_676_n 0.0822527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_X_c_774_n 0.00373262f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=2.2
cc_63 VNB N_X_c_775_n 0.00503584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_817_n 0.0499252f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=2.2
cc_65 VNB N_VGND_c_818_n 0.0415677f $X=-0.19 $Y=-0.24 $X2=2.06 $Y2=2.2
cc_66 VNB N_VGND_c_819_n 0.0154203f $X=-0.19 $Y=-0.24 $X2=0.465 $Y2=2.21
cc_67 VNB N_VGND_c_820_n 0.00639522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_821_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_822_n 0.0148483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_823_n 0.0147312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_824_n 3.41575e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_825_n 0.0402365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_826_n 0.0863125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_827_n 0.00497181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_828_n 0.0225099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_829_n 0.00513431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_830_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_831_n 0.00362205f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_832_n 0.012302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_833_n 0.0043669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_834_n 0.0123057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_835_n 0.00513431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_836_n 0.0170886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_837_n 0.00439458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_838_n 0.0159319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_839_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_840_n 0.0664237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_841_n 0.0182639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_842_n 0.0745763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_843_n 0.525069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_844_n 0.0134401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_845_n 0.459147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_846_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_847_n 0.00978383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 noxref_2 N_LOWLVPWR_c_100_n 0.0309709f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=2.2
cc_96 noxref_2 N_VPWR_c_675_n 0.0228594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 noxref_2 N_VPWR_c_676_n 0.0549811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 N_LOWLVPWR_c_99_n VPB 0.0251748f $X=2.225 $Y=2.2 $X2=-0.19 $Y2=-0.24
cc_99 N_LOWLVPWR_c_99_n N_A_505_297#_M1013_d 0.00144688f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_100 N_LOWLVPWR_M1013_b N_A_505_297#_c_219_n 0.0037173f $X=1.92 $Y=1.305 $X2=0
+ $Y2=0
cc_101 N_LOWLVPWR_c_99_n N_A_505_297#_c_219_n 3.15819e-19 $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_102 N_LOWLVPWR_M1013_b N_A_505_297#_c_220_n 0.00974718f $X=1.92 $Y=1.305
+ $X2=0 $Y2=0
cc_103 N_LOWLVPWR_c_108_p N_A_505_297#_c_220_n 3.29394e-19 $X=2.645 $Y=3.49
+ $X2=0 $Y2=0
cc_104 N_LOWLVPWR_c_99_n N_A_505_297#_c_220_n 0.0372262f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_105 N_LOWLVPWR_c_108_p N_A_505_297#_c_229_n 0.00924483f $X=2.645 $Y=3.49
+ $X2=0 $Y2=0
cc_106 N_LOWLVPWR_c_99_n N_A_505_297#_c_229_n 0.0204768f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_107 N_LOWLVPWR_c_112_p N_A_505_297#_c_229_n 0.0100174f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_108 N_LOWLVPWR_c_108_p N_A_505_297#_c_221_n 0.0678602f $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_109 N_LOWLVPWR_c_114_p N_A_505_297#_c_221_n 0.00525651f $X=2.435 $Y=2.66
+ $X2=0 $Y2=0
cc_110 N_LOWLVPWR_c_108_p N_A_505_297#_c_222_n 0.00169032f $X=2.645 $Y=3.49
+ $X2=0 $Y2=0
cc_111 N_LOWLVPWR_c_99_n N_A_714_47#_c_302_n 5.4797e-19 $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_112 N_LOWLVPWR_c_99_n N_A_714_47#_M1021_g 0.00777495f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_113 N_LOWLVPWR_c_99_n N_A_714_47#_c_297_n 0.0182669f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_114 N_LOWLVPWR_c_99_n N_A_714_47#_c_298_n 0.0104851f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_115 N_LOWLVPWR_c_99_n N_A_714_47#_c_301_n 0.00926075f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_116 N_LOWLVPWR_M1013_b N_A_M1013_g 0.0304234f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_117 N_LOWLVPWR_c_122_p N_A_M1013_g 0.00523247f $X=2.225 $Y=1.79 $X2=0 $Y2=0
cc_118 N_LOWLVPWR_c_108_p N_A_M1013_g 0.0055008f $X=2.645 $Y=3.49 $X2=0 $Y2=0
cc_119 N_LOWLVPWR_c_114_p N_A_M1013_g 0.00938999f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_120 N_LOWLVPWR_c_99_n N_A_M1013_g 0.00645994f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_121 N_LOWLVPWR_c_112_p N_A_M1013_g 0.00218038f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_122 N_LOWLVPWR_M1013_b N_A_c_398_n 0.00316885f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_123 N_LOWLVPWR_M1013_b N_A_c_407_n 0.00111856f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_124 N_LOWLVPWR_c_99_n N_A_c_407_n 0.00229296f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_125 N_LOWLVPWR_c_99_n N_A_620_911#_M1021_s 0.00479759f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_126 N_LOWLVPWR_c_99_n N_A_620_911#_c_469_n 0.0011695f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_127 N_LOWLVPWR_c_99_n N_A_620_911#_c_475_n 0.0174341f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_128 N_LOWLVPWR_c_99_n N_A_1032_911#_c_591_n 0.00737951f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_129 N_LOWLVPWR_c_99_n N_A_1032_911#_M1008_g 0.00870505f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_130 N_LOWLVPWR_c_99_n N_A_1032_911#_M1015_g 0.00715996f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_131 N_LOWLVPWR_c_99_n N_A_1032_911#_M1016_g 0.00712859f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_132 N_LOWLVPWR_c_99_n N_VPWR_M1021_d 0.00413567f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_133 N_LOWLVPWR_c_99_n N_VPWR_M1008_s 0.00463513f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_134 N_LOWLVPWR_c_99_n N_VPWR_M1016_s 0.00454198f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_135 N_LOWLVPWR_c_99_n N_VPWR_c_682_n 0.0221365f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_136 N_LOWLVPWR_c_99_n N_VPWR_c_683_n 0.0172645f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_137 N_LOWLVPWR_c_99_n N_VPWR_c_684_n 0.0200894f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_138 N_LOWLVPWR_c_99_n N_VPWR_c_685_n 0.00466952f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_139 N_LOWLVPWR_c_99_n N_VPWR_c_686_n 0.00411278f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_140 N_LOWLVPWR_c_114_p N_VPWR_c_675_n 0.0123972f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_141 N_LOWLVPWR_c_98_n N_VPWR_c_675_n 5.76636e-19 $X=1.475 $Y=2.2 $X2=0 $Y2=0
cc_142 N_LOWLVPWR_c_100_n N_VPWR_c_675_n 0.00675753f $X=1.36 $Y=2.2 $X2=0 $Y2=0
cc_143 N_LOWLVPWR_c_101_n N_VPWR_c_675_n 0.01865f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_144 N_LOWLVPWR_c_99_n N_VPWR_c_691_n 0.00185735f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_145 N_LOWLVPWR_M1013_b N_VPWR_c_676_n 0.0147849f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_146 N_LOWLVPWR_c_108_p N_VPWR_c_676_n 0.0879787f $X=2.645 $Y=3.49 $X2=0 $Y2=0
cc_147 N_LOWLVPWR_c_114_p N_VPWR_c_676_n 0.02138f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_148 N_LOWLVPWR_c_98_n N_VPWR_c_676_n 0.0948062f $X=1.475 $Y=2.2 $X2=0 $Y2=0
cc_149 N_LOWLVPWR_c_99_n N_VPWR_c_676_n 0.418194f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_150 N_LOWLVPWR_c_100_n N_VPWR_c_676_n 0.116739f $X=1.36 $Y=2.2 $X2=0 $Y2=0
cc_151 N_LOWLVPWR_c_101_n N_VPWR_c_676_n 0.00970859f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_152 N_LOWLVPWR_c_99_n N_X_M1002_d 0.0041104f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_153 N_LOWLVPWR_c_99_n N_X_c_777_n 0.0245217f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_154 N_LOWLVPWR_c_99_n X 0.0251052f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_155 VPB N_A_714_47#_c_302_n 0.0256732f $X=4.25 $Y=1.305 $X2=2.225 $Y2=1.79
cc_156 VPB N_A_714_47#_c_293_n 5.34541e-19 $X=4.25 $Y=1.305 $X2=2.225 $Y2=1.79
cc_157 VPB N_A_714_47#_M1021_g 0.0198732f $X=4.25 $Y=1.305 $X2=2.225 $Y2=2.66
cc_158 VPB N_A_714_47#_c_295_n 0.00466811f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_159 VPB N_A_714_47#_c_298_n 0.0149067f $X=4.25 $Y=1.305 $X2=1.36 $Y2=2.21
cc_160 VPB N_A_714_47#_c_312_n 0.00449536f $X=4.25 $Y=1.305 $X2=2.06 $Y2=2.2
cc_161 VPB N_A_620_911#_c_476_n 0.0169344f $X=4.25 $Y=1.305 $X2=2.225 $Y2=1.79
cc_162 VPB N_A_620_911#_c_464_n 5.21411e-19 $X=4.25 $Y=1.305 $X2=2.225 $Y2=1.79
cc_163 VPB N_A_620_911#_c_478_n 0.0246766f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_620_911#_M1000_g 0.00259316f $X=4.25 $Y=1.305 $X2=2.435 $Y2=2.66
cc_165 VPB N_A_620_911#_c_480_n 0.0249303f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_620_911#_c_481_n 0.0094712f $X=4.25 $Y=1.305 $X2=1.475 $Y2=2.2
cc_167 VPB N_A_620_911#_M1011_g 0.00114838f $X=4.25 $Y=1.305 $X2=2.225 $Y2=2.2
cc_168 VPB N_A_620_911#_M1001_g 0.0064606f $X=4.25 $Y=1.305 $X2=1.36 $Y2=2.21
cc_169 VPB N_A_620_911#_c_484_n 0.00400906f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_620_911#_c_485_n 0.00698872f $X=4.25 $Y=1.305 $X2=0.435 $Y2=2.14
cc_171 VPB N_A_620_911#_c_486_n 0.0141637f $X=4.25 $Y=1.305 $X2=2.06 $Y2=2.2
cc_172 VPB N_A_620_911#_c_467_n 0.0188917f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_620_911#_c_469_n 0.00337762f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_620_911#_c_475_n 0.00324872f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_620_911#_c_472_n 6.57859e-19 $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1032_911#_c_591_n 0.0147881f $X=4.25 $Y=1.305 $X2=2.225 $Y2=1.79
cc_177 VPB N_A_1032_911#_c_582_n 0.00953288f $X=4.25 $Y=1.305 $X2=2.225 $Y2=2.66
cc_178 VPB N_A_1032_911#_M1008_g 0.0277715f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_179 VPB N_A_1032_911#_c_598_n 0.0664838f $X=4.25 $Y=1.305 $X2=2.225 $Y2=2.2
cc_180 VPB N_A_1032_911#_c_599_n 0.0212205f $X=4.25 $Y=1.305 $X2=2.225 $Y2=2.2
cc_181 VPB N_A_1032_911#_M1015_g 0.0202696f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_182 VPB N_A_1032_911#_c_601_n 0.0401913f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1032_911#_c_585_n 0.0223728f $X=4.25 $Y=1.305 $X2=0.465 $Y2=2.21
cc_184 VPB N_A_1032_911#_M1016_g 0.0355931f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1032_911#_c_587_n 0.00747506f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1032_911#_c_605_n 0.00596971f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1032_911#_c_606_n 0.0106787f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1032_911#_c_607_n 0.00808952f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1032_911#_c_588_n 0.00143619f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1032_911#_c_589_n 0.00628335f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1032_911#_c_590_n 0.0238154f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_682_n 0.00429074f $X=4.25 $Y=1.305 $X2=2.435 $Y2=3.49
cc_193 VPB N_VPWR_c_700_n 0.00447924f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_683_n 0.00379002f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_195 VPB N_VPWR_c_684_n 0.00404706f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_703_n 0.00101664f $X=4.25 $Y=1.305 $X2=1.36 $Y2=2.2
cc_197 VPB N_VPWR_c_685_n 0.0107502f $X=4.25 $Y=1.305 $X2=0.435 $Y2=2.14
cc_198 VPB N_VPWR_c_705_n 0.0021751f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_686_n 0.00753446f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_200 VPB N_VPWR_c_707_n 0.00258752f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_691_n 0.0156676f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_676_n 0.0813942f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_X_c_777_n 0.00374381f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_204 VPB X 0.00132567f $X=4.25 $Y=1.305 $X2=1.505 $Y2=2.2
cc_205 N_A_505_297#_c_221_n N_A_714_47#_c_294_n 0.0441264f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_206 N_A_505_297#_c_216_n N_A_714_47#_c_295_n 0.0011083f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_207 N_A_505_297#_c_218_n N_A_714_47#_c_295_n 3.68575e-19 $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_208 N_A_505_297#_c_221_n N_A_714_47#_c_296_n 0.0103626f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_209 N_A_505_297#_c_220_n N_A_714_47#_c_297_n 0.0048486f $X=3.06 $Y=2.25 $X2=0
+ $Y2=0
cc_210 N_A_505_297#_c_221_n N_A_714_47#_c_297_n 9.66994e-19 $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_211 N_A_505_297#_c_220_n N_A_714_47#_c_298_n 0.00327676f $X=3.06 $Y=2.25
+ $X2=0 $Y2=0
cc_212 N_A_505_297#_c_221_n N_A_714_47#_c_298_n 0.00125462f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_213 N_A_505_297#_c_221_n N_A_714_47#_c_301_n 0.0084582f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_214 N_A_505_297#_c_219_n N_A_M1013_g 0.0110528f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_215 N_A_505_297#_c_221_n N_A_M1013_g 0.0027023f $X=3.225 $Y=3.84 $X2=0 $Y2=0
cc_216 N_A_505_297#_c_219_n N_A_c_394_n 0.010267f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_217 N_A_505_297#_c_219_n N_A_c_395_n 0.0218308f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_218 N_A_505_297#_c_219_n N_A_M1004_g 0.00480585f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_219 N_A_505_297#_c_219_n N_A_c_398_n 0.00146935f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_220 N_A_505_297#_c_219_n N_A_c_407_n 0.0360803f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_221 N_A_505_297#_c_220_n N_A_c_407_n 0.00941491f $X=3.06 $Y=2.25 $X2=0 $Y2=0
cc_222 N_A_505_297#_c_216_n N_A_620_911#_c_478_n 0.0155516f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_223 N_A_505_297#_c_216_n N_A_620_911#_M1011_g 0.00777355f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_224 N_A_505_297#_c_211_n N_A_620_911#_c_493_n 0.00968676f $X=3.025 $Y=4.48
+ $X2=0 $Y2=0
cc_225 N_A_505_297#_c_212_n N_A_620_911#_c_493_n 0.00843936f $X=3.455 $Y=4.48
+ $X2=0 $Y2=0
cc_226 N_A_505_297#_c_214_n N_A_620_911#_c_493_n 0.0169132f $X=3.53 $Y=4.405
+ $X2=0 $Y2=0
cc_227 N_A_505_297#_c_215_n N_A_620_911#_c_493_n 2.89638e-19 $X=3.885 $Y=4.48
+ $X2=0 $Y2=0
cc_228 N_A_505_297#_c_214_n N_A_620_911#_c_466_n 0.021891f $X=3.53 $Y=4.405
+ $X2=0 $Y2=0
cc_229 N_A_505_297#_c_222_n N_A_620_911#_c_466_n 0.00420454f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_230 N_A_505_297#_c_221_n N_A_620_911#_c_499_n 0.0226213f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_231 N_A_505_297#_c_222_n N_A_620_911#_c_499_n 0.017913f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_232 N_A_505_297#_c_212_n N_A_620_911#_c_501_n 2.89638e-19 $X=3.455 $Y=4.48
+ $X2=0 $Y2=0
cc_233 N_A_505_297#_c_215_n N_A_620_911#_c_501_n 0.00843936f $X=3.885 $Y=4.48
+ $X2=0 $Y2=0
cc_234 N_A_505_297#_c_216_n N_A_620_911#_c_501_n 0.0149859f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_235 N_A_505_297#_c_217_n N_A_620_911#_c_501_n 0.00985995f $X=4.315 $Y=4.48
+ $X2=0 $Y2=0
cc_236 N_A_505_297#_c_218_n N_A_620_911#_c_501_n 0.00418634f $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_237 N_A_505_297#_c_221_n N_A_620_911#_c_467_n 0.00433954f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_238 N_A_505_297#_c_222_n N_A_620_911#_c_467_n 0.0112331f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_239 N_A_505_297#_c_221_n N_A_620_911#_c_468_n 0.00372705f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_240 N_A_505_297#_c_222_n N_A_620_911#_c_468_n 0.0022314f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_241 N_A_505_297#_c_218_n N_A_620_911#_c_472_n 0.0155516f $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_242 N_A_505_297#_M1013_d N_VPWR_c_676_n 0.00146082f $X=2.525 $Y=1.485 $X2=0
+ $Y2=0
cc_243 N_A_505_297#_c_220_n N_VPWR_c_676_n 0.00782153f $X=3.06 $Y=2.25 $X2=0
+ $Y2=0
cc_244 N_A_505_297#_c_229_n N_VPWR_c_676_n 0.00276885f $X=2.8 $Y=2.25 $X2=0
+ $Y2=0
cc_245 N_A_505_297#_c_221_n N_VPWR_c_676_n 0.0587137f $X=3.225 $Y=3.84 $X2=0
+ $Y2=0
cc_246 N_A_505_297#_c_219_n N_VGND_c_817_n 0.0068636f $X=2.675 $Y=0.62 $X2=0
+ $Y2=0
cc_247 N_A_505_297#_c_211_n N_VGND_c_818_n 0.00414737f $X=3.025 $Y=4.48 $X2=0
+ $Y2=0
cc_248 N_A_505_297#_c_219_n N_VGND_c_819_n 0.0271827f $X=2.675 $Y=0.62 $X2=0
+ $Y2=0
cc_249 N_A_505_297#_c_212_n N_VGND_c_820_n 0.00179869f $X=3.455 $Y=4.48 $X2=0
+ $Y2=0
cc_250 N_A_505_297#_c_213_n N_VGND_c_820_n 0.00240634f $X=3.81 $Y=4.405 $X2=0
+ $Y2=0
cc_251 N_A_505_297#_c_215_n N_VGND_c_820_n 0.00304527f $X=3.885 $Y=4.48 $X2=0
+ $Y2=0
cc_252 N_A_505_297#_c_217_n N_VGND_c_822_n 0.00390324f $X=4.315 $Y=4.48 $X2=0
+ $Y2=0
cc_253 N_A_505_297#_c_219_n N_VGND_c_828_n 0.00966373f $X=2.675 $Y=0.62 $X2=0
+ $Y2=0
cc_254 N_A_505_297#_c_211_n N_VGND_c_830_n 0.0054895f $X=3.025 $Y=4.48 $X2=0
+ $Y2=0
cc_255 N_A_505_297#_c_212_n N_VGND_c_830_n 0.0054895f $X=3.455 $Y=4.48 $X2=0
+ $Y2=0
cc_256 N_A_505_297#_c_215_n N_VGND_c_841_n 0.0054895f $X=3.885 $Y=4.48 $X2=0
+ $Y2=0
cc_257 N_A_505_297#_c_217_n N_VGND_c_841_n 0.0054895f $X=4.315 $Y=4.48 $X2=0
+ $Y2=0
cc_258 N_A_505_297#_c_211_n N_VGND_c_843_n 0.0110264f $X=3.025 $Y=4.48 $X2=0
+ $Y2=0
cc_259 N_A_505_297#_c_212_n N_VGND_c_843_n 0.00972667f $X=3.455 $Y=4.48 $X2=0
+ $Y2=0
cc_260 N_A_505_297#_c_215_n N_VGND_c_843_n 0.00972667f $X=3.885 $Y=4.48 $X2=0
+ $Y2=0
cc_261 N_A_505_297#_c_217_n N_VGND_c_843_n 0.0103929f $X=4.315 $Y=4.48 $X2=0
+ $Y2=0
cc_262 N_A_505_297#_c_219_n N_VGND_c_845_n 0.00857725f $X=2.675 $Y=0.62 $X2=0
+ $Y2=0
cc_263 N_A_714_47#_c_300_n N_A_M1004_g 0.00265062f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_264 N_A_714_47#_c_300_n N_A_c_397_n 0.00391065f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_265 N_A_714_47#_c_297_n N_A_M1005_g 0.00224176f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_266 N_A_714_47#_c_300_n N_A_M1005_g 0.0169165f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_267 N_A_714_47#_c_297_n N_A_c_400_n 0.0205035f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_268 N_A_714_47#_c_300_n N_A_c_400_n 6.96042e-19 $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_269 N_A_714_47#_c_297_n N_A_M1009_g 0.00205104f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_270 N_A_714_47#_c_299_n N_A_M1009_g 0.0169165f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_271 N_A_714_47#_M1021_g N_A_c_402_n 0.0124308f $X=4.78 $Y=1.955 $X2=0 $Y2=0
cc_272 N_A_714_47#_c_299_n N_A_c_402_n 0.00296321f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_273 N_A_714_47#_c_299_n N_A_M1012_g 0.00146631f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_274 N_A_714_47#_c_298_n N_A_c_405_n 0.0062571f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_275 N_A_714_47#_c_302_n N_A_620_911#_c_476_n 0.0315412f $X=4.705 $Y=2.58
+ $X2=0 $Y2=0
cc_276 N_A_714_47#_c_295_n N_A_620_911#_c_476_n 4.83528e-19 $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_277 N_A_714_47#_c_312_n N_A_620_911#_c_476_n 0.00503951f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_278 N_A_714_47#_c_293_n N_A_620_911#_c_464_n 0.0315412f $X=4.27 $Y=2.58 $X2=0
+ $Y2=0
cc_279 N_A_714_47#_c_294_n N_A_620_911#_c_464_n 0.0158995f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_280 N_A_714_47#_c_301_n N_A_620_911#_c_464_n 9.48385e-19 $X=4.105 $Y=2.49
+ $X2=0 $Y2=0
cc_281 N_A_714_47#_c_295_n N_A_620_911#_c_478_n 0.0093238f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_282 N_A_714_47#_c_295_n N_A_620_911#_M1000_g 0.00318484f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_283 N_A_714_47#_c_312_n N_A_620_911#_M1000_g 0.00383717f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_284 N_A_714_47#_c_295_n N_A_620_911#_c_466_n 0.00293645f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_285 N_A_714_47#_c_296_n N_A_620_911#_c_466_n 0.00664702f $X=3.85 $Y=3.555
+ $X2=0 $Y2=0
cc_286 N_A_714_47#_c_294_n N_A_620_911#_c_522_n 0.0272967f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_287 N_A_714_47#_c_295_n N_A_620_911#_c_522_n 0.0121977f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_288 N_A_714_47#_c_312_n N_A_620_911#_c_522_n 0.014378f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_289 N_A_714_47#_c_295_n N_A_620_911#_c_467_n 0.0257916f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_290 N_A_714_47#_c_312_n N_A_620_911#_c_467_n 0.00429612f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_291 N_A_714_47#_c_295_n N_A_620_911#_c_468_n 0.0127974f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_292 N_A_714_47#_c_293_n N_A_620_911#_c_469_n 0.00516777f $X=4.27 $Y=2.58
+ $X2=0 $Y2=0
cc_293 N_A_714_47#_c_295_n N_A_620_911#_c_469_n 0.00294758f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_294 N_A_714_47#_c_312_n N_A_620_911#_c_469_n 0.0174426f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_295 N_A_714_47#_c_293_n N_A_620_911#_c_470_n 9.46557e-19 $X=4.27 $Y=2.58
+ $X2=0 $Y2=0
cc_296 N_A_714_47#_c_294_n N_A_620_911#_c_470_n 0.0121174f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_297 N_A_714_47#_c_301_n N_A_620_911#_c_470_n 0.0118139f $X=4.105 $Y=2.49
+ $X2=0 $Y2=0
cc_298 N_A_714_47#_c_302_n N_A_620_911#_c_475_n 0.0110028f $X=4.705 $Y=2.58
+ $X2=0 $Y2=0
cc_299 N_A_714_47#_M1021_g N_A_620_911#_c_475_n 0.0043455f $X=4.78 $Y=1.955
+ $X2=0 $Y2=0
cc_300 N_A_714_47#_c_294_n N_A_620_911#_c_475_n 0.00251195f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_301 N_A_714_47#_c_297_n N_A_620_911#_c_475_n 0.0372645f $X=4.105 $Y=2.07
+ $X2=0 $Y2=0
cc_302 N_A_714_47#_c_298_n N_A_620_911#_c_475_n 0.00490309f $X=4.105 $Y=2.07
+ $X2=0 $Y2=0
cc_303 N_A_714_47#_c_299_n N_A_620_911#_c_475_n 0.00567249f $X=4.475 $Y=0.855
+ $X2=0 $Y2=0
cc_304 N_A_714_47#_c_301_n N_A_620_911#_c_475_n 0.00754333f $X=4.105 $Y=2.49
+ $X2=0 $Y2=0
cc_305 N_A_714_47#_c_295_n N_A_620_911#_c_471_n 0.00527878f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_306 N_A_714_47#_M1021_g N_A_1032_911#_c_591_n 0.0177359f $X=4.78 $Y=1.955
+ $X2=0 $Y2=0
cc_307 N_A_714_47#_M1021_g N_VPWR_c_682_n 0.00295399f $X=4.78 $Y=1.955 $X2=0
+ $Y2=0
cc_308 N_A_714_47#_c_312_n N_VPWR_c_700_n 0.0145663f $X=4.555 $Y=3.235 $X2=0
+ $Y2=0
cc_309 N_A_714_47#_c_302_n N_VPWR_c_676_n 0.00492007f $X=4.705 $Y=2.58 $X2=0
+ $Y2=0
cc_310 N_A_714_47#_c_293_n N_VPWR_c_676_n 0.00298594f $X=4.27 $Y=2.58 $X2=0
+ $Y2=0
cc_311 N_A_714_47#_M1021_g N_VPWR_c_676_n 0.00197299f $X=4.78 $Y=1.955 $X2=0
+ $Y2=0
cc_312 N_A_714_47#_c_294_n N_VPWR_c_676_n 0.0294373f $X=3.765 $Y=3.47 $X2=0
+ $Y2=0
cc_313 N_A_714_47#_c_295_n N_VPWR_c_676_n 0.0105024f $X=4.39 $Y=3.555 $X2=0
+ $Y2=0
cc_314 N_A_714_47#_c_297_n N_VPWR_c_676_n 2.07821e-19 $X=4.105 $Y=2.07 $X2=0
+ $Y2=0
cc_315 N_A_714_47#_c_298_n N_VPWR_c_676_n 0.00102999f $X=4.105 $Y=2.07 $X2=0
+ $Y2=0
cc_316 N_A_714_47#_c_312_n N_VPWR_c_676_n 0.0118616f $X=4.555 $Y=3.235 $X2=0
+ $Y2=0
cc_317 N_A_714_47#_c_301_n N_VPWR_c_676_n 0.0186535f $X=4.105 $Y=2.49 $X2=0
+ $Y2=0
cc_318 N_A_714_47#_c_299_n N_X_c_775_n 0.00263398f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_319 N_A_714_47#_c_299_n N_VGND_M1005_s 3.36085e-19 $X=4.475 $Y=0.855 $X2=0
+ $Y2=0
cc_320 N_A_714_47#_c_300_n N_VGND_M1005_s 0.00139685f $X=4.19 $Y=0.855 $X2=0
+ $Y2=0
cc_321 N_A_714_47#_c_300_n N_VGND_c_819_n 0.00702407f $X=4.19 $Y=0.855 $X2=0
+ $Y2=0
cc_322 N_A_714_47#_c_300_n N_VGND_c_821_n 0.0168391f $X=4.19 $Y=0.855 $X2=0
+ $Y2=0
cc_323 N_A_714_47#_c_299_n N_VGND_c_823_n 0.00706177f $X=4.475 $Y=0.855 $X2=0
+ $Y2=0
cc_324 N_A_714_47#_c_383_p N_VGND_c_832_n 0.0121541f $X=3.71 $Y=0.42 $X2=0 $Y2=0
cc_325 N_A_714_47#_c_300_n N_VGND_c_832_n 0.00204475f $X=4.19 $Y=0.855 $X2=0
+ $Y2=0
cc_326 N_A_714_47#_c_299_n N_VGND_c_834_n 0.00202943f $X=4.475 $Y=0.855 $X2=0
+ $Y2=0
cc_327 N_A_714_47#_c_386_p N_VGND_c_834_n 0.0124538f $X=4.57 $Y=0.42 $X2=0 $Y2=0
cc_328 N_A_714_47#_M1004_d N_VGND_c_845_n 0.00397884f $X=3.57 $Y=0.235 $X2=0
+ $Y2=0
cc_329 N_A_714_47#_M1009_d N_VGND_c_845_n 0.00400851f $X=4.43 $Y=0.235 $X2=0
+ $Y2=0
cc_330 N_A_714_47#_c_383_p N_VGND_c_845_n 0.00717399f $X=3.71 $Y=0.42 $X2=0
+ $Y2=0
cc_331 N_A_714_47#_c_299_n N_VGND_c_845_n 0.00389716f $X=4.475 $Y=0.855 $X2=0
+ $Y2=0
cc_332 N_A_714_47#_c_300_n N_VGND_c_845_n 0.00522015f $X=4.19 $Y=0.855 $X2=0
+ $Y2=0
cc_333 N_A_714_47#_c_386_p N_VGND_c_845_n 0.00724021f $X=4.57 $Y=0.42 $X2=0
+ $Y2=0
cc_334 N_A_c_402_n N_A_620_911#_c_475_n 0.0037239f $X=4.71 $Y=1.145 $X2=0 $Y2=0
cc_335 N_A_M1012_g N_A_1032_911#_M1006_g 0.00987876f $X=4.785 $Y=0.56 $X2=0
+ $Y2=0
cc_336 N_A_c_402_n N_A_1032_911#_c_587_n 0.00987876f $X=4.71 $Y=1.145 $X2=0
+ $Y2=0
cc_337 N_A_M1013_g N_VPWR_c_676_n 0.00543198f $X=2.45 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A_c_402_n N_X_c_775_n 7.02896e-19 $X=4.71 $Y=1.145 $X2=0 $Y2=0
cc_339 N_A_c_394_n N_VGND_c_817_n 0.0135915f $X=2.46 $Y=1.01 $X2=0 $Y2=0
cc_340 N_A_c_394_n N_VGND_c_819_n 0.00625119f $X=2.46 $Y=1.01 $X2=0 $Y2=0
cc_341 N_A_M1004_g N_VGND_c_819_n 0.0129916f $X=3.495 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A_c_398_n N_VGND_c_819_n 0.00306309f $X=3.63 $Y=1.145 $X2=0 $Y2=0
cc_343 N_A_M1005_g N_VGND_c_819_n 6.36276e-19 $X=3.925 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A_c_407_n N_VGND_c_819_n 0.0150235f $X=3.125 $Y=1.25 $X2=0 $Y2=0
cc_345 N_A_M1004_g N_VGND_c_821_n 5.31107e-19 $X=3.495 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A_M1005_g N_VGND_c_821_n 0.00741971f $X=3.925 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A_M1009_g N_VGND_c_821_n 0.00741971f $X=4.355 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A_M1012_g N_VGND_c_821_n 5.31107e-19 $X=4.785 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A_M1009_g N_VGND_c_823_n 6.33842e-19 $X=4.355 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A_M1012_g N_VGND_c_823_n 0.0112243f $X=4.785 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A_c_394_n N_VGND_c_828_n 0.00585385f $X=2.46 $Y=1.01 $X2=0 $Y2=0
cc_352 N_A_M1004_g N_VGND_c_832_n 0.00486043f $X=3.495 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A_M1005_g N_VGND_c_832_n 0.00364644f $X=3.925 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A_M1009_g N_VGND_c_834_n 0.00364644f $X=4.355 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A_M1012_g N_VGND_c_834_n 0.00486043f $X=4.785 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_c_394_n N_VGND_c_845_n 0.0134051f $X=2.46 $Y=1.01 $X2=0 $Y2=0
cc_357 N_A_M1004_g N_VGND_c_845_n 0.00822531f $X=3.495 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_M1005_g N_VGND_c_845_n 0.00430798f $X=3.925 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_M1009_g N_VGND_c_845_n 0.00430798f $X=4.355 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_M1012_g N_VGND_c_845_n 0.00822531f $X=4.785 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_620_911#_c_480_n N_A_1032_911#_c_591_n 0.00897291f $X=5.16 $Y=2.94
+ $X2=0 $Y2=0
cc_362 N_A_620_911#_c_480_n N_A_1032_911#_M1008_g 0.00835405f $X=5.16 $Y=2.94
+ $X2=0 $Y2=0
cc_363 N_A_620_911#_c_486_n N_A_1032_911#_c_598_n 0.00835405f $X=5.235 $Y=4.045
+ $X2=0 $Y2=0
cc_364 N_A_620_911#_M1001_g N_A_1032_911#_c_605_n 0.00835405f $X=5.235 $Y=3.485
+ $X2=0 $Y2=0
cc_365 N_A_620_911#_M1001_g N_A_1032_911#_c_607_n 0.00763754f $X=5.235 $Y=3.485
+ $X2=0 $Y2=0
cc_366 N_A_620_911#_M1011_g N_A_1032_911#_c_589_n 0.0254294f $X=5.085 $Y=4.88
+ $X2=0 $Y2=0
cc_367 N_A_620_911#_c_486_n N_A_1032_911#_c_589_n 0.00641748f $X=5.235 $Y=4.045
+ $X2=0 $Y2=0
cc_368 N_A_620_911#_M1011_g N_A_1032_911#_c_590_n 0.00384336f $X=5.085 $Y=4.88
+ $X2=0 $Y2=0
cc_369 N_A_620_911#_c_475_n N_VPWR_c_682_n 0.035645f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_370 N_A_620_911#_c_480_n N_VPWR_c_700_n 0.0189101f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_371 N_A_620_911#_c_481_n N_VPWR_c_700_n 0.00521099f $X=5.01 $Y=4.045 $X2=0
+ $Y2=0
cc_372 N_A_620_911#_c_469_n N_VPWR_c_700_n 0.00509169f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_373 N_A_620_911#_c_469_n N_VPWR_c_703_n 0.00305029f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_374 N_A_620_911#_c_475_n N_VPWR_c_703_n 0.00537241f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_375 N_A_620_911#_c_480_n N_VPWR_c_685_n 0.004734f $X=5.16 $Y=2.94 $X2=0 $Y2=0
cc_376 N_A_620_911#_c_476_n N_VPWR_c_676_n 0.0047221f $X=4.705 $Y=2.94 $X2=0
+ $Y2=0
cc_377 N_A_620_911#_c_464_n N_VPWR_c_676_n 0.00442472f $X=4.27 $Y=2.94 $X2=0
+ $Y2=0
cc_378 N_A_620_911#_c_480_n N_VPWR_c_676_n 0.0132723f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_379 N_A_620_911#_c_484_n N_VPWR_c_676_n 0.00736425f $X=4.78 $Y=2.94 $X2=0
+ $Y2=0
cc_380 N_A_620_911#_c_522_n N_VPWR_c_676_n 0.00566481f $X=4.105 $Y=3.135 $X2=0
+ $Y2=0
cc_381 N_A_620_911#_c_469_n N_VPWR_c_676_n 0.0219288f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_382 N_A_620_911#_c_470_n N_VPWR_c_676_n 0.00663704f $X=4.19 $Y=2.83 $X2=0
+ $Y2=0
cc_383 N_A_620_911#_c_475_n N_VPWR_c_676_n 0.0165665f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_384 N_A_620_911#_c_493_n N_VGND_c_818_n 0.0267051f $X=3.24 $Y=4.735 $X2=0
+ $Y2=0
cc_385 N_A_620_911#_c_493_n N_VGND_c_820_n 0.0266323f $X=3.24 $Y=4.735 $X2=0
+ $Y2=0
cc_386 N_A_620_911#_c_466_n N_VGND_c_820_n 0.0146667f $X=3.935 $Y=4.24 $X2=0
+ $Y2=0
cc_387 N_A_620_911#_c_501_n N_VGND_c_820_n 0.0266323f $X=4.1 $Y=4.735 $X2=0
+ $Y2=0
cc_388 N_A_620_911#_c_478_n N_VGND_c_822_n 0.0183082f $X=4.705 $Y=4.045 $X2=0
+ $Y2=0
cc_389 N_A_620_911#_M1011_g N_VGND_c_822_n 0.00390249f $X=5.085 $Y=4.88 $X2=0
+ $Y2=0
cc_390 N_A_620_911#_c_501_n N_VGND_c_822_n 0.025678f $X=4.1 $Y=4.735 $X2=0 $Y2=0
cc_391 N_A_620_911#_c_493_n N_VGND_c_830_n 0.0189253f $X=3.24 $Y=4.735 $X2=0
+ $Y2=0
cc_392 N_A_620_911#_c_501_n N_VGND_c_841_n 0.0189253f $X=4.1 $Y=4.735 $X2=0
+ $Y2=0
cc_393 N_A_620_911#_M1011_g N_VGND_c_842_n 0.00548296f $X=5.085 $Y=4.88 $X2=0
+ $Y2=0
cc_394 N_A_620_911#_M1003_d N_VGND_c_843_n 0.00223231f $X=3.1 $Y=4.555 $X2=0
+ $Y2=0
cc_395 N_A_620_911#_M1019_d N_VGND_c_843_n 0.00223231f $X=3.96 $Y=4.555 $X2=0
+ $Y2=0
cc_396 N_A_620_911#_M1011_g N_VGND_c_843_n 0.0116568f $X=5.085 $Y=4.88 $X2=0
+ $Y2=0
cc_397 N_A_620_911#_c_493_n N_VGND_c_843_n 0.0122674f $X=3.24 $Y=4.735 $X2=0
+ $Y2=0
cc_398 N_A_620_911#_c_501_n N_VGND_c_843_n 0.0122674f $X=4.1 $Y=4.735 $X2=0
+ $Y2=0
cc_399 N_A_1032_911#_c_591_n N_VPWR_c_682_n 0.00897993f $X=5.255 $Y=1.41 $X2=0
+ $Y2=0
cc_400 N_A_1032_911#_M1008_g N_VPWR_c_700_n 0.00163667f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_401 N_A_1032_911#_c_605_n N_VPWR_c_700_n 8.67432e-19 $X=5.775 $Y=3.065 $X2=0
+ $Y2=0
cc_402 N_A_1032_911#_c_607_n N_VPWR_c_700_n 0.00115994f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_403 N_A_1032_911#_M1008_g N_VPWR_c_683_n 0.00377671f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_404 N_A_1032_911#_M1015_g N_VPWR_c_683_n 0.00372221f $X=6.205 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A_1032_911#_c_585_n N_VPWR_c_683_n 0.00228736f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_406 N_A_1032_911#_M1016_g N_VPWR_c_684_n 0.00741785f $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_407 N_A_1032_911#_c_591_n N_VPWR_c_685_n 0.00545125f $X=5.255 $Y=1.41 $X2=0
+ $Y2=0
cc_408 N_A_1032_911#_M1008_g N_VPWR_c_685_n 0.0154662f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_1032_911#_c_607_n N_VPWR_c_685_n 0.00839873f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_410 N_A_1032_911#_c_599_n N_VPWR_c_705_n 0.00325633f $X=6.13 $Y=3.065 $X2=0
+ $Y2=0
cc_411 N_A_1032_911#_M1015_g N_VPWR_c_686_n 0.0132738f $X=6.205 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A_1032_911#_c_601_n N_VPWR_c_686_n 0.00299145f $X=6.56 $Y=3.065 $X2=0
+ $Y2=0
cc_413 N_A_1032_911#_M1016_g N_VPWR_c_686_n 0.0152247f $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A_1032_911#_c_591_n N_VPWR_c_676_n 0.00412295f $X=5.255 $Y=1.41 $X2=0
+ $Y2=0
cc_415 N_A_1032_911#_M1008_g N_VPWR_c_676_n 0.0135788f $X=5.775 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A_1032_911#_c_599_n N_VPWR_c_676_n 0.00282891f $X=6.13 $Y=3.065 $X2=0
+ $Y2=0
cc_417 N_A_1032_911#_M1015_g N_VPWR_c_676_n 0.0112054f $X=6.205 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_A_1032_911#_c_601_n N_VPWR_c_676_n 0.00282891f $X=6.56 $Y=3.065 $X2=0
+ $Y2=0
cc_419 N_A_1032_911#_M1016_g N_VPWR_c_676_n 0.0141754f $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A_1032_911#_c_607_n N_VPWR_c_676_n 0.00687951f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_421 N_A_1032_911#_M1007_g N_X_c_783_n 0.00498668f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_422 N_A_1032_911#_c_582_n N_X_c_784_n 0.00792257f $X=5.7 $Y=1.247 $X2=0 $Y2=0
cc_423 N_A_1032_911#_c_585_n N_X_c_784_n 0.0552661f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_424 N_A_1032_911#_M1016_g N_X_c_777_n 7.94882e-19 $X=6.635 $Y=1.985 $X2=0
+ $Y2=0
cc_425 N_A_1032_911#_M1017_g N_X_c_774_n 0.00496787f $X=6.205 $Y=0.56 $X2=0
+ $Y2=0
cc_426 N_A_1032_911#_M1018_g N_X_c_774_n 0.00458369f $X=6.635 $Y=0.56 $X2=0
+ $Y2=0
cc_427 N_A_1032_911#_c_585_n N_X_c_789_n 0.0308881f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_428 N_A_1032_911#_M1006_g N_X_c_775_n 0.00446469f $X=5.255 $Y=0.56 $X2=0
+ $Y2=0
cc_429 N_A_1032_911#_c_582_n N_X_c_775_n 0.0290305f $X=5.7 $Y=1.247 $X2=0 $Y2=0
cc_430 N_A_1032_911#_M1007_g N_X_c_775_n 0.00667268f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_431 N_A_1032_911#_c_591_n X 0.00308224f $X=5.255 $Y=1.41 $X2=0 $Y2=0
cc_432 N_A_1032_911#_M1008_g X 0.0103699f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_433 N_A_1032_911#_c_589_n N_VGND_c_822_n 0.0259447f $X=5.45 $Y=4.24 $X2=0
+ $Y2=0
cc_434 N_A_1032_911#_M1006_g N_VGND_c_823_n 0.00189452f $X=5.255 $Y=0.56 $X2=0
+ $Y2=0
cc_435 N_A_1032_911#_M1006_g N_VGND_c_824_n 5.88421e-19 $X=5.255 $Y=0.56 $X2=0
+ $Y2=0
cc_436 N_A_1032_911#_M1007_g N_VGND_c_824_n 0.0110235f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_437 N_A_1032_911#_M1017_g N_VGND_c_824_n 0.010662f $X=6.205 $Y=0.56 $X2=0
+ $Y2=0
cc_438 N_A_1032_911#_c_585_n N_VGND_c_824_n 0.00223674f $X=6.635 $Y=1.085 $X2=0
+ $Y2=0
cc_439 N_A_1032_911#_M1018_g N_VGND_c_824_n 6.48459e-19 $X=6.635 $Y=0.56 $X2=0
+ $Y2=0
cc_440 N_A_1032_911#_M1018_g N_VGND_c_825_n 0.00407687f $X=6.635 $Y=0.56 $X2=0
+ $Y2=0
cc_441 N_A_1032_911#_M1006_g N_VGND_c_836_n 0.00585385f $X=5.255 $Y=0.56 $X2=0
+ $Y2=0
cc_442 N_A_1032_911#_M1007_g N_VGND_c_836_n 0.00486043f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_443 N_A_1032_911#_M1017_g N_VGND_c_838_n 0.00486043f $X=6.205 $Y=0.56 $X2=0
+ $Y2=0
cc_444 N_A_1032_911#_M1018_g N_VGND_c_838_n 0.00585385f $X=6.635 $Y=0.56 $X2=0
+ $Y2=0
cc_445 N_A_1032_911#_c_589_n N_VGND_c_842_n 0.0239189f $X=5.45 $Y=4.24 $X2=0
+ $Y2=0
cc_446 N_A_1032_911#_M1011_d N_VGND_c_843_n 0.00214546f $X=5.16 $Y=4.555 $X2=0
+ $Y2=0
cc_447 N_A_1032_911#_c_589_n N_VGND_c_843_n 0.0195213f $X=5.45 $Y=4.24 $X2=0
+ $Y2=0
cc_448 N_A_1032_911#_M1006_g N_VGND_c_845_n 0.010837f $X=5.255 $Y=0.56 $X2=0
+ $Y2=0
cc_449 N_A_1032_911#_M1007_g N_VGND_c_845_n 0.00852643f $X=5.775 $Y=0.56 $X2=0
+ $Y2=0
cc_450 N_A_1032_911#_M1017_g N_VGND_c_845_n 0.00822531f $X=6.205 $Y=0.56 $X2=0
+ $Y2=0
cc_451 N_A_1032_911#_M1018_g N_VGND_c_845_n 0.011676f $X=6.635 $Y=0.56 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_676_n N_X_M1002_d 0.00216609f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_453 N_VPWR_c_676_n N_X_M1015_d 0.00133453f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_c_683_n N_X_c_784_n 0.0121443f $X=5.99 $Y=1.79 $X2=0 $Y2=0
cc_455 N_VPWR_c_683_n N_X_c_777_n 0.0273305f $X=5.99 $Y=1.79 $X2=0 $Y2=0
cc_456 N_VPWR_c_684_n N_X_c_777_n 0.00424153f $X=6.85 $Y=1.79 $X2=0 $Y2=0
cc_457 N_VPWR_c_686_n N_X_c_777_n 0.00966848f $X=6.755 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_676_n N_X_c_777_n 0.00302523f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_459 N_VPWR_c_682_n X 0.0230063f $X=5.005 $Y=1.79 $X2=0 $Y2=0
cc_460 N_VPWR_c_683_n X 0.021786f $X=5.99 $Y=1.79 $X2=0 $Y2=0
cc_461 N_VPWR_c_685_n X 0.0113333f $X=5.905 $Y=2.72 $X2=0 $Y2=0
cc_462 N_VPWR_c_676_n X 0.00302523f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_463 N_X_c_775_n N_VGND_c_823_n 0.001162f $X=5.497 $Y=1.41 $X2=0 $Y2=0
cc_464 N_X_c_783_n N_VGND_c_824_n 0.0406307f $X=5.47 $Y=0.42 $X2=0 $Y2=0
cc_465 N_X_c_784_n N_VGND_c_824_n 0.0165907f $X=6.28 $Y=1.247 $X2=0 $Y2=0
cc_466 N_X_c_775_n N_VGND_c_824_n 0.00106574f $X=5.497 $Y=1.41 $X2=0 $Y2=0
cc_467 N_X_c_774_n N_VGND_c_825_n 0.00274856f $X=6.42 $Y=0.42 $X2=0 $Y2=0
cc_468 N_X_c_783_n N_VGND_c_836_n 0.0191787f $X=5.47 $Y=0.42 $X2=0 $Y2=0
cc_469 N_X_c_774_n N_VGND_c_838_n 0.0135183f $X=6.42 $Y=0.42 $X2=0 $Y2=0
cc_470 N_X_M1006_d N_VGND_c_845_n 0.00542784f $X=5.33 $Y=0.235 $X2=0 $Y2=0
cc_471 N_X_M1017_d N_VGND_c_845_n 0.00431525f $X=6.28 $Y=0.235 $X2=0 $Y2=0
cc_472 N_X_c_783_n N_VGND_c_845_n 0.0114765f $X=5.47 $Y=0.42 $X2=0 $Y2=0
cc_473 N_X_c_774_n N_VGND_c_845_n 0.00839034f $X=6.42 $Y=0.42 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a41o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.075000 4.065000 1.295000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.075000 4.975000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.155000 1.075000 6.185000 1.295000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.495000 1.075000 7.505000 1.295000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135000 1.075000 3.145000 1.280000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.635000 1.605000 0.805000 ;
        RECT 0.150000 0.805000 0.320000 1.575000 ;
        RECT 0.150000 1.575000 1.605000 1.745000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 1.745000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.435000 1.745000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.465000 ;
        RECT 0.935000  0.085000 1.265000 0.465000 ;
        RECT 1.775000  0.085000 2.125000 0.465000 ;
        RECT 2.635000  0.085000 2.965000 0.465000 ;
        RECT 6.615000  0.085000 6.945000 0.465000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.095000 1.915000 0.425000 2.635000 ;
        RECT 0.935000 1.915000 1.265000 2.635000 ;
        RECT 1.775000 1.915000 2.125000 2.635000 ;
        RECT 3.575000 1.915000 3.905000 2.635000 ;
        RECT 4.415000 1.915000 4.745000 2.635000 ;
        RECT 5.345000 1.915000 6.035000 2.635000 ;
        RECT 6.615000 1.915000 6.945000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.490000 1.075000 1.945000 1.245000 ;
      RECT 1.775000 0.645000 3.905000 0.815000 ;
      RECT 1.775000 0.815000 1.945000 1.075000 ;
      RECT 1.775000 1.245000 1.945000 1.455000 ;
      RECT 1.775000 1.455000 2.965000 1.625000 ;
      RECT 2.295000 0.255000 2.465000 0.645000 ;
      RECT 2.375000 1.795000 2.545000 2.295000 ;
      RECT 2.375000 2.295000 3.405000 2.465000 ;
      RECT 2.715000 1.955000 3.045000 2.125000 ;
      RECT 2.795000 1.625000 2.965000 1.955000 ;
      RECT 3.155000 0.295000 4.245000 0.465000 ;
      RECT 3.235000 1.535000 7.370000 1.705000 ;
      RECT 3.235000 1.705000 3.405000 2.295000 ;
      RECT 4.075000 0.465000 4.245000 0.645000 ;
      RECT 4.075000 0.645000 5.165000 0.815000 ;
      RECT 4.075000 1.705000 4.245000 2.465000 ;
      RECT 4.415000 0.295000 6.105000 0.465000 ;
      RECT 4.935000 1.705000 5.105000 2.465000 ;
      RECT 5.355000 0.645000 7.285000 0.815000 ;
      RECT 6.275000 1.705000 6.445000 2.465000 ;
      RECT 7.115000 0.255000 7.285000 0.645000 ;
      RECT 7.115000 1.705000 7.285000 2.465000 ;
  END
END sky130_fd_sc_hd__a41o_4

* NGSPICE file created from sky130_fd_sc_hd__xor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
M1000 a_496_49# a_358_93# a_120_21# VPB phighvt w=840000u l=150000u
+  ad=7.326e+11p pd=5.14e+06u as=3.192e+11p ps=2.44e+06u
M1001 a_919_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.653e+11p pd=1.82e+06u as=8.2505e+11p ps=7.78e+06u
M1002 a_919_297# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.526e+11p pd=2.52e+06u as=1.213e+12p ps=1.048e+07u
M1003 VPWR a_120_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1004 a_1290_49# a_919_297# a_496_49# VNB nshort w=420000u l=150000u
+  ad=5.517e+11p pd=4.37e+06u as=5.401e+11p ps=4.32e+06u
M1005 a_120_21# C a_496_49# VNB nshort w=640000u l=150000u
+  ad=2.56e+11p pd=2.08e+06u as=0p ps=0u
M1006 X a_120_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_358_93# C VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1008 a_496_49# B a_1023_365# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.828e+11p ps=3.78e+06u
M1009 a_120_21# C a_478_325# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=7.592e+11p ps=5.22e+06u
M1010 X a_120_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1011 a_1023_365# a_919_297# a_496_49# VPB phighvt w=840000u l=150000u
+  ad=6.966e+11p pd=5.24e+06u as=0p ps=0u
M1012 a_1290_49# a_1023_365# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=7.57e+11p pd=5.58e+06u as=0p ps=0u
M1013 a_478_325# B a_1290_49# VNB nshort w=640000u l=150000u
+  ad=5.9845e+11p pd=4.47e+06u as=0p ps=0u
M1014 a_496_49# B a_1290_49# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_120_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1290_49# a_919_297# a_478_325# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A a_1023_365# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_478_325# B a_1023_365# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_358_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=0p ps=0u
M1020 a_1290_49# a_1023_365# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_478_325# a_358_93# a_120_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A a_1023_365# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1023_365# a_919_297# a_478_325# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


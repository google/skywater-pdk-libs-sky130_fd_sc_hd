* File: sky130_fd_sc_hd__or2_0.spice
* Created: Thu Aug 27 14:42:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or2_0.spice.pex"
.subckt sky130_fd_sc_hd__or2_0  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_A_68_355#_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_68_355#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0567 PD=0.755 PS=0.69 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_68_355#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.07035 PD=1.36 PS=0.755 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_150_355# N_B_M1005_g N_A_68_355#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_150_355# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0784132 AS=0.0441 PD=0.772642 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8
+ SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_68_355#_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2176 AS=0.119487 PD=1.96 PS=1.17736 NRD=23.0687 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_159 A_150_355# 0 1.0136e-19 $X=0.75 $Y=1.775
*
.include "sky130_fd_sc_hd__or2_0.spice.SKY130_FD_SC_HD__OR2_0.pxi"
*
.ends
*
*

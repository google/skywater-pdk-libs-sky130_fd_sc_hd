* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_8.pex.spice
* Created: Tue Sep  1 19:11:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%A 1 3 4 6 7 9 12 14 16 19 21 23
+ 26 28 30 33 35 37 40 42 44 47 49 51 54 56 58 61 63 65 66 68 69 70 71 72 73 74
+ 75 76 77 112 113
r199 111 113 36.7542 $w=5.75e-07 $l=3.95e-07 $layer=POLY_cond $X=4.7 $Y=1.097
+ $X2=5.095 $Y2=1.097
r200 111 112 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=4.7
+ $Y=1.16 $X2=4.7 $Y2=1.16
r201 109 111 2.32622 $w=5.75e-07 $l=2.5e-08 $layer=POLY_cond $X=4.675 $Y=1.097
+ $X2=4.7 $Y2=1.097
r202 92 93 39.5457 $w=5.75e-07 $l=4.25e-07 $layer=POLY_cond $X=0.89 $Y=1.097
+ $X2=1.315 $Y2=1.097
r203 90 92 25.1231 $w=5.75e-07 $l=2.7e-07 $layer=POLY_cond $X=0.62 $Y=1.097
+ $X2=0.89 $Y2=1.097
r204 87 90 13.9573 $w=5.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.47 $Y=1.097
+ $X2=0.62 $Y2=1.097
r205 77 112 14.688 $w=2.53e-07 $l=3.25e-07 $layer=LI1_cond $X=4.375 $Y=1.162
+ $X2=4.7 $Y2=1.162
r206 76 77 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=3.915 $Y=1.162
+ $X2=4.375 $Y2=1.162
r207 75 76 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=3.455 $Y=1.162
+ $X2=3.915 $Y2=1.162
r208 74 75 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=2.995 $Y=1.162
+ $X2=3.455 $Y2=1.162
r209 73 74 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.162
+ $X2=2.995 $Y2=1.162
r210 72 73 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=2.075 $Y=1.162
+ $X2=2.535 $Y2=1.162
r211 71 72 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=1.615 $Y=1.162
+ $X2=2.075 $Y2=1.162
r212 70 71 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.162
+ $X2=1.615 $Y2=1.162
r213 69 70 24.1787 $w=2.53e-07 $l=5.35e-07 $layer=LI1_cond $X=0.62 $Y=1.162
+ $X2=1.155 $Y2=1.162
r214 69 90 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r215 66 113 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=5.095 $Y=1.385
+ $X2=5.095 $Y2=1.097
r216 66 68 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.095 $Y=1.385
+ $X2=5.095 $Y2=1.985
r217 63 109 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=4.675 $Y=1.385
+ $X2=4.675 $Y2=1.097
r218 63 65 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.675 $Y=1.385
+ $X2=4.675 $Y2=1.985
r219 59 109 23.2622 $w=5.75e-07 $l=2.5e-07 $layer=POLY_cond $X=4.425 $Y=1.097
+ $X2=4.675 $Y2=1.097
r220 59 107 15.8183 $w=5.75e-07 $l=1.7e-07 $layer=POLY_cond $X=4.425 $Y=1.097
+ $X2=4.255 $Y2=1.097
r221 59 61 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=4.425 $Y=0.81
+ $X2=4.425 $Y2=0.445
r222 56 107 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=4.255 $Y=1.385
+ $X2=4.255 $Y2=1.097
r223 56 58 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.255 $Y=1.385
+ $X2=4.255 $Y2=1.985
r224 52 107 24.1926 $w=5.75e-07 $l=2.6e-07 $layer=POLY_cond $X=3.995 $Y=1.097
+ $X2=4.255 $Y2=1.097
r225 52 105 14.8878 $w=5.75e-07 $l=1.6e-07 $layer=POLY_cond $X=3.995 $Y=1.097
+ $X2=3.835 $Y2=1.097
r226 52 54 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.995 $Y=0.81
+ $X2=3.995 $Y2=0.445
r227 49 105 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=3.835 $Y=1.385
+ $X2=3.835 $Y2=1.097
r228 49 51 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.835 $Y=1.385
+ $X2=3.835 $Y2=1.985
r229 45 105 25.1231 $w=5.75e-07 $l=2.7e-07 $layer=POLY_cond $X=3.565 $Y=1.097
+ $X2=3.835 $Y2=1.097
r230 45 103 13.9573 $w=5.75e-07 $l=1.5e-07 $layer=POLY_cond $X=3.565 $Y=1.097
+ $X2=3.415 $Y2=1.097
r231 45 47 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.565 $Y=0.81
+ $X2=3.565 $Y2=0.445
r232 42 103 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=3.415 $Y=1.385
+ $X2=3.415 $Y2=1.097
r233 42 44 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.415 $Y=1.385
+ $X2=3.415 $Y2=1.985
r234 38 103 26.0536 $w=5.75e-07 $l=2.8e-07 $layer=POLY_cond $X=3.135 $Y=1.097
+ $X2=3.415 $Y2=1.097
r235 38 101 13.0268 $w=5.75e-07 $l=1.4e-07 $layer=POLY_cond $X=3.135 $Y=1.097
+ $X2=2.995 $Y2=1.097
r236 38 40 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.135 $Y=0.81
+ $X2=3.135 $Y2=0.445
r237 35 101 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.995 $Y=1.385
+ $X2=2.995 $Y2=1.097
r238 35 37 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.995 $Y=1.385
+ $X2=2.995 $Y2=1.985
r239 31 101 26.9841 $w=5.75e-07 $l=2.9e-07 $layer=POLY_cond $X=2.705 $Y=1.097
+ $X2=2.995 $Y2=1.097
r240 31 99 12.0963 $w=5.75e-07 $l=1.3e-07 $layer=POLY_cond $X=2.705 $Y=1.097
+ $X2=2.575 $Y2=1.097
r241 31 33 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.705 $Y=0.81
+ $X2=2.705 $Y2=0.445
r242 28 99 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.575 $Y=1.385
+ $X2=2.575 $Y2=1.097
r243 28 30 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.575 $Y=1.385
+ $X2=2.575 $Y2=1.985
r244 24 99 27.9146 $w=5.75e-07 $l=3e-07 $layer=POLY_cond $X=2.275 $Y=1.097
+ $X2=2.575 $Y2=1.097
r245 24 97 11.1658 $w=5.75e-07 $l=1.2e-07 $layer=POLY_cond $X=2.275 $Y=1.097
+ $X2=2.155 $Y2=1.097
r246 24 26 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.275 $Y=0.81
+ $X2=2.275 $Y2=0.445
r247 21 97 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.155 $Y=1.385
+ $X2=2.155 $Y2=1.097
r248 21 23 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.155 $Y=1.385
+ $X2=2.155 $Y2=1.985
r249 17 97 28.8451 $w=5.75e-07 $l=3.1e-07 $layer=POLY_cond $X=1.845 $Y=1.097
+ $X2=2.155 $Y2=1.097
r250 17 95 10.2353 $w=5.75e-07 $l=1.1e-07 $layer=POLY_cond $X=1.845 $Y=1.097
+ $X2=1.735 $Y2=1.097
r251 17 19 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.845 $Y=0.81
+ $X2=1.845 $Y2=0.445
r252 14 95 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.097
r253 14 16 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.985
r254 10 95 29.7756 $w=5.75e-07 $l=3.2e-07 $layer=POLY_cond $X=1.415 $Y=1.097
+ $X2=1.735 $Y2=1.097
r255 10 93 9.30486 $w=5.75e-07 $l=1e-07 $layer=POLY_cond $X=1.415 $Y=1.097
+ $X2=1.315 $Y2=1.097
r256 10 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.415 $Y=0.81
+ $X2=1.415 $Y2=0.445
r257 7 93 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=1.315 $Y=1.385
+ $X2=1.315 $Y2=1.097
r258 7 9 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.315 $Y=1.385 $X2=1.315
+ $Y2=1.985
r259 4 92 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=0.89 $Y=1.385
+ $X2=0.89 $Y2=1.097
r260 4 6 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.89 $Y=1.385 $X2=0.89
+ $Y2=1.985
r261 1 87 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=0.47 $Y=1.385
+ $X2=0.47 $Y2=1.097
r262 1 3 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.47 $Y=1.385 $X2=0.47
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%KAPWR 1 2 3 4 5 6 7 38 39 43 44
+ 48 49 53 54 58 59 61 63 65 69 76 81 86 91 96 101
c141 63 0 1.04828e-19 $X=5.195 $Y=2.21
r142 69 72 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=1.965
+ $X2=0.26 $Y2=2.21
r143 65 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.215 $Y=2.21
+ $X2=0.215 $Y2=2.21
r144 62 101 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=5.305 $Y=2.21
+ $X2=5.305 $Y2=1.965
r145 61 63 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=5.34 $Y=2.21
+ $X2=5.195 $Y2=2.21
r146 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.34 $Y=2.21
+ $X2=5.34 $Y2=2.21
r147 59 63 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=4.585 $Y=2.24
+ $X2=5.195 $Y2=2.24
r148 57 96 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=4.465 $Y=2.21
+ $X2=4.465 $Y2=1.965
r149 56 59 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.44 $Y=2.21
+ $X2=4.585 $Y2=2.21
r150 56 58 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.44 $Y=2.21
+ $X2=4.295 $Y2=2.21
r151 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.44 $Y=2.21
+ $X2=4.44 $Y2=2.21
r152 54 58 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=3.725 $Y=2.24
+ $X2=4.295 $Y2=2.24
r153 52 91 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.625 $Y=2.21
+ $X2=3.625 $Y2=1.965
r154 51 54 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.58 $Y=2.21
+ $X2=3.725 $Y2=2.21
r155 51 53 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.58 $Y=2.21
+ $X2=3.435 $Y2=2.21
r156 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.21
+ $X2=3.58 $Y2=2.21
r157 49 53 0.333882 $w=2e-07 $l=4.35e-07 $layer=MET1_cond $X=3 $Y=2.24 $X2=3.435
+ $Y2=2.24
r158 47 86 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.785 $Y=2.21
+ $X2=2.785 $Y2=1.965
r159 46 49 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.855 $Y=2.21
+ $X2=3 $Y2=2.21
r160 46 48 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.855 $Y=2.21
+ $X2=2.71 $Y2=2.21
r161 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.855 $Y=2.21
+ $X2=2.855 $Y2=2.21
r162 44 48 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=2.12 $Y=2.24
+ $X2=2.71 $Y2=2.24
r163 42 81 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.945 $Y=2.21
+ $X2=1.945 $Y2=1.965
r164 41 44 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=2.12 $Y2=2.21
r165 41 43 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=1.83 $Y2=2.21
r166 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.975 $Y=2.21
+ $X2=1.975 $Y2=2.21
r167 39 43 0.468202 $w=2e-07 $l=6.1e-07 $layer=MET1_cond $X=1.22 $Y=2.24
+ $X2=1.83 $Y2=2.24
r168 38 65 0.234171 $w=3.7e-07 $l=5.7e-07 $layer=MET1_cond $X=0.93 $Y=2.24
+ $X2=0.36 $Y2=2.24
r169 37 76 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.105 $Y=2.21
+ $X2=1.105 $Y2=1.965
r170 36 39 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.075 $Y=2.21
+ $X2=1.22 $Y2=2.21
r171 36 38 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.075 $Y=2.21
+ $X2=0.93 $Y2=2.21
r172 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.075 $Y=2.21
+ $X2=1.075 $Y2=2.21
r173 7 101 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=5.17
+ $Y=1.485 $X2=5.305 $Y2=1.965
r174 6 96 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=4.33
+ $Y=1.485 $X2=4.465 $Y2=1.965
r175 5 91 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=1.485 $X2=3.625 $Y2=1.965
r176 4 86 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=2.65
+ $Y=1.485 $X2=2.785 $Y2=1.965
r177 3 81 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=1.485 $X2=1.945 $Y2=1.965
r178 2 76 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.105 $Y2=1.965
r179 1 69 300 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%Y 1 2 3 4 5 6 7 8 9 10 32 33 34
+ 35 36 39 41 45 49 51 53 57 61 63 65 69 73 75 77 81 85 87 89 93 95 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 115 116
c244 116 0 1.04828e-19 $X=5.305 $Y=1.46
r245 109 116 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.305 $Y=1.545
+ $X2=5.305 $Y2=1.46
r246 109 116 0.341465 $w=2.68e-07 $l=8e-09 $layer=LI1_cond $X=5.305 $Y=1.452
+ $X2=5.305 $Y2=1.46
r247 108 109 11.183 $w=2.68e-07 $l=2.62e-07 $layer=LI1_cond $X=5.305 $Y=1.19
+ $X2=5.305 $Y2=1.452
r248 107 115 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.305 $Y=0.78
+ $X2=5.305 $Y2=0.865
r249 107 108 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.305 $Y=0.9
+ $X2=5.305 $Y2=1.19
r250 107 115 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.305 $Y=0.9
+ $X2=5.305 $Y2=0.865
r251 96 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=1.545
+ $X2=4.885 $Y2=1.545
r252 95 109 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.17 $Y=1.545
+ $X2=5.305 $Y2=1.545
r253 95 96 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.17 $Y=1.545
+ $X2=4.97 $Y2=1.545
r254 91 106 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=1.63
+ $X2=4.885 $Y2=1.545
r255 91 93 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.885 $Y=1.63
+ $X2=4.885 $Y2=1.83
r256 90 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.305 $Y=0.78
+ $X2=4.21 $Y2=0.78
r257 89 107 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.17 $Y=0.78
+ $X2=5.305 $Y2=0.78
r258 89 90 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.17 $Y=0.78
+ $X2=4.305 $Y2=0.78
r259 88 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=1.545
+ $X2=4.045 $Y2=1.545
r260 87 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=1.545
+ $X2=4.885 $Y2=1.545
r261 87 88 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.8 $Y=1.545
+ $X2=4.13 $Y2=1.545
r262 83 105 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=0.695
+ $X2=4.21 $Y2=0.78
r263 83 85 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=4.21 $Y=0.695
+ $X2=4.21 $Y2=0.445
r264 79 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=1.63
+ $X2=4.045 $Y2=1.545
r265 79 81 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.045 $Y=1.63
+ $X2=4.045 $Y2=1.83
r266 78 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.445 $Y=0.78
+ $X2=3.35 $Y2=0.78
r267 77 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.115 $Y=0.78
+ $X2=4.21 $Y2=0.78
r268 77 78 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.115 $Y=0.78
+ $X2=3.445 $Y2=0.78
r269 76 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=1.545
+ $X2=3.205 $Y2=1.545
r270 75 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=1.545
+ $X2=4.045 $Y2=1.545
r271 75 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.96 $Y=1.545
+ $X2=3.29 $Y2=1.545
r272 71 103 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.695
+ $X2=3.35 $Y2=0.78
r273 71 73 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.35 $Y=0.695
+ $X2=3.35 $Y2=0.445
r274 67 102 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=1.63
+ $X2=3.205 $Y2=1.545
r275 67 69 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.205 $Y=1.63
+ $X2=3.205 $Y2=1.83
r276 66 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.585 $Y=0.78
+ $X2=2.49 $Y2=0.78
r277 65 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.255 $Y=0.78
+ $X2=3.35 $Y2=0.78
r278 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.255 $Y=0.78
+ $X2=2.585 $Y2=0.78
r279 64 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=1.545
+ $X2=2.365 $Y2=1.545
r280 63 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=1.545
+ $X2=3.205 $Y2=1.545
r281 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.12 $Y=1.545
+ $X2=2.45 $Y2=1.545
r282 59 101 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.695
+ $X2=2.49 $Y2=0.78
r283 59 61 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=2.49 $Y=0.695
+ $X2=2.49 $Y2=0.445
r284 55 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=1.63
+ $X2=2.365 $Y2=1.545
r285 55 57 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.365 $Y=1.63
+ $X2=2.365 $Y2=1.83
r286 54 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=0.78
+ $X2=1.63 $Y2=0.78
r287 53 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.395 $Y=0.78
+ $X2=2.49 $Y2=0.78
r288 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.395 $Y=0.78
+ $X2=1.725 $Y2=0.78
r289 52 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.545
+ $X2=1.525 $Y2=1.545
r290 51 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=1.545
+ $X2=2.365 $Y2=1.545
r291 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.28 $Y=1.545
+ $X2=1.61 $Y2=1.545
r292 47 99 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.695
+ $X2=1.63 $Y2=0.78
r293 47 49 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.63 $Y=0.695
+ $X2=1.63 $Y2=0.445
r294 43 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=1.63
+ $X2=1.525 $Y2=1.545
r295 43 45 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.525 $Y=1.63
+ $X2=1.525 $Y2=1.83
r296 42 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.545
+ $X2=0.68 $Y2=1.545
r297 41 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=1.545
+ $X2=1.525 $Y2=1.545
r298 41 42 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.44 $Y=1.545
+ $X2=0.765 $Y2=1.545
r299 37 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.63
+ $X2=0.68 $Y2=1.545
r300 37 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.68 $Y=1.63 $X2=0.68
+ $Y2=1.93
r301 35 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=1.545
+ $X2=0.68 $Y2=1.545
r302 35 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.595 $Y=1.545
+ $X2=0.285 $Y2=1.545
r303 33 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.535 $Y=0.78
+ $X2=1.63 $Y2=0.78
r304 33 34 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.535 $Y=0.78
+ $X2=0.285 $Y2=0.78
r305 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.46
+ $X2=0.285 $Y2=1.545
r306 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.285 $Y2=0.78
r307 31 32 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.2 $Y2=1.46
r308 10 93 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=4.75
+ $Y=1.485 $X2=4.885 $Y2=1.83
r309 9 81 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=3.91
+ $Y=1.485 $X2=4.045 $Y2=1.83
r310 8 69 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=3.07
+ $Y=1.485 $X2=3.205 $Y2=1.83
r311 7 57 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=2.23
+ $Y=1.485 $X2=2.365 $Y2=1.83
r312 6 45 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=1.39
+ $Y=1.485 $X2=1.525 $Y2=1.83
r313 5 39 300 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.93
r314 4 85 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.235 $X2=4.21 $Y2=0.445
r315 3 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.235 $X2=3.35 $Y2=0.445
r316 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.49 $Y2=0.445
r317 1 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.235 $X2=1.63 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%VGND 1 2 3 4 5 18 22 26 30 34
+ 37 38 40 41 42 44 49 54 70 71 74 77 80 83
r90 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r91 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r93 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r94 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r95 67 70 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r96 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r97 65 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r98 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r99 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r100 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r101 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r102 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.92
+ $Y2=0
r103 59 61 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=3.45 $Y2=0
r104 58 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r105 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r106 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r107 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.06
+ $Y2=0
r108 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.53 $Y2=0
r109 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.92
+ $Y2=0
r110 54 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=2.53 $Y2=0
r111 53 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r112 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r113 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r114 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r115 50 52 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r116 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.06
+ $Y2=0
r117 49 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.61 $Y2=0
r118 47 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r119 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r120 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r121 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r122 42 47 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r123 42 83 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r124 40 64 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r125 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r126 39 67 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.83
+ $Y2=0
r127 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r128 37 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=3.45 $Y2=0
r129 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.78
+ $Y2=0
r130 36 64 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.945 $Y=0
+ $X2=4.37 $Y2=0
r131 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.78
+ $Y2=0
r132 32 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r133 32 34 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.39
r134 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0
r135 28 30 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0.39
r136 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r137 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.39
r138 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0
r139 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0.39
r140 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r141 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r142 5 34 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.5
+ $Y=0.235 $X2=4.64 $Y2=0.39
r143 4 30 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.78 $Y2=0.39
r144 3 26 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.235 $X2=2.92 $Y2=0.39
r145 2 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.235 $X2=2.06 $Y2=0.39
r146 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%VPWR 1 8 9
r80 8 9 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r81 4 8 360.128 $w=1.68e-07 $l=5.52e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=5.75
+ $Y2=2.72
r82 1 9 1.57067 $w=4.8e-07 $l=5.52e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=5.75
+ $Y2=2.72
r83 1 4 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


* File: sky130_fd_sc_hd__lpflow_bleeder_1.spice
* Created: Thu Aug 27 14:23:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_bleeder_1.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_bleeder_1  VNB VPB SHORT VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* SHORT	SHORT
* VPB	VPB
* VNB	VNB
MM1000 A_147_105# N_SHORT_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.36
+ AD=0.0378 AS=0.0936 PD=0.57 PS=1.24 NRD=16.656 NRS=0 M=1 R=2.4 SA=75000.2
+ SB=75001.6 A=0.054 P=1.02 MULT=1
MM1004 A_219_105# N_SHORT_M1004_g A_147_105# VNB NSHORT L=0.15 W=0.36 AD=0.0378
+ AS=0.0378 PD=0.57 PS=0.57 NRD=16.656 NRS=16.656 M=1 R=2.4 SA=75000.5
+ SB=75001.3 A=0.054 P=1.02 MULT=1
MM1001 A_291_105# N_SHORT_M1001_g A_219_105# VNB NSHORT L=0.15 W=0.36 AD=0.0378
+ AS=0.0378 PD=0.57 PS=0.57 NRD=16.656 NRS=16.656 M=1 R=2.4 SA=75000.9
+ SB=75000.9 A=0.054 P=1.02 MULT=1
MM1003 A_363_105# N_SHORT_M1003_g A_291_105# VNB NSHORT L=0.15 W=0.36 AD=0.0378
+ AS=0.0378 PD=0.57 PS=0.57 NRD=16.656 NRS=16.656 M=1 R=2.4 SA=75001.3
+ SB=75000.5 A=0.054 P=1.02 MULT=1
MM1002 N_VPWR_M1002_d N_SHORT_M1002_g A_363_105# VNB NSHORT L=0.15 W=0.36
+ AD=0.0936 AS=0.0378 PD=1.24 PS=0.57 NRD=0 NRS=16.656 M=1 R=2.4 SA=75001.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
DX5_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__lpflow_bleeder_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__and2_4.spice.SKY130_FD_SC_HD__AND2_4.pxi
* Created: Thu Aug 27 14:07:05 2020
* 
x_PM_SKY130_FD_SC_HD__AND2_4%A N_A_M1005_g N_A_M1006_g A N_A_c_57_n N_A_c_58_n
+ N_A_c_59_n PM_SKY130_FD_SC_HD__AND2_4%A
x_PM_SKY130_FD_SC_HD__AND2_4%B N_B_M1000_g N_B_M1010_g B N_B_c_84_n N_B_c_85_n
+ N_B_c_86_n PM_SKY130_FD_SC_HD__AND2_4%B
x_PM_SKY130_FD_SC_HD__AND2_4%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1006_d
+ N_A_27_47#_c_122_n N_A_27_47#_M1002_g N_A_27_47#_M1001_g N_A_27_47#_c_123_n
+ N_A_27_47#_M1003_g N_A_27_47#_M1004_g N_A_27_47#_c_124_n N_A_27_47#_M1007_g
+ N_A_27_47#_M1009_g N_A_27_47#_c_125_n N_A_27_47#_M1008_g N_A_27_47#_M1011_g
+ N_A_27_47#_c_126_n N_A_27_47#_c_140_n N_A_27_47#_c_127_n N_A_27_47#_c_173_p
+ N_A_27_47#_c_151_n N_A_27_47#_c_153_n N_A_27_47#_c_128_n N_A_27_47#_c_135_n
+ N_A_27_47#_c_136_n N_A_27_47#_c_129_n N_A_27_47#_c_130_n
+ PM_SKY130_FD_SC_HD__AND2_4%A_27_47#
x_PM_SKY130_FD_SC_HD__AND2_4%VPWR N_VPWR_M1006_s N_VPWR_M1010_d N_VPWR_M1004_s
+ N_VPWR_M1011_s N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n
+ N_VPWR_c_235_n N_VPWR_c_236_n VPWR N_VPWR_c_237_n N_VPWR_c_238_n
+ N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_230_n
+ PM_SKY130_FD_SC_HD__AND2_4%VPWR
x_PM_SKY130_FD_SC_HD__AND2_4%X N_X_M1002_d N_X_M1007_d N_X_M1001_d N_X_M1009_d
+ N_X_c_312_n N_X_c_289_n N_X_c_292_n N_X_c_296_n N_X_c_332_p N_X_c_316_n
+ N_X_c_298_n N_X_c_287_n N_X_c_302_n N_X_c_304_n N_X_c_306_n X N_X_c_285_n X
+ PM_SKY130_FD_SC_HD__AND2_4%X
x_PM_SKY130_FD_SC_HD__AND2_4%VGND N_VGND_M1000_d N_VGND_M1003_s N_VGND_M1008_s
+ N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n VGND
+ N_VGND_c_347_n N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n
+ N_VGND_c_352_n PM_SKY130_FD_SC_HD__AND2_4%VGND
cc_1 VNB N_A_c_57_n 0.0302805f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_2 VNB N_A_c_58_n 0.0141299f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_3 VNB N_A_c_59_n 0.021624f $X=-0.19 $Y=-0.24 $X2=0.382 $Y2=0.995
cc_4 VNB N_B_c_84_n 0.0213314f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_5 VNB N_B_c_85_n 0.00330631f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_6 VNB N_B_c_86_n 0.0171393f $X=-0.19 $Y=-0.24 $X2=0.382 $Y2=0.995
cc_7 VNB N_A_27_47#_c_122_n 0.0169849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_123_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=0.382 $Y2=1.325
cc_9 VNB N_A_27_47#_c_124_n 0.0160024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_125_n 0.0184169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_126_n 0.0141802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_127_n 0.00929734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_128_n 0.00127837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_129_n 0.00171227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_130_n 0.0667411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_230_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_285_n 0.0108749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0235754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_343_n 0.00501393f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_20 VNB N_VGND_c_344_n 3.21684e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_345_n 0.0115115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_346_n 0.0107852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_347_n 0.0268617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_348_n 0.015947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_349_n 0.0113516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_350_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_351_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_352_n 0.180667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_M1006_g 0.0225934f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_30 VPB N_A_c_57_n 0.00688583f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_31 VPB N_A_c_58_n 0.0116013f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_32 VPB N_B_M1010_g 0.0201094f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_33 VPB N_B_c_84_n 0.00438023f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_34 VPB N_B_c_85_n 0.0017826f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_35 VPB N_A_27_47#_M1001_g 0.0188029f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_36 VPB N_A_27_47#_M1004_g 0.018288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_M1009_g 0.0183103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_M1011_g 0.0210399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_135_n 0.00127073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_136_n 0.00920717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_129_n 4.55278e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_130_n 0.0124075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_231_n 0.0103398f $X=-0.19 $Y=1.305 $X2=0.382 $Y2=0.995
cc_44 VPB N_VPWR_c_232_n 0.0273818f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_45 VPB N_VPWR_c_233_n 0.00431378f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_234_n 3.16049e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_235_n 0.0117752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_236_n 0.0236962f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_237_n 0.0151816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_238_n 0.0152595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_239_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_240_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_241_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_230_n 0.04486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_X_c_287_n 0.0124234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB X 0.0114218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 N_A_M1006_g N_B_M1010_g 0.0245388f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A_c_58_n N_B_M1010_g 0.00129134f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_c_57_n N_B_c_84_n 0.038114f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_c_58_n N_B_c_84_n 2.57313e-19 $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_c_57_n N_B_c_85_n 0.00237503f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_c_58_n N_B_c_85_n 0.0262305f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_c_59_n N_B_c_86_n 0.038114f $X=0.382 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A_c_59_n N_A_27_47#_c_126_n 0.00636458f $X=0.382 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A_c_58_n N_A_27_47#_c_140_n 5.95137e-19 $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_59_n N_A_27_47#_c_140_n 0.0119563f $X=0.382 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A_c_57_n N_A_27_47#_c_127_n 0.00123469f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_c_58_n N_A_27_47#_c_127_n 0.0214429f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_c_59_n N_A_27_47#_c_127_n 7.78534e-19 $X=0.382 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_c_58_n N_VPWR_M1006_s 0.00332814f $X=0.35 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_71 N_A_M1006_g N_VPWR_c_232_n 0.011618f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_c_57_n N_VPWR_c_232_n 6.75944e-19 $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_c_58_n N_VPWR_c_232_n 0.0153825f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_M1006_g N_VPWR_c_237_n 0.00486043f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1006_g N_VPWR_c_230_n 0.00825064f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_c_59_n N_VGND_c_347_n 0.0041289f $X=0.382 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_c_59_n N_VGND_c_352_n 0.00651126f $X=0.382 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B_c_86_n N_A_27_47#_c_122_n 0.0225638f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B_M1010_g N_A_27_47#_M1001_g 0.0204134f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_80 N_B_c_86_n N_A_27_47#_c_126_n 0.00138685f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_84_n N_A_27_47#_c_140_n 0.00354699f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B_c_85_n N_A_27_47#_c_140_n 0.0219556f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B_c_86_n N_A_27_47#_c_140_n 0.0128622f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B_M1010_g N_A_27_47#_c_151_n 0.0154459f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_85 N_B_c_85_n N_A_27_47#_c_151_n 0.00896924f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B_c_84_n N_A_27_47#_c_153_n 6.00846e-19 $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B_c_85_n N_A_27_47#_c_153_n 0.011078f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B_c_85_n N_A_27_47#_c_128_n 0.0018209f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_c_86_n N_A_27_47#_c_128_n 0.00398737f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B_M1010_g N_A_27_47#_c_135_n 0.00498595f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_91 N_B_M1010_g N_A_27_47#_c_129_n 8.45385e-19 $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B_c_84_n N_A_27_47#_c_129_n 0.00243438f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_c_85_n N_A_27_47#_c_129_n 0.025987f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B_c_84_n N_A_27_47#_c_130_n 0.0124263f $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B_c_85_n N_A_27_47#_c_130_n 2.86813e-19 $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B_M1010_g N_VPWR_c_232_n 6.33335e-19 $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B_M1010_g N_VPWR_c_233_n 0.00171766f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B_M1010_g N_VPWR_c_237_n 0.00585385f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_99 N_B_M1010_g N_VPWR_c_230_n 0.0107105f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B_c_86_n N_VGND_c_343_n 0.00441145f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B_c_86_n N_VGND_c_347_n 0.00422112f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B_c_86_n N_VGND_c_352_n 0.00593409f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_151_n N_VPWR_M1010_d 0.00696425f $X=1.15 $Y=1.665 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_135_n N_VPWR_M1010_d 0.00111849f $X=1.255 $Y=1.58 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_M1001_g N_VPWR_c_233_n 0.00170185f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_151_n N_VPWR_c_233_n 0.0193839f $X=1.15 $Y=1.665 $X2=0 $Y2=0
cc_107 N_A_27_47#_M1001_g N_VPWR_c_234_n 6.10667e-19 $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_M1004_g N_VPWR_c_234_n 0.00979109f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1009_g N_VPWR_c_234_n 0.00969908f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_M1011_g N_VPWR_c_234_n 5.94761e-19 $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1009_g N_VPWR_c_236_n 5.94761e-19 $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_M1011_g N_VPWR_c_236_n 0.0107575f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_173_p N_VPWR_c_237_n 0.012099f $X=0.69 $Y=1.96 $X2=0 $Y2=0
cc_114 N_A_27_47#_M1001_g N_VPWR_c_238_n 0.00585385f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1004_g N_VPWR_c_238_n 0.00486043f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_M1009_g N_VPWR_c_239_n 0.00486043f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_M1011_g N_VPWR_c_239_n 0.00486043f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_27_47#_M1006_d N_VPWR_c_230_n 0.00570388f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_M1001_g N_VPWR_c_230_n 0.0106977f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1004_g N_VPWR_c_230_n 0.00822531f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_M1009_g N_VPWR_c_230_n 0.00822531f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_M1011_g N_VPWR_c_230_n 0.00822531f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_173_p N_VPWR_c_230_n 0.00684987f $X=0.69 $Y=1.96 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_123_n N_X_c_289_n 0.011111f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_124_n N_X_c_289_n 0.0110478f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_130_n N_X_c_289_n 0.00231838f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1004_g N_X_c_292_n 0.016114f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1009_g N_X_c_292_n 0.0139045f $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_136_n N_X_c_292_n 0.0417385f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_130_n N_X_c_292_n 6.56764e-19 $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_136_n N_X_c_296_n 0.0147839f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_130_n N_X_c_296_n 7.2697e-19 $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_125_n N_X_c_298_n 0.0160286f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_136_n N_X_c_298_n 0.00590462f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1011_g N_X_c_287_n 0.019007f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_136_n N_X_c_287_n 0.00595992f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_136_n N_X_c_302_n 0.0546247f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_130_n N_X_c_302_n 0.00234013f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_136_n N_X_c_304_n 0.0141519f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_130_n N_X_c_304_n 0.00238051f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_136_n N_X_c_306_n 0.0147839f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_130_n N_X_c_306_n 7.2697e-19 $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_125_n X 0.0240627f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_136_n X 0.0275568f $X=2.52 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_140_n A_110_47# 0.00271764f $X=1.15 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_27_47#_c_140_n N_VGND_M1000_d 0.00919698f $X=1.15 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_27_47#_c_128_n N_VGND_M1000_d 9.90294e-19 $X=1.255 $Y=1.02 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_27_47#_c_122_n N_VGND_c_343_n 0.00296124f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_140_n N_VGND_c_343_n 0.024657f $X=1.15 $Y=0.71 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_122_n N_VGND_c_344_n 0.00109054f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_c_123_n N_VGND_c_344_n 0.00804258f $X=1.84 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_124_n N_VGND_c_344_n 0.00625485f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_125_n N_VGND_c_344_n 4.98572e-19 $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_124_n N_VGND_c_346_n 4.98572e-19 $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_125_n N_VGND_c_346_n 0.00731833f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_126_n N_VGND_c_347_n 0.0207561f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_140_n N_VGND_c_347_n 0.00814185f $X=1.15 $Y=0.71 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_122_n N_VGND_c_348_n 0.00558147f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_123_n N_VGND_c_348_n 0.00351072f $X=1.84 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_140_n N_VGND_c_348_n 9.77174e-19 $X=1.15 $Y=0.71 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_124_n N_VGND_c_349_n 0.00351072f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_125_n N_VGND_c_349_n 0.00351072f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1005_s N_VGND_c_352_n 0.00213418f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_122_n N_VGND_c_352_n 0.0102604f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_123_n N_VGND_c_352_n 0.00411677f $X=1.84 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_124_n N_VGND_c_352_n 0.0040731f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_125_n N_VGND_c_352_n 0.0040731f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_126_n N_VGND_c_352_n 0.0123808f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_140_n N_VGND_c_352_n 0.0176947f $X=1.15 $Y=0.71 $X2=0 $Y2=0
cc_170 N_VPWR_c_230_n N_X_M1001_d 0.00535672f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_171 N_VPWR_c_230_n N_X_M1009_d 0.00535672f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_172 N_VPWR_c_238_n N_X_c_312_n 0.0124538f $X=1.89 $Y=2.72 $X2=0 $Y2=0
cc_173 N_VPWR_c_230_n N_X_c_312_n 0.00724021f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_174 N_VPWR_M1004_s N_X_c_292_n 0.00340327f $X=1.915 $Y=1.485 $X2=0 $Y2=0
cc_175 N_VPWR_c_234_n N_X_c_292_n 0.0170296f $X=2.055 $Y=2.02 $X2=0 $Y2=0
cc_176 N_VPWR_c_239_n N_X_c_316_n 0.0124538f $X=2.75 $Y=2.72 $X2=0 $Y2=0
cc_177 N_VPWR_c_230_n N_X_c_316_n 0.00724021f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_178 N_VPWR_M1011_s N_X_c_287_n 0.00470097f $X=2.775 $Y=1.485 $X2=0 $Y2=0
cc_179 N_VPWR_c_236_n N_X_c_287_n 0.0239152f $X=2.915 $Y=2.02 $X2=0 $Y2=0
cc_180 N_VPWR_M1011_s X 8.60883e-19 $X=2.775 $Y=1.485 $X2=0 $Y2=0
cc_181 N_X_c_289_n N_VGND_M1003_s 0.00327388f $X=2.39 $Y=0.73 $X2=0 $Y2=0
cc_182 N_X_c_298_n N_VGND_M1008_s 0.0010969f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_183 N_X_c_285_n N_VGND_M1008_s 0.00351052f $X=2.995 $Y=0.845 $X2=0 $Y2=0
cc_184 X N_VGND_M1008_s 6.85193e-19 $X=2.99 $Y=0.85 $X2=0 $Y2=0
cc_185 N_X_c_289_n N_VGND_c_344_n 0.0162283f $X=2.39 $Y=0.73 $X2=0 $Y2=0
cc_186 N_X_c_285_n N_VGND_c_345_n 0.00116793f $X=2.995 $Y=0.845 $X2=0 $Y2=0
cc_187 N_X_c_298_n N_VGND_c_346_n 0.00344107f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_188 N_X_c_285_n N_VGND_c_346_n 0.0188167f $X=2.995 $Y=0.845 $X2=0 $Y2=0
cc_189 N_X_c_289_n N_VGND_c_348_n 0.00263122f $X=2.39 $Y=0.73 $X2=0 $Y2=0
cc_190 N_X_c_302_n N_VGND_c_348_n 0.00436709f $X=1.72 $Y=0.68 $X2=0 $Y2=0
cc_191 N_X_c_289_n N_VGND_c_349_n 0.00263122f $X=2.39 $Y=0.73 $X2=0 $Y2=0
cc_192 N_X_c_332_p N_VGND_c_349_n 0.0123333f $X=2.485 $Y=0.42 $X2=0 $Y2=0
cc_193 N_X_c_298_n N_VGND_c_349_n 0.00263122f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_194 N_X_M1002_d N_VGND_c_352_n 0.00434391f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_195 N_X_M1007_d N_VGND_c_352_n 0.00251209f $X=2.345 $Y=0.235 $X2=0 $Y2=0
cc_196 N_X_c_289_n N_VGND_c_352_n 0.0101713f $X=2.39 $Y=0.73 $X2=0 $Y2=0
cc_197 N_X_c_332_p N_VGND_c_352_n 0.00721345f $X=2.485 $Y=0.42 $X2=0 $Y2=0
cc_198 N_X_c_298_n N_VGND_c_352_n 0.00477848f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_199 N_X_c_302_n N_VGND_c_352_n 0.00604783f $X=1.72 $Y=0.68 $X2=0 $Y2=0
cc_200 N_X_c_285_n N_VGND_c_352_n 0.00289812f $X=2.995 $Y=0.845 $X2=0 $Y2=0
cc_201 A_110_47# N_VGND_c_352_n 0.00239227f $X=0.55 $Y=0.235 $X2=1.255 $Y2=0.805

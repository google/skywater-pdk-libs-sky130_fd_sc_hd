* File: sky130_fd_sc_hd__decap_3.pxi.spice
* Created: Tue Sep  1 19:02:08 2020
* 
x_PM_SKY130_FD_SC_HD__DECAP_3%VGND N_VGND_M1001_s N_VGND_c_13_n N_VGND_M1000_g
+ N_VGND_c_14_n VGND N_VGND_c_15_n N_VGND_c_16_n
+ PM_SKY130_FD_SC_HD__DECAP_3%VGND
x_PM_SKY130_FD_SC_HD__DECAP_3%VPWR N_VPWR_M1000_s N_VPWR_c_27_n VPWR
+ N_VPWR_M1001_g N_VPWR_c_31_n N_VPWR_c_29_n PM_SKY130_FD_SC_HD__DECAP_3%VPWR
cc_1 VNB N_VGND_c_13_n 0.0201334f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.76
cc_2 VNB N_VGND_c_14_n 0.0220173f $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=1.29
cc_3 VNB N_VGND_c_15_n 0.0862828f $X=-0.19 $Y=-0.24 $X2=1.12 $Y2=0.485
cc_4 VNB N_VGND_c_16_n 0.102847f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=0
cc_5 VNB N_VPWR_c_27_n 0.0157537f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=2.05
cc_6 VNB N_VPWR_M1001_g 0.0971894f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=-0.085
cc_7 VNB N_VPWR_c_29_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=1.12 $Y2=0.375
cc_8 VPB N_VGND_c_13_n 0.0794504f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.76
cc_9 VPB N_VGND_c_14_n 0.00511056f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.29
cc_10 VPB N_VPWR_c_27_n 0.0113742f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=2.05
cc_11 VPB N_VPWR_c_31_n 0.115327f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.375
cc_12 VPB N_VPWR_c_29_n 0.0418596f $X=-0.19 $Y=1.305 $X2=1.12 $Y2=0.375
cc_13 N_VGND_c_13_n N_VPWR_c_27_n 0.0139364f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_14 N_VGND_c_14_n N_VPWR_c_27_n 0.0329927f $X=0.42 $Y=1.29 $X2=0 $Y2=0
cc_15 N_VGND_c_15_n N_VPWR_c_27_n 0.0460926f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_16 N_VGND_c_13_n N_VPWR_M1001_g 0.03778f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_17 N_VGND_c_14_n N_VPWR_M1001_g 0.0139364f $X=0.42 $Y=1.29 $X2=0 $Y2=0
cc_18 N_VGND_c_15_n N_VPWR_M1001_g 0.0749649f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_19 N_VGND_c_13_n N_VPWR_c_31_n 0.0936943f $X=0.69 $Y=1.76 $X2=0 $Y2=0
cc_20 N_VGND_c_14_n N_VPWR_c_31_n 0.0460926f $X=0.42 $Y=1.29 $X2=0 $Y2=0

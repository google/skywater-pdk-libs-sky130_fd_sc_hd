* File: sky130_fd_sc_hd__and3_1.spice.SKY130_FD_SC_HD__AND3_1.pxi
* Created: Thu Aug 27 14:07:34 2020
* 
x_PM_SKY130_FD_SC_HD__AND3_1%A N_A_M1006_g N_A_M1004_g A N_A_c_54_n N_A_c_55_n
+ PM_SKY130_FD_SC_HD__AND3_1%A
x_PM_SKY130_FD_SC_HD__AND3_1%B N_B_M1002_g N_B_M1000_g N_B_c_80_n B N_B_c_84_n
+ PM_SKY130_FD_SC_HD__AND3_1%B
x_PM_SKY130_FD_SC_HD__AND3_1%C N_C_c_118_n N_C_M1003_g N_C_c_119_n N_C_M1007_g C
+ C N_C_c_122_n PM_SKY130_FD_SC_HD__AND3_1%C
x_PM_SKY130_FD_SC_HD__AND3_1%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1004_s
+ N_A_27_47#_M1000_d N_A_27_47#_M1001_g N_A_27_47#_M1005_g N_A_27_47#_c_164_n
+ N_A_27_47#_c_173_n N_A_27_47#_c_165_n N_A_27_47#_c_166_n N_A_27_47#_c_167_n
+ N_A_27_47#_c_176_n N_A_27_47#_c_168_n N_A_27_47#_c_169_n N_A_27_47#_c_170_n
+ N_A_27_47#_c_171_n PM_SKY130_FD_SC_HD__AND3_1%A_27_47#
x_PM_SKY130_FD_SC_HD__AND3_1%VPWR N_VPWR_M1004_d N_VPWR_M1007_d N_VPWR_c_252_n
+ VPWR N_VPWR_c_253_n N_VPWR_c_254_n N_VPWR_c_251_n N_VPWR_c_256_n
+ N_VPWR_c_257_n PM_SKY130_FD_SC_HD__AND3_1%VPWR
x_PM_SKY130_FD_SC_HD__AND3_1%X N_X_M1001_d N_X_M1005_d N_X_c_287_n N_X_c_284_n
+ N_X_c_285_n X X N_X_c_289_n PM_SKY130_FD_SC_HD__AND3_1%X
x_PM_SKY130_FD_SC_HD__AND3_1%VGND N_VGND_M1003_d N_VGND_c_308_n VGND
+ N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n
+ PM_SKY130_FD_SC_HD__AND3_1%VGND
cc_1 VNB N_A_M1004_g 0.00264232f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.71
cc_2 VNB A 0.0190658f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A_c_54_n 0.064248f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_4 VNB N_A_c_55_n 0.0169709f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=0.73
cc_5 VNB N_B_M1002_g 0.0364558f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_6 VNB N_B_c_80_n 0.00261095f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=0.93
cc_7 VNB N_C_c_118_n 0.0150959f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_8 VNB N_C_c_119_n 0.0427505f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.255
cc_9 VNB N_C_M1007_g 3.96206e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.71
cc_10 VNB C 0.00647375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_C_c_122_n 0.00151102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_164_n 0.00795526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_165_n 0.00339252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_166_n 0.00504859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_167_n 0.0031774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_168_n 0.00330364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_169_n 0.00358757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_170_n 0.0230819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_171_n 0.0204922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_251_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_284_n 0.0251181f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=0.93
cc_22 VNB N_X_c_285_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_23 VNB X 0.0136214f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=0.73
cc_24 VNB N_VGND_c_308_n 0.00237268f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.71
cc_25 VNB N_VGND_c_309_n 0.0413951f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=0.93
cc_26 VNB N_VGND_c_310_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_311_n 0.142297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_312_n 0.00354115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_M1004_g 0.0277804f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.71
cc_30 VPB N_B_M1000_g 0.0164719f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_31 VPB N_B_c_80_n 0.00666805f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=0.93
cc_32 VPB B 0.0107794f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.93
cc_33 VPB N_B_c_84_n 0.0358203f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=1.255
cc_34 VPB N_C_M1007_g 0.0216299f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.71
cc_35 VPB N_A_27_47#_M1005_g 0.0234651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_47#_c_173_n 0.0185069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_c_165_n 0.00279331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_166_n 0.00224001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_176_n 0.00874548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_168_n 0.00682202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_169_n 6.58508e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_170_n 0.00513253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_252_n 0.00248325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_253_n 0.0215577f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=0.73
cc_45 VPB N_VPWR_c_254_n 0.0153939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_251_n 0.0510087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_256_n 0.0593285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_257_n 0.00372629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_X_c_287_n 0.00524127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_X_c_284_n 0.0183925f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=0.93
cc_51 VPB N_X_c_289_n 0.0218575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 A N_B_M1002_g 0.00231842f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_53 N_A_c_55_n N_B_M1002_g 0.0408653f $X=0.335 $Y=0.73 $X2=0 $Y2=0
cc_54 N_A_M1004_g N_B_M1000_g 0.0169206f $X=0.47 $Y=1.71 $X2=0 $Y2=0
cc_55 N_A_c_54_n N_B_c_80_n 0.0408653f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_56 A N_A_27_47#_M1006_s 0.00212885f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_57 A N_A_27_47#_c_164_n 0.0313092f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_58 N_A_c_54_n N_A_27_47#_c_164_n 0.00137178f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_59 N_A_c_55_n N_A_27_47#_c_164_n 0.00744605f $X=0.335 $Y=0.73 $X2=0 $Y2=0
cc_60 N_A_M1004_g N_A_27_47#_c_173_n 0.00363759f $X=0.47 $Y=1.71 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_A_27_47#_c_165_n 0.00833123f $X=0.47 $Y=1.71 $X2=0 $Y2=0
cc_62 A N_A_27_47#_c_165_n 0.021679f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_54_n N_A_27_47#_c_165_n 0.00529802f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_64 A N_A_27_47#_c_166_n 0.0212009f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_c_54_n N_A_27_47#_c_166_n 0.0104883f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_66 A N_A_27_47#_c_167_n 0.0303199f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_A_c_54_n N_A_27_47#_c_167_n 0.00110744f $X=0.26 $Y=0.93 $X2=0 $Y2=0
cc_68 N_A_c_55_n N_A_27_47#_c_167_n 0.00138373f $X=0.335 $Y=0.73 $X2=0 $Y2=0
cc_69 N_A_M1004_g N_A_27_47#_c_168_n 0.00136653f $X=0.47 $Y=1.71 $X2=0 $Y2=0
cc_70 N_A_M1004_g N_VPWR_c_256_n 0.022834f $X=0.47 $Y=1.71 $X2=0 $Y2=0
cc_71 A A_109_47# 5.06513e-19 $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_72 N_A_c_55_n N_VGND_c_309_n 0.00366111f $X=0.335 $Y=0.73 $X2=0 $Y2=0
cc_73 N_A_c_55_n N_VGND_c_311_n 0.00605974f $X=0.335 $Y=0.73 $X2=0 $Y2=0
cc_74 N_B_M1002_g N_C_c_118_n 0.0625976f $X=0.83 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_75 N_B_M1002_g N_C_c_119_n 0.00711137f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_76 N_B_c_80_n N_C_c_119_n 6.15948e-19 $X=0.86 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B_c_80_n N_C_M1007_g 0.0141608f $X=0.86 $Y=1.41 $X2=0 $Y2=0
cc_78 B N_C_M1007_g 0.00201949f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_79 N_B_M1002_g C 2.52771e-19 $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_80 N_B_M1002_g N_C_c_122_n 8.64309e-19 $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_81 B N_A_27_47#_M1005_g 6.22676e-19 $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_82 N_B_c_84_n N_A_27_47#_M1005_g 0.00185069f $X=0.95 $Y=2.295 $X2=0 $Y2=0
cc_83 N_B_M1002_g N_A_27_47#_c_164_n 0.00818238f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_84 N_B_M1002_g N_A_27_47#_c_167_n 0.0158484f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_85 B N_A_27_47#_c_176_n 0.0133235f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_86 N_B_M1002_g N_A_27_47#_c_168_n 0.00495536f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_87 N_B_M1000_g N_A_27_47#_c_168_n 0.00873905f $X=0.89 $Y=1.71 $X2=0 $Y2=0
cc_88 N_B_c_80_n N_A_27_47#_c_168_n 0.00651041f $X=0.86 $Y=1.41 $X2=0 $Y2=0
cc_89 B N_A_27_47#_c_168_n 0.00827708f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_90 N_B_c_84_n N_A_27_47#_c_168_n 4.84666e-19 $X=0.95 $Y=2.295 $X2=0 $Y2=0
cc_91 N_B_M1000_g N_VPWR_c_252_n 8.70215e-19 $X=0.89 $Y=1.71 $X2=0 $Y2=0
cc_92 B N_VPWR_c_252_n 0.0280643f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_93 N_B_c_84_n N_VPWR_c_252_n 7.79965e-19 $X=0.95 $Y=2.295 $X2=0 $Y2=0
cc_94 B N_VPWR_c_253_n 0.0324753f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_95 N_B_c_84_n N_VPWR_c_253_n 0.00329641f $X=0.95 $Y=2.295 $X2=0 $Y2=0
cc_96 B N_VPWR_c_251_n 0.0181571f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_97 N_B_c_84_n N_VPWR_c_251_n 0.00178749f $X=0.95 $Y=2.295 $X2=0 $Y2=0
cc_98 N_B_M1000_g N_VPWR_c_256_n 0.0172349f $X=0.89 $Y=1.71 $X2=0 $Y2=0
cc_99 N_B_c_80_n N_VPWR_c_256_n 2.0902e-19 $X=0.86 $Y=1.41 $X2=0 $Y2=0
cc_100 B N_VPWR_c_256_n 0.0284614f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_101 N_B_M1002_g N_VGND_c_309_n 0.00365976f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_102 N_B_M1002_g N_VGND_c_311_n 0.00500957f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_103 N_C_M1007_g N_A_27_47#_M1005_g 0.0270827f $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_104 N_C_c_118_n N_A_27_47#_c_164_n 0.00107441f $X=1.19 $Y=0.73 $X2=0 $Y2=0
cc_105 N_C_c_122_n N_A_27_47#_c_164_n 0.0128492f $X=1.31 $Y=0.79 $X2=0 $Y2=0
cc_106 N_C_c_118_n N_A_27_47#_c_167_n 0.00349053f $X=1.19 $Y=0.73 $X2=0 $Y2=0
cc_107 N_C_c_122_n N_A_27_47#_c_167_n 0.0536032f $X=1.31 $Y=0.79 $X2=0 $Y2=0
cc_108 N_C_c_119_n N_A_27_47#_c_176_n 0.00496171f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_109 N_C_M1007_g N_A_27_47#_c_176_n 0.0199191f $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_110 C N_A_27_47#_c_176_n 0.0277011f $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_111 N_C_c_119_n N_A_27_47#_c_168_n 0.00112048f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_112 N_C_M1007_g N_A_27_47#_c_168_n 9.77432e-19 $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_113 C N_A_27_47#_c_168_n 0.00221086f $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_114 N_C_c_119_n N_A_27_47#_c_169_n 0.00144494f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_115 N_C_M1007_g N_A_27_47#_c_169_n 8.68757e-19 $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_116 C N_A_27_47#_c_169_n 0.0182304f $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_117 N_C_c_119_n N_A_27_47#_c_170_n 0.0192014f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_118 N_C_M1007_g N_A_27_47#_c_170_n 0.00160999f $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_119 C N_A_27_47#_c_170_n 7.08195e-19 $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_120 N_C_c_118_n N_A_27_47#_c_171_n 0.00877122f $X=1.19 $Y=0.73 $X2=0 $Y2=0
cc_121 N_C_c_119_n N_A_27_47#_c_171_n 0.00621969f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_122 C N_A_27_47#_c_171_n 0.00198953f $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_123 N_C_c_122_n N_A_27_47#_c_171_n 0.00177508f $X=1.31 $Y=0.79 $X2=0 $Y2=0
cc_124 N_C_M1007_g N_VPWR_c_253_n 0.00193172f $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_125 N_C_M1007_g N_VPWR_c_251_n 0.00238657f $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_126 N_C_M1007_g N_VPWR_c_256_n 3.17213e-19 $X=1.355 $Y=1.71 $X2=0 $Y2=0
cc_127 C N_X_c_284_n 0.00665115f $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_128 N_C_c_122_n N_VGND_M1003_d 0.00386934f $X=1.31 $Y=0.79 $X2=-0.19
+ $Y2=-0.24
cc_129 N_C_c_118_n N_VGND_c_308_n 0.00434006f $X=1.19 $Y=0.73 $X2=0 $Y2=0
cc_130 N_C_c_122_n N_VGND_c_308_n 0.0243913f $X=1.31 $Y=0.79 $X2=0 $Y2=0
cc_131 N_C_c_118_n N_VGND_c_309_n 0.00412865f $X=1.19 $Y=0.73 $X2=0 $Y2=0
cc_132 N_C_c_122_n N_VGND_c_309_n 0.00989316f $X=1.31 $Y=0.79 $X2=0 $Y2=0
cc_133 N_C_c_118_n N_VGND_c_311_n 0.00678637f $X=1.19 $Y=0.73 $X2=0 $Y2=0
cc_134 C N_VGND_c_311_n 0.0042617f $X=1.26 $Y=0.85 $X2=0 $Y2=0
cc_135 N_C_c_122_n N_VGND_c_311_n 0.00762473f $X=1.31 $Y=0.79 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_176_n N_VPWR_M1007_d 0.0027927f $X=1.645 $Y=1.635 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_M1005_g N_VPWR_c_252_n 0.0110297f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_176_n N_VPWR_c_252_n 0.0144383f $X=1.645 $Y=1.635 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_M1005_g N_VPWR_c_254_n 0.00525069f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1005_g N_VPWR_c_251_n 0.00987998f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_c_176_n N_VPWR_c_251_n 0.00773634f $X=1.645 $Y=1.635 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_173_n N_VPWR_c_256_n 0.0233778f $X=0.26 $Y=1.645 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_165_n N_VPWR_c_256_n 0.0126037f $X=0.71 $Y=1.275 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_168_n N_VPWR_c_256_n 0.0052698f $X=1.1 $Y=1.635 $X2=0 $Y2=0
cc_145 N_A_27_47#_M1005_g N_X_c_284_n 0.00837861f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_176_n N_X_c_284_n 0.0257002f $X=1.645 $Y=1.635 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_169_n N_X_c_284_n 0.0287806f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_170_n N_X_c_284_n 0.00753248f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_171_n N_X_c_284_n 0.00682852f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_164_n A_109_47# 0.00376423f $X=0.805 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_27_47#_c_164_n A_181_47# 0.0016621f $X=0.805 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_27_47#_c_167_n A_181_47# 0.00156681f $X=0.89 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_27_47#_c_164_n N_VGND_c_308_n 3.41305e-19 $X=0.805 $Y=0.38 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_169_n N_VGND_c_308_n 0.00563404f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_170_n N_VGND_c_308_n 4.70982e-19 $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_171_n N_VGND_c_308_n 0.0108815f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_164_n N_VGND_c_309_n 0.0400798f $X=0.805 $Y=0.38 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_171_n N_VGND_c_310_n 0.0046653f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_27_47#_M1006_s N_VGND_c_311_n 0.00211652f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_164_n N_VGND_c_311_n 0.0311117f $X=0.805 $Y=0.38 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_171_n N_VGND_c_311_n 0.00895857f $X=1.79 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_VPWR_c_251_n N_X_M1005_d 0.00335098f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_c_254_n N_X_c_289_n 0.0185457f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_164 N_VPWR_c_251_n N_X_c_289_n 0.0105168f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_165 X N_VGND_c_310_n 0.0178555f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_166 N_X_M1001_d N_VGND_c_311_n 0.00387172f $X=1.905 $Y=0.235 $X2=0 $Y2=0
cc_167 X N_VGND_c_311_n 0.00990557f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_168 A_109_47# N_VGND_c_311_n 0.0017052f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_169 A_181_47# N_VGND_c_311_n 0.00655254f $X=0.905 $Y=0.235 $X2=0.26 $Y2=0.38

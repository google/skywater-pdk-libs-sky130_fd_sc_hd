* File: sky130_fd_sc_hd__dfbbn_2.spice
* Created: Thu Aug 27 14:14:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dfbbn_2.pex.spice"
.subckt sky130_fd_sc_hd__dfbbn_2  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1038 N_VGND_M1038_d N_CLK_N_M1038_g N_A_27_47#_M1038_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_193_47#_M1025_d N_A_27_47#_M1025_g N_VGND_M1038_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_381_47#_M1011_d N_D_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.1092 PD=0.802308 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1036 N_A_476_47#_M1036_d N_A_193_47#_M1036_g N_A_381_47#_M1011_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0702 AS=0.0609231 PD=0.75 PS=0.687692 NRD=19.992 NRS=16.656
+ M=1 R=2.4 SA=75000.7 SB=75002.7 A=0.054 P=1.02 MULT=1
MM1006 A_584_47# N_A_27_47#_M1006_g N_A_476_47#_M1036_d VNB NSHORT L=0.15 W=0.36
+ AD=0.0618923 AS=0.0702 PD=0.692308 PS=0.75 NRD=38.964 NRS=16.656 M=1 R=2.4
+ SA=75001.2 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1012 N_VGND_M1012_d N_A_650_21#_M1012_g A_584_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.084 AS=0.0722077 PD=0.82 PS=0.807692 NRD=35.712 NRS=33.396 M=1 R=2.8
+ SA=75001.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1037 N_A_790_47#_M1037_d N_SET_B_M1037_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0800377 AS=0.084 PD=0.784528 PS=0.82 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1035 N_A_650_21#_M1035_d N_A_476_47#_M1035_g N_A_790_47#_M1037_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0864 AS=0.121962 PD=0.91 PS=1.19547 NRD=0 NRS=14.052 M=1
+ R=4.26667 SA=75001.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1042 N_A_790_47#_M1042_d N_A_944_21#_M1042_g N_A_650_21#_M1035_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 A_1162_47# N_A_650_21#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.11968 AS=0.1664 PD=1.2352 PS=1.8 NRD=24.744 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1007 N_A_1257_47#_M1007_d N_A_27_47#_M1007_g A_1162_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0711 AS=0.06732 PD=0.755 PS=0.6948 NRD=23.328 NRS=43.992 M=1 R=2.4
+ SA=75000.7 SB=75002.7 A=0.054 P=1.02 MULT=1
MM1004 A_1366_47# N_A_193_47#_M1004_g N_A_1257_47#_M1007_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0711 PD=0.687692 PS=0.755 NRD=38.076 NRS=14.988 M=1
+ R=2.4 SA=75001.2 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1024 N_VGND_M1024_d N_A_1431_21#_M1024_g A_1366_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0710769 PD=0.7 PS=0.802308 NRD=1.428 NRS=32.628 M=1 R=2.8
+ SA=75001.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_1547_47#_M1005_d N_SET_B_M1005_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0950151 AS=0.0588 PD=0.855849 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_1431_21#_M1008_d N_A_1257_47#_M1008_g N_A_1547_47#_M1005_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0864 AS=0.144785 PD=0.91 PS=1.30415 NRD=0 NRS=14.052 M=1
+ R=4.26667 SA=75001.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1016 N_A_1547_47#_M1016_d N_A_944_21#_M1016_g N_A_1431_21#_M1008_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.176 AS=0.0864 PD=1.83 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VGND_M1027_d N_RESET_B_M1027_g N_A_944_21#_M1027_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0787009 AS=0.1113 PD=0.773271 PS=1.37 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1027_d N_A_1431_21#_M1003_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_A_1431_21#_M1022_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.195 AS=0.08775 PD=1.9 PS=0.92 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_A_1431_21#_M1017_g N_A_2236_47#_M1017_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1033 N_Q_M1033_d N_A_2236_47#_M1033_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11785 PD=0.92 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1040 N_Q_M1033_d N_A_2236_47#_M1040_g N_VGND_M1040_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1023 N_VPWR_M1023_d N_CLK_N_M1023_g N_A_27_47#_M1023_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1023_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_381_47#_M1029_d N_D_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06825 AS=0.1092 PD=0.745 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75007 A=0.063 P=1.14 MULT=1
MM1018 N_A_476_47#_M1018_d N_A_27_47#_M1018_g N_A_381_47#_M1029_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.06825 PD=0.69 PS=0.745 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75000.7 SB=75006.5 A=0.063 P=1.14 MULT=1
MM1009 A_560_413# N_A_193_47#_M1009_g N_A_476_47#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0945 AS=0.0567 PD=0.87 PS=0.69 NRD=79.7259 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75006.1 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_650_21#_M1015_g A_560_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0945 PD=0.8 PS=0.87 NRD=21.0987 NRS=79.7259 M=1 R=2.8
+ SA=75001.7 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1041 N_A_650_21#_M1041_d N_SET_B_M1041_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.098 AS=0.0798 PD=0.82 PS=0.8 NRD=53.9386 NRS=25.7873 M=1 R=2.8
+ SA=75002.2 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1020 A_894_329# N_A_476_47#_M1020_g N_A_650_21#_M1041_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.105 AS=0.196 PD=1.09 PS=1.64 NRD=16.4101 NRS=0 M=1 R=5.6
+ SA=75001.5 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1032 N_VPWR_M1032_d N_A_944_21#_M1032_g A_894_329# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2331 AS=0.105 PD=1.395 PS=1.09 NRD=10.5395 NRS=16.4101 M=1 R=5.6
+ SA=75001.9 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1028 A_1115_329# N_A_650_21#_M1028_g N_VPWR_M1032_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2324 AS=0.2331 PD=1.88 PS=1.395 NRD=51.9686 NRS=53.9386 M=1 R=5.6
+ SA=75002.6 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1031 N_A_1257_47#_M1031_d N_A_193_47#_M1031_g A_1115_329# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.1162 PD=0.69 PS=0.94 NRD=0 NRS=103.957 M=1 R=2.8
+ SA=75004.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1019 A_1343_413# N_A_27_47#_M1019_g N_A_1257_47#_M1031_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.0567 PD=0.86 PS=0.69 NRD=77.3816 NRS=0 M=1 R=2.8
+ SA=75005 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1431_21#_M1034_g A_1343_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0924 PD=0.81 PS=0.86 NRD=25.7873 NRS=77.3816 M=1 R=2.8
+ SA=75005.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_1431_21#_M1013_d N_SET_B_M1013_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.78 PS=0.81 NRD=25.7873 NRS=25.7873 M=1 R=2.8
+ SA=75006.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1039 A_1665_329# N_A_1257_47#_M1039_g N_A_1431_21#_M1013_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.1638 PD=1.05 PS=1.56 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75003.4 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1043 N_VPWR_M1043_d N_A_944_21#_M1043_g A_1665_329# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2184 AS=0.0882 PD=2.2 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75003.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_RESET_B_M1001_g N_A_944_21#_M1001_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.120195 AS=0.176 PD=1.04195 PS=1.83 NRD=40.8775 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1014 N_Q_N_M1014_d N_A_1431_21#_M1014_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.187805 PD=1.27 PS=1.62805 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1030 N_Q_N_M1014_d N_A_1431_21#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.3 PD=1.27 PS=2.6 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1026_d N_A_1431_21#_M1026_g N_A_2236_47#_M1026_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1026_d N_A_2236_47#_M1002_g N_Q_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.181707 AS=0.135 PD=1.61585 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_2236_47#_M1010_g N_Q_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX44_noxref VNB VPB NWDIODE A=21.2823 P=29.73
c_262 VPB 0 1.15981e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__dfbbn_2.pxi.spice"
*
.ends
*
*

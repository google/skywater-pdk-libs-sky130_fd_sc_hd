* File: sky130_fd_sc_hd__mux2_1.pxi.spice
* Created: Tue Sep  1 19:14:18 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2_1%A_76_199# N_A_76_199#_M1005_d N_A_76_199#_M1001_d
+ N_A_76_199#_M1010_g N_A_76_199#_M1007_g N_A_76_199#_c_80_n N_A_76_199#_c_141_p
+ N_A_76_199#_c_81_n N_A_76_199#_c_97_p N_A_76_199#_c_100_p N_A_76_199#_c_82_n
+ N_A_76_199#_c_83_n N_A_76_199#_c_84_n N_A_76_199#_c_93_p N_A_76_199#_c_85_n
+ PM_SKY130_FD_SC_HD__MUX2_1%A_76_199#
x_PM_SKY130_FD_SC_HD__MUX2_1%S N_S_M1004_g N_S_M1003_g N_S_M1008_g N_S_M1009_g
+ N_S_c_164_n N_S_c_165_n N_S_c_166_n N_S_c_167_n N_S_c_168_n N_S_c_159_n
+ N_S_c_160_n S S N_S_c_172_n S PM_SKY130_FD_SC_HD__MUX2_1%S
x_PM_SKY130_FD_SC_HD__MUX2_1%A1 N_A1_M1005_g N_A1_M1006_g N_A1_c_250_n
+ N_A1_c_251_n N_A1_c_255_n N_A1_c_256_n A1 A1 N_A1_c_258_n
+ PM_SKY130_FD_SC_HD__MUX2_1%A1
x_PM_SKY130_FD_SC_HD__MUX2_1%A0 N_A0_c_316_n N_A0_M1001_g N_A0_c_317_n
+ N_A0_c_318_n N_A0_M1011_g N_A0_c_313_n A0 N_A0_c_314_n N_A0_c_315_n
+ PM_SKY130_FD_SC_HD__MUX2_1%A0
x_PM_SKY130_FD_SC_HD__MUX2_1%A_505_21# N_A_505_21#_M1008_d N_A_505_21#_M1009_d
+ N_A_505_21#_M1000_g N_A_505_21#_M1002_g N_A_505_21#_c_365_n
+ N_A_505_21#_c_366_n N_A_505_21#_c_367_n N_A_505_21#_c_368_n
+ N_A_505_21#_c_372_n N_A_505_21#_c_369_n PM_SKY130_FD_SC_HD__MUX2_1%A_505_21#
x_PM_SKY130_FD_SC_HD__MUX2_1%X N_X_M1010_s N_X_M1007_s N_X_c_419_n N_X_c_422_n
+ N_X_c_420_n X X X PM_SKY130_FD_SC_HD__MUX2_1%X
x_PM_SKY130_FD_SC_HD__MUX2_1%VPWR N_VPWR_M1007_d N_VPWR_M1002_d N_VPWR_c_440_n
+ N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n VPWR N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_439_n N_VPWR_c_447_n PM_SKY130_FD_SC_HD__MUX2_1%VPWR
x_PM_SKY130_FD_SC_HD__MUX2_1%VGND N_VGND_M1010_d N_VGND_M1000_d N_VGND_c_482_n
+ N_VGND_c_483_n VGND N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n
+ N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n PM_SKY130_FD_SC_HD__MUX2_1%VGND
cc_1 VNB N_A_76_199#_c_80_n 0.0116029f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=0.74
cc_2 VNB N_A_76_199#_c_81_n 0.00447235f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=1.955
cc_3 VNB N_A_76_199#_c_82_n 0.0020543f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_4 VNB N_A_76_199#_c_83_n 0.0229624f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_5 VNB N_A_76_199#_c_84_n 9.59127e-19 $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=0.995
cc_6 VNB N_A_76_199#_c_85_n 0.0196195f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_7 VNB N_S_M1004_g 0.0298002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_S_M1008_g 0.0538388f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_9 VNB N_S_c_159_n 4.01021e-19 $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=1.16
cc_10 VNB N_S_c_160_n 0.0237569f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_11 VNB N_A1_M1005_g 0.0208507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_250_n 0.00376476f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_13 VNB N_A1_c_251_n 0.042985f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_14 VNB A1 0.00703975f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.74
cc_15 VNB N_A0_M1011_g 0.0198887f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_A0_c_313_n 0.0108468f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_17 VNB N_A0_c_314_n 0.0272106f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.995
cc_18 VNB N_A0_c_315_n 0.00762444f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=0.74
cc_19 VNB N_A_505_21#_M1000_g 0.0241214f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_A_505_21#_M1002_g 0.0125644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_505_21#_c_365_n 0.00709026f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.995
cc_22 VNB N_A_505_21#_c_366_n 0.0251039f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=2.04
cc_23 VNB N_A_505_21#_c_367_n 0.0144794f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_24 VNB N_A_505_21#_c_368_n 0.0274406f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_25 VNB N_A_505_21#_c_369_n 0.0496831f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_26 VNB N_X_c_419_n 0.00479254f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_27 VNB N_X_c_420_n 0.0216049f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.825
cc_28 VNB X 0.0169999f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.995
cc_29 VNB N_VPWR_c_439_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_30 VNB N_VGND_c_482_n 0.00281836f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_31 VNB N_VGND_c_483_n 0.00663575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_484_n 0.0151047f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.74
cc_33 VNB N_VGND_c_485_n 0.0506918f $X=-0.19 $Y=-0.24 $X2=2.235 $Y2=2.04
cc_34 VNB N_VGND_c_486_n 0.0262615f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_35 VNB N_VGND_c_487_n 0.229802f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_36 VNB N_VGND_c_488_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_489_n 0.00978572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_76_199#_M1007_g 0.0256335f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB N_A_76_199#_c_81_n 0.0101663f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.955
cc_40 VPB N_A_76_199#_c_82_n 0.00303041f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_41 VPB N_A_76_199#_c_83_n 0.00460251f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_42 VPB N_S_M1003_g 0.0415197f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_43 VPB N_S_M1008_g 0.00441351f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_S_M1009_g 0.0243612f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.995
cc_45 VPB N_S_c_164_n 0.00885822f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=0.825
cc_46 VPB N_S_c_165_n 0.0362312f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.955
cc_47 VPB N_S_c_166_n 0.00241283f $X=-0.19 $Y=1.305 $X2=1.445 $Y2=2.04
cc_48 VPB N_S_c_167_n 0.00210134f $X=-0.19 $Y=1.305 $X2=2.235 $Y2=2.04
cc_49 VPB N_S_c_168_n 0.00169114f $X=-0.19 $Y=1.305 $X2=2.235 $Y2=2.04
cc_50 VPB N_S_c_159_n 8.95108e-19 $X=-0.19 $Y=1.305 $X2=0.557 $Y2=1.16
cc_51 VPB N_S_c_160_n 0.00652915f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_52 VPB S 0.00990495f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=0.54
cc_53 VPB N_S_c_172_n 0.0302448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A1_M1006_g 0.0215074f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_55 VPB N_A1_c_250_n 0.00568866f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_56 VPB N_A1_c_255_n 0.0144573f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.825
cc_57 VPB N_A1_c_256_n 2.22344e-19 $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.995
cc_58 VPB A1 0.00125011f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.74
cc_59 VPB N_A1_c_258_n 0.0301995f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_60 VPB N_A0_c_316_n 0.0186035f $X=-0.19 $Y=1.305 $X2=1.57 $Y2=0.235
cc_61 VPB N_A0_c_317_n 0.0356569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A0_c_318_n 0.00995527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A0_c_313_n 0.019745f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_64 VPB N_A0_c_315_n 0.00291456f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=0.74
cc_65 VPB N_A_505_21#_M1002_g 0.0359247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_505_21#_c_367_n 0.0343287f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_67 VPB N_A_505_21#_c_372_n 0.0232729f $X=-0.19 $Y=1.305 $X2=1.715 $Y2=0.54
cc_68 VPB N_X_c_422_n 0.0065071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_X_c_420_n 0.00903352f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.825
cc_70 VPB X 0.0315701f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=0.74
cc_71 VPB N_VPWR_c_440_n 0.00466757f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_72 VPB N_VPWR_c_441_n 0.0109028f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.995
cc_73 VPB N_VPWR_c_442_n 0.0562811f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=0.825
cc_74 VPB N_VPWR_c_443_n 0.00324402f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.955
cc_75 VPB N_VPWR_c_444_n 0.0178188f $X=-0.19 $Y=1.305 $X2=2.235 $Y2=2.04
cc_76 VPB N_VPWR_c_445_n 0.0253104f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_77 VPB N_VPWR_c_439_n 0.0817053f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_78 VPB N_VPWR_c_447_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 N_A_76_199#_c_80_n N_S_M1004_g 0.0127256f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A_76_199#_c_81_n N_S_M1004_g 0.00169522f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_81 N_A_76_199#_c_84_n N_S_M1004_g 0.0015792f $X=0.557 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_76_199#_c_93_p N_S_M1004_g 0.00658843f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_83 N_A_76_199#_c_85_n N_S_M1004_g 0.0196985f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_76_199#_M1007_g N_S_M1003_g 0.0173935f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_76_199#_c_81_n N_S_M1003_g 0.00320692f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_86 N_A_76_199#_c_97_p N_S_M1003_g 7.01458e-19 $X=1.445 $Y=2.04 $X2=0 $Y2=0
cc_87 N_A_76_199#_M1007_g N_S_c_164_n 0.00184919f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_76_199#_c_97_p N_S_c_165_n 0.011273f $X=1.445 $Y=2.04 $X2=0 $Y2=0
cc_89 N_A_76_199#_c_100_p N_S_c_165_n 0.0635743f $X=2.235 $Y=2.04 $X2=0 $Y2=0
cc_90 N_A_76_199#_c_100_p N_S_c_168_n 0.0073193f $X=2.235 $Y=2.04 $X2=0 $Y2=0
cc_91 N_A_76_199#_c_80_n N_S_c_159_n 0.0147573f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_76_199#_c_81_n N_S_c_159_n 0.0678463f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_93 N_A_76_199#_c_82_n N_S_c_159_n 0.0199828f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_76_199#_c_83_n N_S_c_159_n 3.64005e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_76_199#_c_80_n N_S_c_160_n 0.00319573f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A_76_199#_c_81_n N_S_c_160_n 0.00495531f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_97 N_A_76_199#_c_82_n N_S_c_160_n 0.00197826f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_76_199#_c_83_n N_S_c_160_n 0.0203259f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_76_199#_c_93_p N_A1_M1005_g 0.0212849f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_100 N_A_76_199#_c_100_p N_A1_M1006_g 0.0041715f $X=2.235 $Y=2.04 $X2=0 $Y2=0
cc_101 N_A_76_199#_c_81_n N_A1_c_250_n 0.0570093f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_102 N_A_76_199#_c_93_p N_A1_c_250_n 0.0124631f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_103 N_A_76_199#_c_81_n N_A1_c_251_n 0.00809091f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_104 N_A_76_199#_c_93_p N_A1_c_251_n 0.00213394f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_105 N_A_76_199#_c_100_p N_A1_c_255_n 0.0438796f $X=2.235 $Y=2.04 $X2=0 $Y2=0
cc_106 N_A_76_199#_c_81_n N_A1_c_256_n 0.0137204f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_107 N_A_76_199#_c_100_p N_A1_c_256_n 0.0116475f $X=2.235 $Y=2.04 $X2=0 $Y2=0
cc_108 N_A_76_199#_c_100_p N_A0_c_316_n 0.0161361f $X=2.235 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_76_199#_c_100_p N_A0_c_317_n 0.0123372f $X=2.235 $Y=2.04 $X2=0 $Y2=0
cc_110 N_A_76_199#_c_81_n N_A0_c_318_n 0.00433026f $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_111 N_A_76_199#_c_93_p N_A0_M1011_g 0.00160673f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_112 N_A_76_199#_c_81_n N_A0_c_313_n 2.97582e-19 $X=1.36 $Y=1.955 $X2=0 $Y2=0
cc_113 N_A_76_199#_c_93_p N_A0_c_315_n 0.00589575f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_114 N_A_76_199#_M1007_g N_X_c_422_n 0.00322768f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_76_199#_M1007_g N_X_c_420_n 0.0040804f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_76_199#_c_82_n N_X_c_420_n 0.0243204f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_76_199#_c_83_n N_X_c_420_n 0.00753248f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_76_199#_c_84_n N_X_c_420_n 0.00882561f $X=0.557 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_76_199#_c_85_n N_X_c_420_n 0.00354074f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_76_199#_M1007_g X 0.00877631f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_76_199#_M1007_g N_VPWR_c_440_n 0.00438629f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_76_199#_c_80_n N_VPWR_c_440_n 0.00226749f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_76_199#_c_82_n N_VPWR_c_440_n 0.00756629f $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_124 N_A_76_199#_c_83_n N_VPWR_c_440_n 4.09213e-19 $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_125 N_A_76_199#_M1007_g N_VPWR_c_444_n 0.00541359f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_76_199#_M1007_g N_VPWR_c_439_n 0.0117818f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_76_199#_c_81_n A_218_374# 7.06647e-19 $X=1.36 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_128 N_A_76_199#_c_97_p A_218_374# 0.00277991f $X=1.445 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A_76_199#_c_80_n N_VGND_M1010_d 0.00473865f $X=1.27 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_76_199#_c_141_p N_VGND_M1010_d 8.75693e-19 $X=0.685 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_76_199#_c_84_n N_VGND_M1010_d 8.08664e-19 $X=0.557 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A_76_199#_c_80_n N_VGND_c_482_n 0.01222f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_76_199#_c_141_p N_VGND_c_482_n 0.00929542f $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_134 N_A_76_199#_c_83_n N_VGND_c_482_n 3.09237e-19 $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_76_199#_c_93_p N_VGND_c_482_n 0.00973513f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_136 N_A_76_199#_c_85_n N_VGND_c_482_n 0.00872433f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_A_76_199#_c_85_n N_VGND_c_484_n 0.0046653f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_76_199#_c_80_n N_VGND_c_485_n 0.00714584f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_76_199#_c_93_p N_VGND_c_485_n 0.0320721f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_140 N_A_76_199#_M1005_d N_VGND_c_487_n 0.0096734f $X=1.57 $Y=0.235 $X2=0
+ $Y2=0
cc_141 N_A_76_199#_c_80_n N_VGND_c_487_n 0.0118208f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_76_199#_c_141_p N_VGND_c_487_n 8.0899e-19 $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_76_199#_c_93_p N_VGND_c_487_n 0.019514f $X=1.36 $Y=0.54 $X2=0 $Y2=0
cc_144 N_A_76_199#_c_85_n N_VGND_c_487_n 0.00895857f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_76_199#_c_93_p A_218_47# 0.00606386f $X=1.36 $Y=0.54 $X2=-0.19
+ $Y2=-0.24
cc_146 N_S_M1004_g N_A1_M1005_g 0.0309752f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_147 N_S_c_165_n N_A1_M1006_g 0.0127926f $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_148 N_S_c_160_n N_A1_c_251_n 0.00605477f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_149 N_S_c_165_n N_A1_c_255_n 0.00783263f $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_150 N_S_c_167_n N_A1_c_255_n 0.00133723f $X=2.88 $Y=1.63 $X2=0 $Y2=0
cc_151 N_S_c_168_n N_A1_c_255_n 0.0123063f $X=2.88 $Y=2.295 $X2=0 $Y2=0
cc_152 N_S_c_167_n A1 0.0141868f $X=2.88 $Y=1.63 $X2=0 $Y2=0
cc_153 N_S_c_165_n N_A1_c_258_n 5.84442e-19 $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_154 N_S_c_167_n N_A1_c_258_n 0.00125929f $X=2.88 $Y=1.63 $X2=0 $Y2=0
cc_155 N_S_c_168_n N_A1_c_258_n 0.00939374f $X=2.88 $Y=2.295 $X2=0 $Y2=0
cc_156 N_S_c_164_n N_A0_c_316_n 9.1133e-19 $X=1.02 $Y=2.295 $X2=-0.19 $Y2=-0.24
cc_157 N_S_c_165_n N_A0_c_316_n 0.0108033f $X=2.795 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_158 N_S_M1003_g N_A0_c_318_n 0.0233336f $X=1.015 $Y=2.08 $X2=0 $Y2=0
cc_159 N_S_M1008_g N_A_505_21#_M1000_g 0.00837678f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_160 N_S_M1008_g N_A_505_21#_M1002_g 0.0106395f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_161 N_S_M1009_g N_A_505_21#_M1002_g 0.0106308f $X=3.44 $Y=2.08 $X2=0 $Y2=0
cc_162 N_S_c_165_n N_A_505_21#_M1002_g 0.00406273f $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_163 N_S_c_167_n N_A_505_21#_M1002_g 0.00399688f $X=2.88 $Y=1.63 $X2=0 $Y2=0
cc_164 N_S_c_168_n N_A_505_21#_M1002_g 0.0137565f $X=2.88 $Y=2.295 $X2=0 $Y2=0
cc_165 S N_A_505_21#_M1002_g 0.00746073f $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_166 N_S_c_172_n N_A_505_21#_M1002_g 0.0210687f $X=3.38 $Y=1.545 $X2=0 $Y2=0
cc_167 N_S_M1008_g N_A_505_21#_c_365_n 0.0175175f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_168 N_S_c_167_n N_A_505_21#_c_365_n 0.00591184f $X=2.88 $Y=1.63 $X2=0 $Y2=0
cc_169 S N_A_505_21#_c_365_n 0.0223708f $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_170 N_S_c_172_n N_A_505_21#_c_365_n 0.00248698f $X=3.38 $Y=1.545 $X2=0 $Y2=0
cc_171 N_S_M1008_g N_A_505_21#_c_366_n 0.0101674f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_172 N_S_M1008_g N_A_505_21#_c_367_n 0.0136619f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_173 S N_A_505_21#_c_367_n 0.0166636f $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_174 N_S_c_172_n N_A_505_21#_c_367_n 0.0102485f $X=3.38 $Y=1.545 $X2=0 $Y2=0
cc_175 S N_A_505_21#_c_368_n 4.91502e-19 $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_176 N_S_M1008_g N_A_505_21#_c_369_n 0.0178169f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_177 N_S_c_167_n N_A_505_21#_c_369_n 0.00218549f $X=2.88 $Y=1.63 $X2=0 $Y2=0
cc_178 S N_A_505_21#_c_369_n 0.00237629f $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_179 N_S_c_164_n N_X_c_420_n 0.00478262f $X=1.02 $Y=2.295 $X2=0 $Y2=0
cc_180 N_S_M1003_g N_VPWR_c_440_n 0.00321158f $X=1.015 $Y=2.08 $X2=0 $Y2=0
cc_181 N_S_c_164_n N_VPWR_c_440_n 0.0432455f $X=1.02 $Y=2.295 $X2=0 $Y2=0
cc_182 N_S_c_166_n N_VPWR_c_440_n 0.0141313f $X=1.105 $Y=2.38 $X2=0 $Y2=0
cc_183 N_S_M1009_g N_VPWR_c_441_n 0.00506507f $X=3.44 $Y=2.08 $X2=0 $Y2=0
cc_184 N_S_c_165_n N_VPWR_c_441_n 0.0137894f $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_185 N_S_c_168_n N_VPWR_c_441_n 0.0294585f $X=2.88 $Y=2.295 $X2=0 $Y2=0
cc_186 S N_VPWR_c_441_n 0.010519f $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_187 N_S_c_172_n N_VPWR_c_441_n 0.00145494f $X=3.38 $Y=1.545 $X2=0 $Y2=0
cc_188 N_S_M1003_g N_VPWR_c_442_n 8.50093e-19 $X=1.015 $Y=2.08 $X2=0 $Y2=0
cc_189 N_S_c_165_n N_VPWR_c_442_n 0.121009f $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_190 N_S_c_166_n N_VPWR_c_442_n 0.0121882f $X=1.105 $Y=2.38 $X2=0 $Y2=0
cc_191 N_S_M1009_g N_VPWR_c_445_n 0.00534427f $X=3.44 $Y=2.08 $X2=0 $Y2=0
cc_192 N_S_M1009_g N_VPWR_c_439_n 0.00523659f $X=3.44 $Y=2.08 $X2=0 $Y2=0
cc_193 N_S_c_165_n N_VPWR_c_439_n 0.0694838f $X=2.795 $Y=2.38 $X2=0 $Y2=0
cc_194 N_S_c_166_n N_VPWR_c_439_n 0.006547f $X=1.105 $Y=2.38 $X2=0 $Y2=0
cc_195 N_S_c_168_n A_535_374# 0.00479825f $X=2.88 $Y=2.295 $X2=-0.19 $Y2=-0.24
cc_196 N_S_M1004_g N_VGND_c_482_n 0.00601017f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_197 N_S_M1008_g N_VGND_c_483_n 0.00375687f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_198 N_S_M1004_g N_VGND_c_485_n 0.00428022f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_199 N_S_M1008_g N_VGND_c_486_n 0.00585385f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_200 N_S_M1004_g N_VGND_c_487_n 0.00640514f $X=1.015 $Y=0.445 $X2=0 $Y2=0
cc_201 N_S_M1008_g N_VGND_c_487_n 0.0126275f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A1_M1006_g N_A0_c_317_n 0.00317917f $X=2.6 $Y=2.08 $X2=0 $Y2=0
cc_203 N_A1_c_255_n N_A0_c_317_n 0.012453f $X=2.435 $Y=1.7 $X2=0 $Y2=0
cc_204 N_A1_c_256_n N_A0_c_317_n 0.00733132f $X=1.785 $Y=1.7 $X2=0 $Y2=0
cc_205 N_A1_c_251_n N_A0_c_318_n 0.0102256f $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_206 N_A1_M1005_g N_A0_M1011_g 0.0116149f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_207 A1 N_A0_M1011_g 0.00158356f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_208 N_A1_c_250_n N_A0_c_313_n 0.00586297f $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_209 N_A1_c_255_n N_A0_c_313_n 0.00348659f $X=2.435 $Y=1.7 $X2=0 $Y2=0
cc_210 A1 N_A0_c_313_n 0.0016247f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_211 N_A1_c_258_n N_A0_c_313_n 0.0204691f $X=2.54 $Y=1.545 $X2=0 $Y2=0
cc_212 N_A1_c_250_n N_A0_c_314_n 3.49151e-19 $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_213 N_A1_c_251_n N_A0_c_314_n 0.0209106f $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_214 N_A1_c_255_n N_A0_c_314_n 0.00166378f $X=2.435 $Y=1.7 $X2=0 $Y2=0
cc_215 A1 N_A0_c_314_n 0.00247923f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_216 N_A1_M1005_g N_A0_c_315_n 0.00124204f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A1_c_250_n N_A0_c_315_n 0.0398419f $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_218 N_A1_c_251_n N_A0_c_315_n 0.00209255f $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_219 N_A1_c_255_n N_A0_c_315_n 0.0192865f $X=2.435 $Y=1.7 $X2=0 $Y2=0
cc_220 A1 N_A0_c_315_n 0.0887943f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_221 N_A1_c_258_n N_A0_c_315_n 2.00408e-19 $X=2.54 $Y=1.545 $X2=0 $Y2=0
cc_222 A1 N_A_505_21#_M1000_g 0.0211682f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_223 A1 N_A_505_21#_M1002_g 0.00637504f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_224 N_A1_c_258_n N_A_505_21#_M1002_g 0.0625034f $X=2.54 $Y=1.545 $X2=0 $Y2=0
cc_225 A1 N_A_505_21#_c_365_n 0.0115821f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_226 A1 N_A_505_21#_c_369_n 0.00863073f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_227 N_A1_c_258_n N_A_505_21#_c_369_n 0.00540744f $X=2.54 $Y=1.545 $X2=0 $Y2=0
cc_228 N_A1_M1006_g N_VPWR_c_442_n 8.51345e-19 $X=2.6 $Y=2.08 $X2=0 $Y2=0
cc_229 A1 N_VGND_c_483_n 0.0269885f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_230 N_A1_M1005_g N_VGND_c_485_n 0.00357668f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_231 A1 N_VGND_c_485_n 0.0110225f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_232 N_A1_M1005_g N_VGND_c_487_n 0.00590596f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_233 N_A1_c_251_n N_VGND_c_487_n 8.00495e-19 $X=1.7 $Y=0.98 $X2=0 $Y2=0
cc_234 A1 N_VGND_c_487_n 0.00678747f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_235 A1 A_439_47# 0.00375979f $X=2.45 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_236 N_A0_M1011_g N_A_505_21#_M1000_g 0.0265912f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A0_c_314_n N_A_505_21#_M1000_g 0.0110099f $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_238 N_A0_c_315_n N_A_505_21#_M1000_g 0.00177736f $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_239 N_A0_c_313_n N_A_505_21#_M1002_g 0.0022574f $X=2.12 $Y=1.645 $X2=0 $Y2=0
cc_240 N_A0_c_314_n N_A_505_21#_M1002_g 3.79555e-19 $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_241 N_A0_c_314_n N_A_505_21#_c_369_n 0.00200073f $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_242 N_A0_c_316_n N_VPWR_c_442_n 8.51345e-19 $X=1.53 $Y=1.795 $X2=0 $Y2=0
cc_243 N_A0_M1011_g N_VGND_c_485_n 0.00357668f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_244 N_A0_c_315_n N_VGND_c_485_n 0.0150093f $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_245 N_A0_M1011_g N_VGND_c_487_n 0.00590596f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_246 N_A0_c_314_n N_VGND_c_487_n 0.00116644f $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_247 N_A0_c_315_n N_VGND_c_487_n 0.00982774f $X=2.18 $Y=0.98 $X2=0 $Y2=0
cc_248 N_A0_c_315_n A_439_47# 0.00363136f $X=2.18 $Y=0.98 $X2=-0.19 $Y2=-0.24
cc_249 N_A_505_21#_M1002_g N_VPWR_c_441_n 0.00219666f $X=2.96 $Y=2.08 $X2=0
+ $Y2=0
cc_250 N_A_505_21#_M1002_g N_VPWR_c_442_n 0.00294738f $X=2.96 $Y=2.08 $X2=0
+ $Y2=0
cc_251 N_A_505_21#_c_372_n N_VPWR_c_445_n 0.0157581f $X=3.885 $Y=2.08 $X2=0
+ $Y2=0
cc_252 N_A_505_21#_M1002_g N_VPWR_c_439_n 0.00244374f $X=2.96 $Y=2.08 $X2=0
+ $Y2=0
cc_253 N_A_505_21#_c_372_n N_VPWR_c_439_n 0.017495f $X=3.885 $Y=2.08 $X2=0 $Y2=0
cc_254 N_A_505_21#_M1000_g N_VGND_c_483_n 0.00752592f $X=2.6 $Y=0.445 $X2=0
+ $Y2=0
cc_255 N_A_505_21#_c_365_n N_VGND_c_483_n 0.0272033f $X=3.535 $Y=0.98 $X2=0
+ $Y2=0
cc_256 N_A_505_21#_c_369_n N_VGND_c_483_n 0.00883154f $X=2.96 $Y=0.98 $X2=0
+ $Y2=0
cc_257 N_A_505_21#_M1000_g N_VGND_c_485_n 0.00435091f $X=2.6 $Y=0.445 $X2=0
+ $Y2=0
cc_258 N_A_505_21#_c_366_n N_VGND_c_486_n 0.0129431f $X=3.65 $Y=0.455 $X2=0
+ $Y2=0
cc_259 N_A_505_21#_M1008_d N_VGND_c_487_n 0.0028471f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_260 N_A_505_21#_M1000_g N_VGND_c_487_n 0.00810682f $X=2.6 $Y=0.445 $X2=0
+ $Y2=0
cc_261 N_A_505_21#_c_366_n N_VGND_c_487_n 0.00919761f $X=3.65 $Y=0.455 $X2=0
+ $Y2=0
cc_262 N_A_505_21#_c_369_n N_VGND_c_487_n 0.00264476f $X=2.96 $Y=0.98 $X2=0
+ $Y2=0
cc_263 X N_VPWR_c_444_n 0.0213966f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_264 N_X_M1007_s N_VPWR_c_439_n 0.00209319f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_265 X N_VPWR_c_439_n 0.0126193f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_266 X N_VGND_c_484_n 0.0175724f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_267 N_X_M1010_s N_VGND_c_487_n 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_268 X N_VGND_c_487_n 0.00972866f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_269 N_VGND_c_487_n A_218_47# 0.00335872f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_270 N_VGND_c_487_n A_439_47# 0.00746861f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

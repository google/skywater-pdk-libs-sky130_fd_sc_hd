* File: sky130_fd_sc_hd__ebufn_4.pxi.spice
* Created: Tue Sep  1 19:07:19 2020
* 
x_PM_SKY130_FD_SC_HD__EBUFN_4%A N_A_M1018_g N_A_M1013_g A A N_A_c_101_n
+ N_A_c_102_n PM_SKY130_FD_SC_HD__EBUFN_4%A
x_PM_SKY130_FD_SC_HD__EBUFN_4%TE_B N_TE_B_M1014_g N_TE_B_c_136_n N_TE_B_M1002_g
+ N_TE_B_c_137_n N_TE_B_c_134_n N_TE_B_c_139_n N_TE_B_M1000_g N_TE_B_c_140_n
+ N_TE_B_c_141_n N_TE_B_M1011_g N_TE_B_c_142_n N_TE_B_c_143_n N_TE_B_M1016_g
+ N_TE_B_c_144_n N_TE_B_c_145_n N_TE_B_M1019_g N_TE_B_c_146_n N_TE_B_c_147_n
+ N_TE_B_c_148_n TE_B PM_SKY130_FD_SC_HD__EBUFN_4%TE_B
x_PM_SKY130_FD_SC_HD__EBUFN_4%A_214_47# N_A_214_47#_M1014_d N_A_214_47#_M1002_d
+ N_A_214_47#_c_217_n N_A_214_47#_M1003_g N_A_214_47#_c_218_n
+ N_A_214_47#_c_219_n N_A_214_47#_c_220_n N_A_214_47#_M1004_g
+ N_A_214_47#_c_221_n N_A_214_47#_c_222_n N_A_214_47#_M1005_g
+ N_A_214_47#_c_223_n N_A_214_47#_M1006_g N_A_214_47#_c_224_n
+ N_A_214_47#_c_225_n N_A_214_47#_c_226_n N_A_214_47#_c_233_n
+ N_A_214_47#_c_227_n N_A_214_47#_c_228_n N_A_214_47#_c_229_n
+ N_A_214_47#_c_230_n N_A_214_47#_c_231_n N_A_214_47#_c_232_n
+ PM_SKY130_FD_SC_HD__EBUFN_4%A_214_47#
x_PM_SKY130_FD_SC_HD__EBUFN_4%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1013_s
+ N_A_27_47#_M1007_g N_A_27_47#_M1001_g N_A_27_47#_M1008_g N_A_27_47#_M1009_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1012_g N_A_27_47#_M1015_g N_A_27_47#_M1017_g
+ N_A_27_47#_c_329_n N_A_27_47#_c_330_n N_A_27_47#_c_319_n N_A_27_47#_c_320_n
+ N_A_27_47#_c_321_n N_A_27_47#_c_322_n N_A_27_47#_c_333_n N_A_27_47#_c_323_n
+ N_A_27_47#_c_324_n PM_SKY130_FD_SC_HD__EBUFN_4%A_27_47#
x_PM_SKY130_FD_SC_HD__EBUFN_4%VPWR N_VPWR_M1013_d N_VPWR_M1000_d N_VPWR_M1016_d
+ N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n VPWR N_VPWR_c_414_n
+ N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_410_n N_VPWR_c_419_n
+ N_VPWR_c_420_n N_VPWR_c_421_n PM_SKY130_FD_SC_HD__EBUFN_4%VPWR
x_PM_SKY130_FD_SC_HD__EBUFN_4%A_320_309# N_A_320_309#_M1000_s
+ N_A_320_309#_M1011_s N_A_320_309#_M1019_s N_A_320_309#_M1009_d
+ N_A_320_309#_M1017_d N_A_320_309#_c_485_n N_A_320_309#_c_512_n
+ N_A_320_309#_c_486_n N_A_320_309#_c_519_n N_A_320_309#_c_487_n
+ N_A_320_309#_c_493_n PM_SKY130_FD_SC_HD__EBUFN_4%A_320_309#
x_PM_SKY130_FD_SC_HD__EBUFN_4%Z N_Z_M1007_d N_Z_M1010_d N_Z_M1001_s N_Z_M1012_s
+ N_Z_c_556_n Z Z Z Z Z Z Z Z Z Z N_Z_c_540_n N_Z_c_537_n
+ PM_SKY130_FD_SC_HD__EBUFN_4%Z
x_PM_SKY130_FD_SC_HD__EBUFN_4%VGND N_VGND_M1018_d N_VGND_M1003_d N_VGND_M1005_d
+ N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n VGND N_VGND_c_605_n
+ N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n N_VGND_c_609_n N_VGND_c_610_n
+ N_VGND_c_611_n N_VGND_c_612_n PM_SKY130_FD_SC_HD__EBUFN_4%VGND
x_PM_SKY130_FD_SC_HD__EBUFN_4%A_393_47# N_A_393_47#_M1003_s N_A_393_47#_M1004_s
+ N_A_393_47#_M1006_s N_A_393_47#_M1008_s N_A_393_47#_M1015_s
+ N_A_393_47#_c_681_n N_A_393_47#_c_686_n N_A_393_47#_c_682_n
+ N_A_393_47#_c_729_n N_A_393_47#_c_692_n N_A_393_47#_c_736_n
+ N_A_393_47#_c_683_n N_A_393_47#_c_697_n PM_SKY130_FD_SC_HD__EBUFN_4%A_393_47#
cc_1 VNB A 0.00215563f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_2 VNB N_A_c_101_n 0.0269023f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_3 VNB N_A_c_102_n 0.019414f $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=0.995
cc_4 VNB N_TE_B_M1014_g 0.0226981f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_5 VNB N_TE_B_c_134_n 0.0406042f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_6 VNB TE_B 0.00130093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_214_47#_c_217_n 0.0175571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_214_47#_c_218_n 0.00893548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_214_47#_c_219_n 0.00846217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_214_47#_c_220_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.16
cc_11 VNB N_A_214_47#_c_221_n 0.00893472f $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=0.995
cc_12 VNB N_A_214_47#_c_222_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.85
cc_13 VNB N_A_214_47#_c_223_n 0.0126529f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_14 VNB N_A_214_47#_c_224_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_214_47#_c_225_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_214_47#_c_226_n 0.0111771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_214_47#_c_227_n 0.0122386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_214_47#_c_228_n 0.00105691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_214_47#_c_229_n 0.0236972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_214_47#_c_230_n 0.00159906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_214_47#_c_231_n 0.0338621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_214_47#_c_232_n 0.0150954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1007_g 0.0185496f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_24 VNB N_A_27_47#_M1001_g 7.20477e-19 $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_25 VNB N_A_27_47#_M1008_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.85
cc_26 VNB N_A_27_47#_M1009_g 4.13757e-19 $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.53
cc_27 VNB N_A_27_47#_M1010_g 0.0175045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_M1012_g 4.5009e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_M1015_g 0.0210785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_M1017_g 5.06554e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_319_n 0.0150059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_320_n 0.00828112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_321_n 0.0113098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_322_n 0.023363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_323_n 0.00588605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_324_n 0.0646544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_410_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB Z 0.0228337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Z_c_537_n 0.0136094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_602_n 5.72709e-19 $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.16
cc_41 VNB N_VGND_c_603_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.325
cc_42 VNB N_VGND_c_604_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_43 VNB N_VGND_c_605_n 0.0151734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_606_n 0.0336478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_607_n 0.0110833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_608_n 0.0582981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_609_n 0.307493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_610_n 0.00558939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_611_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_612_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_393_47#_c_681_n 0.00521061f $X=-0.19 $Y=-0.24 $X2=0.552 $Y2=1.325
cc_52 VNB N_A_393_47#_c_682_n 0.00281657f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_53 VNB N_A_393_47#_c_683_n 0.00812227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VPB N_A_M1013_g 0.0221199f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_55 VPB A 0.00131181f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_56 VPB N_A_c_101_n 0.00605063f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_57 VPB N_TE_B_c_136_n 0.0179427f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_58 VPB N_TE_B_c_137_n 0.0180786f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_59 VPB N_TE_B_c_134_n 0.0265907f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_60 VPB N_TE_B_c_139_n 0.0167523f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_TE_B_c_140_n 0.0127572f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_62 VPB N_TE_B_c_141_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0.552 $Y2=0.995
cc_63 VPB N_TE_B_c_142_n 0.0113042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_TE_B_c_143_n 0.0133656f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_65 VPB N_TE_B_c_144_n 0.0238745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_TE_B_c_145_n 0.0172196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_TE_B_c_146_n 0.00612638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_TE_B_c_147_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_TE_B_c_148_n 0.0049211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB TE_B 0.00297755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_214_47#_c_233_n 0.00715433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_214_47#_c_228_n 0.0123134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_M1001_g 0.0267252f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_74 VPB N_A_27_47#_M1009_g 0.0191885f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.53
cc_75 VPB N_A_27_47#_M1012_g 0.01917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_M1017_g 0.0233497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_329_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_330_n 0.0219831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_321_n 0.00158633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_322_n 0.0194644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_333_n 0.00136192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_411_n 5.72709e-19 $X=-0.19 $Y=1.305 $X2=0.552 $Y2=1.16
cc_83 VPB N_VPWR_c_412_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.552 $Y2=1.325
cc_84 VPB N_VPWR_c_413_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_85 VPB N_VPWR_c_414_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_415_n 0.0260256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_416_n 0.0111333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_417_n 0.0656674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_410_n 0.0550152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_419_n 0.00558939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_420_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_421_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_320_309#_c_485_n 0.0034618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_320_309#_c_486_n 0.00179358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_320_309#_c_487_n 0.0298921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB Z 0.00750198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB Z 0.0150079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Z_c_540_n 0.0148687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 A N_TE_B_M1014_g 0.00729568f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A_c_101_n N_TE_B_M1014_g 0.0215008f $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_c_102_n N_TE_B_M1014_g 0.0220615f $X=0.552 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_M1013_g N_TE_B_c_134_n 0.0280837f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_103 A TE_B 0.049885f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A_c_101_n TE_B 4.16903e-19 $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_c_102_n TE_B 2.00312e-19 $X=0.552 $Y=0.995 $X2=0 $Y2=0
cc_106 A N_A_214_47#_c_228_n 0.00489798f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_107 A N_A_27_47#_c_320_n 0.0194626f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_108 N_A_c_101_n N_A_27_47#_c_320_n 0.00964443f $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_109 A N_A_27_47#_c_321_n 0.00274795f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_110 N_A_c_101_n N_A_27_47#_c_321_n 0.00262964f $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_111 A N_A_27_47#_c_322_n 0.0667582f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_112 N_A_c_102_n N_A_27_47#_c_322_n 0.0274299f $X=0.552 $Y=0.995 $X2=0 $Y2=0
cc_113 A N_VPWR_M1013_d 0.00489945f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_114 N_A_M1013_g N_VPWR_c_411_n 0.0132693f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_115 A N_VPWR_c_411_n 0.0179123f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_116 N_A_c_101_n N_VPWR_c_411_n 5.35719e-19 $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_M1013_g N_VPWR_c_414_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_M1013_g N_VPWR_c_410_n 0.008846f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_119 A N_VGND_M1018_d 0.00304146f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_120 A N_VGND_c_602_n 0.0172572f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_121 N_A_c_101_n N_VGND_c_602_n 6.62542e-19 $X=0.575 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_102_n N_VGND_c_602_n 0.0116256f $X=0.552 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_102_n N_VGND_c_605_n 0.0046653f $X=0.552 $Y=0.995 $X2=0 $Y2=0
cc_124 A N_VGND_c_609_n 0.00190664f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_125 N_A_c_102_n N_VGND_c_609_n 0.00818925f $X=0.552 $Y=0.995 $X2=0 $Y2=0
cc_126 TE_B N_A_214_47#_M1014_d 0.0030848f $X=1.07 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_127 N_TE_B_c_147_n N_A_214_47#_c_218_n 0.0133811f $X=2.355 $Y=1.395 $X2=0
+ $Y2=0
cc_128 N_TE_B_c_140_n N_A_214_47#_c_219_n 0.0133811f $X=2.28 $Y=1.395 $X2=0
+ $Y2=0
cc_129 N_TE_B_c_148_n N_A_214_47#_c_221_n 0.0133811f $X=2.775 $Y=1.395 $X2=0
+ $Y2=0
cc_130 N_TE_B_c_142_n N_A_214_47#_c_224_n 0.0133811f $X=2.7 $Y=1.395 $X2=0 $Y2=0
cc_131 N_TE_B_c_144_n N_A_214_47#_c_225_n 0.0133811f $X=3.12 $Y=1.395 $X2=0
+ $Y2=0
cc_132 N_TE_B_c_134_n N_A_214_47#_c_226_n 0.00398079f $X=1.595 $Y=1.395 $X2=0
+ $Y2=0
cc_133 TE_B N_A_214_47#_c_226_n 0.0121175f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_134 N_TE_B_c_139_n N_A_214_47#_c_233_n 0.00457052f $X=1.935 $Y=1.47 $X2=0
+ $Y2=0
cc_135 N_TE_B_M1014_g N_A_214_47#_c_227_n 0.00569329f $X=0.995 $Y=0.56 $X2=0
+ $Y2=0
cc_136 TE_B N_A_214_47#_c_227_n 0.0211308f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_137 N_TE_B_c_136_n N_A_214_47#_c_228_n 0.00255621f $X=0.995 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_TE_B_c_137_n N_A_214_47#_c_228_n 0.0132701f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_134_n N_A_214_47#_c_228_n 0.0172417f $X=1.595 $Y=1.395 $X2=0
+ $Y2=0
cc_140 N_TE_B_c_139_n N_A_214_47#_c_228_n 0.00683098f $X=1.935 $Y=1.47 $X2=0
+ $Y2=0
cc_141 TE_B N_A_214_47#_c_228_n 0.0243073f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_142 N_TE_B_c_137_n N_A_214_47#_c_229_n 0.022517f $X=1.86 $Y=1.395 $X2=0 $Y2=0
cc_143 N_TE_B_c_134_n N_A_214_47#_c_230_n 0.00912967f $X=1.595 $Y=1.395 $X2=0
+ $Y2=0
cc_144 TE_B N_A_214_47#_c_230_n 0.0189956f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_145 N_TE_B_c_134_n N_A_27_47#_c_320_n 0.00906049f $X=1.595 $Y=1.395 $X2=0
+ $Y2=0
cc_146 TE_B N_A_27_47#_c_320_n 0.0271555f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_147 N_TE_B_c_136_n N_VPWR_c_411_n 0.021108f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_148 N_TE_B_c_139_n N_VPWR_c_412_n 0.00812573f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_149 N_TE_B_c_141_n N_VPWR_c_412_n 0.00643377f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_150 N_TE_B_c_143_n N_VPWR_c_412_n 5.02907e-19 $X=2.775 $Y=1.47 $X2=0 $Y2=0
cc_151 N_TE_B_c_141_n N_VPWR_c_413_n 5.02907e-19 $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_152 N_TE_B_c_143_n N_VPWR_c_413_n 0.00643498f $X=2.775 $Y=1.47 $X2=0 $Y2=0
cc_153 N_TE_B_c_145_n N_VPWR_c_413_n 0.00815483f $X=3.195 $Y=1.47 $X2=0 $Y2=0
cc_154 N_TE_B_c_136_n N_VPWR_c_415_n 0.00544582f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_155 N_TE_B_c_139_n N_VPWR_c_415_n 0.00336882f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_156 N_TE_B_c_141_n N_VPWR_c_416_n 0.00336882f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_157 N_TE_B_c_143_n N_VPWR_c_416_n 0.00337001f $X=2.775 $Y=1.47 $X2=0 $Y2=0
cc_158 N_TE_B_c_145_n N_VPWR_c_417_n 0.00337001f $X=3.195 $Y=1.47 $X2=0 $Y2=0
cc_159 N_TE_B_c_136_n N_VPWR_c_410_n 0.0104464f $X=0.995 $Y=1.41 $X2=0 $Y2=0
cc_160 N_TE_B_c_139_n N_VPWR_c_410_n 0.00522984f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_161 N_TE_B_c_141_n N_VPWR_c_410_n 0.00390377f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_162 N_TE_B_c_143_n N_VPWR_c_410_n 0.00390568f $X=2.775 $Y=1.47 $X2=0 $Y2=0
cc_163 N_TE_B_c_145_n N_VPWR_c_410_n 0.0053254f $X=3.195 $Y=1.47 $X2=0 $Y2=0
cc_164 N_TE_B_c_137_n N_A_320_309#_c_486_n 0.0021044f $X=1.86 $Y=1.395 $X2=0
+ $Y2=0
cc_165 N_TE_B_c_139_n N_A_320_309#_c_486_n 0.014832f $X=1.935 $Y=1.47 $X2=0
+ $Y2=0
cc_166 N_TE_B_c_140_n N_A_320_309#_c_486_n 3.68533e-19 $X=2.28 $Y=1.395 $X2=0
+ $Y2=0
cc_167 N_TE_B_c_141_n N_A_320_309#_c_486_n 0.0128906f $X=2.355 $Y=1.47 $X2=0
+ $Y2=0
cc_168 N_TE_B_c_142_n N_A_320_309#_c_486_n 4.01342e-19 $X=2.7 $Y=1.395 $X2=0
+ $Y2=0
cc_169 N_TE_B_c_143_n N_A_320_309#_c_493_n 0.012893f $X=2.775 $Y=1.47 $X2=0
+ $Y2=0
cc_170 N_TE_B_c_144_n N_A_320_309#_c_493_n 3.68277e-19 $X=3.12 $Y=1.395 $X2=0
+ $Y2=0
cc_171 N_TE_B_c_145_n N_A_320_309#_c_493_n 0.0154967f $X=3.195 $Y=1.47 $X2=0
+ $Y2=0
cc_172 N_TE_B_c_139_n N_Z_c_540_n 0.00874586f $X=1.935 $Y=1.47 $X2=0 $Y2=0
cc_173 N_TE_B_c_140_n N_Z_c_540_n 0.00450614f $X=2.28 $Y=1.395 $X2=0 $Y2=0
cc_174 N_TE_B_c_141_n N_Z_c_540_n 0.0115096f $X=2.355 $Y=1.47 $X2=0 $Y2=0
cc_175 N_TE_B_c_142_n N_Z_c_540_n 0.0043665f $X=2.7 $Y=1.395 $X2=0 $Y2=0
cc_176 N_TE_B_c_143_n N_Z_c_540_n 0.0115275f $X=2.775 $Y=1.47 $X2=0 $Y2=0
cc_177 N_TE_B_c_144_n N_Z_c_540_n 0.00643784f $X=3.12 $Y=1.395 $X2=0 $Y2=0
cc_178 N_TE_B_c_145_n N_Z_c_540_n 0.0146945f $X=3.195 $Y=1.47 $X2=0 $Y2=0
cc_179 N_TE_B_c_146_n N_Z_c_540_n 0.00154844f $X=1.935 $Y=1.395 $X2=0 $Y2=0
cc_180 N_TE_B_c_147_n N_Z_c_540_n 0.00146804f $X=2.355 $Y=1.395 $X2=0 $Y2=0
cc_181 N_TE_B_c_148_n N_Z_c_540_n 0.00146804f $X=2.775 $Y=1.395 $X2=0 $Y2=0
cc_182 N_TE_B_M1014_g N_VGND_c_602_n 0.0142944f $X=0.995 $Y=0.56 $X2=0 $Y2=0
cc_183 N_TE_B_M1014_g N_VGND_c_606_n 0.00544582f $X=0.995 $Y=0.56 $X2=0 $Y2=0
cc_184 N_TE_B_M1014_g N_VGND_c_609_n 0.00681521f $X=0.995 $Y=0.56 $X2=0 $Y2=0
cc_185 TE_B N_VGND_c_609_n 0.005623f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_186 N_A_214_47#_c_231_n N_A_27_47#_M1007_g 0.0221173f $X=3.645 $Y=1.035 $X2=0
+ $Y2=0
cc_187 N_A_214_47#_c_232_n N_A_27_47#_M1007_g 0.0143373f $X=3.645 $Y=0.96 $X2=0
+ $Y2=0
cc_188 N_A_214_47#_c_226_n N_A_27_47#_c_320_n 0.00655698f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_189 N_A_214_47#_c_228_n N_A_27_47#_c_320_n 0.00778923f $X=1.587 $Y=1.595
+ $X2=0 $Y2=0
cc_190 N_A_214_47#_c_229_n N_A_27_47#_c_320_n 0.0890663f $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_214_47#_c_230_n N_A_27_47#_c_320_n 0.0291445f $X=1.587 $Y=1.15 $X2=0
+ $Y2=0
cc_192 N_A_214_47#_c_231_n N_A_27_47#_c_320_n 7.09467e-19 $X=3.645 $Y=1.035
+ $X2=0 $Y2=0
cc_193 N_A_214_47#_c_229_n N_A_27_47#_c_333_n 2.5595e-19 $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_194 N_A_214_47#_c_229_n N_A_27_47#_c_323_n 0.0192917f $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_214_47#_c_231_n N_A_27_47#_c_323_n 8.01321e-19 $X=3.645 $Y=1.035
+ $X2=0 $Y2=0
cc_196 N_A_214_47#_c_229_n N_A_27_47#_c_324_n 3.70419e-19 $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_197 N_A_214_47#_c_233_n N_VPWR_c_415_n 0.0169526f $X=1.205 $Y=1.96 $X2=0
+ $Y2=0
cc_198 N_A_214_47#_M1002_d N_VPWR_c_410_n 0.00313466f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_A_214_47#_c_233_n N_VPWR_c_410_n 0.00975095f $X=1.205 $Y=1.96 $X2=0
+ $Y2=0
cc_200 N_A_214_47#_c_228_n N_A_320_309#_M1000_s 0.00472796f $X=1.587 $Y=1.595
+ $X2=-0.19 $Y2=-0.24
cc_201 N_A_214_47#_c_233_n N_A_320_309#_c_485_n 0.0247516f $X=1.205 $Y=1.96
+ $X2=0 $Y2=0
cc_202 N_A_214_47#_c_233_n N_A_320_309#_c_486_n 0.0140932f $X=1.205 $Y=1.96
+ $X2=0 $Y2=0
cc_203 N_A_214_47#_c_228_n N_A_320_309#_c_486_n 0.0128275f $X=1.587 $Y=1.595
+ $X2=0 $Y2=0
cc_204 N_A_214_47#_c_229_n N_A_320_309#_c_486_n 0.00415949f $X=3.645 $Y=1.16
+ $X2=0 $Y2=0
cc_205 N_A_214_47#_c_219_n N_Z_c_540_n 7.87147e-19 $X=2.375 $Y=1.035 $X2=0 $Y2=0
cc_206 N_A_214_47#_c_223_n N_Z_c_540_n 0.00103061f $X=3.48 $Y=1.035 $X2=0 $Y2=0
cc_207 N_A_214_47#_c_228_n N_Z_c_540_n 0.0232389f $X=1.587 $Y=1.595 $X2=0 $Y2=0
cc_208 N_A_214_47#_c_229_n N_Z_c_540_n 0.133896f $X=3.645 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_214_47#_c_231_n N_Z_c_540_n 0.00830267f $X=3.645 $Y=1.035 $X2=0 $Y2=0
cc_210 N_A_214_47#_c_217_n N_VGND_c_603_n 0.00856801f $X=2.3 $Y=0.96 $X2=0 $Y2=0
cc_211 N_A_214_47#_c_220_n N_VGND_c_603_n 0.00699289f $X=2.72 $Y=0.96 $X2=0
+ $Y2=0
cc_212 N_A_214_47#_c_222_n N_VGND_c_603_n 6.07018e-19 $X=3.14 $Y=0.96 $X2=0
+ $Y2=0
cc_213 N_A_214_47#_c_220_n N_VGND_c_604_n 6.07018e-19 $X=2.72 $Y=0.96 $X2=0
+ $Y2=0
cc_214 N_A_214_47#_c_222_n N_VGND_c_604_n 0.00699289f $X=3.14 $Y=0.96 $X2=0
+ $Y2=0
cc_215 N_A_214_47#_c_232_n N_VGND_c_604_n 0.00810839f $X=3.645 $Y=0.96 $X2=0
+ $Y2=0
cc_216 N_A_214_47#_c_217_n N_VGND_c_606_n 0.00341689f $X=2.3 $Y=0.96 $X2=0 $Y2=0
cc_217 N_A_214_47#_c_226_n N_VGND_c_606_n 0.0422474f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_218 N_A_214_47#_c_220_n N_VGND_c_607_n 0.00341689f $X=2.72 $Y=0.96 $X2=0
+ $Y2=0
cc_219 N_A_214_47#_c_222_n N_VGND_c_607_n 0.00341689f $X=3.14 $Y=0.96 $X2=0
+ $Y2=0
cc_220 N_A_214_47#_c_232_n N_VGND_c_608_n 0.00341689f $X=3.645 $Y=0.96 $X2=0
+ $Y2=0
cc_221 N_A_214_47#_M1014_d N_VGND_c_609_n 0.00225448f $X=1.07 $Y=0.235 $X2=0
+ $Y2=0
cc_222 N_A_214_47#_c_217_n N_VGND_c_609_n 0.00540327f $X=2.3 $Y=0.96 $X2=0 $Y2=0
cc_223 N_A_214_47#_c_220_n N_VGND_c_609_n 0.0040262f $X=2.72 $Y=0.96 $X2=0 $Y2=0
cc_224 N_A_214_47#_c_222_n N_VGND_c_609_n 0.0040262f $X=3.14 $Y=0.96 $X2=0 $Y2=0
cc_225 N_A_214_47#_c_226_n N_VGND_c_609_n 0.0238257f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_226 N_A_214_47#_c_232_n N_VGND_c_609_n 0.00433138f $X=3.645 $Y=0.96 $X2=0
+ $Y2=0
cc_227 N_A_214_47#_c_226_n N_A_393_47#_c_681_n 0.0295289f $X=1.45 $Y=0.425 $X2=0
+ $Y2=0
cc_228 N_A_214_47#_c_227_n N_A_393_47#_c_681_n 0.00478569f $X=1.587 $Y=1.025
+ $X2=0 $Y2=0
cc_229 N_A_214_47#_c_217_n N_A_393_47#_c_686_n 0.0122116f $X=2.3 $Y=0.96 $X2=0
+ $Y2=0
cc_230 N_A_214_47#_c_218_n N_A_393_47#_c_686_n 0.00186586f $X=2.645 $Y=1.035
+ $X2=0 $Y2=0
cc_231 N_A_214_47#_c_220_n N_A_393_47#_c_686_n 0.0113204f $X=2.72 $Y=0.96 $X2=0
+ $Y2=0
cc_232 N_A_214_47#_c_229_n N_A_393_47#_c_686_n 0.0379559f $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_233 N_A_214_47#_c_227_n N_A_393_47#_c_682_n 0.0174646f $X=1.587 $Y=1.025
+ $X2=0 $Y2=0
cc_234 N_A_214_47#_c_229_n N_A_393_47#_c_682_n 0.02155f $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_235 N_A_214_47#_c_222_n N_A_393_47#_c_692_n 0.0113204f $X=3.14 $Y=0.96 $X2=0
+ $Y2=0
cc_236 N_A_214_47#_c_223_n N_A_393_47#_c_692_n 0.00186586f $X=3.48 $Y=1.035
+ $X2=0 $Y2=0
cc_237 N_A_214_47#_c_229_n N_A_393_47#_c_692_n 0.0466922f $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_238 N_A_214_47#_c_231_n N_A_393_47#_c_692_n 0.00311914f $X=3.645 $Y=1.035
+ $X2=0 $Y2=0
cc_239 N_A_214_47#_c_232_n N_A_393_47#_c_692_n 0.0116005f $X=3.645 $Y=0.96 $X2=0
+ $Y2=0
cc_240 N_A_214_47#_c_221_n N_A_393_47#_c_697_n 0.00193161f $X=3.065 $Y=1.035
+ $X2=0 $Y2=0
cc_241 N_A_214_47#_c_229_n N_A_393_47#_c_697_n 0.0119538f $X=3.645 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_320_n N_VPWR_c_411_n 0.00627922f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_330_n N_VPWR_c_414_n 0.0180037f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_244 N_A_27_47#_M1001_g N_VPWR_c_417_n 0.00357877f $X=4.1 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_27_47#_M1009_g N_VPWR_c_417_n 0.00357877f $X=4.52 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_M1012_g N_VPWR_c_417_n 0.00357877f $X=4.94 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_M1017_g N_VPWR_c_417_n 0.00357877f $X=5.36 $Y=1.985 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1013_s N_VPWR_c_410_n 0.00382897f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1001_g N_VPWR_c_410_n 0.00655123f $X=4.1 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1009_g N_VPWR_c_410_n 0.00522516f $X=4.52 $Y=1.985 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1012_g N_VPWR_c_410_n 0.00522516f $X=4.94 $Y=1.985 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1017_g N_VPWR_c_410_n 0.00629538f $X=5.36 $Y=1.985 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_330_n N_VPWR_c_410_n 0.00993674f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_254 N_A_27_47#_M1001_g N_A_320_309#_c_487_n 0.0179753f $X=4.1 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1009_g N_A_320_309#_c_487_n 0.0179713f $X=4.52 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1012_g N_A_320_309#_c_487_n 0.0179753f $X=4.94 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1017_g N_A_320_309#_c_487_n 0.0179753f $X=5.36 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1007_g N_Z_c_556_n 0.00331535f $X=4.1 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1008_g N_Z_c_556_n 0.0101668f $X=4.52 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_27_47#_M1010_g N_Z_c_556_n 0.0102073f $X=4.94 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_27_47#_M1015_g N_Z_c_556_n 0.0127239f $X=5.36 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_320_n N_Z_c_556_n 6.36393e-19 $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_333_n N_Z_c_556_n 0.00193698f $X=4.395 $Y=1.19 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_323_n N_Z_c_556_n 0.0828592f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_324_n N_Z_c_556_n 0.00585817f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_27_47#_M1015_g Z 0.00557285f $X=5.36 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_323_n Z 0.0213183f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_324_n Z 0.0071668f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1001_g N_Z_c_540_n 0.0151477f $X=4.1 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_27_47#_M1009_g N_Z_c_540_n 0.0116868f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_27_47#_M1012_g N_Z_c_540_n 0.0117437f $X=4.94 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_27_47#_M1017_g N_Z_c_540_n 0.0146833f $X=5.36 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_320_n N_Z_c_540_n 0.0216421f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_333_n N_Z_c_540_n 0.00792175f $X=4.395 $Y=1.19 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_323_n N_Z_c_540_n 0.10964f $X=5.27 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_324_n N_Z_c_540_n 0.00559408f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_320_n N_VGND_c_602_n 0.00667101f $X=4.25 $Y=1.19 $X2=0 $Y2=0
cc_278 N_A_27_47#_M1007_g N_VGND_c_604_n 0.00107009f $X=4.1 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_319_n N_VGND_c_605_n 0.0154729f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_27_47#_M1007_g N_VGND_c_608_n 0.00357877f $X=4.1 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A_27_47#_M1008_g N_VGND_c_608_n 0.00357877f $X=4.52 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_27_47#_M1010_g N_VGND_c_608_n 0.00357877f $X=4.94 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_27_47#_M1015_g N_VGND_c_608_n 0.00357877f $X=5.36 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_27_47#_M1018_s N_VGND_c_609_n 0.00388065f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1007_g N_VGND_c_609_n 0.00556923f $X=4.1 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_27_47#_M1008_g N_VGND_c_609_n 0.00522516f $X=4.52 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_27_47#_M1010_g N_VGND_c_609_n 0.00522516f $X=4.94 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_27_47#_M1015_g N_VGND_c_609_n 0.00629538f $X=5.36 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_319_n N_VGND_c_609_n 0.00980171f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_320_n N_A_393_47#_c_686_n 0.00400213f $X=4.25 $Y=1.19 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_320_n N_A_393_47#_c_682_n 0.00189895f $X=4.25 $Y=1.19 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_320_n N_A_393_47#_c_692_n 0.00974424f $X=4.25 $Y=1.19 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1007_g N_A_393_47#_c_683_n 0.0111875f $X=4.1 $Y=0.56 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1008_g N_A_393_47#_c_683_n 0.00814603f $X=4.52 $Y=0.56 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1010_g N_A_393_47#_c_683_n 0.00814603f $X=4.94 $Y=0.56 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1015_g N_A_393_47#_c_683_n 0.00814603f $X=5.36 $Y=0.56 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_323_n N_A_393_47#_c_683_n 0.00382597f $X=5.27 $Y=1.16 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_320_n N_A_393_47#_c_697_n 0.00114955f $X=4.25 $Y=1.19 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_410_n N_A_320_309#_M1000_s 0.00382897f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_300 N_VPWR_c_410_n N_A_320_309#_M1011_s 0.0040445f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_410_n N_A_320_309#_M1019_s 0.00628971f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_410_n N_A_320_309#_M1009_d 0.00215227f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_410_n N_A_320_309#_M1017_d 0.00225742f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_415_n N_A_320_309#_c_485_n 0.0166237f $X=1.98 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_410_n N_A_320_309#_c_485_n 0.00929827f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_416_n N_A_320_309#_c_512_n 0.0112554f $X=2.82 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_410_n N_A_320_309#_c_512_n 0.00644035f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_M1000_d N_A_320_309#_c_486_n 0.0031368f $X=2.01 $Y=1.545 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_412_n N_A_320_309#_c_486_n 0.0161728f $X=2.145 $Y=2.36 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_415_n N_A_320_309#_c_486_n 0.00207669f $X=1.98 $Y=2.72 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_416_n N_A_320_309#_c_486_n 0.00208431f $X=2.82 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_410_n N_A_320_309#_c_486_n 0.00729963f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_417_n N_A_320_309#_c_519_n 0.160759f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_410_n N_A_320_309#_c_519_n 0.0956142f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_M1016_d N_A_320_309#_c_493_n 0.00314385f $X=2.85 $Y=1.545 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_413_n N_A_320_309#_c_493_n 0.0160815f $X=2.985 $Y=2.36 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_416_n N_A_320_309#_c_493_n 0.00259065f $X=2.82 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_417_n N_A_320_309#_c_493_n 0.00259065f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_410_n N_A_320_309#_c_493_n 0.0101931f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_410_n N_Z_M1001_s 0.00216833f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_321 N_VPWR_c_410_n N_Z_M1012_s 0.00216833f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_M1000_d N_Z_c_540_n 0.00168399f $X=2.01 $Y=1.545 $X2=0 $Y2=0
cc_323 N_VPWR_M1016_d N_Z_c_540_n 0.0016881f $X=2.85 $Y=1.545 $X2=0 $Y2=0
cc_324 N_A_320_309#_c_487_n N_Z_M1001_s 0.00314062f $X=5.57 $Y=2.02 $X2=0 $Y2=0
cc_325 N_A_320_309#_c_487_n N_Z_M1012_s 0.00316076f $X=5.57 $Y=2.02 $X2=0 $Y2=0
cc_326 N_A_320_309#_M1017_d Z 9.75102e-19 $X=5.435 $Y=1.485 $X2=0 $Y2=0
cc_327 N_A_320_309#_c_487_n Z 0.020022f $X=5.57 $Y=2.02 $X2=0 $Y2=0
cc_328 N_A_320_309#_M1011_s N_Z_c_540_n 0.00168399f $X=2.43 $Y=1.545 $X2=0 $Y2=0
cc_329 N_A_320_309#_M1019_s N_Z_c_540_n 0.0121617f $X=3.27 $Y=1.545 $X2=0 $Y2=0
cc_330 N_A_320_309#_M1009_d N_Z_c_540_n 0.0016881f $X=4.595 $Y=1.485 $X2=0 $Y2=0
cc_331 N_A_320_309#_M1017_d N_Z_c_540_n 0.00274995f $X=5.435 $Y=1.485 $X2=0
+ $Y2=0
cc_332 N_A_320_309#_c_486_n N_Z_c_540_n 0.0440435f $X=2.65 $Y=2 $X2=0 $Y2=0
cc_333 N_A_320_309#_c_493_n N_Z_c_540_n 0.185742f $X=3.32 $Y=2.18 $X2=0 $Y2=0
cc_334 N_Z_c_537_n N_VGND_c_608_n 0.00338803f $X=5.785 $Y=0.855 $X2=0 $Y2=0
cc_335 N_Z_M1007_d N_VGND_c_609_n 0.00216833f $X=4.175 $Y=0.235 $X2=0 $Y2=0
cc_336 N_Z_M1010_d N_VGND_c_609_n 0.00216833f $X=5.015 $Y=0.235 $X2=0 $Y2=0
cc_337 N_Z_c_537_n N_VGND_c_609_n 0.00504335f $X=5.785 $Y=0.855 $X2=0 $Y2=0
cc_338 N_Z_c_556_n N_A_393_47#_M1008_s 0.00308199f $X=5.675 $Y=0.735 $X2=0 $Y2=0
cc_339 N_Z_c_556_n N_A_393_47#_M1015_s 0.00592387f $X=5.675 $Y=0.735 $X2=0 $Y2=0
cc_340 Z N_A_393_47#_M1015_s 4.28177e-19 $X=5.69 $Y=0.765 $X2=0 $Y2=0
cc_341 N_Z_c_537_n N_A_393_47#_M1015_s 9.56518e-19 $X=5.785 $Y=0.855 $X2=0 $Y2=0
cc_342 N_Z_c_540_n N_A_393_47#_c_692_n 0.00225779f $X=5.675 $Y=1.585 $X2=0 $Y2=0
cc_343 N_Z_M1007_d N_A_393_47#_c_683_n 0.00305132f $X=4.175 $Y=0.235 $X2=0 $Y2=0
cc_344 N_Z_M1010_d N_A_393_47#_c_683_n 0.00305132f $X=5.015 $Y=0.235 $X2=0 $Y2=0
cc_345 N_Z_c_556_n N_A_393_47#_c_683_n 0.0777916f $X=5.675 $Y=0.735 $X2=0 $Y2=0
cc_346 N_Z_c_537_n N_A_393_47#_c_683_n 0.0046867f $X=5.785 $Y=0.855 $X2=0 $Y2=0
cc_347 N_VGND_c_609_n N_A_393_47#_M1003_s 0.00229009f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_348 N_VGND_c_609_n N_A_393_47#_M1004_s 0.00255104f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_609_n N_A_393_47#_M1006_s 0.00332861f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_609_n N_A_393_47#_M1008_s 0.00215227f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_609_n N_A_393_47#_M1015_s 0.00225742f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_606_n N_A_393_47#_c_681_n 0.0192583f $X=2.345 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_609_n N_A_393_47#_c_681_n 0.0106713f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_M1003_d N_A_393_47#_c_686_n 0.00288179f $X=2.375 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_VGND_c_603_n N_A_393_47#_c_686_n 0.0162338f $X=2.51 $Y=0.36 $X2=0 $Y2=0
cc_356 N_VGND_c_606_n N_A_393_47#_c_686_n 0.00234306f $X=2.345 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_607_n N_A_393_47#_c_686_n 0.00234306f $X=3.185 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_609_n N_A_393_47#_c_686_n 0.00978207f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_359 N_VGND_c_607_n N_A_393_47#_c_729_n 0.00998989f $X=3.185 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_609_n N_A_393_47#_c_729_n 0.00637943f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_M1005_d N_A_393_47#_c_692_n 0.00296184f $X=3.215 $Y=0.235 $X2=0
+ $Y2=0
cc_362 N_VGND_c_604_n N_A_393_47#_c_692_n 0.0162338f $X=3.35 $Y=0.36 $X2=0 $Y2=0
cc_363 N_VGND_c_607_n N_A_393_47#_c_692_n 0.00234306f $X=3.185 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_608_n N_A_393_47#_c_692_n 0.00234306f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_609_n N_A_393_47#_c_692_n 0.00978207f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_608_n N_A_393_47#_c_736_n 0.0197284f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_609_n N_A_393_47#_c_736_n 0.011132f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_608_n N_A_393_47#_c_683_n 0.0983668f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_609_n N_A_393_47#_c_683_n 0.0627626f $X=5.75 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a22oi_1.spice
* Created: Thu Aug 27 14:02:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a22oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a22oi_1  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1007 A_109_47# N_B2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.169 PD=0.88 PS=1.82 NRD=11.076 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.07475 PD=1.82 PS=0.88 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 A_381_47# N_A1_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.169 PD=0.86 PS=1.82 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g A_381_47# VNB NSHORT L=0.15 W=0.65 AD=0.234
+ AS=0.06825 PD=2.02 PS=0.86 NRD=11.988 NRS=9.228 M=1 R=4.33333 SA=75000.5
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 N_A_109_297#_M1004_d N_B2_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_109_297#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_109_297#_M1006_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_109_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.3 AS=0.135 PD=2.6 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__a22oi_1.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__o2bb2ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 3.505000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 1.825000 1.285000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.045000 1.075000 10.005000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.075000 7.875000 1.285000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415000 0.645000 6.155000 0.905000 ;
        RECT 4.425000 1.455000 7.715000 1.625000 ;
        RECT 4.425000 1.625000 4.675000 2.465000 ;
        RECT 5.265000 1.625000 5.515000 2.465000 ;
        RECT 5.875000 0.905000 6.155000 1.455000 ;
        RECT 6.625000 1.625000 6.875000 2.125000 ;
        RECT 7.465000 1.625000 7.715000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 2.295000  0.085000  2.465000 0.555000 ;
        RECT 3.135000  0.085000  3.305000 0.555000 ;
        RECT 6.665000  0.085000  6.835000 0.555000 ;
        RECT 7.505000  0.085000  7.675000 0.555000 ;
        RECT 8.345000  0.085000  8.515000 0.555000 ;
        RECT 9.185000  0.085000  9.355000 0.555000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
        RECT 9.805000 -0.085000 9.975000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.155000 1.795000  0.405000 2.635000 ;
        RECT 0.995000 1.795000  1.245000 2.635000 ;
        RECT 1.835000 1.795000  2.085000 2.635000 ;
        RECT 2.675000 1.795000  2.925000 2.635000 ;
        RECT 3.515000 1.795000  4.255000 2.635000 ;
        RECT 4.845000 1.795000  5.095000 2.635000 ;
        RECT 5.685000 1.795000  5.935000 2.635000 ;
        RECT 8.305000 1.795000  8.555000 2.635000 ;
        RECT 9.145000 1.795000  9.395000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
        RECT 9.805000 2.635000 9.975000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.645000 1.705000 0.905000 ;
      RECT 0.085000 0.905000 0.255000 1.455000 ;
      RECT 0.085000 1.455000 3.915000 1.625000 ;
      RECT 0.100000 0.255000 2.125000 0.475000 ;
      RECT 0.575000 1.625000 0.825000 2.465000 ;
      RECT 1.415000 1.625000 1.665000 2.465000 ;
      RECT 1.875000 0.475000 2.125000 0.725000 ;
      RECT 1.875000 0.725000 3.805000 0.905000 ;
      RECT 2.255000 1.625000 2.505000 2.465000 ;
      RECT 2.635000 0.255000 2.965000 0.725000 ;
      RECT 3.095000 1.625000 3.345000 2.465000 ;
      RECT 3.475000 0.255000 3.805000 0.725000 ;
      RECT 3.745000 1.075000 5.705000 1.285000 ;
      RECT 3.745000 1.285000 3.915000 1.455000 ;
      RECT 4.060000 0.255000 6.495000 0.475000 ;
      RECT 4.060000 0.475000 4.245000 0.835000 ;
      RECT 6.175000 1.795000 6.455000 2.295000 ;
      RECT 6.175000 2.295000 8.135000 2.465000 ;
      RECT 6.325000 0.475000 6.495000 0.735000 ;
      RECT 6.325000 0.735000 9.855000 0.905000 ;
      RECT 7.005000 0.255000 7.335000 0.725000 ;
      RECT 7.005000 0.725000 9.855000 0.735000 ;
      RECT 7.045000 1.795000 7.295000 2.295000 ;
      RECT 7.845000 0.255000 8.175000 0.725000 ;
      RECT 7.885000 1.455000 9.875000 1.625000 ;
      RECT 7.885000 1.625000 8.135000 2.295000 ;
      RECT 8.685000 0.255000 9.015000 0.725000 ;
      RECT 8.725000 1.625000 8.975000 2.465000 ;
      RECT 9.525000 0.255000 9.855000 0.725000 ;
      RECT 9.565000 1.625000 9.875000 2.465000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_4

* File: sky130_fd_sc_hd__o2bb2a_2.pex.spice
* Created: Thu Aug 27 14:38:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%A_84_21# 1 2 7 9 12 14 16 19 23 24 27 28 29
+ 38 41 44 45 47 49
c114 19 0 1.14156e-19 $X=0.915 $Y=1.985
r115 51 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.915 $Y2=1.16
r116 45 47 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.715 $Y=1.245
+ $X2=2.715 $Y2=1.495
r117 44 45 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.705 $Y=1.075
+ $X2=2.705 $Y2=1.245
r118 43 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.695 $Y=0.69
+ $X2=2.695 $Y2=1.075
r119 41 43 10.7341 $w=2.43e-07 $l=2.05e-07 $layer=LI1_cond $X=2.657 $Y=0.485
+ $X2=2.657 $Y2=0.69
r120 36 38 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.96 $Y=1.53
+ $X2=1.185 $Y2=1.53
r121 28 49 0.646529 $w=5.53e-07 $l=3e-08 $layer=LI1_cond $X=2.907 $Y=1.97
+ $X2=2.907 $Y2=2
r122 28 47 16.5449 $w=5.53e-07 $l=4.75e-07 $layer=LI1_cond $X=2.907 $Y=1.97
+ $X2=2.907 $Y2=1.495
r123 28 29 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.63 $Y=1.97
+ $X2=1.27 $Y2=1.97
r124 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.185 $Y=1.885
+ $X2=1.27 $Y2=1.97
r125 26 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.615
+ $X2=1.185 $Y2=1.53
r126 26 27 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.185 $Y=1.615
+ $X2=1.185 $Y2=1.885
r127 24 53 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=0.96 $Y=1.16
+ $X2=0.915 $Y2=1.16
r128 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.16 $X2=0.96 $Y2=1.16
r129 21 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=1.445
+ $X2=0.96 $Y2=1.53
r130 21 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.96 $Y=1.445
+ $X2=0.96 $Y2=1.16
r131 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.325
+ $X2=0.915 $Y2=1.16
r132 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.915 $Y=1.325
+ $X2=0.915 $Y2=1.985
r133 14 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=0.995
+ $X2=0.915 $Y2=1.16
r134 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.915 $Y=0.995
+ $X2=0.915 $Y2=0.56
r135 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r136 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.985
r137 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=1.16
r138 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=0.56
r139 2 49 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.885
+ $Y=1.845 $X2=3.02 $Y2=2
r140 1 41 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.62 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%A1_N 3 7 9 12
c38 9 0 1.58869e-19 $X=1.6 $Y=1.19
r39 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.16
+ $X2=1.44 $Y2=1.325
r40 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.16
+ $X2=1.44 $Y2=0.995
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.44
+ $Y=1.16 $X2=1.44 $Y2=1.16
r42 9 13 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=1.6 $Y=1.175 $X2=1.44
+ $Y2=1.175
r43 7 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.4 $Y=2.165 $X2=1.4
+ $Y2=1.325
r44 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.395 $Y=0.445
+ $X2=1.395 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%A2_N 3 6 8 12 13 16
c44 12 0 1.58869e-19 $X=1.94 $Y=0.935
r45 12 17 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=0.935
+ $X2=1.93 $Y2=1.1
r46 12 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=0.935
+ $X2=1.93 $Y2=0.77
r47 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=0.935 $X2=1.94 $Y2=0.935
r48 9 13 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.625 $Y=0.735
+ $X2=1.625 $Y2=0.51
r49 8 11 16.4231 $w=2.34e-07 $l=3.15e-07 $layer=LI1_cond $X=1.625 $Y=0.905
+ $X2=1.94 $Y2=0.905
r50 8 9 1.08988 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=1.625 $Y=0.905
+ $X2=1.625 $Y2=0.735
r51 6 17 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=1.95 $Y=2.165
+ $X2=1.95 $Y2=1.1
r52 3 16 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.86 $Y=0.445
+ $X2=1.86 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%A_295_369# 1 2 9 13 15 16 17 21 28 30
c67 17 0 1.14156e-19 $X=2.195 $Y=1.605
r68 28 30 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.327 $Y=1.52
+ $X2=2.327 $Y2=1.355
r69 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.52 $X2=2.375 $Y2=1.52
r70 25 30 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.28 $Y=0.565
+ $X2=2.28 $Y2=1.355
r71 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.195 $Y=0.48
+ $X2=2.28 $Y2=0.565
r72 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=0.48
+ $X2=2.07 $Y2=0.48
r73 17 28 3.69652 $w=2.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.327 $Y=1.605
+ $X2=2.327 $Y2=1.52
r74 17 19 27.2396 $w=2.18e-07 $l=5.2e-07 $layer=LI1_cond $X=2.195 $Y=1.605
+ $X2=1.675 $Y2=1.605
r75 15 29 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.735 $Y=1.52
+ $X2=2.375 $Y2=1.52
r76 15 16 5.03009 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=2.735 $Y=1.52
+ $X2=2.82 $Y2=1.52
r77 11 16 37.0704 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.83 $Y=1.355
+ $X2=2.82 $Y2=1.52
r78 11 13 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.83 $Y=1.355
+ $X2=2.83 $Y2=0.445
r79 7 16 37.0704 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.81 $Y=1.685
+ $X2=2.82 $Y2=1.52
r80 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.81 $Y=1.685 $X2=2.81
+ $Y2=2.165
r81 2 19 600 $w=1.7e-07 $l=2.98706e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=1.845 $X2=1.675 $Y2=1.63
r82 1 23 182 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.235 $X2=2.07 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%B2 3 7 9 12 14
r50 13 14 14.7118 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.44 $Y=1.325
+ $X2=3.44 $Y2=1.53
r51 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.16 $X2=3.25 $Y2=1.16
r52 9 13 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.355 $Y=1.2
+ $X2=3.44 $Y2=1.325
r53 9 11 5.124 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.355 $Y=1.2 $X2=3.25
+ $Y2=1.2
r54 5 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.16
r55 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.25 $Y=1.325 $X2=3.25
+ $Y2=2.165
r56 1 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=1.16
r57 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.25 $Y=0.995 $X2=3.25
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%B1 3 7 9 10 16
r27 13 16 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.67 $Y=1.16
+ $X2=3.865 $Y2=1.16
r28 9 10 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.872 $Y=1.16
+ $X2=3.872 $Y2=1.53
r29 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.865
+ $Y=1.16 $X2=3.865 $Y2=1.16
r30 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r31 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.67 $Y=1.325 $X2=3.67
+ $Y2=2.165
r32 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r33 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.67 $Y=0.995 $X2=3.67
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%VPWR 1 2 3 4 13 15 21 23 25 27 29 34 39 48
+ 51 59 63
r61 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 45 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 43 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 43 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r66 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 40 42 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 39 58 4.63403 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.935 $Y2=2.72
r69 39 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 38 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r73 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=2.72
+ $X2=1.125 $Y2=2.72
r74 35 37 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.29 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 34 40 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=2.362 $Y=2.72
+ $X2=2.565 $Y2=2.72
r76 34 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 34 51 11.3822 $w=4.03e-07 $l=4e-07 $layer=LI1_cond $X=2.362 $Y=2.72
+ $X2=2.362 $Y2=2.32
r78 34 37 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=2.72 $X2=2.07
+ $Y2=2.72
r79 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r80 33 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 30 45 4.06635 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r83 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.69 $Y2=2.72
r84 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=1.125 $Y2=2.72
r85 29 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.96 $Y=2.72 $X2=0.69
+ $Y2=2.72
r86 27 63 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 23 58 3.00647 $w=3.15e-07 $l=1.06325e-07 $layer=LI1_cond $X=3.887 $Y=2.635
+ $X2=3.935 $Y2=2.72
r88 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=3.887 $Y=2.635
+ $X2=3.887 $Y2=2
r89 19 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=2.635
+ $X2=1.125 $Y2=2.72
r90 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.125 $Y=2.635
+ $X2=1.125 $Y2=2.32
r91 15 18 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.237 $Y=1.62
+ $X2=0.237 $Y2=2.3
r92 13 45 3.11087 $w=2.55e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.182 $Y2=2.72
r93 13 18 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.237 $Y2=2.3
r94 4 25 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.845 $X2=3.88 $Y2=2
r95 3 51 600 $w=1.7e-07 $l=6.22194e-07 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.845 $X2=2.365 $Y2=2.32
r96 2 21 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.485 $X2=1.125 $Y2=2.32
r97 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r98 1 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%X 1 2 9 13 14 15 16 19
r29 16 19 11.2985 $w=2.53e-07 $l=2.5e-07 $layer=LI1_cond $X=0.662 $Y=2.21
+ $X2=0.662 $Y2=1.96
r30 14 19 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=0.662 $Y=1.922
+ $X2=0.662 $Y2=1.96
r31 14 15 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=0.662 $Y=1.922
+ $X2=0.662 $Y2=1.795
r32 13 15 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.62 $Y=0.825
+ $X2=0.62 $Y2=1.795
r33 7 13 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=0.702 $Y=0.658
+ $X2=0.702 $Y2=0.825
r34 7 9 9.90757 $w=3.33e-07 $l=2.88e-07 $layer=LI1_cond $X=0.702 $Y=0.658
+ $X2=0.702 $Y2=0.37
r35 2 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.485 $X2=0.705 $Y2=1.96
r36 1 9 91 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.705 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
+ 51
r60 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r61 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 40 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r63 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r64 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r65 34 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=0 $X2=3.46
+ $Y2=0
r66 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.545 $Y=0 $X2=3.91
+ $Y2=0
r67 33 47 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r68 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r69 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r70 30 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.15
+ $Y2=0
r71 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.61
+ $Y2=0
r72 29 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.46
+ $Y2=0
r73 29 32 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=3.375 $Y=0 $X2=1.61
+ $Y2=0
r74 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r75 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r76 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r77 25 40 4.06635 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r78 25 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r79 24 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.15
+ $Y2=0
r80 24 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.69
+ $Y2=0
r81 22 51 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=0 $X2=0.23
+ $Y2=0
r82 18 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0
r83 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0.39
r84 14 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r85 14 16 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.525
r86 10 40 3.11087 $w=2.55e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.182 $Y2=0
r87 10 12 12.8802 $w=2.53e-07 $l=2.85e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.37
r88 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.39
r89 2 16 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.235 $X2=1.15 $Y2=0.525
r90 1 12 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_2%A_581_47# 1 2 9 11 12 15
r32 13 15 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.88 $Y=0.725
+ $X2=3.88 $Y2=0.435
r33 11 13 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.715 $Y=0.815
+ $X2=3.88 $Y2=0.725
r34 11 12 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=3.715 $Y=0.815
+ $X2=3.185 $Y2=0.815
r35 7 12 6.94918 $w=1.8e-07 $l=1.53542e-07 $layer=LI1_cond $X=3.07 $Y=0.725
+ $X2=3.185 $Y2=0.815
r36 7 9 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.07 $Y=0.725 $X2=3.07
+ $Y2=0.485
r37 2 15 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.435
r38 1 9 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.04 $Y2=0.485
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o32ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.075000 5.865000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 1.075000 4.480000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 3.065000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.075000 1.705000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.845000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 2.045000 0.905000 ;
        RECT 0.515000 1.495000 3.105000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.095000 ;
        RECT 1.875000 0.905000 2.045000 1.105000 ;
        RECT 1.875000 1.105000 2.170000 1.495000 ;
        RECT 2.775000 1.665000 3.105000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 2.620000  0.085000 2.950000 0.545000 ;
        RECT 3.635000  0.085000 3.805000 0.545000 ;
        RECT 4.905000  0.085000 5.235000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 1.435000 2.175000 1.605000 2.635000 ;
        RECT 4.620000 1.835000 4.825000 2.635000 ;
        RECT 5.495000 1.495000 5.715000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 2.405000 0.485000 ;
      RECT 0.090000 0.485000 0.345000 0.905000 ;
      RECT 0.090000 1.495000 0.345000 2.295000 ;
      RECT 0.090000 2.295000 1.265000 2.465000 ;
      RECT 1.015000 1.835000 2.105000 2.005000 ;
      RECT 1.015000 2.005000 1.265000 2.295000 ;
      RECT 1.775000 2.005000 2.105000 2.455000 ;
      RECT 2.235000 0.485000 2.405000 0.715000 ;
      RECT 2.235000 0.715000 5.755000 0.905000 ;
      RECT 2.335000 1.835000 2.585000 2.255000 ;
      RECT 2.335000 2.255000 4.385000 2.445000 ;
      RECT 3.135000 0.255000 3.465000 0.715000 ;
      RECT 3.275000 1.495000 3.445000 2.255000 ;
      RECT 3.615000 1.495000 5.325000 1.665000 ;
      RECT 3.615000 1.665000 3.945000 2.085000 ;
      RECT 4.055000 0.255000 4.725000 0.715000 ;
      RECT 4.135000 1.835000 4.385000 2.255000 ;
      RECT 4.995000 1.665000 5.325000 2.460000 ;
      RECT 5.425000 0.255000 5.755000 0.715000 ;
  END
END sky130_fd_sc_hd__o32ai_2

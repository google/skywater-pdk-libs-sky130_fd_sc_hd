* File: sky130_fd_sc_hd__or2_0.spice.pex
* Created: Thu Aug 27 14:42:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR2_0%B 1 3 6 8 12 15
r25 14 15 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.615 $Y=1.16
+ $X2=0.675 $Y2=1.16
r26 11 14 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.415 $Y=1.16
+ $X2=0.615 $Y2=1.16
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.16 $X2=0.415 $Y2=1.16
r28 8 12 3.56894 $w=6.18e-07 $l=1.85e-07 $layer=LI1_cond $X=0.23 $Y=1.305
+ $X2=0.415 $Y2=1.305
r29 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=1.325
+ $X2=0.675 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.675 $Y=1.325
+ $X2=0.675 $Y2=1.985
r31 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=1.16
r32 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_0%A 3 6 8 9 13 15
r32 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.16
+ $X2=1.095 $Y2=1.325
r33 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.16
+ $X2=1.095 $Y2=0.995
r34 8 9 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.172 $Y=1.16
+ $X2=1.172 $Y2=1.53
r35 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.16 $X2=1.095 $Y2=1.16
r36 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.035 $Y=1.985
+ $X2=1.035 $Y2=1.325
r37 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.035 $Y=0.675
+ $X2=1.035 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_0%A_68_355# 1 2 9 12 15 16 17 20 21 27 31
c60 20 0 9.5905e-20 $X=1.61 $Y=1.16
c61 15 0 1.0136e-19 $X=0.755 $Y=1.785
r62 27 29 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0.66
+ $X2=0.81 $Y2=0.825
r63 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.61 $Y2=1.325
r64 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.61 $Y2=0.995
r65 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r66 18 20 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.61 $Y=1.785
+ $X2=1.61 $Y2=1.16
r67 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.87
+ $X2=1.61 $Y2=1.785
r68 16 17 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.525 $Y=1.87
+ $X2=0.84 $Y2=1.87
r69 15 17 5.63966 $w=2.89e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.84 $Y2=1.87
r70 15 24 12.2422 $w=2.89e-07 $l=3.66033e-07 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.465 $Y2=1.957
r71 15 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.755 $Y2=0.825
r72 12 32 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.52 $Y=2.095
+ $X2=1.52 $Y2=1.325
r73 9 31 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.52 $Y=0.675
+ $X2=1.52 $Y2=0.995
r74 2 24 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.775 $X2=0.465 $Y2=1.95
r75 1 27 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.465 $X2=0.825 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_0%VPWR 1 6 8 10 17 18 21
r23 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r26 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.31 $Y2=2.72
r27 15 17 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=2.07 $Y2=2.72
r28 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=2.72
+ $X2=1.31 $Y2=2.72
r29 10 12 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.145 $Y=2.72
+ $X2=0.23 $Y2=2.72
r30 8 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r31 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r32 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=2.635 $X2=1.31
+ $Y2=2.72
r33 4 6 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.31 $Y=2.635
+ $X2=1.31 $Y2=2.21
r34 1 6 600 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.775 $X2=1.31 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_0%X 1 2 10 16 19
c21 2 0 9.5905e-20 $X=1.595 $Y=1.775
r22 17 19 9.69516 $w=3.13e-07 $l=2.65e-07 $layer=LI1_cond $X=2.022 $Y=2.135
+ $X2=2.022 $Y2=1.87
r23 16 17 1.01705 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=2.022 $Y=2.3
+ $X2=2.022 $Y2=2.135
r24 14 16 7.40357 $w=3.28e-07 $l=2.12e-07 $layer=LI1_cond $X=1.81 $Y=2.3
+ $X2=2.022 $Y2=2.3
r25 11 19 38.2318 $w=3.13e-07 $l=1.045e-06 $layer=LI1_cond $X=2.022 $Y=0.825
+ $X2=2.022 $Y2=1.87
r26 10 11 0.437101 $w=3.15e-07 $l=1.5e-07 $layer=LI1_cond $X=2.022 $Y=0.675
+ $X2=2.022 $Y2=0.825
r27 8 10 11.2171 $w=2.98e-07 $l=2.92e-07 $layer=LI1_cond $X=1.73 $Y=0.675
+ $X2=2.022 $Y2=0.675
r28 2 14 600 $w=1.7e-07 $l=5.41941e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.775 $X2=1.81 $Y2=2.22
r29 1 8 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.465 $X2=1.73 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_0%VGND 1 2 7 9 13 16 17 18 25 26
r26 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r27 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r28 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r29 20 29 3.81131 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=0 $X2=0.245
+ $Y2=0
r30 20 22 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=0.49 $Y=0 $X2=1.15
+ $Y2=0
r31 18 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r32 18 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r33 16 22 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.15
+ $Y2=0
r34 16 17 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.287
+ $Y2=0
r35 15 25 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=2.07
+ $Y2=0
r36 15 17 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.287
+ $Y2=0
r37 11 17 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.287 $Y=0.085
+ $X2=1.287 $Y2=0
r38 11 13 30.8211 $w=2.13e-07 $l=5.75e-07 $layer=LI1_cond $X=1.287 $Y=0.085
+ $X2=1.287 $Y2=0.66
r39 7 29 3.26684 $w=2.4e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.245 $Y2=0
r40 7 9 27.6106 $w=2.38e-07 $l=5.75e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.66
r41 2 13 182 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.465 $X2=1.305 $Y2=0.66
r42 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.28
+ $Y=0.465 $X2=0.405 $Y2=0.66
.ends


* File: sky130_fd_sc_hd__o2111ai_1.spice
* Created: Thu Aug 27 14:34:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2111ai_1.pex.spice"
.subckt sky130_fd_sc_hd__o2111ai_1  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1002 A_163_47# N_D1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.17225 PD=0.86 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75002.2
+ A=0.0975 P=1.6 MULT=1
MM1003 A_235_47# N_C1_M1003_g A_163_47# VNB NSHORT L=0.15 W=0.65 AD=0.12675
+ AS=0.06825 PD=1.04 PS=0.86 NRD=25.836 NRS=9.228 M=1 R=4.33333 SA=75000.5
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_343_47#_M1005_d N_B1_M1005_g A_235_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.131625 AS=0.12675 PD=1.055 PS=1.04 NRD=13.836 NRS=25.836 M=1 R=4.33333
+ SA=75001.1 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_343_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.131625 PD=1.04 PS=1.055 NRD=7.38 NRS=9.228 M=1 R=4.33333
+ SA=75001.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1000 N_A_343_47#_M1000_d N_A1_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.12675 PD=1.83 PS=1.04 NRD=0 NRS=12.912 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_D1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.14 PD=1.39 PS=1.28 NRD=11.8003 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001.8
+ A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1 AD=0.2025
+ AS=0.195 PD=1.405 PS=1.39 NRD=14.7553 NRS=9.8303 M=1 R=6.66667 SA=75001.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1008 A_454_297# N_A2_M1008_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.2025 PD=1.39 PS=1.405 NRD=27.5603 NRS=9.8303 M=1 R=6.66667 SA=75001.7
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_454_297# VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.195 PD=2.53 PS=1.39 NRD=0 NRS=27.5603 M=1 R=6.66667 SA=75002.3 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_29 VNB 0 1.59109e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__o2111ai_1.pxi.spice"
*
.ends
*
*

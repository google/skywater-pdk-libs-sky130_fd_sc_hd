* NGSPICE file created from sky130_fd_sc_hd__clkbuf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=5.85e+11p ps=5.17e+06u
M1001 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=1.113e+11p ps=1.37e+06u
M1002 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1003 X a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1004 VGND a_27_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_27_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


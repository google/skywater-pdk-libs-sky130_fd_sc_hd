* File: sky130_fd_sc_hd__or4_4.spice
* Created: Tue Sep  1 19:28:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4_4.pex.spice"
.subckt sky130_fd_sc_hd__or4_4  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_A_32_297#_M1004_d N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.169 PD=1.03 PS=1.82 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_C_M1012_g N_A_32_297#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=4.608 M=1 R=4.33333 SA=75000.7
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1014 N_A_32_297#_M1014_d N_B_M1014_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_32_297#_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=17.532 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_32_297#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75002.1
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1001_d N_A_32_297#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_32_297#_M1006_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1006_d N_A_32_297#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.17875 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 A_114_297# N_D_M1002_g N_A_32_297#_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.19
+ AS=0.26 PD=1.38 PS=2.52 NRD=26.5753 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75003.4
+ A=0.15 P=2.3 MULT=1
MM1009 A_220_297# N_C_M1009_g A_114_297# VPB PHIGHVT L=0.15 W=1 AD=0.135 AS=0.19
+ PD=1.27 PS=1.38 NRD=15.7403 NRS=26.5753 M=1 R=6.66667 SA=75000.7 SB=75002.8
+ A=0.15 P=2.3 MULT=1
MM1008 A_304_297# N_B_M1008_g A_220_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_304_297# VPB PHIGHVT L=0.15 W=1 AD=0.19
+ AS=0.135 PD=1.38 PS=1.27 NRD=9.8303 NRS=15.7403 M=1 R=6.66667 SA=75001.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1005_d N_A_32_297#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.19 AS=0.135 PD=1.38 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75002.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_32_297#_M1010_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1010_d N_A_32_297#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_32_297#_M1013_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.135 PD=2.54 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__or4_4.pxi.spice"
*
.ends
*
*

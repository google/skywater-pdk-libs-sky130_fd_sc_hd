* File: sky130_fd_sc_hd__nor3b_1.spice
* Created: Tue Sep  1 19:18:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor3b_1.pex.spice"
.subckt sky130_fd_sc_hd__nor3b_1  VNB VPB B A C_N Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* C_N	C_N
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_91_199#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.221 PD=0.92 PS=1.98 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75000.3
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1004 N_A_91_199#_M1004_d N_C_N_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0787009 PD=1.36 PS=0.773271 NRD=0 NRS=17.856 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_161_297# N_A_91_199#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.32 PD=1.27 PS=2.64 NRD=15.7403 NRS=10.8153 M=1 R=6.66667
+ SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1002 A_245_297# N_B_M1002_g A_161_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.7
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_245_297# VPB PHIGHVT L=0.15 W=1 AD=0.205282
+ AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75000.4 A=0.15 P=2.3 MULT=1
MM1001 N_A_91_199#_M1001_d N_C_N_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0862183 PD=1.36 PS=0.789718 NRD=0 NRS=70.4866 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__nor3b_1.pxi.spice"
*
.ends
*
*

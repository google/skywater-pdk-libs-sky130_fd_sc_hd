* File: sky130_fd_sc_hd__a21boi_4.spice
* Created: Tue Sep  1 18:51:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21boi_4.pex.spice"
.subckt sky130_fd_sc_hd__a21boi_4  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_B1_N_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.26975 PD=1.03 PS=2.13 NRD=11.076 NRS=23.988 M=1 R=4.33333
+ SA=75000.3 SB=75005.8 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1016_d N_A_27_47#_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.091 PD=1.03 PS=0.93 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_27_47#_M1009_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.3
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1009_d N_A_27_47#_M1018_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A_27_47#_M1019_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.091 PD=1.27 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1019_d N_A2_M1007_g N_A_658_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.091 PD=1.27 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_658_47#_M1007_s N_A1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.4
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1011 N_A_658_47#_M1011_d N_A1_M1011_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.8
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1021 N_A_658_47#_M1011_d N_A1_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1022 N_A_658_47#_M1022_d N_A1_M1022_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.6
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A2_M1014_g N_A_658_47#_M1022_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.1
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1014_d N_A2_M1015_g N_A_658_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_A2_M1024_g N_A_658_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1025 N_VPWR_M1025_d N_B1_N_M1025_g N_A_27_47#_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_223_297#_M1000_d N_A_27_47#_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005 A=0.15 P=2.3 MULT=1
MM1005 N_A_223_297#_M1005_d N_A_27_47#_M1005_g N_Y_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1010 N_A_223_297#_M1005_d N_A_27_47#_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1020 N_A_223_297#_M1020_d N_A_27_47#_M1020_g N_Y_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.155 AS=0.14 PD=1.31 PS=1.28 NRD=5.8903 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_223_297#_M1020_d VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.155 PD=1.29 PS=1.31 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1002_d N_A1_M1003_g N_A_223_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.14 PD=1.29 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_223_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1008_d N_A1_M1012_g N_A_223_297#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_A1_M1023_g N_A_223_297#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.7
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1023_d N_A2_M1004_g N_A_223_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A2_M1013_g N_A_223_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1013_d N_A2_M1017_g N_A_223_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75005 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=11.6844 P=17.77
c_52 VNB 0 9.67612e-20 $X=0.145 $Y=-0.085
c_100 VPB 0 3.12905e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a21boi_4.pxi.spice"
*
.ends
*
*

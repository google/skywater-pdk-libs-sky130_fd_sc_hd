* File: sky130_fd_sc_hd__o22a_1.spice
* Created: Tue Sep  1 19:23:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o22a_1.pex.spice"
.subckt sky130_fd_sc_hd__o22a_1  VNB VPB B1 B2 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_78_199#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_78_199#_M1004_d N_B1_M1004_g N_A_215_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1001 N_A_215_47#_M1001_d N_B2_M1001_g N_A_78_199#_M1004_d VNB NSHORT L=0.15
+ W=0.65 AD=0.11375 AS=0.08775 PD=1 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_215_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1005 N_A_215_47#_M1005_d N_A1_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_78_199#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3725 AS=0.28 PD=1.745 PS=2.56 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1006 A_292_297# N_B1_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.1175
+ AS=0.3725 PD=1.235 PS=1.745 NRD=12.2928 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1002 N_A_78_199#_M1002_d N_B2_M1002_g A_292_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.235 AS=0.1175 PD=1.47 PS=1.235 NRD=0 NRS=12.2928 M=1 R=6.66667 SA=75001.5
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1007 A_493_297# N_A2_M1007_g N_A_78_199#_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.235 PD=1.21 PS=1.47 NRD=9.8303 NRS=38.3953 M=1 R=6.66667
+ SA=75002.1 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_493_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_31 VNB 0 9.14711e-20 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__o22a_1.pxi.spice"
*
.ends
*
*

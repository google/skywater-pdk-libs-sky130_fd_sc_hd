* File: sky130_fd_sc_hd__nand2b_1.pex.spice
* Created: Thu Aug 27 14:29:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2B_1%A_N 1 3 6 8 14
c27 8 0 1.91765e-19 $X=0.235 $Y=1.19
r28 11 14 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r30 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r31 4 6 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r32 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r33 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_1%B 3 6 8 11 12 13
c34 11 0 1.91765e-19 $X=0.92 $Y=1.16
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=1.325
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.92
+ $Y=1.16 $X2=0.92 $Y2=1.16
r38 8 12 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=0.695 $Y=1.195
+ $X2=0.92 $Y2=1.195
r39 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.985
+ $X2=0.955 $Y2=1.325
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.56
+ $X2=0.955 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_1%A_27_93# 1 2 9 12 14 16 19 21 23 27 35 36
+ 39
r71 36 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.16
+ $X2=1.465 $Y2=1.325
r72 36 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.16
+ $X2=1.465 $Y2=0.995
r73 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.16 $X2=1.465 $Y2=1.16
r74 32 35 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=1.2
+ $X2=1.465 $Y2=1.2
r75 27 30 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=0.23 $Y=1.58 $X2=0.23
+ $Y2=1.66
r76 23 25 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.225 $Y=0.69
+ $X2=0.225 $Y2=0.82
r77 20 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.2
r78 20 21 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.495
r79 19 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=1.075
+ $X2=1.34 $Y2=1.2
r80 18 19 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.34 $Y=0.905
+ $X2=1.34 $Y2=1.075
r81 17 27 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.37 $Y=1.58 $X2=0.23
+ $Y2=1.58
r82 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.255 $Y=1.58
+ $X2=1.34 $Y2=1.495
r83 16 17 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.255 $Y=1.58
+ $X2=0.37 $Y2=1.58
r84 15 25 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.36 $Y=0.82
+ $X2=0.225 $Y2=0.82
r85 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.255 $Y=0.82
+ $X2=1.34 $Y2=0.905
r86 14 15 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.255 $Y=0.82
+ $X2=0.36 $Y2=0.82
r87 12 40 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.375 $Y=1.985
+ $X2=1.375 $Y2=1.325
r88 9 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.375 $Y=0.56
+ $X2=1.375 $Y2=0.995
r89 2 30 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r90 1 23 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r30 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r32 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 27 36 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.715 $Y=2.72
+ $X2=1.607 $Y2=2.72
r35 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.715 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.83 $Y=2.72
+ $X2=0.705 $Y2=2.72
r40 23 25 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=2.72 $X2=1.15
+ $Y2=2.72
r41 22 36 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.5 $Y=2.72
+ $X2=1.607 $Y2=2.72
r42 22 25 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.5 $Y=2.72 $X2=1.15
+ $Y2=2.72
r43 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.705 $Y2=2.72
r44 17 19 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.23 $Y2=2.72
r45 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 11 36 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.72
r48 11 13 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.34
r49 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r50 7 9 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2
r51 2 13 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.585 $Y2=2.34
r52 1 9 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.745 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_1%Y 1 2 9 11 16 17 18 19 20 21 29 30
r43 21 30 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.92
+ $X2=1.985 $Y2=1.835
r44 21 30 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.985 $Y=1.81
+ $X2=1.985 $Y2=1.835
r45 20 21 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.985 $Y=1.53
+ $X2=1.985 $Y2=1.81
r46 19 20 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.985 $Y=1.19
+ $X2=1.985 $Y2=1.53
r47 18 19 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.985 $Y=0.85
+ $X2=1.985 $Y2=1.19
r48 17 29 3.05272 $w=3.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.985 $Y=0.4
+ $X2=1.985 $Y2=0.545
r49 17 18 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.985 $Y=0.57
+ $X2=1.985 $Y2=0.85
r50 17 29 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.985 $Y=0.57
+ $X2=1.985 $Y2=0.545
r51 11 17 3.89485 $w=2.9e-07 $l=1.85e-07 $layer=LI1_cond $X=1.8 $Y=0.4 $X2=1.985
+ $Y2=0.4
r52 11 13 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.8 $Y=0.4
+ $X2=1.585 $Y2=0.4
r53 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=1.92
+ $X2=1.165 $Y2=1.92
r54 9 21 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.8 $Y=1.92 $X2=1.985
+ $Y2=1.92
r55 9 10 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.8 $Y=1.92 $X2=1.33
+ $Y2=1.92
r56 2 16 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=2
r57 1 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.585 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_1%VGND 1 6 8 10 20 21 24
r28 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r29 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r30 18 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r31 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r32 17 20 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r33 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r34 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.745
+ $Y2=0
r35 15 17 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.15
+ $Y2=0
r36 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.745
+ $Y2=0
r37 10 12 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.23
+ $Y2=0
r38 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r39 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r40 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r41 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.38
r42 1 6 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.745 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__nand3b_2.pex.spice
* Created: Thu Aug 27 14:29:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND3B_2%A_N 3 7 9 12
c27 12 0 1.90991e-19 $X=0.595 $Y=1.16
r28 12 15 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=1.325
r29 12 14 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=0.995
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r31 9 13 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.595 $Y2=1.175
r32 7 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r33 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%C 3 7 11 15 17 18 26
c46 26 0 1.37483e-19 $X=1.435 $Y=1.16
c47 18 0 1.90991e-19 $X=1.53 $Y=1.105
r48 24 26 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.225 $Y=1.16
+ $X2=1.435 $Y2=1.16
r49 21 24 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.015 $Y=1.16
+ $X2=1.225 $Y2=1.16
r50 17 18 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.615 $Y2=1.175
r51 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.16 $X2=1.225 $Y2=1.16
r52 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.435 $Y=1.295
+ $X2=1.435 $Y2=1.16
r53 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.435 $Y=1.295
+ $X2=1.435 $Y2=1.985
r54 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.435 $Y=1.025
+ $X2=1.435 $Y2=1.16
r55 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.435 $Y=1.025
+ $X2=1.435 $Y2=0.56
r56 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.015 $Y=1.295
+ $X2=1.015 $Y2=1.16
r57 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.015 $Y=1.295
+ $X2=1.015 $Y2=1.985
r58 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.015 $Y=1.025
+ $X2=1.015 $Y2=1.16
r59 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.015 $Y=1.025
+ $X2=1.015 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%B 3 7 11 15 17 18 19 30
c46 19 0 1.37483e-19 $X=2.93 $Y=1.105
c47 15 0 1.52405e-19 $X=2.795 $Y=0.56
r48 28 30 71.0956 $w=2.7e-07 $l=3.2e-07 $layer=POLY_cond $X=2.475 $Y=1.16
+ $X2=2.795 $Y2=1.16
r49 26 28 22.2174 $w=2.7e-07 $l=1e-07 $layer=POLY_cond $X=2.375 $Y=1.16
+ $X2=2.475 $Y2=1.16
r50 25 26 22.2174 $w=2.7e-07 $l=1e-07 $layer=POLY_cond $X=2.275 $Y=1.16
+ $X2=2.375 $Y2=1.16
r51 23 25 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=2.275 $Y2=1.16
r52 18 19 29.9455 $w=1.98e-07 $l=5.4e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=3.015 $Y2=1.175
r53 18 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.475
+ $Y=1.16 $X2=2.475 $Y2=1.16
r54 17 18 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=2.475 $Y2=1.175
r55 13 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.795 $Y=1.025
+ $X2=2.795 $Y2=1.16
r56 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.795 $Y=1.025
+ $X2=2.795 $Y2=0.56
r57 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.375 $Y=1.025
+ $X2=2.375 $Y2=1.16
r58 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.375 $Y=1.025
+ $X2=2.375 $Y2=0.56
r59 5 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.275 $Y=1.295
+ $X2=2.275 $Y2=1.16
r60 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.275 $Y=1.295
+ $X2=2.275 $Y2=1.985
r61 1 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.855 $Y=1.295
+ $X2=1.855 $Y2=1.16
r62 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.855 $Y=1.295
+ $X2=1.855 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%A_27_47# 1 2 9 13 17 21 24 27 31 35 38 40
+ 41 46
c84 31 0 9.80354e-20 $X=3.485 $Y=1.16
c85 9 0 1.52405e-19 $X=3.215 $Y=0.56
r86 40 41 10.9812 $w=3.18e-07 $l=2.35e-07 $layer=LI1_cond $X=0.25 $Y=2.3
+ $X2=0.25 $Y2=2.065
r87 35 37 10.9812 $w=3.18e-07 $l=2.35e-07 $layer=LI1_cond $X=0.25 $Y=0.42
+ $X2=0.25 $Y2=0.655
r88 32 46 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.485 $Y=1.16
+ $X2=3.635 $Y2=1.16
r89 32 43 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=3.485 $Y=1.16
+ $X2=3.215 $Y2=1.16
r90 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=1.16 $X2=3.485 $Y2=1.16
r91 29 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.485 $Y=1.445
+ $X2=3.485 $Y2=1.16
r92 28 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.53
+ $X2=0.175 $Y2=1.53
r93 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.32 $Y=1.53
+ $X2=3.485 $Y2=1.445
r94 27 28 199.636 $w=1.68e-07 $l=3.06e-06 $layer=LI1_cond $X=3.32 $Y=1.53
+ $X2=0.26 $Y2=1.53
r95 25 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1.615
+ $X2=0.175 $Y2=1.53
r96 25 41 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.175 $Y=1.615
+ $X2=0.175 $Y2=2.065
r97 24 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=1.445
+ $X2=0.175 $Y2=1.53
r98 24 37 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.175 $Y=1.445
+ $X2=0.175 $Y2=0.655
r99 19 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.635 $Y=1.295
+ $X2=3.635 $Y2=1.16
r100 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.635 $Y=1.295
+ $X2=3.635 $Y2=1.985
r101 15 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.635 $Y=1.025
+ $X2=3.635 $Y2=1.16
r102 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.635 $Y=1.025
+ $X2=3.635 $Y2=0.56
r103 11 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.215 $Y=1.295
+ $X2=3.215 $Y2=1.16
r104 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.215 $Y=1.295
+ $X2=3.215 $Y2=1.985
r105 7 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.215 $Y=1.025
+ $X2=3.215 $Y2=1.16
r106 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.215 $Y=1.025
+ $X2=3.215 $Y2=0.56
r107 2 40 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r108 1 35 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%VPWR 1 2 3 4 5 18 20 24 28 30 34 36 38 40
+ 42 47 52 58 61 64 67 71
r71 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 65 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 56 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 56 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r80 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 53 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=2.72
+ $X2=2.965 $Y2=2.72
r82 53 55 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.09 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 52 70 4.41622 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.76 $Y=2.72 $X2=3.95
+ $Y2=2.72
r84 52 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 51 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r86 51 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r87 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 48 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=2.72
+ $X2=1.645 $Y2=2.72
r89 48 50 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.73 $Y=2.72
+ $X2=2.07 $Y2=2.72
r90 47 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.4 $Y=2.72
+ $X2=2.525 $Y2=2.72
r91 47 50 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.4 $Y=2.72 $X2=2.07
+ $Y2=2.72
r92 42 58 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.735 $Y2=2.72
r93 42 44 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.23 $Y2=2.72
r94 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 40 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r96 36 70 3.02162 $w=2.9e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.905 $Y=2.635
+ $X2=3.95 $Y2=2.72
r97 36 38 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.905 $Y=2.635
+ $X2=3.905 $Y2=2.34
r98 32 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=2.635
+ $X2=2.965 $Y2=2.72
r99 32 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.965 $Y=2.635
+ $X2=2.965 $Y2=2.34
r100 31 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.65 $Y=2.72
+ $X2=2.525 $Y2=2.72
r101 30 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.84 $Y=2.72
+ $X2=2.965 $Y2=2.72
r102 30 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.84 $Y=2.72
+ $X2=2.65 $Y2=2.72
r103 26 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.635
+ $X2=2.525 $Y2=2.72
r104 26 28 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.525 $Y=2.635
+ $X2=2.525 $Y2=2.34
r105 22 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.72
r106 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.34
r107 21 58 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.89 $Y=2.72
+ $X2=0.735 $Y2=2.72
r108 20 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=2.72
+ $X2=1.645 $Y2=2.72
r109 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.56 $Y=2.72
+ $X2=0.89 $Y2=2.72
r110 16 58 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=2.635
+ $X2=0.735 $Y2=2.72
r111 16 18 23.6065 $w=3.08e-07 $l=6.35e-07 $layer=LI1_cond $X=0.735 $Y=2.635
+ $X2=0.735 $Y2=2
r112 5 38 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.485 $X2=3.845 $Y2=2.34
r113 4 34 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.485 $X2=3.005 $Y2=2.34
r114 3 28 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.485 $X2=2.485 $Y2=2.34
r115 2 24 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.485 $X2=1.645 $Y2=2.34
r116 1 18 300 $w=1.7e-07 $l=2.30217e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=2.065 $X2=0.745 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%Y 1 2 3 4 15 19 21 27 30 32 34 37 38
r65 37 38 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.95 $Y=1.19
+ $X2=3.95 $Y2=1.53
r66 36 38 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.95 $Y=1.785
+ $X2=3.95 $Y2=1.53
r67 35 37 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=3.95 $Y=0.905
+ $X2=3.95 $Y2=1.19
r68 28 34 6.31926 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=3.51 $Y=1.895
+ $X2=3.385 $Y2=1.895
r69 27 36 6.83662 $w=2.2e-07 $l=1.51987e-07 $layer=LI1_cond $X=3.85 $Y=1.895
+ $X2=3.95 $Y2=1.785
r70 27 28 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=3.85 $Y=1.895
+ $X2=3.51 $Y2=1.895
r71 21 35 7.01501 $w=2.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=3.85 $Y=0.77
+ $X2=3.95 $Y2=0.905
r72 21 23 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.85 $Y=0.77
+ $X2=3.425 $Y2=0.77
r73 20 32 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.23 $Y=1.87
+ $X2=2.065 $Y2=1.895
r74 19 34 6.31926 $w=1.95e-07 $l=1.36931e-07 $layer=LI1_cond $X=3.26 $Y=1.87
+ $X2=3.385 $Y2=1.895
r75 19 20 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.26 $Y=1.87
+ $X2=2.23 $Y2=1.87
r76 16 30 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.895
+ $X2=1.225 $Y2=1.895
r77 15 32 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=1.895
+ $X2=2.065 $Y2=1.895
r78 15 16 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=1.9 $Y=1.895
+ $X2=1.39 $Y2=1.895
r79 4 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=1.485 $X2=3.425 $Y2=1.96
r80 3 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.485 $X2=2.065 $Y2=2
r81 2 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.485 $X2=1.225 $Y2=2
r82 1 23 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.235 $X2=3.425 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%VGND 1 2 9 11 15 17 19 29 30 33 36
r54 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r56 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r58 27 30 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r59 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r60 26 29 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r61 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r62 24 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.685
+ $Y2=0
r63 24 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=2.07
+ $Y2=0
r64 19 33 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.735
+ $Y2=0
r65 19 21 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.23
+ $Y2=0
r66 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r67 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r68 13 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0
r69 13 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0.38
r70 12 33 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.735
+ $Y2=0
r71 11 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.685
+ $Y2=0
r72 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=0.89
+ $Y2=0
r73 7 33 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r74 7 9 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.38
r75 2 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.235 $X2=1.645 $Y2=0.38
r76 1 9 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.745 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%A_218_47# 1 2 9 12 13 15 17
r34 13 17 6.78806 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.135 $Y=0.77 $X2=2
+ $Y2=0.77
r35 13 15 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.135 $Y=0.77
+ $X2=2.585 $Y2=0.77
r36 12 17 35.6077 $w=1.88e-07 $l=6.1e-07 $layer=LI1_cond $X=1.39 $Y=0.81 $X2=2
+ $Y2=0.81
r37 7 12 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.225 $Y=0.715
+ $X2=1.39 $Y2=0.81
r38 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.225 $Y=0.715
+ $X2=1.225 $Y2=0.38
r39 2 15 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.235 $X2=2.585 $Y2=0.72
r40 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.235 $X2=1.225 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_2%A_408_47# 1 2 3 10 16 20 23
c28 16 0 3.0481e-19 $X=3.005 $Y=0.72
r29 18 23 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=0.36 $X2=3.005
+ $Y2=0.36
r30 18 20 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.09 $Y=0.36
+ $X2=3.845 $Y2=0.36
r31 14 23 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.005 $Y=0.465
+ $X2=3.005 $Y2=0.36
r32 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.005 $Y=0.465
+ $X2=3.005 $Y2=0.72
r33 10 23 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.36 $X2=3.005
+ $Y2=0.36
r34 10 12 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=2.92 $Y=0.36
+ $X2=2.165 $Y2=0.36
r35 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.235 $X2=3.845 $Y2=0.38
r36 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.005 $Y2=0.38
r37 2 16 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.005 $Y2=0.72
r38 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.165 $Y2=0.38
.ends


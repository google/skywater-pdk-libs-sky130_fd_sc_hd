* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
M1000 Z a_27_47# a_383_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.15e+11p pd=2.63e+06u as=9.5e+11p ps=3.9e+06u
M1001 a_193_369# TE_B VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=4.428e+11p ps=4.36e+06u
M1002 a_531_47# a_193_369# VGND VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=4.2375e+11p ps=4.01e+06u
M1003 VPWR A a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1004 a_383_297# TE_B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1006 Z a_27_47# a_531_47# VNB nshort w=650000u l=150000u
+  ad=2.86e+11p pd=2.18e+06u as=0p ps=0u
M1007 a_193_369# TE_B VGND VNB nshort w=420000u l=150000u
+  ad=2.583e+11p pd=2.07e+06u as=0p ps=0u
.ends

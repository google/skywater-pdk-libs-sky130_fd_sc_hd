* File: sky130_fd_sc_hd__o31ai_1.spice.pex
* Created: Thu Aug 27 14:40:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O31AI_1%A1 1 3 6 8 14
r24 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.255 $Y=1.16
+ $X2=0.47 $Y2=1.16
r25 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r26 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r27 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r28 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r29 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%A2 1 3 6 8 9 10 11 17 18
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r39 10 11 8.80518 $w=4.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.832 $Y=1.87
+ $X2=0.832 $Y2=2.21
r40 9 10 8.80518 $w=4.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.832 $Y=1.53
+ $X2=0.832 $Y2=1.87
r41 8 9 8.80518 $w=4.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.832 $Y=1.19
+ $X2=0.832 $Y2=1.53
r42 8 18 0.776928 $w=4.43e-07 $l=3e-08 $layer=LI1_cond $X=0.832 $Y=1.19
+ $X2=0.832 $Y2=1.16
r43 4 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r44 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r45 1 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%A3 3 6 10 13 15 19
r35 14 19 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=1.46 $Y=1.2 $X2=1.58
+ $Y2=1.2
r36 13 16 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.43 $Y2=1.325
r37 13 15 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.43 $Y2=0.995
r38 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.46
+ $Y=1.16 $X2=1.46 $Y2=1.16
r39 10 19 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=1.615 $Y=1.2
+ $X2=1.58 $Y2=1.2
r40 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=1.325
r41 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.56 $X2=1.31
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%B1 3 6 8 10 12 15
r28 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.16 $X2=2.51 $Y2=1.16
r29 9 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.32 $Y=1.16 $X2=2.51
+ $Y2=1.16
r30 8 11 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.157 $Y=1.16
+ $X2=2.157 $Y2=1.325
r31 8 10 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.157 $Y=1.16
+ $X2=2.157 $Y2=0.995
r32 8 9 2.462 $w=3.3e-07 $l=1.63e-07 $layer=POLY_cond $X=2.157 $Y=1.16 $X2=2.32
+ $Y2=1.16
r33 6 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.245 $Y=1.985
+ $X2=2.245 $Y2=1.325
r34 3 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.07 $Y=0.56 $X2=2.07
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%VPWR 1 2 7 9 13 15 19 21 34
r32 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r33 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r34 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r35 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 22 30 4.98888 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=2.72 $X2=0.22
+ $Y2=2.72
r39 22 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.44 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 21 33 4.94809 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.33 $Y=2.72
+ $X2=2.545 $Y2=2.72
r41 21 27 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.33 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 19 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 19 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r44 15 18 22.7148 $w=3.43e-07 $l=6.8e-07 $layer=LI1_cond $X=2.502 $Y=1.66
+ $X2=2.502 $Y2=2.34
r45 13 33 2.94584 $w=3.45e-07 $l=1.04307e-07 $layer=LI1_cond $X=2.502 $Y=2.635
+ $X2=2.545 $Y2=2.72
r46 13 18 9.85422 $w=3.43e-07 $l=2.95e-07 $layer=LI1_cond $X=2.502 $Y=2.635
+ $X2=2.502 $Y2=2.34
r47 9 12 22.3903 $w=3.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.265 $Y=1.66
+ $X2=0.265 $Y2=2.34
r48 7 30 2.94797 $w=3.5e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.22 $Y2=2.72
r49 7 12 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.34
r50 2 18 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.485 $X2=2.495 $Y2=2.34
r51 2 15 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.485 $X2=2.495 $Y2=1.66
r52 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r53 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%Y 1 2 7 9 10 11 12 13 24
r24 22 37 6.46626 $w=2.15e-07 $l=2.83e-07 $layer=LI1_cond $X=2.052 $Y=0.825
+ $X2=2.052 $Y2=0.542
r25 22 24 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.052 $Y=0.825
+ $X2=2.052 $Y2=0.85
r26 13 42 4.12806 $w=5.63e-07 $l=1.95e-07 $layer=LI1_cond $X=2.535 $Y=0.542
+ $X2=2.34 $Y2=0.542
r27 11 12 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.052 $Y=1.87
+ $X2=2.052 $Y2=2.21
r28 11 31 12.5965 $w=2.13e-07 $l=2.35e-07 $layer=LI1_cond $X=2.052 $Y=1.87
+ $X2=2.052 $Y2=1.635
r29 10 31 5.62821 $w=2.13e-07 $l=1.05e-07 $layer=LI1_cond $X=2.052 $Y=1.53
+ $X2=2.052 $Y2=1.635
r30 9 10 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.052 $Y=1.19
+ $X2=2.052 $Y2=1.53
r31 7 42 5.60993 $w=5.63e-07 $l=2.65e-07 $layer=LI1_cond $X=2.075 $Y=0.542
+ $X2=2.34 $Y2=0.542
r32 7 37 0.486899 $w=5.63e-07 $l=2.3e-08 $layer=LI1_cond $X=2.075 $Y=0.542
+ $X2=2.052 $Y2=0.542
r33 7 9 16.6166 $w=2.13e-07 $l=3.1e-07 $layer=LI1_cond $X=2.052 $Y=0.88
+ $X2=2.052 $Y2=1.19
r34 7 24 1.60806 $w=2.13e-07 $l=3e-08 $layer=LI1_cond $X=2.052 $Y=0.88 $X2=2.052
+ $Y2=0.85
r35 2 31 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=2.03 $Y2=1.635
r36 1 42 182 $w=1.7e-07 $l=5.94559e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.34 $Y2=0.74
r37 1 42 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.34 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%VGND 1 2 7 9 13 15 17 24 25 31
r35 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r36 25 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.15
+ $Y2=0
r37 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r38 22 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r39 22 24 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=2.53 $Y2=0
r40 21 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r41 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r42 18 28 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r43 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r44 17 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r45 17 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.69
+ $Y2=0
r46 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r47 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r48 11 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r49 11 13 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.4
r50 7 28 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r51 7 9 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r52 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r53 1 9 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_1%A_109_47# 1 2 9 11 12 15
r32 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0.735
+ $X2=1.535 $Y2=0.4
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.37 $Y=0.82
+ $X2=1.535 $Y2=0.735
r34 11 12 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.37 $Y=0.82
+ $X2=0.845 $Y2=0.82
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.68 $Y=0.735
+ $X2=0.845 $Y2=0.82
r36 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.735 $X2=0.68
+ $Y2=0.4
r37 2 15 91 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.535 $Y2=0.4
r38 1 9 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__dlclkp_4.spice
* Created: Tue Sep  1 19:04:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlclkp_4.pex.spice"
.subckt sky130_fd_sc_hd__dlclkp_4  VNB VPB CLK GATE VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* GATE	GATE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_CLK_M1022_g N_A_27_47#_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_193_47#_M1011_d N_A_27_47#_M1011_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_381_47# N_GATE_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0827077 AS=0.1092 PD=0.866923 PS=1.36 NRD=40.548 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_477_413#_M1025_d N_A_27_47#_M1025_g A_381_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0513 AS=0.0708923 PD=0.645 PS=0.743077 NRD=0 NRS=47.304 M=1 R=2.4
+ SA=75000.7 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1003 A_575_47# N_A_193_47#_M1003_g N_A_477_413#_M1025_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0513 PD=0.687692 PS=0.645 NRD=38.076 NRS=1.656 M=1
+ R=2.4 SA=75001.2 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1009 N_VGND_M1009_d N_A_627_153#_M1009_g A_575_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_477_413#_M1007_g N_A_627_153#_M1007_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1020 A_1046_47# N_A_627_153#_M1020_g N_A_953_297#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=14.76 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_CLK_M1018_g A_1046_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1018_d N_A_953_297#_M1004_g N_GCLK_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.117 PD=0.92 PS=1.01 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_953_297#_M1013_g N_GCLK_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.117 PD=0.92 PS=1.01 NRD=0 NRS=15.684 M=1 R=4.33333
+ SA=75001.5 SB=75001 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1013_d N_A_953_297#_M1021_g N_GCLK_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A_953_297#_M1023_g N_GCLK_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 A_381_369# N_GATE_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116891 AS=0.1664 PD=1.17132 PS=1.8 NRD=39.2818 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_477_413#_M1006_d N_A_193_47#_M1006_g A_381_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0767094 PD=0.81 PS=0.768679 NRD=53.9386 NRS=59.8683 M=1
+ R=2.8 SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 A_585_413# N_A_27_47#_M1012_g N_A_477_413#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.2 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_627_153#_M1016_g A_585_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_477_413#_M1017_g N_A_627_153#_M1017_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.175 AS=0.26 PD=1.35 PS=2.52 NRD=1.9503 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1024 N_A_953_297#_M1024_d N_A_627_153#_M1024_g N_VPWR_M1017_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.3375 AS=0.175 PD=1.675 PS=1.35 NRD=8.8453 NRS=11.8003 M=1
+ R=6.66667 SA=75000.7 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_CLK_M1008_g N_A_953_297#_M1024_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.3375 PD=1.33 PS=1.675 NRD=4.9053 NRS=68.95 M=1 R=6.66667
+ SA=75001.5 SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_GCLK_M1001_d N_A_953_297#_M1001_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.165 PD=1.36 PS=1.33 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75002
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1002 N_GCLK_M1001_d N_A_953_297#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.135 PD=1.36 PS=1.27 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75002.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1015 N_GCLK_M1015_d N_A_953_297#_M1015_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1019 N_GCLK_M1015_d N_A_953_297#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=13.161 P=19.61
c_82 VNB 0 7.84261e-20 $X=0.15 $Y=-0.085
c_163 VPB 0 1.43275e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__dlclkp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__dfstp_1.spice.pex
* Created: Thu Aug 27 14:15:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFSTP_1%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.265 $Y=1.19
+ $X2=0.265 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_27_47# 1 2 9 13 15 17 20 24 28 31 35 36 37
+ 40 42 46 47 50 51 52 54 55 59 61 62 63 64 73 78 85 86 92 93 96
c275 92 0 3.09108e-19 $X=5.175 $Y=1.74
c276 73 0 1.6788e-19 $X=5.335 $Y=1.87
c277 52 0 3.02058e-20 $X=5.07 $Y=0.81
c278 47 0 9.71454e-20 $X=2.435 $Y=0.87
c279 46 0 1.76471e-19 $X=2.435 $Y=0.87
c280 40 0 1.81794e-19 $X=0.725 $Y=1.795
c281 37 0 3.29888e-20 $X=0.61 $Y=1.88
c282 24 0 7.39505e-20 $X=5.085 $Y=2.275
r283 93 104 7.06336 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.175 $Y=1.81
+ $X2=4.985 $Y2=1.81
r284 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.74 $X2=5.175 $Y2=1.74
r285 89 92 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.085 $Y=1.74
+ $X2=5.175 $Y2=1.74
r286 85 88 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.74
+ $X2=2.765 $Y2=1.875
r287 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.74 $X2=2.765 $Y2=1.74
r288 73 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.335 $Y=1.87
+ $X2=5.335 $Y2=1.87
r289 71 86 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=2.555 $Y=1.765
+ $X2=2.765 $Y2=1.765
r290 71 99 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.555 $Y=1.765
+ $X2=2.46 $Y2=1.765
r291 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.87
+ $X2=2.555 $Y2=1.87
r292 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.87
+ $X2=0.695 $Y2=1.87
r293 64 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.7 $Y=1.87
+ $X2=2.555 $Y2=1.87
r294 63 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.19 $Y=1.87
+ $X2=5.335 $Y2=1.87
r295 63 64 3.08168 $w=1.4e-07 $l=2.49e-06 $layer=MET1_cond $X=5.19 $Y=1.87
+ $X2=2.7 $Y2=1.87
r296 62 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.87
+ $X2=0.695 $Y2=1.87
r297 61 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=2.555 $Y2=1.87
r298 61 62 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=0.84 $Y2=1.87
r299 59 96 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=0.93
+ $X2=5.985 $Y2=0.765
r300 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=0.93 $X2=5.985 $Y2=0.93
r301 55 58 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.985 $Y=0.81
+ $X2=5.985 $Y2=0.93
r302 51 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.985 $Y2=0.81
r303 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.07 $Y2=0.81
r304 50 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=1.655
+ $X2=4.985 $Y2=1.81
r305 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.985 $Y=0.895
+ $X2=5.07 $Y2=0.81
r306 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.985 $Y=0.895
+ $X2=4.985 $Y2=1.655
r307 47 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.435 $Y=0.87
+ $X2=2.305 $Y2=0.87
r308 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=0.87 $X2=2.435 $Y2=0.87
r309 44 99 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=1.765
r310 44 46 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=0.87
r311 43 78 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r312 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r313 40 67 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r314 40 42 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r315 39 42 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r316 38 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r317 37 67 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r318 37 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r319 35 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r320 35 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r321 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r322 29 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r323 28 96 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.045 $Y=0.445
+ $X2=6.045 $Y2=0.765
r324 22 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.085 $Y=1.875
+ $X2=5.085 $Y2=1.74
r325 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.085 $Y=1.875
+ $X2=5.085 $Y2=2.275
r326 20 88 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.875
r327 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r328 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r329 11 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r330 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r331 7 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r332 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r333 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r334 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%D 3 7 9 10 14 15
c39 14 0 1.34441e-19 $X=1.855 $Y=1.17
c40 7 0 1.76471e-19 $X=1.83 $Y=2.065
r41 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.335
r42 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.005
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.17 $X2=1.855 $Y2=1.17
r44 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.53
r45 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.17
r46 7 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.83 $Y=2.065
+ $X2=1.83 $Y2=1.335
r47 3 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.83 $Y=0.555
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_193_47# 1 2 9 11 12 15 18 21 23 25 28 29
+ 30 32 33 34 41 45 46 53 54 58
c195 46 0 4.49853e-20 $X=5.335 $Y=1.19
c196 45 0 2.33963e-19 $X=5.335 $Y=1.19
c197 33 0 1.51904e-19 $X=5.19 $Y=1.19
c198 32 0 9.71454e-20 $X=3.052 $Y=1.12
c199 25 0 1.80017e-19 $X=5.625 $Y=2.275
c200 9 0 4.43992e-20 $X=2.315 $Y=2.275
r201 53 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=1.095
r202 53 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=0.765
r203 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=0.93 $X2=2.915 $Y2=0.93
r204 46 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.335
+ $Y=1.26 $X2=5.335 $Y2=1.26
r205 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.335 $Y=1.19
+ $X2=5.335 $Y2=1.19
r206 41 43 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=3.015 $Y=0.85
+ $X2=3.015 $Y2=0.965
r207 41 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=0.85
+ $X2=3.015 $Y2=0.85
r208 37 62 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r209 37 58 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r210 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=0.85
+ $X2=1.155 $Y2=0.85
r211 33 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.19 $Y=1.19
+ $X2=5.335 $Y2=1.19
r212 33 34 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=5.19 $Y=1.19
+ $X2=3.16 $Y2=1.19
r213 32 34 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.052 $Y=1.12
+ $X2=3.16 $Y2=1.19
r214 32 43 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=3.052 $Y=1.12
+ $X2=3.052 $Y2=0.965
r215 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=0.85
+ $X2=1.155 $Y2=0.85
r216 29 41 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=0.85
+ $X2=3.015 $Y2=0.85
r217 29 30 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.87 $Y=0.85
+ $X2=1.3 $Y2=0.85
r218 28 49 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=5.49 $Y=1.26
+ $X2=5.335 $Y2=1.26
r219 23 28 54.3623 $w=1.77e-07 $l=2.09464e-07 $layer=POLY_cond $X=5.625 $Y=1.455
+ $X2=5.595 $Y2=1.26
r220 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.625 $Y=1.455
+ $X2=5.625 $Y2=2.275
r221 19 28 38.0233 $w=1.77e-07 $l=1.49248e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.595 $Y2=1.26
r222 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.565 $Y2=0.445
r223 18 56 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.855 $Y=1.245
+ $X2=2.855 $Y2=1.095
r224 15 55 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.855 $Y=0.415
+ $X2=2.855 $Y2=0.765
r225 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.855 $Y2=1.245
r226 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.39 $Y2=1.32
r227 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.39 $Y2=1.32
r228 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.315 $Y2=2.275
r229 2 62 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r230 1 58 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_652_21# 1 2 9 13 15 19 21 25 28 30 31 35
+ 38
c115 38 0 1.31911e-19 $X=4.635 $Y=0.895
c116 35 0 2.11834e-19 $X=4.075 $Y=1.96
c117 28 0 3.26119e-19 $X=4.635 $Y=1.835
c118 21 0 1.80719e-19 $X=4.54 $Y=1.96
r119 36 38 6.77908 $w=3.38e-07 $l=2e-07 $layer=LI1_cond $X=4.435 $Y=0.895
+ $X2=4.635 $Y2=0.895
r120 31 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.905
r121 31 41 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.575
r122 30 33 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=3.485 $Y=1.74
+ $X2=3.485 $Y2=1.96
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.74 $X2=3.445 $Y2=1.74
r124 27 38 4.14298 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=4.635 $Y=1.065
+ $X2=4.635 $Y2=0.895
r125 27 28 44.9474 $w=1.88e-07 $l=7.7e-07 $layer=LI1_cond $X=4.635 $Y=1.065
+ $X2=4.635 $Y2=1.835
r126 23 36 2.53954 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.895
r127 23 25 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.46
r128 22 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.96
+ $X2=4.075 $Y2=1.96
r129 21 28 6.98266 $w=2.5e-07 $l=1.65831e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.635 $Y2=1.835
r130 21 22 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.16 $Y2=1.96
r131 17 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=1.96
r132 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=2.21
r133 16 33 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.61 $Y=1.96
+ $X2=3.485 $Y2=1.96
r134 15 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=4.075 $Y2=1.96
r135 15 16 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=3.61 $Y2=1.96
r136 13 42 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.335 $Y=2.275
+ $X2=3.335 $Y2=1.905
r137 9 41 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.335 $Y=0.445
+ $X2=3.335 $Y2=1.575
r138 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.065 $X2=4.075 $Y2=2.21
r139 1 25 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.235 $X2=4.475 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%SET_B 1 3 7 11 17 19 20 24 26 27 29 30 36 37
c135 36 0 1.54133e-19 $X=7.195 $Y=0.85
c136 29 0 2.74106e-19 $X=7.05 $Y=0.85
c137 26 0 1.49785e-19 $X=7.01 $Y=0.9
c138 19 0 1.13471e-19 $X=6.915 $Y=1.535
c139 1 0 9.38739e-20 $X=3.865 $Y=1.145
r140 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.195 $Y=0.85
+ $X2=7.195 $Y2=0.85
r141 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.08 $Y=0.85
+ $X2=3.935 $Y2=0.85
r142 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.05 $Y=0.85
+ $X2=7.195 $Y2=0.85
r143 29 30 3.67574 $w=1.4e-07 $l=2.97e-06 $layer=MET1_cond $X=7.05 $Y=0.85
+ $X2=4.08 $Y2=0.85
r144 27 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=0.98 $X2=3.775 $Y2=0.98
r145 27 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=0.85
+ $X2=3.935 $Y2=0.85
r146 26 37 7.89637 $w=2.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.01 $Y=0.87
+ $X2=7.195 $Y2=0.87
r147 24 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=0.98
+ $X2=6.845 $Y2=1.145
r148 24 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=0.98
+ $X2=6.845 $Y2=0.815
r149 23 26 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=0.9
+ $X2=7.01 $Y2=0.9
r150 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.845
+ $Y=0.98 $X2=6.845 $Y2=0.98
r151 19 20 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=6.915 $Y=1.535
+ $X2=6.915 $Y2=1.685
r152 19 44 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.905 $Y=1.535
+ $X2=6.905 $Y2=1.145
r153 17 20 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.925 $Y=2.275
+ $X2=6.925 $Y2=1.685
r154 11 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.785 $Y=0.445
+ $X2=6.785 $Y2=0.815
r155 5 40 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.81 $Y2=0.98
r156 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.905 $Y2=0.445
r157 1 40 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.81 $Y2=0.98
r158 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.865 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_476_47# 1 2 7 9 11 14 16 20 22 24 25 26 30
+ 35 37 38 43 44 53
c158 53 0 1.57127e-19 $X=4.705 $Y=1.4
c159 43 0 4.43992e-20 $X=3.44 $Y=1.3
c160 22 0 3.80375e-20 $X=5.205 $Y=0.735
c161 16 0 1.05575e-19 $X=5.13 $Y=0.825
c162 7 0 3.02058e-20 $X=4.265 $Y=0.735
r163 48 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.705 $Y2=1.4
r164 48 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.265 $Y2=1.4
r165 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.4 $X2=4.285 $Y2=1.4
r166 44 47 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.245 $Y=1.32
+ $X2=4.245 $Y2=1.4
r167 42 43 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=1.3
+ $X2=3.44 $Y2=1.3
r168 40 42 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=3.105 $Y=1.3
+ $X2=3.355 $Y2=1.3
r169 38 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=4.245 $Y2=1.32
r170 38 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=3.44 $Y2=1.32
r171 37 42 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.355 $Y=1.195
+ $X2=3.355 $Y2=1.3
r172 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.355 $Y=0.465
+ $X2=3.355 $Y2=1.195
r173 34 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=1.3
r174 34 35 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=2.25
r175 30 36 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=3.355 $Y2=0.465
r176 30 32 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=2.59 $Y2=0.365
r177 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=3.105 $Y2=2.25
r178 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=2.525 $Y2=2.335
r179 22 24 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.205 $Y=0.735
+ $X2=5.205 $Y2=0.445
r180 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=1.4
r181 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=2.275
r182 17 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.34 $Y=0.825
+ $X2=4.265 $Y2=0.825
r183 16 22 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=5.205 $Y2=0.735
r184 16 17 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=4.34 $Y2=0.825
r185 12 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=1.4
r186 12 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=2.275
r187 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.235
+ $X2=4.265 $Y2=1.4
r188 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=0.825
r189 10 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=1.235
r190 7 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.825
r191 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.445
r192 2 28 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.065 $X2=2.525 $Y2=2.335
r193 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_1182_261# 1 2 9 13 18 21 25 29 32 36 39 40
c80 39 0 1.80017e-19 $X=7.53 $Y=1.67
c81 32 0 1.13471e-19 $X=7.755 $Y=1.575
c82 18 0 6.36548e-20 $X=6.405 $Y=1.38
r83 38 40 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=7.615 $Y=1.67
+ $X2=7.755 $Y2=1.67
r84 38 39 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=1.67
+ $X2=7.53 $Y2=1.67
r85 34 36 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.615 $Y=0.515
+ $X2=7.755 $Y2=0.515
r86 32 40 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=7.755 $Y=1.575
+ $X2=7.755 $Y2=1.67
r87 31 36 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=0.68
+ $X2=7.755 $Y2=0.515
r88 31 32 52.244 $w=1.88e-07 $l=8.95e-07 $layer=LI1_cond $X=7.755 $Y=0.68
+ $X2=7.755 $Y2=1.575
r89 27 38 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.615 $Y=1.765
+ $X2=7.615 $Y2=1.67
r90 27 29 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.615 $Y=1.765
+ $X2=7.615 $Y2=1.87
r91 24 39 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=6.095 $Y=1.66
+ $X2=7.53 $Y2=1.66
r92 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.095
+ $Y=1.66 $X2=6.095 $Y2=1.66
r93 20 25 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=6.07 $Y=1.665
+ $X2=6.07 $Y2=1.66
r94 20 21 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=6.07 $Y=1.665
+ $X2=6.07 $Y2=1.825
r95 16 25 36.9668 $w=3.2e-07 $l=2.05e-07 $layer=POLY_cond $X=6.07 $Y=1.455
+ $X2=6.07 $Y2=1.66
r96 16 18 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.07 $Y=1.38
+ $X2=6.405 $Y2=1.38
r97 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=1.38
r98 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=0.445
r99 9 21 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.985 $Y=2.275
+ $X2=5.985 $Y2=1.825
r100 2 29 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=7.48
+ $Y=1.645 $X2=7.615 $Y2=1.87
r101 1 34 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=7.48
+ $Y=0.235 $X2=7.615 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_1032_413# 1 2 3 12 16 18 22 26 28 29 34 35
+ 39 40 41 44 49 51 54 56 57 58
c164 54 0 9.39049e-20 $X=6.405 $Y=1.32
c165 34 0 7.39505e-20 $X=5.675 $Y=1.915
r166 56 58 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.325 $Y=1.29
+ $X2=7.16 $Y2=1.29
r167 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.325
+ $Y=1.26 $X2=7.325 $Y2=1.26
r168 47 49 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=6.68 $Y=2.085
+ $X2=6.68 $Y2=2.21
r169 46 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=6.405 $Y2=1.32
r170 46 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=7.16 $Y2=1.32
r171 44 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.235
+ $X2=6.405 $Y2=1.32
r172 43 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.405 $Y=0.475
+ $X2=6.405 $Y2=1.235
r173 42 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2 $X2=5.675
+ $Y2=2
r174 41 47 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=6.56 $Y=2
+ $X2=6.68 $Y2=2.085
r175 41 42 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.56 $Y=2 $X2=5.76
+ $Y2=2
r176 39 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=6.405 $Y2=1.32
r177 39 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=5.76 $Y2=1.32
r178 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=6.405 $Y2=0.475
r179 35 37 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=5.805 $Y2=0.39
r180 34 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.915
+ $X2=5.675 $Y2=2
r181 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=1.405
+ $X2=5.76 $Y2=1.32
r182 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.675 $Y=1.405
+ $X2=5.675 $Y2=1.915
r183 29 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.675 $Y=2.29
+ $X2=5.675 $Y2=2
r184 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.59 $Y=2.29
+ $X2=5.295 $Y2=2.29
r185 24 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.345 $Y=1.425
+ $X2=8.345 $Y2=1.26
r186 24 26 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.345 $Y=1.425
+ $X2=8.345 $Y2=2.165
r187 20 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.345 $Y=1.095
+ $X2=8.345 $Y2=1.26
r188 20 22 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=8.345 $Y=1.095
+ $X2=8.345 $Y2=0.445
r189 19 57 5.03009 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.48 $Y=1.26
+ $X2=7.335 $Y2=1.26
r190 18 28 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.27 $Y=1.26
+ $X2=8.345 $Y2=1.26
r191 18 19 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=8.27 $Y=1.26
+ $X2=7.48 $Y2=1.26
r192 14 57 37.0704 $w=1.5e-07 $l=1.96914e-07 $layer=POLY_cond $X=7.405 $Y=1.425
+ $X2=7.335 $Y2=1.26
r193 14 16 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.405 $Y=1.425
+ $X2=7.405 $Y2=2.065
r194 10 57 37.0704 $w=1.5e-07 $l=1.96914e-07 $layer=POLY_cond $X=7.405 $Y=1.095
+ $X2=7.335 $Y2=1.26
r195 10 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.405 $Y=1.095
+ $X2=7.405 $Y2=0.505
r196 3 49 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.59
+ $Y=2.065 $X2=6.715 $Y2=2.21
r197 2 31 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=5.16
+ $Y=2.065 $X2=5.295 $Y2=2.33
r198 1 37 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.805 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_1602_47# 1 2 9 12 18 24 25 28 29 30 32
r56 28 29 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.135 $Y=2 $X2=8.135
+ $Y2=1.915
r57 25 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=1.16
+ $X2=8.765 $Y2=1.325
r58 25 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=1.16
+ $X2=8.765 $Y2=0.995
r59 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.765
+ $Y=1.16 $X2=8.765 $Y2=1.16
r60 22 30 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=8.3 $Y=1.16
+ $X2=8.175 $Y2=1.16
r61 22 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.3 $Y=1.16
+ $X2=8.765 $Y2=1.16
r62 20 30 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=1.325
+ $X2=8.175 $Y2=1.16
r63 20 29 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=8.175 $Y=1.325
+ $X2=8.175 $Y2=1.915
r64 16 30 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=0.995
+ $X2=8.175 $Y2=1.16
r65 16 18 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=8.175 $Y=0.995
+ $X2=8.175 $Y2=0.51
r66 12 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.82 $Y=1.985
+ $X2=8.82 $Y2=1.325
r67 9 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.82 $Y=0.56 $X2=8.82
+ $Y2=0.995
r68 2 28 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=8.01
+ $Y=1.845 $X2=8.135 $Y2=2
r69 1 18 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=8.01
+ $Y=0.235 $X2=8.135 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%VPWR 1 2 3 4 5 6 7 24 28 30 34 38 42 44 46
+ 48 54 59 64 72 77 84 85 88 91 94 101 104 111 114
c165 85 0 1.81794e-19 $X=9.43 $Y=2.72
c166 1 0 3.29888e-20 $X=0.545 $Y=1.815
r167 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r168 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r169 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r170 104 107 10.4269 $w=4.18e-07 $l=3.8e-07 $layer=LI1_cond $X=6.15 $Y=2.34
+ $X2=6.15 $Y2=2.72
r171 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r172 98 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r173 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r174 94 97 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.62 $Y=2.34
+ $X2=3.62 $Y2=2.72
r175 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r176 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r177 85 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.51 $Y2=2.72
r178 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r179 82 114 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=8.765 $Y=2.72
+ $X2=8.622 $Y2=2.72
r180 82 84 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.765 $Y=2.72
+ $X2=9.43 $Y2=2.72
r181 81 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r182 81 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r183 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r184 78 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.36 $Y=2.72
+ $X2=7.195 $Y2=2.72
r185 78 80 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.36 $Y=2.72
+ $X2=7.59 $Y2=2.72
r186 77 114 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=8.48 $Y=2.72
+ $X2=8.622 $Y2=2.72
r187 77 80 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=8.48 $Y=2.72
+ $X2=7.59 $Y2=2.72
r188 76 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r189 76 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r190 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r191 73 107 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.15 $Y2=2.72
r192 73 75 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.67 $Y2=2.72
r193 72 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.03 $Y=2.72
+ $X2=7.195 $Y2=2.72
r194 72 75 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.03 $Y=2.72
+ $X2=6.67 $Y2=2.72
r195 71 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r196 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r197 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r198 68 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r199 67 70 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r200 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r201 65 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.495 $Y2=2.72
r202 65 67 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.83 $Y2=2.72
r203 64 107 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.94 $Y=2.72
+ $X2=6.15 $Y2=2.72
r204 64 70 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.94 $Y=2.72
+ $X2=5.75 $Y2=2.72
r205 63 98 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r206 63 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r207 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r208 60 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r209 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r210 59 97 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=3.62 $Y2=2.72
r211 59 62 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=2.07 $Y2=2.72
r212 58 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r213 58 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r214 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r215 55 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r216 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r217 54 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r218 54 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r219 48 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r220 46 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r221 44 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r222 44 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r223 40 114 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.622 $Y=2.635
+ $X2=8.622 $Y2=2.72
r224 40 42 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=8.622 $Y=2.635
+ $X2=8.622 $Y2=2
r225 36 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=2.635
+ $X2=7.195 $Y2=2.72
r226 36 38 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.195 $Y=2.635
+ $X2=7.195 $Y2=2.21
r227 32 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.72
r228 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.34
r229 31 97 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.81 $Y=2.72
+ $X2=3.62 $Y2=2.72
r230 30 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=4.495 $Y2=2.72
r231 30 31 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=3.81 $Y2=2.72
r232 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r233 26 28 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.22
r234 22 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r235 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r236 7 42 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=8.42
+ $Y=1.845 $X2=8.61 $Y2=2
r237 6 38 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=7
+ $Y=2.065 $X2=7.195 $Y2=2.21
r238 5 104 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.06
+ $Y=2.065 $X2=6.195 $Y2=2.34
r239 4 34 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.065 $X2=4.495 $Y2=2.34
r240 3 94 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.065 $X2=3.595 $Y2=2.34
r241 2 28 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.645 $X2=1.62 $Y2=2.22
r242 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%A_381_47# 1 2 8 9 10 11 12 15 20
c59 20 0 1.34441e-19 $X=2.04 $Y=1.96
r60 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r61 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.88
r62 11 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.6 $Y2=1.88
r63 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r64 9 10 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.6 $Y2=0.73
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.795
+ $X2=1.6 $Y2=1.88
r66 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.6 $Y2=0.73
r67 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.515 $Y2=1.795
r68 2 20 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.645 $X2=2.04 $Y2=1.96
r69 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%Q 1 2 10 11 12 13 14 15
r16 14 15 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=9.072 $Y=1.82
+ $X2=9.072 $Y2=2.21
r17 13 23 5.42326 $w=2.53e-07 $l=1.2e-07 $layer=LI1_cond $X=9.072 $Y=0.51
+ $X2=9.072 $Y2=0.63
r18 11 14 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=9.072 $Y=1.782
+ $X2=9.072 $Y2=1.82
r19 11 12 6.75127 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=9.072 $Y=1.782
+ $X2=9.072 $Y2=1.655
r20 10 12 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=9.11 $Y=0.795
+ $X2=9.11 $Y2=1.655
r21 9 23 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=9.072 $Y=0.668
+ $X2=9.072 $Y2=0.63
r22 9 10 6.75127 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=9.072 $Y=0.668
+ $X2=9.072 $Y2=0.795
r23 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=8.895
+ $Y=1.485 $X2=9.03 $Y2=1.82
r24 1 23 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=8.895
+ $Y=0.235 $X2=9.03 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_1%VGND 1 2 3 4 5 6 21 25 29 31 35 39 41 43 45
+ 51 56 72 79 80 83 86 89 92 96 100 102
c148 96 0 1.49785e-19 $X=6.69 $Y=0.24
c149 80 0 2.71124e-20 $X=9.43 $Y=0
r150 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r151 98 100 11.494 $w=6.48e-07 $l=2.2e-07 $layer=LI1_cond $X=7.13 $Y=0.24
+ $X2=7.35 $Y2=0.24
r152 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r153 95 98 0.644042 $w=6.48e-07 $l=3.5e-08 $layer=LI1_cond $X=7.095 $Y=0.24
+ $X2=7.13 $Y2=0.24
r154 95 96 14.8982 $w=6.48e-07 $l=4.05e-07 $layer=LI1_cond $X=7.095 $Y=0.24
+ $X2=6.69 $Y2=0.24
r155 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r156 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r157 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r158 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r159 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r160 80 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.51 $Y2=0
r161 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r162 77 102 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=8.765 $Y=0
+ $X2=8.622 $Y2=0
r163 77 79 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.765 $Y=0 $X2=9.43
+ $Y2=0
r164 76 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r165 76 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r166 75 100 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.59 $Y=0 $X2=7.35
+ $Y2=0
r167 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r168 72 102 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=8.48 $Y=0
+ $X2=8.622 $Y2=0
r169 72 75 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=8.48 $Y=0 $X2=7.59
+ $Y2=0
r170 71 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r171 70 96 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.69
+ $Y2=0
r172 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r173 68 71 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r174 68 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r175 67 70 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=6.67
+ $Y2=0
r176 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r177 65 92 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.92
+ $Y2=0
r178 65 67 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.29
+ $Y2=0
r179 63 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r180 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r181 60 63 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r182 60 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r183 59 62 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r184 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r185 57 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r186 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r187 56 89 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.815
+ $Y2=0
r188 56 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.45
+ $Y2=0
r189 55 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r190 55 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r191 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r192 52 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r193 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r194 51 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r195 51 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r196 45 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r197 43 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r198 41 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r199 41 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r200 37 102 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.622 $Y=0.085
+ $X2=8.622 $Y2=0
r201 37 39 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=8.622 $Y=0.085
+ $X2=8.622 $Y2=0.38
r202 33 92 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=0.085
+ $X2=4.92 $Y2=0
r203 33 35 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=4.92 $Y=0.085
+ $X2=4.92 $Y2=0.38
r204 32 89 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=3.815
+ $Y2=0
r205 31 92 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.76 $Y=0 $X2=4.92
+ $Y2=0
r206 31 32 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.76 $Y=0 $X2=4.02
+ $Y2=0
r207 27 89 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r208 27 29 7.7298 $w=4.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.36
r209 23 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r210 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.38
r211 19 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r212 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r213 6 39 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=8.42
+ $Y=0.235 $X2=8.61 $Y2=0.38
r214 5 95 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=6.86
+ $Y=0.235 $X2=7.095 $Y2=0.48
r215 4 35 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=4.995 $Y2=0.38
r216 3 29 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.235 $X2=3.695 $Y2=0.36
r217 2 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r218 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__and4b_4.pex.spice
* Created: Tue Sep  1 18:58:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4B_4%A_N 3 7 9 10 11 16
c34 7 0 1.68659e-19 $X=0.47 $Y=2.275
c35 3 0 1.33943e-19 $X=0.47 $Y=0.445
r36 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.16
+ $X2=0.525 $Y2=1.325
r37 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.16
+ $X2=0.525 $Y2=0.995
r38 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.16 $X2=0.525 $Y2=1.16
r39 10 11 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.615 $Y=1.19
+ $X2=0.615 $Y2=1.53
r40 10 17 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.615 $Y=1.19
+ $X2=0.615 $Y2=1.16
r41 9 17 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.615 $Y=0.85
+ $X2=0.615 $Y2=1.16
r42 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r43 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%A_174_21# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 45 47 49 50 51 52 56 59 60 61 62
r145 71 72 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.785 $Y=1.16
+ $X2=2.205 $Y2=1.16
r146 67 69 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.945 $Y=1.16
+ $X2=1.365 $Y2=1.16
r147 60 61 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=4.39 $Y=0.385
+ $X2=2.965 $Y2=0.385
r148 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.88 $Y=0.47
+ $X2=2.965 $Y2=0.385
r149 58 59 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.88 $Y=0.47
+ $X2=2.88 $Y2=0.615
r150 54 56 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.22 $Y=1.63
+ $X2=4.38 $Y2=1.63
r151 52 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.55 $Y=1.63
+ $X2=3.22 $Y2=1.63
r152 50 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.795 $Y=0.7
+ $X2=2.88 $Y2=0.615
r153 50 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.795 $Y=0.7
+ $X2=2.55 $Y2=0.7
r154 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=1.545
+ $X2=2.55 $Y2=1.63
r155 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.245
+ $X2=2.465 $Y2=1.16
r156 48 49 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.465 $Y=1.245
+ $X2=2.465 $Y2=1.545
r157 47 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.075
+ $X2=2.465 $Y2=1.16
r158 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=0.785
+ $X2=2.55 $Y2=0.7
r159 46 47 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.465 $Y=0.785
+ $X2=2.465 $Y2=1.075
r160 45 72 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.285 $Y=1.16
+ $X2=2.205 $Y2=1.16
r161 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=1.16 $X2=2.285 $Y2=1.16
r162 41 71 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.605 $Y=1.16
+ $X2=1.785 $Y2=1.16
r163 41 69 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.605 $Y=1.16
+ $X2=1.365 $Y2=1.16
r164 40 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=1.16
+ $X2=2.285 $Y2=1.16
r165 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.16 $X2=1.605 $Y2=1.16
r166 38 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=1.16
+ $X2=2.465 $Y2=1.16
r167 38 44 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.38 $Y=1.16
+ $X2=2.285 $Y2=1.16
r168 34 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.325
+ $X2=2.205 $Y2=1.16
r169 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.205 $Y=1.325
+ $X2=2.205 $Y2=1.985
r170 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=0.995
+ $X2=2.205 $Y2=1.16
r171 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.205 $Y=0.995
+ $X2=2.205 $Y2=0.56
r172 27 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.16
r173 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.985
r174 24 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=0.995
+ $X2=1.785 $Y2=1.16
r175 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.785 $Y=0.995
+ $X2=1.785 $Y2=0.56
r176 20 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.16
r177 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.985
r178 17 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=1.16
r179 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=0.56
r180 13 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.325
+ $X2=0.945 $Y2=1.16
r181 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.945 $Y=1.325
+ $X2=0.945 $Y2=1.985
r182 10 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=1.16
r183 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r184 3 56 600 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=4.075
+ $Y=1.485 $X2=4.38 $Y2=1.63
r185 2 54 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.63
r186 1 60 91 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=2 $X=4.665
+ $Y=0.235 $X2=4.8 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%D 3 6 8 11 13
c42 8 0 1.34065e-19 $X=2.995 $Y=1.19
r43 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.16
+ $X2=2.95 $Y2=1.325
r44 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.16
+ $X2=2.95 $Y2=0.995
r45 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r46 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.985
+ $X2=3.01 $Y2=1.325
r47 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.56 $X2=3.01
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%C 1 3 6 8 9 13
r35 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.16 $X2=3.43 $Y2=1.16
r36 8 9 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=3.45 $Y=0.85 $X2=3.45
+ $Y2=1.16
r37 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r38 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325 $X2=3.43
+ $Y2=1.985
r39 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995 $X2=3.43
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%B 3 6 8 9 13 15
r36 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.16
+ $X2=4.06 $Y2=1.325
r37 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.16
+ $X2=4.06 $Y2=0.995
r38 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.16 $X2=4.06 $Y2=1.16
r39 9 14 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.98 $Y=1.19 $X2=3.98
+ $Y2=1.16
r40 8 14 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.98 $Y=0.85 $X2=3.98
+ $Y2=1.16
r41 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4 $Y=1.985 $X2=4
+ $Y2=1.325
r42 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4 $Y=0.56 $X2=4
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%A_27_47# 1 2 7 9 12 15 18 20 24 25 28 31
r76 28 30 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.42
+ $X2=0.215 $Y2=0.585
r77 25 32 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.815 $Y=1.16
+ $X2=4.59 $Y2=1.16
r78 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.815
+ $Y=1.16 $X2=4.815 $Y2=1.16
r79 22 24 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.815 $Y=1.915
+ $X2=4.815 $Y2=1.16
r80 21 31 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.215
+ $Y2=2
r81 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.73 $Y=2
+ $X2=4.815 $Y2=1.915
r82 20 21 286.08 $w=1.68e-07 $l=4.385e-06 $layer=LI1_cond $X=4.73 $Y=2 $X2=0.345
+ $Y2=2
r83 16 31 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2
r84 16 18 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2.3
r85 15 31 4.18896 $w=2.17e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.215 $Y2=2
r86 15 30 84.2909 $w=1.73e-07 $l=1.33e-06 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.172 $Y2=0.585
r87 10 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.16
r88 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.985
r89 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=1.16
r90 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.59 $Y=0.995 $X2=4.59
+ $Y2=0.56
r91 2 18 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r92 1 28 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%VPWR 1 2 3 4 5 18 22 26 30 32 34 37 38 39 41
+ 46 51 60 65 68 71 75
r79 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r80 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r81 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r82 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 63 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 60 74 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=4.635 $Y=2.72
+ $X2=4.847 $Y2=2.72
r86 60 62 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.635 $Y=2.72
+ $X2=4.37 $Y2=2.72
r87 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r88 59 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r90 56 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=2.72
+ $X2=2.415 $Y2=2.72
r91 56 58 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.58 $Y=2.72
+ $X2=3.45 $Y2=2.72
r92 55 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r93 55 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r95 52 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=1.575 $Y2=2.72
r96 52 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=2.07 $Y2=2.72
r97 51 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.415 $Y2=2.72
r98 51 54 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.07 $Y2=2.72
r99 50 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r100 50 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r101 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r103 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r104 46 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.575 $Y2=2.72
r105 46 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 41 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r107 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r108 39 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r109 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r110 37 58 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.45 $Y2=2.72
r111 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.64 $Y2=2.72
r112 36 62 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=4.37 $Y2=2.72
r113 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.64 $Y2=2.72
r114 32 74 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=4.8 $Y=2.635
+ $X2=4.847 $Y2=2.72
r115 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.8 $Y=2.635
+ $X2=4.8 $Y2=2.34
r116 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.635
+ $X2=3.64 $Y2=2.72
r117 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.64 $Y=2.635
+ $X2=3.64 $Y2=2.34
r118 24 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.72
r119 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.34
r120 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.72
r121 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.34
r122 16 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r123 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r124 5 34 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=1.485 $X2=4.8 $Y2=2.34
r125 4 30 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=2.34
r126 3 26 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.485 $X2=2.415 $Y2=2.34
r127 2 22 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.485 $X2=1.575 $Y2=2.34
r128 1 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%X 1 2 3 4 15 17 21 25 27 28 29 36 38 44
c46 38 0 3.02602e-19 $X=1.155 $Y=0.85
r47 36 44 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.12 $Y=1.545
+ $X2=1.12 $Y2=1.53
r48 35 38 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=1.12 $Y=0.82 $X2=1.12
+ $Y2=0.85
r49 29 36 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.63 $X2=1.12
+ $Y2=1.545
r50 29 44 1.44055 $w=2.78e-07 $l=3.5e-08 $layer=LI1_cond $X=1.12 $Y=1.495
+ $X2=1.12 $Y2=1.53
r51 28 29 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=1.19
+ $X2=1.12 $Y2=1.495
r52 27 35 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.735
+ $X2=1.12 $Y2=0.82
r53 27 28 12.8827 $w=2.78e-07 $l=3.13e-07 $layer=LI1_cond $X=1.12 $Y=0.877
+ $X2=1.12 $Y2=1.19
r54 27 38 1.11128 $w=2.78e-07 $l=2.7e-08 $layer=LI1_cond $X=1.12 $Y=0.877
+ $X2=1.12 $Y2=0.85
r55 23 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.995 $Y=0.65
+ $X2=1.995 $Y2=0.42
r56 19 29 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.26 $Y=1.63 $X2=1.12
+ $Y2=1.63
r57 19 21 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.26 $Y=1.63
+ $X2=1.995 $Y2=1.63
r58 18 27 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.26 $Y=0.735
+ $X2=1.12 $Y2=0.735
r59 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.91 $Y=0.735
+ $X2=1.995 $Y2=0.65
r60 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.91 $Y=0.735
+ $X2=1.26 $Y2=0.735
r61 13 27 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=1.155 $Y=0.65
+ $X2=1.12 $Y2=0.735
r62 13 15 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.155 $Y=0.65
+ $X2=1.155 $Y2=0.42
r63 4 21 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.485 $X2=1.995 $Y2=1.63
r64 3 29 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.485 $X2=1.155 $Y2=1.63
r65 2 25 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=1.995 $Y2=0.42
r66 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_4%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r79 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r80 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r81 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r82 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r83 42 45 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=4.83
+ $Y2=0
r84 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r85 41 44 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.83
+ $Y2=0
r86 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r87 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.45
+ $Y2=0
r88 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.99
+ $Y2=0
r89 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r90 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r91 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.575
+ $Y2=0
r93 35 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=2.07
+ $Y2=0
r94 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.45
+ $Y2=0
r95 34 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.07
+ $Y2=0
r96 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r97 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r98 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r99 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.735
+ $Y2=0
r100 30 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.15
+ $Y2=0
r101 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.575
+ $Y2=0
r102 29 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.15
+ $Y2=0
r103 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.735
+ $Y2=0
r104 24 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.23
+ $Y2=0
r105 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r106 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r107 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0
r108 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.36
r109 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0
r110 14 16 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0.385
r111 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r112 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.38
r113 3 20 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.45 $Y2=0.36
r114 2 16 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.575 $Y2=0.385
r115 1 12 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.735 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__decap_3.pex.spice
* Created: Thu Aug 27 14:13:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DECAP_3%VGND 1 7 9 12 15 25 28
r14 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r15 25 27 0.442563 $w=8.27e-07 $l=3e-08 $layer=LI1_cond $X=1.12 $Y=0.375
+ $X2=1.15 $Y2=0.375
r16 23 25 11.4329 $w=8.27e-07 $l=7.75e-07 $layer=LI1_cond $X=0.345 $Y=0.375
+ $X2=1.12 $Y2=0.375
r17 22 23 1.25393 $w=8.27e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.375
+ $X2=0.345 $Y2=0.375
r18 19 22 0.442563 $w=8.27e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.375
+ $X2=0.26 $Y2=0.375
r19 15 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r20 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r21 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.29 $X2=0.42 $Y2=1.29
r22 10 23 3.45185 $w=5.2e-07 $l=4.6e-07 $layer=LI1_cond $X=0.345 $Y=0.835
+ $X2=0.345 $Y2=0.375
r23 10 12 10.4657 $w=5.18e-07 $l=4.55e-07 $layer=LI1_cond $X=0.345 $Y=0.835
+ $X2=0.345 $Y2=1.29
r24 7 13 41.3046 $w=5.9e-07 $l=5.89746e-07 $layer=POLY_cond $X=0.69 $Y=1.76
+ $X2=0.42 $Y2=1.29
r25 7 9 23.6915 $w=5.9e-07 $l=2.9e-07 $layer=POLY_cond $X=0.69 $Y=1.76 $X2=0.69
+ $Y2=2.05
r26 1 25 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.485
r27 1 22 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=0.26 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__DECAP_3%VPWR 1 9 12 15 21 24
r14 21 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r15 18 21 8.46672 $w=1.232e-06 $l=8.55e-07 $layer=LI1_cond $X=0.69 $Y=1.865
+ $X2=0.69 $Y2=2.72
r16 12 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r17 12 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r18 10 15 54.7084 $w=5.11e-07 $l=6.72607e-07 $layer=POLY_cond $X=0.96 $Y=1.09
+ $X2=0.76 $Y2=0.51
r19 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.09 $X2=0.96 $Y2=1.09
r20 7 18 7.3378 $w=1.232e-06 $l=4.78983e-07 $layer=LI1_cond $X=1.035 $Y=1.545
+ $X2=0.69 $Y2=1.865
r21 7 9 10.4657 $w=5.18e-07 $l=4.55e-07 $layer=LI1_cond $X=1.035 $Y=1.545
+ $X2=1.035 $Y2=1.09
r22 1 18 300 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.615 $X2=1.12 $Y2=1.865
r23 1 18 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.615 $X2=0.26 $Y2=1.865
.ends


* File: sky130_fd_sc_hd__lpflow_decapkapwr_4.pex.spice
* Created: Thu Aug 27 14:24:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%VGND 1 7 10 13 24 27
r11 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r12 24 26 0.338889 $w=1.08e-06 $l=3e-08 $layer=LI1_cond $X=1.58 $Y=0.645
+ $X2=1.61 $Y2=0.645
r13 22 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r14 21 24 10.0537 $w=1.08e-06 $l=8.9e-07 $layer=LI1_cond $X=0.69 $Y=0.645
+ $X2=1.58 $Y2=0.645
r15 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r16 15 18 0.338889 $w=1.08e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.645
+ $X2=0.26 $Y2=0.645
r17 11 21 4.74444 $w=1.08e-06 $l=4.2e-07 $layer=LI1_cond $X=0.27 $Y=0.645
+ $X2=0.69 $Y2=0.645
r18 11 18 0.112963 $w=1.08e-06 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=0.645
+ $X2=0.26 $Y2=0.645
r19 10 13 41.1323 $w=9.62e-07 $l=7.6e-07 $layer=POLY_cond $X=0.775 $Y=1.29
+ $X2=0.775 $Y2=2.05
r20 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.29 $X2=0.27 $Y2=1.29
r21 7 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r22 7 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r23 1 24 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.51
r24 1 18 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%KAPWR 1 9 13 24 27 28 30
c14 27 0 7.9696e-20 $X=1.61 $Y=2.21
r15 28 30 0.0085136 $w=2.6e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.21
+ $X2=0.23 $Y2=2.21
r16 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.21
+ $X2=1.61 $Y2=2.21
r17 24 26 0.317433 $w=1.153e-06 $l=3e-08 $layer=LI1_cond $X=1.58 $Y=1.745
+ $X2=1.61 $Y2=1.745
r18 18 21 0.317433 $w=1.153e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=1.745
+ $X2=0.26 $Y2=1.745
r19 18 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r20 16 24 0.105811 $w=1.153e-06 $l=1e-08 $layer=LI1_cond $X=1.57 $Y=1.745
+ $X2=1.58 $Y2=1.745
r21 16 21 13.8612 $w=1.153e-06 $l=1.31e-06 $layer=LI1_cond $X=1.57 $Y=1.745
+ $X2=0.26 $Y2=1.745
r22 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.11 $X2=1.57 $Y2=1.11
r23 13 15 38.6501 $w=8.18e-07 $l=8.33966e-07 $layer=POLY_cond $X=0.92 $Y=0.69
+ $X2=1.57 $Y2=1.11
r24 9 28 0.0120192 $w=2.6e-07 $l=2.5e-08 $layer=MET1_cond $X=0.19 $Y=2.21
+ $X2=0.215 $Y2=2.21
r25 9 27 0.756575 $w=2.6e-07 $l=1.333e-06 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=1.61 $Y2=2.21
r26 9 30 0.0266759 $w=2.6e-07 $l=4.7e-08 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=0.23 $Y2=2.21
r27 1 24 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.615 $X2=1.58 $Y2=1.83
r28 1 21 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%VPWR 1 8 9
c10 8 0 7.9696e-20 $X=1.61 $Y=2.72
r11 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72 $X2=1.61
+ $Y2=2.72
r12 4 8 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=1.61
+ $Y2=2.72
r13 1 9 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r14 1 4 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends


* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1.pxi.spice
* Created: Tue Sep  1 19:13:10 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VGND N_VGND_M1010_s
+ N_VGND_M1004_s N_VGND_M1005_s N_VGND_M1007_s N_VGND_M1006_s N_VGND_M1014_s
+ N_VGND_M1012_s N_VGND_M1010_b N_VGND_c_30_p N_VGND_c_9_p N_VGND_c_31_p
+ N_VGND_c_13_p N_VGND_c_52_p N_VGND_c_25_p N_VGND_c_83_p N_VGND_c_32_p
+ N_VGND_c_10_p N_VGND_c_39_p N_VGND_c_48_p N_VGND_c_124_p N_VGND_c_103_p VGND
+ VGND N_VGND_c_21_p N_VGND_c_33_p N_VGND_c_11_p
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPB N_VPB_X16_noxref_D1
+ N_VPB_M1015_b N_VPB_c_214_p N_VPB_c_140_n VPB N_VPB_c_141_n N_VPB_c_142_n VPB
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPB
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPWRIN N_VPWRIN_M1009_s
+ N_VPWRIN_M1009_b N_VPWRIN_c_245_p N_VPWRIN_c_224_n N_VPWRIN_c_237_p
+ N_VPWRIN_c_219_n N_VPWRIN_c_220_n N_VPWRIN_c_235_p N_VPWRIN_c_221_n VPWRIN
+ N_VPWRIN_c_222_n PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPWRIN
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_505_297#
+ N_A_505_297#_M1010_d N_A_505_297#_M1009_d N_A_505_297#_c_274_n
+ N_A_505_297#_M1004_g N_A_505_297#_c_278_n N_A_505_297#_M1007_g
+ N_A_505_297#_c_282_n N_A_505_297#_c_284_n N_A_505_297#_c_285_n
+ N_A_505_297#_M1013_g N_A_505_297#_c_289_n N_A_505_297#_c_290_n
+ N_A_505_297#_M1014_g N_A_505_297#_c_294_n N_A_505_297#_c_295_n
+ N_A_505_297#_c_300_n N_A_505_297#_c_311_n N_A_505_297#_c_301_n
+ N_A_505_297#_c_302_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_505_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_714_58#
+ N_A_714_58#_M1005_d N_A_714_58#_M1011_d N_A_714_58#_M1001_s
+ N_A_714_58#_c_381_n N_A_714_58#_c_358_n N_A_714_58#_M1015_g
+ N_A_714_58#_c_359_n N_A_714_58#_c_362_n N_A_714_58#_c_363_n
+ N_A_714_58#_c_364_n N_A_714_58#_c_365_n N_A_714_58#_c_366_n
+ N_A_714_58#_c_367_n N_A_714_58#_c_371_n N_A_714_58#_c_388_n
+ N_A_714_58#_c_376_n N_A_714_58#_c_377_n N_A_714_58#_c_380_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_714_58#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A N_A_M1009_g N_A_c_463_n
+ N_A_M1010_g N_A_c_468_n N_A_M1005_g N_A_c_474_n N_A_c_475_n N_A_M1006_g
+ N_A_c_482_n N_A_M1011_g N_A_c_488_n N_A_M1012_g N_A_c_494_n N_A_c_495_n
+ N_A_c_496_n A N_A_c_497_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_620_911#
+ N_A_620_911#_M1004_d N_A_620_911#_M1013_d N_A_620_911#_M1015_s
+ N_A_620_911#_c_557_n N_A_620_911#_c_535_n N_A_620_911#_c_536_n
+ N_A_620_911#_M1001_g N_A_620_911#_c_563_n N_A_620_911#_c_564_n
+ N_A_620_911#_M1008_g N_A_620_911#_M1002_g N_A_620_911#_c_568_n
+ N_A_620_911#_c_569_n N_A_620_911#_c_570_n N_A_620_911#_c_541_n
+ N_A_620_911#_c_545_n N_A_620_911#_c_572_n N_A_620_911#_c_547_n
+ N_A_620_911#_c_573_n N_A_620_911#_c_551_n N_A_620_911#_c_552_n
+ N_A_620_911#_c_553_n N_A_620_911#_c_554_n N_A_620_911#_c_579_n
+ N_A_620_911#_c_555_n N_A_620_911#_c_556_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_620_911#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_1028_32#
+ N_A_1028_32#_M1008_d N_A_1028_32#_M1002_d N_A_1028_32#_c_660_n
+ N_A_1028_32#_M1003_g N_A_1028_32#_M1000_g N_A_1028_32#_c_673_n
+ N_A_1028_32#_c_674_n N_A_1028_32#_c_675_n N_A_1028_32#_c_676_n
+ N_A_1028_32#_c_664_n N_A_1028_32#_c_680_n N_A_1028_32#_c_681_n
+ N_A_1028_32#_c_665_n N_A_1028_32#_c_666_n N_A_1028_32#_c_670_n
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_1028_32#
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPWR N_VPWR_M1015_d
+ N_VPWR_M1001_d N_VPWR_c_730_n N_VPWR_c_731_n N_VPWR_c_733_n VPWR
+ N_VPWR_c_727_n N_VPWR_c_736_n N_VPWR_c_728_n VPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%X N_X_M1003_d N_X_M1000_d
+ N_X_c_808_n X X X PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%X
cc_1 N_VGND_M1010_b N_VPB_c_140_n 0.0790644f $X=-0.19 $Y=-0.24 $X2=5.87 $Y2=3.57
cc_2 N_VGND_M1010_b N_VPB_c_141_n 0.0100791f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=3.29
cc_3 N_VGND_M1010_b N_VPB_c_142_n 0.00243231f $X=-0.19 $Y=-0.24 $X2=6.01
+ $Y2=3.29
cc_4 N_VGND_M1010_b N_VPWRIN_c_219_n 0.00447854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 N_VGND_M1010_b N_VPWRIN_c_220_n 0.0244366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 N_VGND_M1010_b N_VPWRIN_c_221_n 0.0306316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 N_VGND_M1010_b N_VPWRIN_c_222_n 0.0344347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 N_VGND_M1010_b N_A_505_297#_c_274_n 0.0179052f $X=-0.19 $Y=-0.24 $X2=-0.19
+ $Y2=1.305
cc_9 N_VGND_c_9_p N_A_505_297#_c_274_n 0.00414737f $X=2.81 $Y=4.7 $X2=-0.19
+ $Y2=1.305
cc_10 N_VGND_c_10_p N_A_505_297#_c_274_n 0.0054895f $X=3.575 $Y=5.44 $X2=-0.19
+ $Y2=1.305
cc_11 N_VGND_c_11_p N_A_505_297#_c_274_n 0.0110264f $X=6.21 $Y=5.44 $X2=-0.19
+ $Y2=1.305
cc_12 N_VGND_M1010_b N_A_505_297#_c_278_n 0.0140848f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_13 N_VGND_c_13_p N_A_505_297#_c_278_n 0.00179869f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_14 N_VGND_c_10_p N_A_505_297#_c_278_n 0.0054895f $X=3.575 $Y=5.44 $X2=0 $Y2=0
cc_15 N_VGND_c_11_p N_A_505_297#_c_278_n 0.00972667f $X=6.21 $Y=5.44 $X2=0 $Y2=0
cc_16 N_VGND_M1010_b N_A_505_297#_c_282_n 0.0130779f $X=-0.19 $Y=-0.24 $X2=0.225
+ $Y2=3.57
cc_17 N_VGND_c_13_p N_A_505_297#_c_282_n 0.00240634f $X=3.67 $Y=4.735 $X2=0.225
+ $Y2=3.57
cc_18 N_VGND_M1010_b N_A_505_297#_c_284_n 0.0294363f $X=-0.19 $Y=-0.24 $X2=0.225
+ $Y2=3.57
cc_19 N_VGND_M1010_b N_A_505_297#_c_285_n 0.0140848f $X=-0.19 $Y=-0.24 $X2=5.87
+ $Y2=3.57
cc_20 N_VGND_c_13_p N_A_505_297#_c_285_n 0.00304527f $X=3.67 $Y=4.735 $X2=5.87
+ $Y2=3.57
cc_21 N_VGND_c_21_p N_A_505_297#_c_285_n 0.0054895f $X=4.445 $Y=5.44 $X2=5.87
+ $Y2=3.57
cc_22 N_VGND_c_11_p N_A_505_297#_c_285_n 0.00972667f $X=6.21 $Y=5.44 $X2=5.87
+ $Y2=3.57
cc_23 N_VGND_M1010_b N_A_505_297#_c_289_n 0.0195784f $X=-0.19 $Y=-0.24 $X2=6.015
+ $Y2=3.57
cc_24 N_VGND_M1010_b N_A_505_297#_c_290_n 0.0162763f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_25 N_VGND_c_25_p N_A_505_297#_c_290_n 0.00390324f $X=4.87 $Y=4.735 $X2=0
+ $Y2=0
cc_26 N_VGND_c_21_p N_A_505_297#_c_290_n 0.0054895f $X=4.445 $Y=5.44 $X2=0 $Y2=0
cc_27 N_VGND_c_11_p N_A_505_297#_c_290_n 0.0103929f $X=6.21 $Y=5.44 $X2=0 $Y2=0
cc_28 N_VGND_M1010_b N_A_505_297#_c_294_n 0.00569361f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_29 N_VGND_M1010_b N_A_505_297#_c_295_n 0.00997858f $X=-0.19 $Y=-0.24
+ $X2=0.557 $Y2=3.57
cc_30 N_VGND_c_30_p N_A_505_297#_c_295_n 0.0068636f $X=2.245 $Y=0.62 $X2=0.557
+ $Y2=3.57
cc_31 N_VGND_c_31_p N_A_505_297#_c_295_n 0.0271827f $X=3.28 $Y=0.475 $X2=0.557
+ $Y2=3.57
cc_32 N_VGND_c_32_p N_A_505_297#_c_295_n 0.00966373f $X=3.115 $Y=0 $X2=0.557
+ $Y2=3.57
cc_33 N_VGND_c_33_p N_A_505_297#_c_295_n 0.00857725f $X=6.21 $Y=0 $X2=0.557
+ $Y2=3.57
cc_34 N_VGND_M1010_b N_A_505_297#_c_300_n 0.016089f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_35 N_VGND_M1010_b N_A_505_297#_c_301_n 0.034685f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_36 N_VGND_M1010_b N_A_505_297#_c_302_n 0.0845171f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_37 N_VGND_M1010_b N_A_714_58#_c_358_n 0.0129761f $X=-0.19 $Y=-0.24 $X2=0.37
+ $Y2=3.57
cc_38 N_VGND_M1010_b N_A_714_58#_c_359_n 0.00127602f $X=-0.19 $Y=-0.24 $X2=0.49
+ $Y2=3.5
cc_39 N_VGND_c_39_p N_A_714_58#_c_359_n 0.00988313f $X=3.975 $Y=0 $X2=0.49
+ $Y2=3.5
cc_40 N_VGND_c_33_p N_A_714_58#_c_359_n 0.00702789f $X=6.21 $Y=0 $X2=0.49
+ $Y2=3.5
cc_41 N_VGND_M1010_b N_A_714_58#_c_362_n 0.0175549f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.29
cc_42 N_VGND_M1010_b N_A_714_58#_c_363_n 0.00209323f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_43 N_VGND_M1010_b N_A_714_58#_c_364_n 0.00298088f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.57
cc_44 N_VGND_M1010_b N_A_714_58#_c_365_n 0.0397033f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_45 N_VGND_M1010_b N_A_714_58#_c_366_n 0.0516547f $X=-0.19 $Y=-0.24 $X2=6.01
+ $Y2=3.57
cc_46 N_VGND_M1006_s N_A_714_58#_c_367_n 3.36085e-19 $X=4 $Y=0.29 $X2=0 $Y2=0
cc_47 N_VGND_M1010_b N_A_714_58#_c_367_n 0.00479086f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_48 N_VGND_c_48_p N_A_714_58#_c_367_n 0.00202943f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_49 N_VGND_c_33_p N_A_714_58#_c_367_n 0.00393502f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_50 N_VGND_M1006_s N_A_714_58#_c_371_n 0.00139685f $X=4 $Y=0.29 $X2=0.557
+ $Y2=3.57
cc_51 N_VGND_M1010_b N_A_714_58#_c_371_n 0.00744058f $X=-0.19 $Y=-0.24 $X2=0.557
+ $Y2=3.57
cc_52 N_VGND_c_52_p N_A_714_58#_c_371_n 0.0168391f $X=4.14 $Y=0.475 $X2=0.557
+ $Y2=3.57
cc_53 N_VGND_c_39_p N_A_714_58#_c_371_n 0.00204475f $X=3.975 $Y=0 $X2=0.557
+ $Y2=3.57
cc_54 N_VGND_c_33_p N_A_714_58#_c_371_n 0.00525801f $X=6.21 $Y=0 $X2=0.557
+ $Y2=3.57
cc_55 N_VGND_M1010_b N_A_714_58#_c_376_n 0.00351628f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_56 N_VGND_M1010_b N_A_714_58#_c_377_n 0.00128614f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_57 N_VGND_c_48_p N_A_714_58#_c_377_n 0.0101829f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_58 N_VGND_c_33_p N_A_714_58#_c_377_n 0.00711893f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_59 N_VGND_M1010_b N_A_714_58#_c_380_n 0.00576889f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_60 N_VGND_M1010_b N_A_M1009_g 0.00675179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 N_VGND_M1010_b N_A_c_463_n 0.0408343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 N_VGND_c_30_p N_A_c_463_n 0.0135915f $X=2.245 $Y=0.62 $X2=0 $Y2=0
cc_63 N_VGND_c_31_p N_A_c_463_n 0.00625119f $X=3.28 $Y=0.475 $X2=0 $Y2=0
cc_64 N_VGND_c_32_p N_A_c_463_n 0.00585385f $X=3.115 $Y=0 $X2=0 $Y2=0
cc_65 N_VGND_c_33_p N_A_c_463_n 0.0134051f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_66 N_VGND_M1010_b N_A_c_468_n 0.0352506f $X=-0.19 $Y=-0.24 $X2=4.25 $Y2=1.305
cc_67 N_VGND_M1010_b N_A_M1005_g 0.0208571f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=3.57
cc_68 N_VGND_c_31_p N_A_M1005_g 0.0122275f $X=3.28 $Y=0.475 $X2=0.225 $Y2=3.57
cc_69 N_VGND_c_52_p N_A_M1005_g 4.84532e-19 $X=4.14 $Y=0.475 $X2=0.225 $Y2=3.57
cc_70 N_VGND_c_39_p N_A_M1005_g 0.00441152f $X=3.975 $Y=0 $X2=0.225 $Y2=3.57
cc_71 N_VGND_c_33_p N_A_M1005_g 0.00802014f $X=6.21 $Y=0 $X2=0.225 $Y2=3.57
cc_72 N_VGND_M1010_b N_A_c_474_n 0.0168496f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=3.57
cc_73 N_VGND_M1010_b N_A_c_475_n 0.0656946f $X=-0.19 $Y=-0.24 $X2=5.87 $Y2=3.57
cc_74 N_VGND_c_31_p N_A_c_475_n 0.00306309f $X=3.28 $Y=0.475 $X2=5.87 $Y2=3.57
cc_75 N_VGND_M1010_b N_A_M1006_g 0.0168071f $X=-0.19 $Y=-0.24 $X2=6.015 $Y2=3.57
cc_76 N_VGND_c_31_p N_A_M1006_g 5.35342e-19 $X=3.28 $Y=0.475 $X2=6.015 $Y2=3.57
cc_77 N_VGND_c_52_p N_A_M1006_g 0.00698688f $X=4.14 $Y=0.475 $X2=6.015 $Y2=3.57
cc_78 N_VGND_c_39_p N_A_M1006_g 0.00327003f $X=3.975 $Y=0 $X2=6.015 $Y2=3.57
cc_79 N_VGND_c_33_p N_A_M1006_g 0.00407147f $X=6.21 $Y=0 $X2=6.015 $Y2=3.57
cc_80 N_VGND_M1010_b N_A_c_482_n 0.0149976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 N_VGND_M1010_b N_A_M1011_g 0.0168094f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=3.57
cc_82 N_VGND_c_52_p N_A_M1011_g 0.00698688f $X=4.14 $Y=0.475 $X2=0.23 $Y2=3.57
cc_83 N_VGND_c_83_p N_A_M1011_g 5.32908e-19 $X=5 $Y=0.475 $X2=0.23 $Y2=3.57
cc_84 N_VGND_c_48_p N_A_M1011_g 0.00327003f $X=4.835 $Y=0 $X2=0.23 $Y2=3.57
cc_85 N_VGND_c_33_p N_A_M1011_g 0.00407147f $X=6.21 $Y=0 $X2=0.23 $Y2=3.57
cc_86 N_VGND_M1010_b N_A_c_488_n 0.0253117f $X=-0.19 $Y=-0.24 $X2=6.01 $Y2=3.29
cc_87 N_VGND_M1010_b N_A_M1012_g 0.0174292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 N_VGND_c_52_p N_A_M1012_g 4.84532e-19 $X=4.14 $Y=0.475 $X2=0 $Y2=0
cc_89 N_VGND_c_83_p N_A_M1012_g 0.0104329f $X=5 $Y=0.475 $X2=0 $Y2=0
cc_90 N_VGND_c_48_p N_A_M1012_g 0.00441152f $X=4.835 $Y=0 $X2=0 $Y2=0
cc_91 N_VGND_c_33_p N_A_M1012_g 0.00802014f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_92 N_VGND_M1010_b N_A_c_494_n 0.017446f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=3.57
cc_93 N_VGND_M1010_b N_A_c_495_n 0.00933068f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=3.57
cc_94 N_VGND_M1010_b N_A_c_496_n 0.0106787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 N_VGND_M1010_b N_A_c_497_n 0.0169952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 N_VGND_c_31_p N_A_c_497_n 0.014754f $X=3.28 $Y=0.475 $X2=0 $Y2=0
cc_97 N_VGND_c_11_p N_A_620_911#_M1004_d 0.00223231f $X=6.21 $Y=5.44 $X2=0.145
+ $Y2=3.04
cc_98 N_VGND_c_11_p N_A_620_911#_M1013_d 0.00223231f $X=6.21 $Y=5.44 $X2=5.925
+ $Y2=3.04
cc_99 N_VGND_M1010_b N_A_620_911#_c_535_n 0.0127228f $X=-0.19 $Y=-0.24 $X2=0.37
+ $Y2=3.57
cc_100 N_VGND_c_25_p N_A_620_911#_c_536_n 0.0183082f $X=4.87 $Y=4.735 $X2=0.225
+ $Y2=3.57
cc_101 N_VGND_M1010_b N_A_620_911#_M1008_g 0.0484682f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.57
cc_102 N_VGND_c_25_p N_A_620_911#_M1008_g 0.00390249f $X=4.87 $Y=4.735 $X2=0.23
+ $Y2=3.57
cc_103 N_VGND_c_103_p N_A_620_911#_M1008_g 0.00548296f $X=5.865 $Y=5.44 $X2=0.23
+ $Y2=3.57
cc_104 N_VGND_c_11_p N_A_620_911#_M1008_g 0.0116568f $X=6.21 $Y=5.44 $X2=0.23
+ $Y2=3.57
cc_105 N_VGND_c_9_p N_A_620_911#_c_541_n 0.0267051f $X=2.81 $Y=4.7 $X2=0 $Y2=0
cc_106 N_VGND_c_13_p N_A_620_911#_c_541_n 0.0266323f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_107 N_VGND_c_10_p N_A_620_911#_c_541_n 0.0189253f $X=3.575 $Y=5.44 $X2=0
+ $Y2=0
cc_108 N_VGND_c_11_p N_A_620_911#_c_541_n 0.0122674f $X=6.21 $Y=5.44 $X2=0 $Y2=0
cc_109 N_VGND_M1010_b N_A_620_911#_c_545_n 0.0128475f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_110 N_VGND_c_13_p N_A_620_911#_c_545_n 0.0146667f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_111 N_VGND_c_13_p N_A_620_911#_c_547_n 0.0266323f $X=3.67 $Y=4.735 $X2=0
+ $Y2=0
cc_112 N_VGND_c_25_p N_A_620_911#_c_547_n 0.025678f $X=4.87 $Y=4.735 $X2=0 $Y2=0
cc_113 N_VGND_c_21_p N_A_620_911#_c_547_n 0.0189253f $X=4.445 $Y=5.44 $X2=0
+ $Y2=0
cc_114 N_VGND_c_11_p N_A_620_911#_c_547_n 0.0122674f $X=6.21 $Y=5.44 $X2=0 $Y2=0
cc_115 N_VGND_M1010_b N_A_620_911#_c_551_n 0.0561622f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_116 N_VGND_M1010_b N_A_620_911#_c_552_n 0.0016479f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_117 N_VGND_M1010_b N_A_620_911#_c_553_n 7.55444e-19 $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_118 N_VGND_M1010_b N_A_620_911#_c_554_n 9.83343e-19 $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_119 N_VGND_M1010_b N_A_620_911#_c_555_n 0.00835191f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_120 N_VGND_M1010_b N_A_620_911#_c_556_n 0.0133087f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_121 N_VGND_c_11_p N_A_1028_32#_M1008_d 0.00214546f $X=6.21 $Y=5.44 $X2=0.145
+ $Y2=3.04
cc_122 N_VGND_M1010_b N_A_1028_32#_c_660_n 0.0202016f $X=-0.19 $Y=-0.24
+ $X2=-0.19 $Y2=1.305
cc_123 N_VGND_c_83_p N_A_1028_32#_c_660_n 0.0134873f $X=5 $Y=0.475 $X2=-0.19
+ $Y2=1.305
cc_124 N_VGND_c_124_p N_A_1028_32#_c_660_n 0.00441152f $X=5.865 $Y=0 $X2=-0.19
+ $Y2=1.305
cc_125 N_VGND_c_33_p N_A_1028_32#_c_660_n 0.00881995f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=1.305
cc_126 N_VGND_M1010_b N_A_1028_32#_c_664_n 0.0702068f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.29
cc_127 N_VGND_M1010_b N_A_1028_32#_c_665_n 0.0216787f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_128 N_VGND_M1010_b N_A_1028_32#_c_666_n 0.067692f $X=-0.19 $Y=-0.24 $X2=0.56
+ $Y2=3.57
cc_129 N_VGND_c_25_p N_A_1028_32#_c_666_n 0.0259447f $X=4.87 $Y=4.735 $X2=0.56
+ $Y2=3.57
cc_130 N_VGND_c_103_p N_A_1028_32#_c_666_n 0.0239189f $X=5.865 $Y=5.44 $X2=0.56
+ $Y2=3.57
cc_131 N_VGND_c_11_p N_A_1028_32#_c_666_n 0.0195213f $X=6.21 $Y=5.44 $X2=0.56
+ $Y2=3.57
cc_132 N_VGND_M1010_b N_A_1028_32#_c_670_n 0.0379295f $X=-0.19 $Y=-0.24 $X2=0
+ $Y2=0
cc_133 N_VGND_M1010_b N_VPWR_c_727_n 0.0363208f $X=-0.19 $Y=-0.24 $X2=0.23
+ $Y2=3.57
cc_134 N_VGND_M1010_b N_VPWR_c_728_n 0.0368329f $X=-0.19 $Y=-0.24 $X2=0.56
+ $Y2=3.57
cc_135 N_VGND_M1010_b N_X_c_808_n 0.0439478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 N_VGND_c_124_p N_X_c_808_n 0.0168697f $X=5.865 $Y=0 $X2=0 $Y2=0
cc_137 N_VGND_c_33_p N_X_c_808_n 0.0112798f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_138 N_VGND_M1010_b X 0.00616885f $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=3.57
cc_139 N_VGND_M1010_b X 0.00156813f $X=-0.19 $Y=-0.24 $X2=6.015 $Y2=3.57
cc_140 N_VPB_c_140_n N_VPWRIN_M1009_b 0.0152996f $X=5.87 $Y=3.57 $X2=4.86
+ $Y2=0.29
cc_141 N_VPB_c_140_n N_VPWRIN_c_224_n 0.0727088f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_142 N_VPB_M1015_b N_VPWRIN_c_220_n 0.0283959f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_143 N_VPB_X16_noxref_D1 N_VPWRIN_c_221_n 0.0309709f $X=-0.19 $Y=1.305 $X2=0
+ $Y2=0
cc_144 N_VPB_c_140_n N_A_505_297#_c_301_n 0.0247683f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_145 N_VPB_c_140_n N_A_505_297#_c_302_n 6.63876e-19 $X=5.87 $Y=3.57 $X2=0.23
+ $Y2=0.085
cc_146 N_VPB_M1015_b N_A_714_58#_c_381_n 0.0255327f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_147 N_VPB_M1015_b N_A_714_58#_c_358_n 5.34541e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_148 N_VPB_M1015_b N_A_714_58#_M1015_g 0.0196228f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_149 N_VPB_M1015_b N_A_714_58#_c_363_n 0.0045246f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_150 N_VPB_c_140_n N_A_714_58#_c_363_n 0.0451176f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_151 N_VPB_c_140_n N_A_714_58#_c_364_n 0.010882f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_152 N_VPB_M1015_b N_A_714_58#_c_366_n 0.0149067f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_153 N_VPB_M1015_b N_A_714_58#_c_388_n 0.00449536f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_154 N_VPB_M1015_b N_A_620_911#_c_557_n 0.0169344f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_155 N_VPB_M1015_b N_A_620_911#_c_535_n 5.21411e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_156 N_VPB_M1015_b N_A_620_911#_c_536_n 0.0246766f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_157 N_VPB_c_140_n N_A_620_911#_c_536_n 5.78421e-19 $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_158 N_VPB_M1015_b N_A_620_911#_M1001_g 0.00259316f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_159 N_VPB_c_140_n N_A_620_911#_M1001_g 0.00720206f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_160 N_VPB_M1015_b N_A_620_911#_c_563_n 0.0243277f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_161 N_VPB_M1015_b N_A_620_911#_c_564_n 0.0094712f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_162 N_VPB_M1015_b N_A_620_911#_M1008_g 0.00114838f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_163 N_VPB_M1015_b N_A_620_911#_M1002_g 0.00645643f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_164 N_VPB_c_140_n N_A_620_911#_M1002_g 0.00821798f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_165 N_VPB_M1015_b N_A_620_911#_c_568_n 0.00400906f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_166 N_VPB_M1015_b N_A_620_911#_c_569_n 0.00698872f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_167 N_VPB_M1015_b N_A_620_911#_c_570_n 0.0141637f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_168 N_VPB_c_140_n N_A_620_911#_c_545_n 0.0118014f $X=5.87 $Y=3.57 $X2=0.23
+ $Y2=0.085
cc_169 N_VPB_c_140_n N_A_620_911#_c_572_n 0.00154646f $X=5.87 $Y=3.57 $X2=0.23
+ $Y2=0.64
cc_170 N_VPB_c_140_n N_A_620_911#_c_573_n 7.52174e-19 $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_171 N_VPB_M1015_b N_A_620_911#_c_551_n 0.0188917f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_172 N_VPB_c_140_n N_A_620_911#_c_551_n 0.00519139f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_173 N_VPB_c_140_n N_A_620_911#_c_552_n 0.00368761f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_174 N_VPB_M1015_b N_A_620_911#_c_553_n 0.00337762f $X=4.25 $Y=1.305 $X2=2.81
+ $Y2=4.7
cc_175 N_VPB_c_140_n N_A_620_911#_c_553_n 8.12088e-19 $X=5.87 $Y=3.57 $X2=2.81
+ $Y2=4.7
cc_176 N_VPB_M1015_b N_A_620_911#_c_579_n 0.00324872f $X=4.25 $Y=1.305 $X2=3.28
+ $Y2=0.475
cc_177 N_VPB_c_140_n N_A_620_911#_c_555_n 0.00167232f $X=5.87 $Y=3.57 $X2=3.67
+ $Y2=5.355
cc_178 N_VPB_M1015_b N_A_620_911#_c_556_n 6.57859e-19 $X=4.25 $Y=1.305 $X2=3.67
+ $Y2=4.735
cc_179 N_VPB_c_140_n N_A_1028_32#_M1002_d 0.00329366f $X=5.87 $Y=3.57 $X2=2.685
+ $Y2=4.555
cc_180 N_VPB_M1015_b N_A_1028_32#_M1000_g 0.00952509f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_181 N_VPB_M1015_b N_A_1028_32#_c_673_n 0.0246441f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_182 N_VPB_M1015_b N_A_1028_32#_c_674_n 0.00607427f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_183 N_VPB_M1015_b N_A_1028_32#_c_675_n 0.0805674f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_184 N_VPB_M1015_b N_A_1028_32#_c_676_n 0.0884656f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_185 N_VPB_c_140_n N_A_1028_32#_c_676_n 0.00776237f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_186 N_VPB_c_142_n N_A_1028_32#_c_676_n 0.0261557f $X=6.01 $Y=3.29 $X2=0 $Y2=0
cc_187 N_VPB_M1015_b N_A_1028_32#_c_664_n 0.037361f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_188 N_VPB_M1015_b N_A_1028_32#_c_680_n 0.00738594f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_189 N_VPB_M1015_b N_A_1028_32#_c_681_n 0.00744458f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_190 N_VPB_c_140_n N_A_1028_32#_c_681_n 0.0227f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_191 N_VPB_c_142_n N_A_1028_32#_c_681_n 0.0419493f $X=6.01 $Y=3.29 $X2=0 $Y2=0
cc_192 N_VPB_M1015_b N_A_1028_32#_c_665_n 6.19031e-19 $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_193 N_VPB_c_140_n N_A_1028_32#_c_665_n 0.00369231f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_194 N_VPB_c_142_n N_A_1028_32#_c_665_n 0.0174681f $X=6.01 $Y=3.29 $X2=0 $Y2=0
cc_195 N_VPB_M1015_b N_A_1028_32#_c_666_n 0.00293548f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_196 N_VPB_c_140_n N_A_1028_32#_c_666_n 0.00771994f $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_197 N_VPB_M1015_b N_A_1028_32#_c_670_n 0.0181697f $X=4.25 $Y=1.305 $X2=0
+ $Y2=0
cc_198 N_VPB_c_140_n N_A_1028_32#_c_670_n 3.47599e-19 $X=5.87 $Y=3.57 $X2=0
+ $Y2=0
cc_199 N_VPB_c_142_n N_A_1028_32#_c_670_n 0.005123f $X=6.01 $Y=3.29 $X2=0 $Y2=0
cc_200 N_VPB_c_140_n N_VPWR_M1001_d 0.00370825f $X=5.87 $Y=3.57 $X2=2.685
+ $Y2=4.555
cc_201 N_VPB_M1015_b N_VPWR_c_730_n 0.00616116f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_202 N_VPB_M1015_b N_VPWR_c_731_n 0.00447924f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_203 N_VPB_c_140_n N_VPWR_c_731_n 0.0205244f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_204 N_VPB_M1015_b N_VPWR_c_733_n 9.70405e-19 $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_205 N_VPB_X16_noxref_D1 N_VPWR_c_727_n 0.0202024f $X=-0.19 $Y=1.305 $X2=0
+ $Y2=0
cc_206 N_VPB_c_141_n N_VPWR_c_727_n 0.0194225f $X=0.23 $Y=3.29 $X2=0 $Y2=0
cc_207 N_VPB_M1015_b N_VPWR_c_736_n 0.0235549f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_208 N_VPB_c_142_n N_VPWR_c_736_n 0.0194225f $X=6.01 $Y=3.29 $X2=0 $Y2=0
cc_209 N_VPB_X16_noxref_D1 N_VPWR_c_728_n 0.0368104f $X=-0.19 $Y=1.305 $X2=0
+ $Y2=0
cc_210 N_VPB_M1015_b N_VPWR_c_728_n 0.0550446f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_211 N_VPB_c_214_p N_VPWR_c_728_n 0.0152864f $X=0.37 $Y=3.57 $X2=0 $Y2=0
cc_212 N_VPB_c_140_n N_VPWR_c_728_n 0.279538f $X=5.87 $Y=3.57 $X2=0 $Y2=0
cc_213 N_VPB_c_141_n N_VPWR_c_728_n 0.00501853f $X=0.23 $Y=3.29 $X2=0 $Y2=0
cc_214 N_VPB_c_142_n N_VPWR_c_728_n 0.00501853f $X=6.01 $Y=3.29 $X2=0 $Y2=0
cc_215 N_VPB_M1015_b X 0.0157781f $X=4.25 $Y=1.305 $X2=0 $Y2=0
cc_216 N_VPWRIN_c_220_n N_A_505_297#_M1009_d 0.00144688f $X=2.225 $Y=2.2
+ $X2=2.685 $Y2=4.555
cc_217 N_VPWRIN_M1009_b N_A_505_297#_c_295_n 0.0037173f $X=1.92 $Y=1.305 $X2=0
+ $Y2=0
cc_218 N_VPWRIN_c_220_n N_A_505_297#_c_295_n 3.15819e-19 $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_219 N_VPWRIN_M1009_b N_A_505_297#_c_300_n 0.00974718f $X=1.92 $Y=1.305 $X2=0
+ $Y2=0
cc_220 N_VPWRIN_c_224_n N_A_505_297#_c_300_n 3.29394e-19 $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_221 N_VPWRIN_c_220_n N_A_505_297#_c_300_n 0.0372262f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_222 N_VPWRIN_c_224_n N_A_505_297#_c_311_n 0.00924483f $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_223 N_VPWRIN_c_220_n N_A_505_297#_c_311_n 0.0204768f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_224 N_VPWRIN_c_235_p N_A_505_297#_c_311_n 0.0100174f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_225 N_VPWRIN_c_224_n N_A_505_297#_c_301_n 0.0654251f $X=2.645 $Y=3.49 $X2=0
+ $Y2=0
cc_226 N_VPWRIN_c_237_p N_A_505_297#_c_301_n 0.00525651f $X=2.435 $Y=2.66 $X2=0
+ $Y2=0
cc_227 N_VPWRIN_c_224_n N_A_505_297#_c_302_n 0.00169032f $X=2.645 $Y=3.49
+ $X2=0.23 $Y2=0.085
cc_228 N_VPWRIN_c_220_n N_A_714_58#_c_381_n 5.4797e-19 $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_229 N_VPWRIN_c_220_n N_A_714_58#_M1015_g 0.00777495f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_230 N_VPWRIN_c_220_n N_A_714_58#_c_365_n 0.0182669f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_231 N_VPWRIN_c_220_n N_A_714_58#_c_366_n 0.0104851f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_232 N_VPWRIN_c_220_n N_A_714_58#_c_380_n 0.00926075f $X=2.225 $Y=2.2 $X2=0.23
+ $Y2=4.8
cc_233 N_VPWRIN_M1009_b N_A_M1009_g 0.0304234f $X=1.92 $Y=1.305 $X2=3.135
+ $Y2=0.29
cc_234 N_VPWRIN_c_245_p N_A_M1009_g 0.00523247f $X=2.225 $Y=1.79 $X2=3.135
+ $Y2=0.29
cc_235 N_VPWRIN_c_224_n N_A_M1009_g 0.0055008f $X=2.645 $Y=3.49 $X2=3.135
+ $Y2=0.29
cc_236 N_VPWRIN_c_237_p N_A_M1009_g 0.00938999f $X=2.435 $Y=2.66 $X2=3.135
+ $Y2=0.29
cc_237 N_VPWRIN_c_220_n N_A_M1009_g 0.00645994f $X=2.225 $Y=2.2 $X2=3.135
+ $Y2=0.29
cc_238 N_VPWRIN_c_235_p N_A_M1009_g 0.00218038f $X=2.225 $Y=2.2 $X2=3.135
+ $Y2=0.29
cc_239 N_VPWRIN_M1009_b N_A_c_475_n 0.00316885f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_240 N_VPWRIN_M1009_b N_A_c_497_n 0.00111856f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_241 N_VPWRIN_c_220_n N_A_c_497_n 0.00229296f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_242 N_VPWRIN_c_220_n N_A_620_911#_M1015_s 0.00479759f $X=2.225 $Y=2.2
+ $X2=3.135 $Y2=0.29
cc_243 N_VPWRIN_c_220_n N_A_620_911#_c_553_n 0.0011695f $X=2.225 $Y=2.2 $X2=2.81
+ $Y2=4.7
cc_244 N_VPWRIN_c_220_n N_A_620_911#_c_579_n 0.0174341f $X=2.225 $Y=2.2 $X2=3.28
+ $Y2=0.475
cc_245 N_VPWRIN_c_220_n N_A_1028_32#_M1000_g 0.00737951f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_246 N_VPWRIN_c_220_n N_A_1028_32#_c_675_n 0.0108557f $X=2.225 $Y=2.2 $X2=0
+ $Y2=0
cc_247 N_VPWRIN_c_220_n N_VPWR_M1015_d 0.00296071f $X=2.225 $Y=2.2 $X2=2.12
+ $Y2=0.41
cc_248 N_VPWRIN_c_220_n N_VPWR_c_730_n 0.0222006f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_249 N_VPWRIN_c_237_p N_VPWR_c_727_n 0.0123972f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_250 N_VPWRIN_c_219_n N_VPWR_c_727_n 5.76636e-19 $X=1.475 $Y=2.2 $X2=0 $Y2=0
cc_251 N_VPWRIN_c_221_n N_VPWR_c_727_n 0.00675753f $X=1.36 $Y=2.2 $X2=0 $Y2=0
cc_252 N_VPWRIN_c_222_n N_VPWR_c_727_n 0.01865f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_253 N_VPWRIN_c_220_n N_VPWR_c_736_n 0.00711378f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_254 N_VPWRIN_M1009_b N_VPWR_c_728_n 0.00623335f $X=1.92 $Y=1.305 $X2=0 $Y2=0
cc_255 N_VPWRIN_c_224_n N_VPWR_c_728_n 0.0659883f $X=2.645 $Y=3.49 $X2=0 $Y2=0
cc_256 N_VPWRIN_c_237_p N_VPWR_c_728_n 0.02138f $X=2.435 $Y=2.66 $X2=0 $Y2=0
cc_257 N_VPWRIN_c_219_n N_VPWR_c_728_n 0.0948062f $X=1.475 $Y=2.2 $X2=0 $Y2=0
cc_258 N_VPWRIN_c_220_n N_VPWR_c_728_n 0.32456f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_259 N_VPWRIN_c_221_n N_VPWR_c_728_n 0.116739f $X=1.36 $Y=2.2 $X2=0 $Y2=0
cc_260 N_VPWRIN_c_222_n N_VPWR_c_728_n 0.00970859f $X=2.06 $Y=2.2 $X2=0 $Y2=0
cc_261 N_VPWRIN_c_220_n N_X_M1000_d 0.00229479f $X=2.225 $Y=2.2 $X2=2.685
+ $Y2=4.555
cc_262 N_VPWRIN_c_220_n X 0.0277336f $X=2.225 $Y=2.2 $X2=0 $Y2=0
cc_263 N_A_505_297#_c_301_n N_A_714_58#_c_362_n 0.0441264f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_264 N_A_505_297#_c_289_n N_A_714_58#_c_363_n 6.95188e-19 $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_265 N_A_505_297#_c_294_n N_A_714_58#_c_363_n 3.7852e-19 $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_266 N_A_505_297#_c_301_n N_A_714_58#_c_364_n 0.00788518f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_267 N_A_505_297#_c_300_n N_A_714_58#_c_365_n 0.0048486f $X=3.06 $Y=2.25 $X2=0
+ $Y2=0
cc_268 N_A_505_297#_c_301_n N_A_714_58#_c_365_n 9.66994e-19 $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_269 N_A_505_297#_c_300_n N_A_714_58#_c_366_n 0.00327676f $X=3.06 $Y=2.25
+ $X2=0 $Y2=0
cc_270 N_A_505_297#_c_301_n N_A_714_58#_c_366_n 0.00125462f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_271 N_A_505_297#_c_301_n N_A_714_58#_c_380_n 0.0084582f $X=3.225 $Y=3.84
+ $X2=0.23 $Y2=4.8
cc_272 N_A_505_297#_c_295_n N_A_M1009_g 0.0110528f $X=2.675 $Y=0.62 $X2=3.135
+ $Y2=0.29
cc_273 N_A_505_297#_c_301_n N_A_M1009_g 0.0027023f $X=3.225 $Y=3.84 $X2=3.135
+ $Y2=0.29
cc_274 N_A_505_297#_c_295_n N_A_c_463_n 0.010267f $X=2.675 $Y=0.62 $X2=4
+ $Y2=0.29
cc_275 N_A_505_297#_c_295_n N_A_c_468_n 0.0218308f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_276 N_A_505_297#_c_295_n N_A_M1005_g 0.00336998f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_277 N_A_505_297#_c_295_n N_A_c_475_n 0.00146935f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_278 N_A_505_297#_c_295_n N_A_c_497_n 0.0360803f $X=2.675 $Y=0.62 $X2=0 $Y2=0
cc_279 N_A_505_297#_c_300_n N_A_c_497_n 0.00941491f $X=3.06 $Y=2.25 $X2=0 $Y2=0
cc_280 N_A_505_297#_c_289_n N_A_620_911#_c_536_n 0.0155516f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_281 N_A_505_297#_c_289_n N_A_620_911#_M1008_g 0.00777355f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_282 N_A_505_297#_c_274_n N_A_620_911#_c_541_n 0.00968676f $X=3.025 $Y=4.48
+ $X2=-0.19 $Y2=-0.24
cc_283 N_A_505_297#_c_278_n N_A_620_911#_c_541_n 0.00843936f $X=3.455 $Y=4.48
+ $X2=-0.19 $Y2=-0.24
cc_284 N_A_505_297#_c_284_n N_A_620_911#_c_541_n 0.0169132f $X=3.53 $Y=4.405
+ $X2=-0.19 $Y2=-0.24
cc_285 N_A_505_297#_c_285_n N_A_620_911#_c_541_n 2.89638e-19 $X=3.885 $Y=4.48
+ $X2=-0.19 $Y2=-0.24
cc_286 N_A_505_297#_c_284_n N_A_620_911#_c_545_n 0.021891f $X=3.53 $Y=4.405
+ $X2=0.23 $Y2=0.085
cc_287 N_A_505_297#_c_302_n N_A_620_911#_c_545_n 0.00420454f $X=3.225 $Y=3.84
+ $X2=0.23 $Y2=0.085
cc_288 N_A_505_297#_c_301_n N_A_620_911#_c_572_n 0.0218015f $X=3.225 $Y=3.84
+ $X2=0.23 $Y2=0.64
cc_289 N_A_505_297#_c_302_n N_A_620_911#_c_572_n 0.0175078f $X=3.225 $Y=3.84
+ $X2=0.23 $Y2=0.64
cc_290 N_A_505_297#_c_278_n N_A_620_911#_c_547_n 2.89638e-19 $X=3.455 $Y=4.48
+ $X2=0 $Y2=0
cc_291 N_A_505_297#_c_285_n N_A_620_911#_c_547_n 0.00843936f $X=3.885 $Y=4.48
+ $X2=0 $Y2=0
cc_292 N_A_505_297#_c_289_n N_A_620_911#_c_547_n 0.0149859f $X=4.24 $Y=4.405
+ $X2=0 $Y2=0
cc_293 N_A_505_297#_c_290_n N_A_620_911#_c_547_n 0.00985995f $X=4.315 $Y=4.48
+ $X2=0 $Y2=0
cc_294 N_A_505_297#_c_294_n N_A_620_911#_c_547_n 0.00418634f $X=3.885 $Y=4.405
+ $X2=0 $Y2=0
cc_295 N_A_505_297#_c_301_n N_A_620_911#_c_551_n 0.00421035f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_296 N_A_505_297#_c_302_n N_A_620_911#_c_551_n 0.0112331f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_297 N_A_505_297#_c_301_n N_A_620_911#_c_552_n 0.00372705f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_298 N_A_505_297#_c_302_n N_A_620_911#_c_552_n 0.0022314f $X=3.225 $Y=3.84
+ $X2=0 $Y2=0
cc_299 N_A_505_297#_c_294_n N_A_620_911#_c_556_n 0.0155516f $X=3.885 $Y=4.405
+ $X2=3.67 $Y2=4.735
cc_300 N_A_505_297#_M1009_d N_VPWR_c_728_n 0.00146082f $X=2.525 $Y=1.485 $X2=0
+ $Y2=0
cc_301 N_A_505_297#_c_300_n N_VPWR_c_728_n 0.00782153f $X=3.06 $Y=2.25 $X2=0
+ $Y2=0
cc_302 N_A_505_297#_c_311_n N_VPWR_c_728_n 0.00276885f $X=2.8 $Y=2.25 $X2=0
+ $Y2=0
cc_303 N_A_505_297#_c_301_n N_VPWR_c_728_n 0.0490709f $X=3.225 $Y=3.84 $X2=0
+ $Y2=0
cc_304 N_A_714_58#_c_371_n N_A_M1005_g 0.00122167f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_305 N_A_714_58#_c_371_n N_A_c_474_n 0.00391065f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_306 N_A_714_58#_c_365_n N_A_M1006_g 0.00224176f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_307 N_A_714_58#_c_371_n N_A_M1006_g 0.0163574f $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_308 N_A_714_58#_c_365_n N_A_c_482_n 0.0205035f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_309 N_A_714_58#_c_371_n N_A_c_482_n 6.96042e-19 $X=4.19 $Y=0.855 $X2=0 $Y2=0
cc_310 N_A_714_58#_c_365_n N_A_M1011_g 0.00205104f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_311 N_A_714_58#_c_367_n N_A_M1011_g 0.0163574f $X=4.475 $Y=0.855 $X2=0 $Y2=0
cc_312 N_A_714_58#_M1015_g N_A_c_488_n 0.0124308f $X=4.78 $Y=1.955 $X2=0 $Y2=0
cc_313 N_A_714_58#_c_376_n N_A_c_488_n 0.00295241f $X=4.57 $Y=0.73 $X2=0 $Y2=0
cc_314 N_A_714_58#_c_376_n N_A_M1012_g 6.61267e-19 $X=4.57 $Y=0.73 $X2=0 $Y2=0
cc_315 N_A_714_58#_c_366_n N_A_c_495_n 0.0062571f $X=4.105 $Y=2.07 $X2=0 $Y2=0
cc_316 N_A_714_58#_c_381_n N_A_620_911#_c_557_n 0.0315412f $X=4.705 $Y=2.58
+ $X2=0 $Y2=0
cc_317 N_A_714_58#_c_363_n N_A_620_911#_c_557_n 4.83528e-19 $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_318 N_A_714_58#_c_388_n N_A_620_911#_c_557_n 0.00503951f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_319 N_A_714_58#_c_358_n N_A_620_911#_c_535_n 0.0315412f $X=4.27 $Y=2.58 $X2=0
+ $Y2=0
cc_320 N_A_714_58#_c_362_n N_A_620_911#_c_535_n 0.0158995f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_321 N_A_714_58#_c_380_n N_A_620_911#_c_535_n 9.48385e-19 $X=4.105 $Y=2.49
+ $X2=0 $Y2=0
cc_322 N_A_714_58#_c_363_n N_A_620_911#_c_536_n 0.00905183f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_323 N_A_714_58#_c_363_n N_A_620_911#_M1001_g 0.00273734f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_324 N_A_714_58#_c_388_n N_A_620_911#_M1001_g 0.00383717f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_325 N_A_714_58#_c_363_n N_A_620_911#_c_545_n 0.00177263f $X=4.39 $Y=3.555
+ $X2=0.23 $Y2=0.085
cc_326 N_A_714_58#_c_364_n N_A_620_911#_c_545_n 0.0036785f $X=3.85 $Y=3.555
+ $X2=0.23 $Y2=0.085
cc_327 N_A_714_58#_c_362_n N_A_620_911#_c_573_n 0.0272967f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_328 N_A_714_58#_c_363_n N_A_620_911#_c_573_n 0.0109877f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_329 N_A_714_58#_c_388_n N_A_620_911#_c_573_n 0.014378f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_330 N_A_714_58#_c_363_n N_A_620_911#_c_551_n 0.0241447f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_331 N_A_714_58#_c_388_n N_A_620_911#_c_551_n 0.00429612f $X=4.555 $Y=3.235
+ $X2=0 $Y2=0
cc_332 N_A_714_58#_c_363_n N_A_620_911#_c_552_n 0.0112348f $X=4.39 $Y=3.555
+ $X2=0 $Y2=0
cc_333 N_A_714_58#_c_358_n N_A_620_911#_c_553_n 0.00516777f $X=4.27 $Y=2.58
+ $X2=2.81 $Y2=4.7
cc_334 N_A_714_58#_c_363_n N_A_620_911#_c_553_n 0.00294758f $X=4.39 $Y=3.555
+ $X2=2.81 $Y2=4.7
cc_335 N_A_714_58#_c_388_n N_A_620_911#_c_553_n 0.0174384f $X=4.555 $Y=3.235
+ $X2=2.81 $Y2=4.7
cc_336 N_A_714_58#_c_358_n N_A_620_911#_c_554_n 9.46557e-19 $X=4.27 $Y=2.58
+ $X2=0 $Y2=0
cc_337 N_A_714_58#_c_362_n N_A_620_911#_c_554_n 0.0121174f $X=3.765 $Y=3.47
+ $X2=0 $Y2=0
cc_338 N_A_714_58#_c_380_n N_A_620_911#_c_554_n 0.0118139f $X=4.105 $Y=2.49
+ $X2=0 $Y2=0
cc_339 N_A_714_58#_c_381_n N_A_620_911#_c_579_n 0.0110028f $X=4.705 $Y=2.58
+ $X2=3.28 $Y2=0.475
cc_340 N_A_714_58#_M1015_g N_A_620_911#_c_579_n 0.0043455f $X=4.78 $Y=1.955
+ $X2=3.28 $Y2=0.475
cc_341 N_A_714_58#_c_362_n N_A_620_911#_c_579_n 0.00251195f $X=3.765 $Y=3.47
+ $X2=3.28 $Y2=0.475
cc_342 N_A_714_58#_c_365_n N_A_620_911#_c_579_n 0.0372645f $X=4.105 $Y=2.07
+ $X2=3.28 $Y2=0.475
cc_343 N_A_714_58#_c_366_n N_A_620_911#_c_579_n 0.00490309f $X=4.105 $Y=2.07
+ $X2=3.28 $Y2=0.475
cc_344 N_A_714_58#_c_376_n N_A_620_911#_c_579_n 0.005679f $X=4.57 $Y=0.73
+ $X2=3.28 $Y2=0.475
cc_345 N_A_714_58#_c_380_n N_A_620_911#_c_579_n 0.00754333f $X=4.105 $Y=2.49
+ $X2=3.28 $Y2=0.475
cc_346 N_A_714_58#_c_363_n N_A_620_911#_c_555_n 0.00345728f $X=4.39 $Y=3.555
+ $X2=3.67 $Y2=5.355
cc_347 N_A_714_58#_c_381_n N_A_1028_32#_M1000_g 0.0107884f $X=4.705 $Y=2.58
+ $X2=0 $Y2=0
cc_348 N_A_714_58#_M1015_g N_A_1028_32#_c_664_n 0.0107884f $X=4.78 $Y=1.955
+ $X2=0 $Y2=0
cc_349 N_A_714_58#_M1015_g N_VPWR_c_730_n 0.00284928f $X=4.78 $Y=1.955 $X2=0
+ $Y2=0
cc_350 N_A_714_58#_c_363_n N_VPWR_c_731_n 0.0121345f $X=4.39 $Y=3.555 $X2=0
+ $Y2=0
cc_351 N_A_714_58#_c_388_n N_VPWR_c_731_n 0.0145663f $X=4.555 $Y=3.235 $X2=0
+ $Y2=0
cc_352 N_A_714_58#_c_381_n N_VPWR_c_728_n 0.00485266f $X=4.705 $Y=2.58 $X2=0
+ $Y2=0
cc_353 N_A_714_58#_c_358_n N_VPWR_c_728_n 0.00298594f $X=4.27 $Y=2.58 $X2=0
+ $Y2=0
cc_354 N_A_714_58#_M1015_g N_VPWR_c_728_n 0.00196242f $X=4.78 $Y=1.955 $X2=0
+ $Y2=0
cc_355 N_A_714_58#_c_362_n N_VPWR_c_728_n 0.0244983f $X=3.765 $Y=3.47 $X2=0
+ $Y2=0
cc_356 N_A_714_58#_c_363_n N_VPWR_c_728_n 0.0055128f $X=4.39 $Y=3.555 $X2=0
+ $Y2=0
cc_357 N_A_714_58#_c_365_n N_VPWR_c_728_n 2.07821e-19 $X=4.105 $Y=2.07 $X2=0
+ $Y2=0
cc_358 N_A_714_58#_c_366_n N_VPWR_c_728_n 0.00102999f $X=4.105 $Y=2.07 $X2=0
+ $Y2=0
cc_359 N_A_714_58#_c_388_n N_VPWR_c_728_n 0.00647659f $X=4.555 $Y=3.235 $X2=0
+ $Y2=0
cc_360 N_A_714_58#_c_380_n N_VPWR_c_728_n 0.0186535f $X=4.105 $Y=2.49 $X2=0
+ $Y2=0
cc_361 N_A_714_58#_c_376_n X 0.00128222f $X=4.57 $Y=0.73 $X2=0 $Y2=0
cc_362 N_A_714_58#_M1015_g X 0.00145345f $X=4.78 $Y=1.955 $X2=0 $Y2=0
cc_363 N_A_c_488_n N_A_620_911#_c_579_n 0.0037239f $X=4.71 $Y=1.145 $X2=3.28
+ $Y2=0.475
cc_364 N_A_M1012_g N_A_1028_32#_c_660_n 0.0104298f $X=4.785 $Y=0.615 $X2=4.86
+ $Y2=0.29
cc_365 N_A_c_488_n N_A_1028_32#_c_664_n 0.0104298f $X=4.71 $Y=1.145 $X2=0 $Y2=0
cc_366 N_A_M1009_g N_VPWR_c_728_n 0.00543198f $X=2.45 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A_M1012_g X 9.61814e-19 $X=4.785 $Y=0.615 $X2=0 $Y2=0
cc_368 N_A_620_911#_c_563_n N_A_1028_32#_c_674_n 0.0106294f $X=5.16 $Y=2.94
+ $X2=0 $Y2=0
cc_369 N_A_620_911#_c_563_n N_A_1028_32#_c_676_n 0.0121261f $X=5.16 $Y=2.94
+ $X2=0 $Y2=0
cc_370 N_A_620_911#_M1002_g N_A_1028_32#_c_681_n 0.00786959f $X=5.235 $Y=3.485
+ $X2=0 $Y2=0
cc_371 N_A_620_911#_M1008_g N_A_1028_32#_c_666_n 0.0254294f $X=5.085 $Y=4.88
+ $X2=0 $Y2=0
cc_372 N_A_620_911#_c_570_n N_A_1028_32#_c_666_n 0.00641748f $X=5.235 $Y=4.045
+ $X2=0 $Y2=0
cc_373 N_A_620_911#_M1008_g N_A_1028_32#_c_670_n 0.00384336f $X=5.085 $Y=4.88
+ $X2=0 $Y2=0
cc_374 N_A_620_911#_M1002_g N_A_1028_32#_c_670_n 0.0121261f $X=5.235 $Y=3.485
+ $X2=0 $Y2=0
cc_375 N_A_620_911#_c_579_n N_VPWR_c_730_n 0.035645f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_376 N_A_620_911#_c_563_n N_VPWR_c_731_n 0.0189101f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_377 N_A_620_911#_c_564_n N_VPWR_c_731_n 0.00521099f $X=5.01 $Y=4.045 $X2=0
+ $Y2=0
cc_378 N_A_620_911#_c_553_n N_VPWR_c_731_n 0.00509169f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_379 N_A_620_911#_c_553_n N_VPWR_c_733_n 0.00305029f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_380 N_A_620_911#_c_579_n N_VPWR_c_733_n 0.00537241f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_381 N_A_620_911#_c_563_n N_VPWR_c_736_n 0.00433894f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_382 N_A_620_911#_c_557_n N_VPWR_c_728_n 0.00365797f $X=4.705 $Y=2.94 $X2=0
+ $Y2=0
cc_383 N_A_620_911#_c_535_n N_VPWR_c_728_n 0.00398455f $X=4.27 $Y=2.94 $X2=0
+ $Y2=0
cc_384 N_A_620_911#_c_563_n N_VPWR_c_728_n 0.0064951f $X=5.16 $Y=2.94 $X2=0
+ $Y2=0
cc_385 N_A_620_911#_c_568_n N_VPWR_c_728_n 0.00339161f $X=4.78 $Y=2.94 $X2=0
+ $Y2=0
cc_386 N_A_620_911#_c_573_n N_VPWR_c_728_n 0.00622378f $X=4.105 $Y=3.135 $X2=0
+ $Y2=0
cc_387 N_A_620_911#_c_553_n N_VPWR_c_728_n 0.0219288f $X=4.47 $Y=2.83 $X2=0
+ $Y2=0
cc_388 N_A_620_911#_c_554_n N_VPWR_c_728_n 0.00663704f $X=4.19 $Y=2.83 $X2=0
+ $Y2=0
cc_389 N_A_620_911#_c_579_n N_VPWR_c_728_n 0.0165665f $X=4.555 $Y=1.79 $X2=0
+ $Y2=0
cc_390 N_A_1028_32#_M1000_g N_VPWR_c_730_n 0.00707023f $X=5.23 $Y=1.955 $X2=0
+ $Y2=0
cc_391 N_A_1028_32#_c_676_n N_VPWR_c_731_n 0.00238815f $X=5.775 $Y=4.015 $X2=0
+ $Y2=0
cc_392 N_A_1028_32#_c_681_n N_VPWR_c_731_n 0.00470553f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_393 N_A_1028_32#_c_673_n N_VPWR_c_736_n 0.0123843f $X=5.7 $Y=2.58 $X2=0 $Y2=0
cc_394 N_A_1028_32#_c_674_n N_VPWR_c_736_n 0.00491588f $X=5.305 $Y=2.58 $X2=0
+ $Y2=0
cc_395 N_A_1028_32#_c_676_n N_VPWR_c_736_n 0.0126975f $X=5.775 $Y=4.015 $X2=0
+ $Y2=0
cc_396 N_A_1028_32#_c_680_n N_VPWR_c_736_n 0.00431658f $X=5.775 $Y=2.58 $X2=0
+ $Y2=0
cc_397 N_A_1028_32#_c_681_n N_VPWR_c_736_n 0.00839796f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_398 N_A_1028_32#_M1000_g N_VPWR_c_728_n 0.00179018f $X=5.23 $Y=1.955 $X2=0
+ $Y2=0
cc_399 N_A_1028_32#_c_673_n N_VPWR_c_728_n 0.00231984f $X=5.7 $Y=2.58 $X2=0
+ $Y2=0
cc_400 N_A_1028_32#_c_674_n N_VPWR_c_728_n 0.00100275f $X=5.305 $Y=2.58 $X2=0
+ $Y2=0
cc_401 N_A_1028_32#_c_675_n N_VPWR_c_728_n 0.00204024f $X=5.775 $Y=2.505 $X2=0
+ $Y2=0
cc_402 N_A_1028_32#_c_676_n N_VPWR_c_728_n 0.00689358f $X=5.775 $Y=4.015 $X2=0
+ $Y2=0
cc_403 N_A_1028_32#_c_680_n N_VPWR_c_728_n 0.00208775f $X=5.775 $Y=2.58 $X2=0
+ $Y2=0
cc_404 N_A_1028_32#_c_681_n N_VPWR_c_728_n 0.00327036f $X=5.455 $Y=3.235 $X2=0
+ $Y2=0
cc_405 N_A_1028_32#_c_660_n X 0.00117381f $X=5.215 $Y=1.015 $X2=0 $Y2=0
cc_406 N_A_1028_32#_c_664_n X 0.0013393f $X=5.23 $Y=1.25 $X2=0 $Y2=0
cc_407 N_A_1028_32#_c_660_n X 0.00137501f $X=5.215 $Y=1.015 $X2=0 $Y2=0
cc_408 N_A_1028_32#_M1000_g X 6.87819e-19 $X=5.23 $Y=1.955 $X2=0 $Y2=0
cc_409 N_A_1028_32#_c_673_n X 0.00413561f $X=5.7 $Y=2.58 $X2=0 $Y2=0
cc_410 N_A_1028_32#_c_675_n X 0.02096f $X=5.775 $Y=2.505 $X2=0 $Y2=0
cc_411 N_A_1028_32#_c_664_n X 0.0569333f $X=5.23 $Y=1.25 $X2=0 $Y2=0
cc_412 N_VPWR_c_730_n X 0.00475824f $X=5.005 $Y=1.79 $X2=0 $Y2=0
cc_413 N_VPWR_c_736_n X 0.0113211f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_728_n X 0.00302523f $X=6.21 $Y=2.72 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=2.0496e+12p ps=1.849e+07u
M1001 Q_N a_1887_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.1888e+12p ps=1.291e+07u
M1002 Q a_2596_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1003 VGND a_1887_21# a_1822_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1004 a_1241_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=3.705e+11p pd=3.79e+06u as=0p ps=0u
M1005 VPWR RESET_B a_1396_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1006 a_2004_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=4.041e+11p pd=3.95e+06u as=0p ps=0u
M1007 a_381_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_1887_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.457e+11p pd=2.34e+06u as=0p ps=0u
M1009 VGND a_1102_21# a_1030_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.467e+11p ps=1.56e+06u
M1010 a_1714_47# a_27_47# a_1614_47# VNB nshort w=360000u l=150000u
+  ad=1.404e+11p pd=1.5e+06u as=1.96e+11p ps=1.98e+06u
M1011 a_1017_413# a_193_47# a_917_47# VPB phighvt w=420000u l=150000u
+  ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u
M1012 a_1102_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.94e+11p pd=2.46e+06u as=0p ps=0u
M1013 a_453_47# SCE a_381_47# VNB nshort w=420000u l=150000u
+  ad=2.559e+11p pd=2.92e+06u as=0p ps=0u
M1014 a_917_47# a_193_47# a_453_47# VNB nshort w=360000u l=150000u
+  ad=1.494e+11p pd=1.55e+06u as=0p ps=0u
M1015 VGND RESET_B a_1396_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1016 a_1614_47# a_1102_21# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_453_47# D a_752_413# VPB phighvt w=420000u l=150000u
+  ad=3.071e+11p pd=3.31e+06u as=1.134e+11p ps=1.38e+06u
M1018 Q a_2596_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1019 a_1800_413# a_27_47# a_1714_47# VPB phighvt w=420000u l=150000u
+  ad=1.848e+11p pd=1.72e+06u as=1.134e+11p ps=1.38e+06u
M1020 a_1887_21# a_1714_47# a_2004_47# VNB nshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1021 a_752_413# SCE VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1887_21# a_2596_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1023 a_2122_329# a_1714_47# a_1887_21# VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1024 a_1822_47# a_193_47# a_1714_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR CLK_N a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1026 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1027 a_453_47# D a_735_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1028 VPWR a_1396_21# a_2122_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_2004_47# a_1396_21# a_1887_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1396_21# a_1351_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1031 a_1714_47# a_193_47# a_1572_329# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.486e+11p ps=2.82e+06u
M1032 a_1241_47# a_1396_21# a_1102_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1033 a_381_363# SCD VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1034 VPWR SCE a_423_315# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1035 VPWR a_1102_21# a_1017_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1351_329# a_917_47# a_1102_21# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q_N a_1887_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1038 a_453_47# a_423_315# a_381_363# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_917_47# a_27_47# a_453_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1102_21# a_917_47# a_1241_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND SCE a_423_315# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1042 a_735_47# a_423_315# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_1887_21# a_1800_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1030_47# a_27_47# a_917_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND CLK_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1046 VGND a_1887_21# a_2596_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1047 a_1572_329# a_1102_21# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

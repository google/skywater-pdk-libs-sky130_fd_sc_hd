* File: sky130_fd_sc_hd__a2bb2o_2.pxi.spice
* Created: Thu Aug 27 14:03:17 2020
* 
x_PM_SKY130_FD_SC_HD__A2BB2O_2%A_82_21# N_A_82_21#_M1001_d N_A_82_21#_M1009_s
+ N_A_82_21#_c_76_n N_A_82_21#_M1007_g N_A_82_21#_M1002_g N_A_82_21#_c_77_n
+ N_A_82_21#_M1008_g N_A_82_21#_M1012_g N_A_82_21#_c_85_n N_A_82_21#_c_95_p
+ N_A_82_21#_c_136_p N_A_82_21#_c_86_n N_A_82_21#_c_87_n N_A_82_21#_c_88_n
+ N_A_82_21#_c_78_n N_A_82_21#_c_79_n N_A_82_21#_c_80_n N_A_82_21#_c_81_n
+ N_A_82_21#_c_91_n N_A_82_21#_c_82_n PM_SKY130_FD_SC_HD__A2BB2O_2%A_82_21#
x_PM_SKY130_FD_SC_HD__A2BB2O_2%A1_N N_A1_N_M1011_g N_A1_N_M1005_g A1_N A1_N
+ N_A1_N_c_191_n N_A1_N_c_192_n PM_SKY130_FD_SC_HD__A2BB2O_2%A1_N
x_PM_SKY130_FD_SC_HD__A2BB2O_2%A2_N N_A2_N_c_227_n N_A2_N_M1006_g N_A2_N_M1000_g
+ A2_N PM_SKY130_FD_SC_HD__A2BB2O_2%A2_N
x_PM_SKY130_FD_SC_HD__A2BB2O_2%A_313_47# N_A_313_47#_M1011_d N_A_313_47#_M1006_d
+ N_A_313_47#_c_258_n N_A_313_47#_M1001_g N_A_313_47#_c_259_n
+ N_A_313_47#_M1009_g N_A_313_47#_c_310_p N_A_313_47#_c_260_n
+ N_A_313_47#_c_261_n N_A_313_47#_c_264_n N_A_313_47#_c_265_n
+ N_A_313_47#_c_280_n PM_SKY130_FD_SC_HD__A2BB2O_2%A_313_47#
x_PM_SKY130_FD_SC_HD__A2BB2O_2%B2 N_B2_M1004_g N_B2_M1013_g B2 N_B2_c_320_n
+ N_B2_c_321_n PM_SKY130_FD_SC_HD__A2BB2O_2%B2
x_PM_SKY130_FD_SC_HD__A2BB2O_2%B1 N_B1_M1003_g N_B1_M1010_g B1 B1 B1
+ N_B1_c_366_n PM_SKY130_FD_SC_HD__A2BB2O_2%B1
x_PM_SKY130_FD_SC_HD__A2BB2O_2%VPWR N_VPWR_M1002_s N_VPWR_M1012_s N_VPWR_M1013_d
+ N_VPWR_c_394_n N_VPWR_c_395_n VPWR VPWR N_VPWR_c_397_n N_VPWR_c_398_n
+ N_VPWR_c_399_n N_VPWR_c_393_n N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n
+ VPWR PM_SKY130_FD_SC_HD__A2BB2O_2%VPWR
x_PM_SKY130_FD_SC_HD__A2BB2O_2%X N_X_M1007_s N_X_M1002_d N_X_c_457_n N_X_c_459_n
+ N_X_c_455_n X X X N_X_c_469_n PM_SKY130_FD_SC_HD__A2BB2O_2%X
x_PM_SKY130_FD_SC_HD__A2BB2O_2%A_574_369# N_A_574_369#_M1009_d
+ N_A_574_369#_M1010_d N_A_574_369#_c_483_n N_A_574_369#_c_481_n
+ N_A_574_369#_c_482_n N_A_574_369#_c_506_n N_A_574_369#_c_494_n
+ PM_SKY130_FD_SC_HD__A2BB2O_2%A_574_369#
x_PM_SKY130_FD_SC_HD__A2BB2O_2%VGND N_VGND_M1007_d N_VGND_M1008_d N_VGND_M1000_d
+ N_VGND_M1003_d N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n VGND VGND
+ N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n N_VGND_c_517_n N_VGND_c_518_n
+ N_VGND_c_519_n N_VGND_c_520_n VGND PM_SKY130_FD_SC_HD__A2BB2O_2%VGND
cc_1 VNB N_A_82_21#_c_76_n 0.0203464f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_A_82_21#_c_77_n 0.017306f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_A_82_21#_c_78_n 0.00168749f $X=-0.19 $Y=-0.24 $X2=2.765 $Y2=1.895
cc_4 VNB N_A_82_21#_c_79_n 0.00126207f $X=-0.19 $Y=-0.24 $X2=2.945 $Y2=0.445
cc_5 VNB N_A_82_21#_c_80_n 0.00405192f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_6 VNB N_A_82_21#_c_81_n 0.0477328f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_7 VNB N_A_82_21#_c_82_n 0.00849818f $X=-0.19 $Y=-0.24 $X2=2.945 $Y2=0.785
cc_8 VNB N_A1_N_M1011_g 0.0314275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A1_N_c_191_n 0.0208395f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_10 VNB N_A1_N_c_192_n 0.00632248f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_11 VNB N_A2_N_c_227_n 0.0213219f $X=-0.19 $Y=-0.24 $X2=2.81 $Y2=0.235
cc_12 VNB N_A2_N_M1000_g 0.0292979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A2_N 0.00262102f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.56
cc_14 VNB N_A_313_47#_c_258_n 0.0183385f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_15 VNB N_A_313_47#_c_259_n 0.061271f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.325
cc_16 VNB N_A_313_47#_c_260_n 0.0112681f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_17 VNB N_A_313_47#_c_261_n 0.00674176f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_18 VNB N_B2_M1004_g 0.0449337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B2_c_320_n 0.00452196f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_20 VNB N_B2_c_321_n 0.0100943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B1_M1003_g 0.0328058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB B1 0.0236663f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.56
cc_23 VNB N_B1_c_366_n 0.0395916f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_24 VNB N_VPWR_c_393_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_25 VNB N_X_c_455_n 0.00103298f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.985
cc_26 VNB N_VGND_c_510_n 0.00263482f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_27 VNB N_VGND_c_511_n 0.0128438f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.325
cc_28 VNB N_VGND_c_512_n 0.0192404f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_29 VNB VGND 0.0113688f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.325
cc_30 VNB N_VGND_c_514_n 0.0153157f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=2.2
cc_31 VNB N_VGND_c_515_n 0.0246972f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=1.16
cc_32 VNB N_VGND_c_516_n 0.00699789f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_33 VNB N_VGND_c_517_n 0.0148665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_518_n 0.0137885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_519_n 0.221737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_520_n 0.00868793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_A_82_21#_M1002_g 0.0242689f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_38 VPB N_A_82_21#_M1012_g 0.0204978f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_39 VPB N_A_82_21#_c_85_n 0.00111481f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.805
cc_40 VPB N_A_82_21#_c_86_n 6.73913e-19 $X=-0.19 $Y=1.305 $X2=1.625 $Y2=2.2
cc_41 VPB N_A_82_21#_c_87_n 0.0182324f $X=-0.19 $Y=1.305 $X2=2.44 $Y2=2.285
cc_42 VPB N_A_82_21#_c_88_n 0.0024581f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=2.285
cc_43 VPB N_A_82_21#_c_78_n 0.00450287f $X=-0.19 $Y=1.305 $X2=2.765 $Y2=1.895
cc_44 VPB N_A_82_21#_c_81_n 0.00810031f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_45 VPB N_A_82_21#_c_91_n 0.00489497f $X=-0.19 $Y=1.305 $X2=2.585 $Y2=2.275
cc_46 VPB N_A1_N_M1005_g 0.0181122f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.995
cc_47 VPB N_A1_N_c_191_n 0.0046179f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.995
cc_48 VPB N_A1_N_c_192_n 0.00267071f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.56
cc_49 VPB N_A2_N_c_227_n 0.0270662f $X=-0.19 $Y=1.305 $X2=2.81 $Y2=0.235
cc_50 VPB A2_N 0.00183417f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_51 VPB N_A_313_47#_c_259_n 0.0255619f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.325
cc_52 VPB N_A_313_47#_M1009_g 0.0391128f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_53 VPB N_A_313_47#_c_264_n 0.0103697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_313_47#_c_265_n 0.00191553f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=1.975
cc_55 VPB N_B2_M1013_g 0.0219077f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.995
cc_56 VPB B2 0.00846849f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_57 VPB N_B2_c_320_n 0.0249797f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.995
cc_58 VPB N_B2_c_321_n 8.181e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B1_M1010_g 0.0487316f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.995
cc_60 VPB B1 0.0161044f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_61 VPB N_B1_c_366_n 0.00754525f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.56
cc_62 VPB N_VPWR_c_394_n 0.00907939f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_63 VPB N_VPWR_c_395_n 0.00232023f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.56
cc_64 VPB VPWR 0.0113429f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_65 VPB N_VPWR_c_397_n 0.0153157f $X=-0.19 $Y=1.305 $X2=1.54 $Y2=1.89
cc_66 VPB N_VPWR_c_398_n 0.0523121f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=2.285
cc_67 VPB N_VPWR_c_399_n 0.0152513f $X=-0.19 $Y=1.305 $X2=0.992 $Y2=1.16
cc_68 VPB N_VPWR_c_393_n 0.0585297f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_69 VPB N_VPWR_c_401_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_402_n 0.0035381f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.16
cc_71 VPB N_VPWR_c_403_n 0.00845764f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=1.16
cc_72 VPB N_X_c_455_n 0.00108005f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_73 VPB N_A_574_369#_c_481_n 0.00483152f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_74 VPB N_A_574_369#_c_482_n 0.00148243f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.325
cc_75 N_A_82_21#_c_77_n N_A1_N_M1011_g 0.0182272f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_82_21#_M1012_g N_A1_N_M1005_g 0.0206265f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_82_21#_c_85_n N_A1_N_M1005_g 0.00451623f $X=1.035 $Y=1.805 $X2=0 $Y2=0
cc_78 N_A_82_21#_c_95_p N_A1_N_M1005_g 0.0109485f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_79 N_A_82_21#_c_86_n N_A1_N_M1005_g 0.00553351f $X=1.625 $Y=2.2 $X2=0 $Y2=0
cc_80 N_A_82_21#_c_88_n N_A1_N_M1005_g 0.00194344f $X=1.71 $Y=2.285 $X2=0 $Y2=0
cc_81 N_A_82_21#_c_95_p N_A1_N_c_191_n 0.00156259f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_82 N_A_82_21#_c_80_n N_A1_N_c_191_n 0.00197826f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_82_21#_c_81_n N_A1_N_c_191_n 0.0204271f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_82_21#_M1012_g N_A1_N_c_192_n 8.79726e-19 $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_85 N_A_82_21#_c_95_p N_A1_N_c_192_n 0.0156175f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_86 N_A_82_21#_c_80_n N_A1_N_c_192_n 0.0392215f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_82_21#_c_81_n N_A1_N_c_192_n 3.57546e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_82_21#_c_95_p N_A2_N_c_227_n 0.003006f $X=1.54 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_82_21#_c_86_n N_A2_N_c_227_n 0.00505208f $X=1.625 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_82_21#_c_87_n N_A2_N_c_227_n 0.0116667f $X=2.44 $Y=2.285 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_82_21#_c_91_n N_A2_N_c_227_n 0.00762679f $X=2.585 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_82_21#_c_79_n N_A_313_47#_c_258_n 4.8064e-19 $X=2.945 $Y=0.445 $X2=0
+ $Y2=0
cc_93 N_A_82_21#_c_82_n N_A_313_47#_c_258_n 0.00476835f $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_94 N_A_82_21#_c_78_n N_A_313_47#_c_259_n 0.0220074f $X=2.765 $Y=1.895 $X2=0
+ $Y2=0
cc_95 N_A_82_21#_c_91_n N_A_313_47#_c_259_n 0.0058762f $X=2.585 $Y=2.275 $X2=0
+ $Y2=0
cc_96 N_A_82_21#_c_82_n N_A_313_47#_c_259_n 0.00503935f $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_97 N_A_82_21#_c_78_n N_A_313_47#_M1009_g 0.0162553f $X=2.765 $Y=1.895 $X2=0
+ $Y2=0
cc_98 N_A_82_21#_c_91_n N_A_313_47#_M1009_g 0.00936639f $X=2.585 $Y=2.275 $X2=0
+ $Y2=0
cc_99 N_A_82_21#_c_79_n N_A_313_47#_c_260_n 0.00227074f $X=2.945 $Y=0.445 $X2=0
+ $Y2=0
cc_100 N_A_82_21#_c_82_n N_A_313_47#_c_260_n 0.010242f $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_101 N_A_82_21#_c_87_n N_A_313_47#_c_264_n 0.0110871f $X=2.44 $Y=2.285 $X2=0
+ $Y2=0
cc_102 N_A_82_21#_c_78_n N_A_313_47#_c_264_n 0.013656f $X=2.765 $Y=1.895 $X2=0
+ $Y2=0
cc_103 N_A_82_21#_c_91_n N_A_313_47#_c_264_n 0.00605907f $X=2.585 $Y=2.275 $X2=0
+ $Y2=0
cc_104 N_A_82_21#_c_78_n N_A_313_47#_c_265_n 0.04654f $X=2.765 $Y=1.895 $X2=0
+ $Y2=0
cc_105 N_A_82_21#_c_82_n N_A_313_47#_c_265_n 0.00313949f $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_106 N_A_82_21#_c_87_n N_A_313_47#_c_280_n 0.00792284f $X=2.44 $Y=2.285 $X2=0
+ $Y2=0
cc_107 N_A_82_21#_c_78_n N_A_313_47#_c_280_n 0.00501479f $X=2.765 $Y=1.895 $X2=0
+ $Y2=0
cc_108 N_A_82_21#_c_91_n N_A_313_47#_c_280_n 5.37178e-19 $X=2.585 $Y=2.275 $X2=0
+ $Y2=0
cc_109 N_A_82_21#_c_78_n N_B2_M1004_g 0.00238194f $X=2.765 $Y=1.895 $X2=0 $Y2=0
cc_110 N_A_82_21#_c_79_n N_B2_M1004_g 0.00111676f $X=2.945 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_82_21#_c_82_n N_B2_M1004_g 0.00266107f $X=2.945 $Y=0.785 $X2=0 $Y2=0
cc_112 N_A_82_21#_c_78_n N_B2_M1013_g 0.00115651f $X=2.765 $Y=1.895 $X2=0 $Y2=0
cc_113 N_A_82_21#_c_78_n B2 0.0206288f $X=2.765 $Y=1.895 $X2=0 $Y2=0
cc_114 N_A_82_21#_c_78_n N_B2_c_320_n 3.22868e-19 $X=2.765 $Y=1.895 $X2=0 $Y2=0
cc_115 N_A_82_21#_c_78_n N_B2_c_321_n 0.0187734f $X=2.765 $Y=1.895 $X2=0 $Y2=0
cc_116 N_A_82_21#_c_82_n N_B2_c_321_n 0.00673007f $X=2.945 $Y=0.785 $X2=0 $Y2=0
cc_117 N_A_82_21#_c_85_n N_VPWR_M1012_s 0.00369532f $X=1.035 $Y=1.805 $X2=0
+ $Y2=0
cc_118 N_A_82_21#_c_95_p N_VPWR_M1012_s 0.0117288f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_119 N_A_82_21#_c_136_p N_VPWR_M1012_s 0.00106957f $X=1.12 $Y=1.89 $X2=0 $Y2=0
cc_120 N_A_82_21#_M1002_g N_VPWR_c_394_n 6.18893e-19 $X=0.485 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_82_21#_M1012_g N_VPWR_c_394_n 0.00825406f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_82_21#_c_95_p N_VPWR_c_394_n 0.00862919f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_123 N_A_82_21#_c_136_p N_VPWR_c_394_n 0.00642951f $X=1.12 $Y=1.89 $X2=0 $Y2=0
cc_124 N_A_82_21#_c_88_n N_VPWR_c_394_n 0.00877693f $X=1.71 $Y=2.285 $X2=0 $Y2=0
cc_125 N_A_82_21#_M1002_g N_VPWR_c_397_n 0.00533769f $X=0.485 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_82_21#_M1012_g N_VPWR_c_397_n 0.0046653f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_82_21#_c_95_p N_VPWR_c_398_n 0.00309642f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_128 N_A_82_21#_c_87_n N_VPWR_c_398_n 0.0294488f $X=2.44 $Y=2.285 $X2=0 $Y2=0
cc_129 N_A_82_21#_c_88_n N_VPWR_c_398_n 0.00749299f $X=1.71 $Y=2.285 $X2=0 $Y2=0
cc_130 N_A_82_21#_c_91_n N_VPWR_c_398_n 0.0168205f $X=2.585 $Y=2.275 $X2=0 $Y2=0
cc_131 N_A_82_21#_M1009_s N_VPWR_c_393_n 0.00231177f $X=2.46 $Y=1.845 $X2=0
+ $Y2=0
cc_132 N_A_82_21#_M1002_g N_VPWR_c_393_n 0.0103364f $X=0.485 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_82_21#_M1012_g N_VPWR_c_393_n 0.00796766f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_82_21#_c_95_p N_VPWR_c_393_n 0.00736589f $X=1.54 $Y=1.89 $X2=0 $Y2=0
cc_135 N_A_82_21#_c_136_p N_VPWR_c_393_n 8.6225e-19 $X=1.12 $Y=1.89 $X2=0 $Y2=0
cc_136 N_A_82_21#_c_87_n N_VPWR_c_393_n 0.0255669f $X=2.44 $Y=2.285 $X2=0 $Y2=0
cc_137 N_A_82_21#_c_88_n N_VPWR_c_393_n 0.00618211f $X=1.71 $Y=2.285 $X2=0 $Y2=0
cc_138 N_A_82_21#_c_91_n N_VPWR_c_393_n 0.0133196f $X=2.585 $Y=2.275 $X2=0 $Y2=0
cc_139 N_A_82_21#_M1002_g N_VPWR_c_403_n 0.0039228f $X=0.485 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_82_21#_c_76_n N_X_c_457_n 0.00192423f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_82_21#_c_81_n N_X_c_457_n 0.00190599f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_82_21#_M1002_g N_X_c_459_n 0.00179207f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_82_21#_c_81_n N_X_c_459_n 0.00193622f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_82_21#_c_76_n N_X_c_455_n 0.00523711f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_82_21#_M1002_g N_X_c_455_n 0.00714657f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_82_21#_c_77_n N_X_c_455_n 0.00395119f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_82_21#_M1012_g N_X_c_455_n 0.00136611f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_82_21#_c_85_n N_X_c_455_n 0.0104644f $X=1.035 $Y=1.805 $X2=0 $Y2=0
cc_149 N_A_82_21#_c_80_n N_X_c_455_n 0.0230865f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_82_21#_c_81_n N_X_c_455_n 0.024289f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_82_21#_c_76_n X 0.00610081f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_82_21#_M1002_g N_X_c_469_n 0.0105532f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_82_21#_c_95_p A_313_297# 0.00411397f $X=1.54 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_82_21#_c_86_n A_313_297# 0.00164129f $X=1.625 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_82_21#_c_91_n N_A_574_369#_c_483_n 0.00420617f $X=2.585 $Y=2.275
+ $X2=0 $Y2=0
cc_156 N_A_82_21#_c_78_n N_A_574_369#_c_482_n 0.00442235f $X=2.765 $Y=1.895
+ $X2=0 $Y2=0
cc_157 N_A_82_21#_c_91_n N_A_574_369#_c_482_n 0.00867828f $X=2.585 $Y=2.275
+ $X2=0 $Y2=0
cc_158 N_A_82_21#_c_76_n N_VGND_c_510_n 6.58943e-19 $X=0.485 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_82_21#_c_77_n N_VGND_c_510_n 0.00849001f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_82_21#_c_80_n N_VGND_c_510_n 0.00551674f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_82_21#_c_81_n N_VGND_c_510_n 4.58244e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_82_21#_c_76_n N_VGND_c_514_n 0.00533769f $X=0.485 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_82_21#_c_77_n N_VGND_c_514_n 0.0046653f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_82_21#_c_79_n N_VGND_c_515_n 0.0110645f $X=2.945 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_82_21#_c_82_n N_VGND_c_515_n 0.00251982f $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_166 N_A_82_21#_c_82_n N_VGND_c_518_n 5.80399e-19 $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_167 N_A_82_21#_M1001_d N_VGND_c_519_n 0.00413042f $X=2.81 $Y=0.235 $X2=0
+ $Y2=0
cc_168 N_A_82_21#_c_76_n N_VGND_c_519_n 0.0103364f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_82_21#_c_77_n N_VGND_c_519_n 0.00796766f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_82_21#_c_79_n N_VGND_c_519_n 0.00640047f $X=2.945 $Y=0.445 $X2=0
+ $Y2=0
cc_171 N_A_82_21#_c_82_n N_VGND_c_519_n 0.00407678f $X=2.945 $Y=0.785 $X2=0
+ $Y2=0
cc_172 N_A_82_21#_c_76_n N_VGND_c_520_n 0.00403247f $X=0.485 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A1_N_c_191_n N_A2_N_c_227_n 0.0736355f $X=1.43 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A1_N_c_192_n N_A2_N_c_227_n 0.00506264f $X=1.43 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A1_N_M1011_g N_A2_N_M1000_g 0.0240597f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A1_N_c_191_n A2_N 3.51879e-19 $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A1_N_c_192_n A2_N 0.0297809f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A1_N_M1011_g N_A_313_47#_c_261_n 0.00536216f $X=1.49 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A1_N_c_192_n N_A_313_47#_c_261_n 0.00541889f $X=1.43 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_A1_N_c_192_n N_A_313_47#_c_265_n 0.00486283f $X=1.43 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A1_N_c_192_n N_VPWR_M1012_s 0.00147965f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A1_N_M1005_g N_VPWR_c_398_n 0.0029384f $X=1.49 $Y=1.805 $X2=0 $Y2=0
cc_183 N_A1_N_M1005_g N_VPWR_c_393_n 0.00395811f $X=1.49 $Y=1.805 $X2=0 $Y2=0
cc_184 N_A1_N_c_192_n A_313_297# 0.0022125f $X=1.43 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_185 N_A1_N_M1011_g N_VGND_c_510_n 0.00364237f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A1_N_c_191_n N_VGND_c_510_n 0.00176065f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A1_N_c_192_n N_VGND_c_510_n 8.57019e-19 $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A1_N_M1011_g N_VGND_c_517_n 0.00585385f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A1_N_M1011_g N_VGND_c_518_n 5.89496e-19 $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A1_N_M1011_g N_VGND_c_519_n 0.0110737f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A2_N_M1000_g N_A_313_47#_c_258_n 0.00378302f $X=1.91 $Y=0.445 $X2=0
+ $Y2=0
cc_192 N_A2_N_c_227_n N_A_313_47#_c_259_n 0.0235992f $X=1.85 $Y=1.375 $X2=0
+ $Y2=0
cc_193 N_A2_N_M1000_g N_A_313_47#_c_259_n 0.0102385f $X=1.91 $Y=0.445 $X2=0
+ $Y2=0
cc_194 A2_N N_A_313_47#_c_259_n 0.00265567f $X=1.965 $Y=1.105 $X2=0 $Y2=0
cc_195 N_A2_N_c_227_n N_A_313_47#_c_260_n 0.00377055f $X=1.85 $Y=1.375 $X2=0
+ $Y2=0
cc_196 N_A2_N_M1000_g N_A_313_47#_c_260_n 0.0122585f $X=1.91 $Y=0.445 $X2=0
+ $Y2=0
cc_197 A2_N N_A_313_47#_c_260_n 0.0218033f $X=1.965 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A2_N_c_227_n N_A_313_47#_c_261_n 3.76221e-19 $X=1.85 $Y=1.375 $X2=0
+ $Y2=0
cc_199 N_A2_N_c_227_n N_A_313_47#_c_265_n 0.00214962f $X=1.85 $Y=1.375 $X2=0
+ $Y2=0
cc_200 N_A2_N_M1000_g N_A_313_47#_c_265_n 9.47693e-19 $X=1.91 $Y=0.445 $X2=0
+ $Y2=0
cc_201 A2_N N_A_313_47#_c_265_n 0.0246561f $X=1.965 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A2_N_c_227_n N_A_313_47#_c_280_n 7.48305e-19 $X=1.85 $Y=1.375 $X2=0
+ $Y2=0
cc_203 A2_N N_A_313_47#_c_280_n 0.013002f $X=1.965 $Y=1.105 $X2=0 $Y2=0
cc_204 N_A2_N_c_227_n N_VPWR_c_398_n 6.45813e-19 $X=1.85 $Y=1.375 $X2=0 $Y2=0
cc_205 N_A2_N_M1000_g N_VGND_c_517_n 0.00341689f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A2_N_M1000_g N_VGND_c_518_n 0.00817983f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A2_N_M1000_g N_VGND_c_519_n 0.0040385f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A_313_47#_c_258_n N_B2_M1004_g 0.0249353f $X=2.735 $Y=0.765 $X2=0 $Y2=0
cc_209 N_A_313_47#_c_259_n N_B2_M1004_g 0.0179776f $X=2.795 $Y=1.435 $X2=0 $Y2=0
cc_210 N_A_313_47#_M1009_g N_B2_M1013_g 0.0252052f $X=2.795 $Y=2.165 $X2=0 $Y2=0
cc_211 N_A_313_47#_c_259_n B2 0.00178503f $X=2.795 $Y=1.435 $X2=0 $Y2=0
cc_212 N_A_313_47#_M1009_g N_B2_c_320_n 0.0179776f $X=2.795 $Y=2.165 $X2=0 $Y2=0
cc_213 N_A_313_47#_M1009_g N_VPWR_c_398_n 0.00448878f $X=2.795 $Y=2.165 $X2=0
+ $Y2=0
cc_214 N_A_313_47#_M1009_g N_VPWR_c_393_n 0.00798716f $X=2.795 $Y=2.165 $X2=0
+ $Y2=0
cc_215 N_A_313_47#_M1009_g N_A_574_369#_c_483_n 0.00148209f $X=2.795 $Y=2.165
+ $X2=0 $Y2=0
cc_216 N_A_313_47#_M1009_g N_A_574_369#_c_482_n 0.00118382f $X=2.795 $Y=2.165
+ $X2=0 $Y2=0
cc_217 N_A_313_47#_c_260_n N_VGND_M1000_d 0.00182057f $X=2.34 $Y=0.74 $X2=0
+ $Y2=0
cc_218 N_A_313_47#_c_258_n N_VGND_c_515_n 0.0034676f $X=2.735 $Y=0.765 $X2=0
+ $Y2=0
cc_219 N_A_313_47#_c_310_p N_VGND_c_517_n 0.0112554f $X=1.7 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_313_47#_c_260_n N_VGND_c_517_n 0.00273399f $X=2.34 $Y=0.74 $X2=0
+ $Y2=0
cc_221 N_A_313_47#_c_258_n N_VGND_c_518_n 0.00995519f $X=2.735 $Y=0.765 $X2=0
+ $Y2=0
cc_222 N_A_313_47#_c_259_n N_VGND_c_518_n 0.00636187f $X=2.795 $Y=1.435 $X2=0
+ $Y2=0
cc_223 N_A_313_47#_c_260_n N_VGND_c_518_n 0.0414636f $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_313_47#_M1011_d N_VGND_c_519_n 0.00412745f $X=1.565 $Y=0.235 $X2=0
+ $Y2=0
cc_225 N_A_313_47#_c_258_n N_VGND_c_519_n 0.00412709f $X=2.735 $Y=0.765 $X2=0
+ $Y2=0
cc_226 N_A_313_47#_c_310_p N_VGND_c_519_n 0.00644035f $X=1.7 $Y=0.445 $X2=0
+ $Y2=0
cc_227 N_A_313_47#_c_260_n N_VGND_c_519_n 0.00660739f $X=2.34 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_B2_M1004_g N_B1_M1003_g 0.0464258f $X=3.155 $Y=0.445 $X2=0 $Y2=0
cc_229 N_B2_c_321_n N_B1_M1003_g 0.00547864f $X=3.4 $Y=1.505 $X2=0 $Y2=0
cc_230 N_B2_M1013_g N_B1_M1010_g 0.0307678f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_231 B2 N_B1_M1010_g 0.00229097f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_232 B2 B1 0.0212548f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_233 N_B2_c_320_n B1 2.55263e-19 $X=3.215 $Y=1.47 $X2=0 $Y2=0
cc_234 N_B2_c_321_n B1 0.0391911f $X=3.4 $Y=1.505 $X2=0 $Y2=0
cc_235 N_B2_M1004_g N_B1_c_366_n 0.00402935f $X=3.155 $Y=0.445 $X2=0 $Y2=0
cc_236 N_B2_c_320_n N_B1_c_366_n 0.0158489f $X=3.215 $Y=1.47 $X2=0 $Y2=0
cc_237 N_B2_c_321_n N_B1_c_366_n 0.00649814f $X=3.4 $Y=1.505 $X2=0 $Y2=0
cc_238 N_B2_M1013_g N_VPWR_c_395_n 0.00279634f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_239 N_B2_M1013_g N_VPWR_c_398_n 0.00422411f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_240 N_B2_M1013_g N_VPWR_c_393_n 0.00583767f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_241 N_B2_M1013_g N_A_574_369#_c_483_n 0.00524398f $X=3.25 $Y=2.165 $X2=0
+ $Y2=0
cc_242 N_B2_M1013_g N_A_574_369#_c_481_n 0.00844573f $X=3.25 $Y=2.165 $X2=0
+ $Y2=0
cc_243 B2 N_A_574_369#_c_481_n 0.0235455f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_244 N_B2_M1013_g N_A_574_369#_c_482_n 0.00222048f $X=3.25 $Y=2.165 $X2=0
+ $Y2=0
cc_245 B2 N_A_574_369#_c_482_n 0.0123423f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_246 N_B2_c_320_n N_A_574_369#_c_482_n 6.67241e-19 $X=3.215 $Y=1.47 $X2=0
+ $Y2=0
cc_247 N_B2_M1013_g N_A_574_369#_c_494_n 0.00214984f $X=3.25 $Y=2.165 $X2=0
+ $Y2=0
cc_248 N_B2_M1004_g N_VGND_c_512_n 0.00224511f $X=3.155 $Y=0.445 $X2=0 $Y2=0
cc_249 N_B2_M1004_g N_VGND_c_515_n 0.00585385f $X=3.155 $Y=0.445 $X2=0 $Y2=0
cc_250 N_B2_M1004_g N_VGND_c_518_n 0.00126121f $X=3.155 $Y=0.445 $X2=0 $Y2=0
cc_251 N_B2_M1004_g N_VGND_c_519_n 0.0108681f $X=3.155 $Y=0.445 $X2=0 $Y2=0
cc_252 N_B2_c_321_n N_VGND_c_519_n 0.0104262f $X=3.4 $Y=1.505 $X2=0 $Y2=0
cc_253 N_B1_M1010_g N_VPWR_c_395_n 0.00884045f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_254 N_B1_M1010_g N_VPWR_c_399_n 0.00348405f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_255 N_B1_M1010_g N_VPWR_c_393_n 0.00513647f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_256 N_B1_M1010_g N_A_574_369#_c_483_n 4.53479e-19 $X=3.67 $Y=2.165 $X2=0
+ $Y2=0
cc_257 N_B1_M1010_g N_A_574_369#_c_481_n 0.0170411f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_258 B1 N_A_574_369#_c_481_n 0.0202429f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_259 N_B1_c_366_n N_A_574_369#_c_481_n 0.00237269f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B1_M1003_g N_VGND_c_512_n 0.0157597f $X=3.575 $Y=0.445 $X2=0 $Y2=0
cc_261 B1 N_VGND_c_512_n 0.0230984f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_262 N_B1_c_366_n N_VGND_c_512_n 0.00301045f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_M1003_g N_VGND_c_515_n 0.00407992f $X=3.575 $Y=0.445 $X2=0 $Y2=0
cc_264 N_B1_M1003_g N_VGND_c_519_n 0.00618209f $X=3.575 $Y=0.445 $X2=0 $Y2=0
cc_265 B1 N_VGND_c_519_n 0.00104546f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_266 N_VPWR_c_393_n N_X_M1002_d 0.00393857f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_267 N_VPWR_c_403_n N_X_c_455_n 0.0380133f $X=0.27 $Y=1.64 $X2=0 $Y2=0
cc_268 N_VPWR_c_397_n N_X_c_469_n 0.0155235f $X=0.95 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_c_393_n N_X_c_469_n 0.00958799f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_393_n N_A_574_369#_M1009_d 0.00242787f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_271 N_VPWR_c_393_n N_A_574_369#_M1010_d 0.00375766f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_272 N_VPWR_M1013_d N_A_574_369#_c_481_n 0.00161592f $X=3.325 $Y=1.845 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_395_n N_A_574_369#_c_481_n 0.014257f $X=3.46 $Y=2.34 $X2=0 $Y2=0
cc_274 N_VPWR_c_398_n N_A_574_369#_c_481_n 0.0020257f $X=3.375 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_399_n N_A_574_369#_c_481_n 0.00203142f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_393_n N_A_574_369#_c_481_n 0.00878585f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_399_n N_A_574_369#_c_506_n 0.0115413f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_393_n N_A_574_369#_c_506_n 0.00645703f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_398_n N_A_574_369#_c_494_n 0.0142246f $X=3.375 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_393_n N_A_574_369#_c_494_n 0.0117845f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_403_n N_VGND_c_520_n 0.00726759f $X=0.27 $Y=1.64 $X2=0 $Y2=0
cc_282 X N_VGND_c_514_n 0.0154428f $X=0.585 $Y=0.425 $X2=0 $Y2=0
cc_283 N_X_M1007_s N_VGND_c_519_n 0.00393857f $X=0.56 $Y=0.235 $X2=0 $Y2=0
cc_284 X N_VGND_c_519_n 0.00957098f $X=0.585 $Y=0.425 $X2=0 $Y2=0
cc_285 X N_VGND_c_520_n 0.0256705f $X=0.585 $Y=0.425 $X2=0 $Y2=0
cc_286 N_VGND_c_519_n A_646_47# 0.00486328f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__nand4_1.spice
* Created: Tue Sep  1 19:16:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4_1.pex.spice"
.subckt sky130_fd_sc_hd__nand4_1  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1007 A_109_47# N_D_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.5
+ A=0.0975 P=1.6 MULT=1
MM1002 A_193_47# N_C_M1002_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=14.76 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 A_277_47# N_B_M1004_g A_193_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=14.76 M=1 R=4.33333 SA=75001
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g A_277_47# VNB NSHORT L=0.15 W=0.65 AD=0.195
+ AS=0.10725 PD=1.9 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333 SA=75001.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_D_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.5 A=0.15
+ P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1 AD=0.3
+ AS=0.165 PD=2.6 PS=1.33 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75001.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_295 A_277_47# 0 1.04363e-19 $X=1.385 $Y=0.235
*
.include "sky130_fd_sc_hd__nand4_1.pxi.spice"
*
.ends
*
*

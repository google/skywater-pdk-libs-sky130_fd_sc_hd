* File: sky130_fd_sc_hd__dlxtp_1.pex.spice
* Created: Tue Sep  1 19:06:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLXTP_1%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39414e-20 $X=0.21 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.21 $Y=1.19
+ $X2=0.21 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%A_27_47# 1 2 9 13 17 19 20 23 27 30 34 35 36
+ 41 44 46 49 50 53 56 57 60 64
c146 57 0 7.63528e-20 $X=2.555 $Y=1.53
c147 13 0 2.69707e-20 $X=0.89 $Y=2.135
c148 9 0 2.69707e-20 $X=0.89 $Y=0.445
r149 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r150 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.53
+ $X2=2.555 $Y2=1.53
r151 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r152 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r153 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.53
+ $X2=2.555 $Y2=1.53
r154 49 50 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.41 $Y=1.53
+ $X2=0.84 $Y2=1.53
r155 48 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r156 47 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r157 45 64 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r158 44 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r159 44 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r160 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r161 38 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r162 37 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r163 36 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r164 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r165 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r166 34 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r167 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r168 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r169 26 60 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r170 26 27 40.8463 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r171 25 60 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r172 21 23 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.22 $Y=1.245
+ $X2=3.22 $Y2=0.415
r173 20 25 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r174 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=3.22 $Y2=1.245
r175 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=2.805 $Y2=1.32
r176 17 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.725 $Y=2.275
+ $X2=2.725 $Y2=1.685
r177 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r178 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r179 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r180 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r181 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r182 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 34 0 1.98767e-19 $X=2.255 $Y=0.765
c84 32 0 1.12109e-19 $X=2.255 $Y=0.93
c85 18 0 7.13094e-20 $X=1.97 $Y=0.7
r86 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r87 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r88 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r89 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r90 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r91 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r92 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r93 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r94 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r95 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r96 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r97 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r98 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r99 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r100 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r101 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r102 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%A_193_47# 1 2 9 12 16 20 24 26 28 29 32 35
+ 39 42 43 50
c124 42 0 7.63528e-20 $X=3.18 $Y=1.74
c125 26 0 1.98767e-19 $X=3.01 $Y=0.87
r126 43 50 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=1.74
+ $X2=3.095 $Y2=1.575
r127 42 45 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.18 $Y2=1.875
r128 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r129 35 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.87
+ $X2=3.015 $Y2=1.87
r130 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r131 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r132 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.87
+ $X2=3.015 $Y2=1.87
r133 28 29 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.87 $Y=1.87
+ $X2=1.3 $Y2=1.87
r134 24 39 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=2.792 $Y=0.87
+ $X2=2.792 $Y2=0.705
r135 23 26 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0.87
+ $X2=3.01 $Y2=0.87
r136 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=0.87 $X2=2.8 $Y2=0.87
r137 20 32 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r138 20 21 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r139 18 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=0.87
r140 18 50 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.575
r141 16 21 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r142 12 45 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.145 $Y=2.275
+ $X2=3.145 $Y2=1.875
r143 9 39 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.725 $Y=0.415
+ $X2=2.725 $Y2=0.705
r144 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r145 1 16 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%A_713_21# 1 2 9 13 17 20 22 25 29 32 34 37
+ 38 41 45 46 52
c77 38 0 1.01102e-19 $X=5.01 $Y=1.16
r78 41 43 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=0.58
+ $X2=4.405 $Y2=0.745
r79 38 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.01 $Y=1.16
+ $X2=5.01 $Y2=1.325
r80 38 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.01 $Y=1.16
+ $X2=5.01 $Y2=0.995
r81 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.16 $X2=5.01 $Y2=1.16
r82 35 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.515 $Y=1.16
+ $X2=4.43 $Y2=1.16
r83 35 37 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.515 $Y=1.16
+ $X2=5.01 $Y2=1.16
r84 34 45 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.43 $Y=1.535
+ $X2=4.405 $Y2=1.7
r85 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=1.325
+ $X2=4.43 $Y2=1.16
r86 33 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.43 $Y=1.325
+ $X2=4.43 $Y2=1.535
r87 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=1.16
r88 32 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=0.745
r89 27 45 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=1.865
+ $X2=4.405 $Y2=1.7
r90 27 29 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.405 $Y=1.865
+ $X2=4.405 $Y2=2.27
r91 25 47 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.64 $Y2=1.7
r92 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r93 22 45 0.463323 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.295 $Y=1.7
+ $X2=4.405 $Y2=1.7
r94 22 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.295 $Y=1.7
+ $X2=3.925 $Y2=1.7
r95 20 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.025 $Y=1.985
+ $X2=5.025 $Y2=1.325
r96 17 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.025 $Y=0.56
+ $X2=5.025 $Y2=0.995
r97 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.865
+ $X2=3.64 $Y2=1.7
r98 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.64 $Y=1.865
+ $X2=3.64 $Y2=2.275
r99 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.535
+ $X2=3.64 $Y2=1.7
r100 7 9 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=3.64 $Y=1.535
+ $X2=3.64 $Y2=0.415
r101 2 45 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.485 $X2=4.38 $Y2=1.755
r102 2 29 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.485 $X2=4.38 $Y2=2.27
r103 1 41 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.255
+ $Y=0.235 $X2=4.38 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%A_560_47# 1 2 7 9 12 14 15 16 20 25 27 30 33
c83 33 0 1.54137e-19 $X=3.33 $Y=0.995
c84 30 0 1.01102e-19 $X=4.09 $Y=1.16
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.16 $X2=4.09 $Y2=1.16
r86 28 33 0.89609 $w=3.3e-07 $l=3.47851e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=3.33 $Y2=0.995
r87 28 30 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=4.09 $Y2=1.16
r88 26 33 8.61065 $w=1.7e-07 $l=4.14246e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.33 $Y2=0.995
r89 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=2.255
r90 25 33 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=0.995
+ $X2=3.33 $Y2=0.995
r91 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=0.995
r92 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r93 20 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.005 $Y2=0.45
r94 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.435 $Y=2.34
+ $X2=3.52 $Y2=2.255
r95 16 18 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.435 $Y=2.34
+ $X2=2.935 $Y2=2.34
r96 14 31 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=4.515 $Y=1.16
+ $X2=4.09 $Y2=1.16
r97 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.515 $Y=1.16
+ $X2=4.59 $Y2=1.16
r98 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.16
r99 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.985
r100 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=1.16
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=0.56
r102 2 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=2.065 $X2=2.935 $Y2=2.34
r103 1 22 182 $w=1.7e-07 $l=3.005e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=3.005 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 42 58 59 62 65
r87 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r90 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r91 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r92 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r93 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r94 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r95 50 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r96 49 52 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r97 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 47 65 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r99 47 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r100 46 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r101 46 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r102 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r103 43 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r104 43 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r105 42 65 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r106 42 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 37 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r108 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r109 35 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r110 35 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r111 33 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.695 $Y=2.72
+ $X2=4.37 $Y2=2.72
r112 33 34 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.695 $Y=2.72
+ $X2=4.797 $Y2=2.72
r113 32 58 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.9 $Y=2.72
+ $X2=5.29 $Y2=2.72
r114 32 34 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=4.9 $Y=2.72
+ $X2=4.797 $Y2=2.72
r115 30 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.775 $Y=2.72
+ $X2=3.45 $Y2=2.72
r116 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=2.72
+ $X2=3.86 $Y2=2.72
r117 29 55 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.945 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=2.72
+ $X2=3.86 $Y2=2.72
r119 25 34 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.797 $Y=2.635
+ $X2=4.797 $Y2=2.72
r120 25 27 48.6918 $w=2.03e-07 $l=9e-07 $layer=LI1_cond $X=4.797 $Y=2.635
+ $X2=4.797 $Y2=1.735
r121 21 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=2.635
+ $X2=3.86 $Y2=2.72
r122 21 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.86 $Y=2.635
+ $X2=3.86 $Y2=2.3
r123 17 65 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r124 17 19 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r125 13 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r126 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r127 4 27 300 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=1.485 $X2=4.815 $Y2=1.735
r128 3 23 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=2.065 $X2=3.86 $Y2=2.3
r129 2 19 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r130 1 15 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%Q 1 2 9 10 11 19 30
r15 28 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.35 $Y=0.745
+ $X2=5.35 $Y2=1.67
r16 16 19 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=5.292 $Y=1.812
+ $X2=5.292 $Y2=1.835
r17 10 16 0.566112 $w=2.83e-07 $l=1.4e-08 $layer=LI1_cond $X=5.292 $Y=1.798
+ $X2=5.292 $Y2=1.812
r18 10 30 7.03738 $w=2.83e-07 $l=1.28e-07 $layer=LI1_cond $X=5.292 $Y=1.798
+ $X2=5.292 $Y2=1.67
r19 10 11 13.2228 $w=2.83e-07 $l=3.27e-07 $layer=LI1_cond $X=5.292 $Y=1.883
+ $X2=5.292 $Y2=2.21
r20 10 19 1.94096 $w=2.83e-07 $l=4.8e-08 $layer=LI1_cond $X=5.292 $Y=1.883
+ $X2=5.292 $Y2=1.835
r21 9 28 11.3641 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=5.292 $Y=0.51
+ $X2=5.292 $Y2=0.745
r22 2 19 300 $w=1.7e-07 $l=4.22493e-07 $layer=licon1_PDIFF $count=2 $X=5.1
+ $Y=1.485 $X2=5.26 $Y2=1.835
r23 1 9 182 $w=1.7e-07 $l=4.17403e-07 $layer=licon1_NDIFF $count=1 $X=5.1
+ $Y=0.235 $X2=5.26 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTP_1%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 44
+ 57 58 61 64 67
c88 58 0 2.71124e-20 $X=5.29 $Y=0
c89 2 0 7.13094e-20 $X=1.905 $Y=0.235
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r91 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r93 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r94 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r95 55 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r96 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r97 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.85
+ $Y2=0
r98 52 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.37
+ $Y2=0
r99 51 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r100 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r101 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r102 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r103 47 50 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r104 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r105 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r106 45 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r107 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.85
+ $Y2=0
r108 44 50 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.685 $Y=0
+ $X2=3.45 $Y2=0
r109 43 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r110 43 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r111 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r112 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r113 40 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r114 39 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r115 39 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r116 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r117 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r118 32 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 30 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=4.37 $Y2=0
r121 30 31 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.695 $Y=0
+ $X2=4.797 $Y2=0
r122 29 57 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.9 $Y=0 $X2=5.29
+ $Y2=0
r123 29 31 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=4.9 $Y=0 $X2=4.797
+ $Y2=0
r124 25 31 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.797 $Y=0.085
+ $X2=4.797 $Y2=0
r125 25 27 25.1574 $w=2.03e-07 $l=4.65e-07 $layer=LI1_cond $X=4.797 $Y=0.085
+ $X2=4.797 $Y2=0.55
r126 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0
r127 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0.445
r128 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r129 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r130 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r131 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r132 4 27 182 $w=1.7e-07 $l=3.82721e-07 $layer=licon1_NDIFF $count=1 $X=4.665
+ $Y=0.235 $X2=4.815 $Y2=0.55
r133 3 23 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.715
+ $Y=0.235 $X2=3.85 $Y2=0.445
r134 2 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r135 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


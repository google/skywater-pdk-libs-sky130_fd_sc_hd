* File: sky130_fd_sc_hd__inv_8.pex.spice
* Created: Tue Sep  1 19:10:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_8%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 57 58 59 60 61 62 83
r160 81 83 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.365 $Y=1.16
+ $X2=3.575 $Y2=1.16
r161 79 81 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.155 $Y=1.16
+ $X2=3.365 $Y2=1.16
r162 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=3.155 $Y2=1.16
r163 77 78 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.315 $Y=1.16
+ $X2=2.735 $Y2=1.16
r164 76 77 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.895 $Y=1.16
+ $X2=2.315 $Y2=1.16
r165 75 76 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.475 $Y=1.16
+ $X2=1.895 $Y2=1.16
r166 74 75 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=1.475 $Y2=1.16
r167 72 74 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.845 $Y=1.16
+ $X2=1.055 $Y2=1.16
r168 72 73 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.845
+ $Y=1.16 $X2=0.845 $Y2=1.16
r169 69 72 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.635 $Y=1.16
+ $X2=0.845 $Y2=1.16
r170 62 81 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.365
+ $Y=1.16 $X2=3.365 $Y2=1.16
r171 61 62 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=2.99 $Y=1.2
+ $X2=3.365 $Y2=1.2
r172 60 61 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=1.2 $X2=2.99
+ $Y2=1.2
r173 59 60 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=1.2 $X2=2.53
+ $Y2=1.2
r174 58 59 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=2.07
+ $Y2=1.2
r175 57 58 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.61
+ $Y2=1.2
r176 57 73 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=1.15 $Y=1.2
+ $X2=0.845 $Y2=1.2
r177 53 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.325
+ $X2=3.575 $Y2=1.16
r178 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.575 $Y=1.325
+ $X2=3.575 $Y2=1.985
r179 50 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=1.16
r180 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=0.56
r181 46 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=1.325
+ $X2=3.155 $Y2=1.16
r182 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.155 $Y=1.325
+ $X2=3.155 $Y2=1.985
r183 43 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=0.995
+ $X2=3.155 $Y2=1.16
r184 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.155 $Y=0.995
+ $X2=3.155 $Y2=0.56
r185 39 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.325
+ $X2=2.735 $Y2=1.16
r186 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.735 $Y=1.325
+ $X2=2.735 $Y2=1.985
r187 36 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=1.16
r188 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=0.56
r189 32 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.16
r190 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.985
r191 29 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=1.16
r192 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=0.56
r193 25 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.325
+ $X2=1.895 $Y2=1.16
r194 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.895 $Y=1.325
+ $X2=1.895 $Y2=1.985
r195 22 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=1.16
r196 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=0.56
r197 18 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.325
+ $X2=1.475 $Y2=1.16
r198 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.475 $Y=1.325
+ $X2=1.475 $Y2=1.985
r199 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=1.16
r200 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.56
r201 11 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.325
+ $X2=1.055 $Y2=1.16
r202 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.055 $Y=1.325
+ $X2=1.055 $Y2=1.985
r203 8 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=1.16
r204 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r205 4 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=1.325
+ $X2=0.635 $Y2=1.16
r206 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.635 $Y=1.325
+ $X2=0.635 $Y2=1.985
r207 1 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=1.16
r208 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_8%VPWR 1 2 3 4 5 16 18 22 24 28 32 34 36 38 39
+ 41 42 43 53 61 65
c64 5 0 1.47581e-19 $X=3.65 $Y=1.485
c65 1 0 1.50838e-19 $X=0.3 $Y=1.485
r66 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 56 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 53 64 4.41037 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.92
+ $Y2=2.72
r71 53 55 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.45
+ $Y2=2.72
r72 52 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 52 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 49 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.72
+ $X2=2.105 $Y2=2.72
r76 49 51 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 48 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r78 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 45 58 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=0.255 $Y2=2.72
r80 45 47 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=2.72 $X2=1.15
+ $Y2=2.72
r81 43 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r82 43 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r83 41 51 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.86 $Y=2.72
+ $X2=2.53 $Y2=2.72
r84 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=2.72
+ $X2=2.945 $Y2=2.72
r85 40 55 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.03 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 40 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.72
+ $X2=2.945 $Y2=2.72
r87 38 47 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=2.72 $X2=1.15
+ $Y2=2.72
r88 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.72
+ $X2=1.265 $Y2=2.72
r89 34 64 3.1073 $w=3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.92 $Y2=2.72
r90 34 36 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2
r91 30 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2.72
r92 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2
r93 26 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2.72
r94 26 28 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2
r95 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=2.72
+ $X2=1.265 $Y2=2.72
r96 24 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=2.72
+ $X2=2.105 $Y2=2.72
r97 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.02 $Y=2.72
+ $X2=1.35 $Y2=2.72
r98 20 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2.72
r99 20 22 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.265 $Y=2.635
+ $X2=1.265 $Y2=2
r100 16 58 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.255 $Y2=2.72
r101 16 18 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.382 $Y2=2
r102 5 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.65
+ $Y=1.485 $X2=3.785 $Y2=2
r103 4 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.485 $X2=2.945 $Y2=2
r104 3 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=1.485 $X2=2.105 $Y2=2
r105 2 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.485 $X2=1.265 $Y2=2
r106 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=1.485 $X2=0.425 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__INV_8%Y 1 2 3 4 5 6 7 8 25 26 27 28 31 35 37 39 43
+ 47 49 51 55 59 61 63 67 71 73 75 79 81 82 84 85 87 88 90 93 94
c174 94 0 1.47581e-19 $X=3.91 $Y=1.19
c175 93 0 1.50838e-19 $X=0.23 $Y=1.19
r176 92 94 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=3.895 $Y=1.495
+ $X2=3.895 $Y2=1.19
r177 91 94 10.2639 $w=3.18e-07 $l=2.85e-07 $layer=LI1_cond $X=3.895 $Y=0.905
+ $X2=3.895 $Y2=1.19
r178 78 93 10.1883 $w=3.43e-07 $l=3.05e-07 $layer=LI1_cond $X=0.257 $Y=1.495
+ $X2=0.257 $Y2=1.19
r179 77 93 9.52018 $w=3.43e-07 $l=2.85e-07 $layer=LI1_cond $X=0.257 $Y=0.905
+ $X2=0.257 $Y2=1.19
r180 76 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=1.58
+ $X2=3.365 $Y2=1.58
r181 75 92 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=3.735 $Y=1.58
+ $X2=3.895 $Y2=1.495
r182 75 76 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.735 $Y=1.58
+ $X2=3.53 $Y2=1.58
r183 74 88 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=0.81
+ $X2=3.365 $Y2=0.81
r184 73 91 7.40893 $w=1.9e-07 $l=2.0199e-07 $layer=LI1_cond $X=3.735 $Y=0.81
+ $X2=3.895 $Y2=0.905
r185 73 74 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=3.735 $Y=0.81
+ $X2=3.53 $Y2=0.81
r186 69 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=1.665
+ $X2=3.365 $Y2=1.58
r187 69 71 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.365 $Y=1.665
+ $X2=3.365 $Y2=2.34
r188 65 88 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.365 $Y=0.715
+ $X2=3.365 $Y2=0.81
r189 65 67 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.365 $Y=0.715
+ $X2=3.365 $Y2=0.38
r190 64 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.58
+ $X2=2.525 $Y2=1.58
r191 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=1.58
+ $X2=3.365 $Y2=1.58
r192 63 64 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.2 $Y=1.58
+ $X2=2.69 $Y2=1.58
r193 62 85 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.81
+ $X2=2.525 $Y2=0.81
r194 61 88 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=0.81
+ $X2=3.365 $Y2=0.81
r195 61 62 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=3.2 $Y=0.81
+ $X2=2.69 $Y2=0.81
r196 57 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.665
+ $X2=2.525 $Y2=1.58
r197 57 59 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.525 $Y=1.665
+ $X2=2.525 $Y2=2.34
r198 53 85 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.525 $Y=0.715
+ $X2=2.525 $Y2=0.81
r199 53 55 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.525 $Y=0.715
+ $X2=2.525 $Y2=0.38
r200 52 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=1.58
+ $X2=1.685 $Y2=1.58
r201 51 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=1.58
+ $X2=2.525 $Y2=1.58
r202 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.36 $Y=1.58
+ $X2=1.85 $Y2=1.58
r203 50 82 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0.81
+ $X2=1.685 $Y2=0.81
r204 49 85 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0.81
+ $X2=2.525 $Y2=0.81
r205 49 50 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=2.36 $Y=0.81
+ $X2=1.85 $Y2=0.81
r206 45 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.58
r207 45 47 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.34
r208 41 82 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=1.685 $Y=0.715
+ $X2=1.685 $Y2=0.81
r209 41 43 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.685 $Y=0.715
+ $X2=1.685 $Y2=0.38
r210 40 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.58
+ $X2=0.845 $Y2=1.58
r211 39 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=1.685 $Y2=1.58
r212 39 40 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=1.01 $Y2=1.58
r213 38 79 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0.81
+ $X2=0.845 $Y2=0.81
r214 37 82 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0.81
+ $X2=1.685 $Y2=0.81
r215 37 38 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=1.52 $Y=0.81
+ $X2=1.01 $Y2=0.81
r216 33 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=1.665
+ $X2=0.845 $Y2=1.58
r217 33 35 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.845 $Y=1.665
+ $X2=0.845 $Y2=2.34
r218 29 79 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=0.845 $Y=0.715
+ $X2=0.845 $Y2=0.81
r219 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.845 $Y=0.715
+ $X2=0.845 $Y2=0.38
r220 28 78 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.43 $Y=1.58
+ $X2=0.257 $Y2=1.495
r221 27 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.58
+ $X2=0.845 $Y2=1.58
r222 27 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.68 $Y=1.58
+ $X2=0.43 $Y2=1.58
r223 26 77 7.58838 $w=1.9e-07 $l=2.15323e-07 $layer=LI1_cond $X=0.43 $Y=0.81
+ $X2=0.257 $Y2=0.905
r224 25 79 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.81
+ $X2=0.845 $Y2=0.81
r225 25 26 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=0.68 $Y=0.81
+ $X2=0.43 $Y2=0.81
r226 8 90 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.485 $X2=3.365 $Y2=1.66
r227 8 71 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.485 $X2=3.365 $Y2=2.34
r228 7 87 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.525 $Y2=1.66
r229 7 59 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.525 $Y2=2.34
r230 6 84 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.685 $Y2=1.66
r231 6 47 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.685 $Y2=2.34
r232 5 81 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.485 $X2=0.845 $Y2=1.66
r233 5 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.485 $X2=0.845 $Y2=2.34
r234 4 67 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.23
+ $Y=0.235 $X2=3.365 $Y2=0.38
r235 3 55 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.39
+ $Y=0.235 $X2=2.525 $Y2=0.38
r236 2 43 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.235 $X2=1.685 $Y2=0.38
r237 1 31 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.71
+ $Y=0.235 $X2=0.845 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__INV_8%VGND 1 2 3 4 5 16 18 22 24 28 32 34 36 38 39
+ 41 42 43 53 61 65
r79 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r80 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r81 56 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r82 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r83 53 64 4.45794 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.92
+ $Y2=0
r84 53 55 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.45
+ $Y2=0
r85 52 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r86 52 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r87 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r88 49 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.105
+ $Y2=0
r89 49 51 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.53
+ $Y2=0
r90 48 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r91 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r92 45 58 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r93 45 47 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=1.15
+ $Y2=0
r94 43 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r95 43 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r96 41 51 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.53
+ $Y2=0
r97 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.945
+ $Y2=0
r98 40 55 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.45
+ $Y2=0
r99 40 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.945
+ $Y2=0
r100 38 47 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.15
+ $Y2=0
r101 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.265
+ $Y2=0
r102 34 64 3.1003 $w=3.05e-07 $l=1.14039e-07 $layer=LI1_cond $X=3.852 $Y=0.085
+ $X2=3.92 $Y2=0
r103 34 36 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=3.852 $Y=0.085
+ $X2=3.852 $Y2=0.38
r104 30 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0
r105 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.38
r106 26 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r107 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.38
r108 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.265
+ $Y2=0
r109 24 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0 $X2=2.105
+ $Y2=0
r110 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=1.35
+ $Y2=0
r111 20 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=0.085
+ $X2=1.265 $Y2=0
r112 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.265 $Y=0.085
+ $X2=1.265 $Y2=0.38
r113 16 58 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.255 $Y2=0
r114 16 18 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.382 $Y2=0.38
r115 5 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.785 $Y2=0.38
r116 4 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.945 $Y2=0.38
r117 3 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.105 $Y2=0.38
r118 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.265 $Y2=0.38
r119 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.38
.ends


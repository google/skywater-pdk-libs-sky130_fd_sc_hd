* File: sky130_fd_sc_hd__a2bb2o_1.spice
* Created: Thu Aug 27 14:03:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2bb2o_1.spice.pex"
.subckt sky130_fd_sc_hd__a2bb2o_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_76_199#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.145916 AS=0.169 PD=1.31822 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1009 N_A_226_47#_M1009_d N_A1_N_M1009_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0942841 PD=0.69 PS=0.851776 NRD=0 NRS=45.708 M=1 R=2.8
+ SA=75000.8 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A2_N_M1007_g N_A_226_47#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1386 AS=0.0567 PD=1.08 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_76_199#_M1001_d N_A_226_47#_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1386 PD=0.69 PS=1.08 NRD=0 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_556_47# N_B2_M1004_g N_A_76_199#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=22.848 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g A_556_47# VNB NSHORT L=0.15 W=0.42 AD=0.1092
+ AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_76_199#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.234859 AS=0.26 PD=2.02113 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 A_226_297# N_A1_N_M1010_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0986408 PD=0.63 PS=0.848873 NRD=23.443 NRS=84.3554 M=1 R=2.8
+ SA=75000.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_226_47#_M1000_d N_A2_N_M1000_g A_226_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_489_413#_M1002_d N_A_226_47#_M1002_g N_A_76_199#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_B2_M1008_g N_A_489_413#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_489_413#_M1006_d N_B1_M1006_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_79 VPB 0 1.32536e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__a2bb2o_1.spice.SKY130_FD_SC_HD__A2BB2O_1.pxi"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__or4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755000 1.075000 2.320000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 2.125000 2.670000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.550000 1.075000 3.550000 1.275000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.435000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.675000 1.250000 0.680000 ;
        RECT 0.935000 0.680000 1.245000 0.790000 ;
        RECT 0.935000 0.790000 1.105000 1.495000 ;
        RECT 0.935000 1.495000 1.250000 1.825000 ;
        RECT 0.970000 0.260000 1.250000 0.675000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.630000  0.085000 0.800000 0.565000 ;
        RECT 1.435000  0.085000 1.815000 0.485000 ;
        RECT 2.385000  0.085000 2.715000 0.485000 ;
        RECT 3.225000  0.085000 3.555000 0.585000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.515000 2.335000 0.845000 2.635000 ;
        RECT 1.480000 2.335000 1.815000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.325000 0.350000 0.735000 ;
      RECT 0.085000 0.735000 0.765000 0.905000 ;
      RECT 0.085000 1.605000 0.765000 1.890000 ;
      RECT 0.510000 1.890000 0.765000 1.995000 ;
      RECT 0.510000 1.995000 1.715000 2.165000 ;
      RECT 0.595000 0.905000 0.765000 1.605000 ;
      RECT 1.290000 0.995000 1.585000 1.325000 ;
      RECT 1.415000 0.735000 3.055000 0.905000 ;
      RECT 1.415000 0.905000 1.585000 0.995000 ;
      RECT 1.415000 1.325000 1.585000 1.355000 ;
      RECT 1.415000 1.355000 1.600000 1.370000 ;
      RECT 1.415000 1.370000 1.610000 1.380000 ;
      RECT 1.415000 1.380000 1.620000 1.390000 ;
      RECT 1.415000 1.390000 1.625000 1.400000 ;
      RECT 1.415000 1.400000 1.630000 1.410000 ;
      RECT 1.415000 1.410000 1.645000 1.420000 ;
      RECT 1.415000 1.420000 1.655000 1.425000 ;
      RECT 1.415000 1.425000 1.665000 1.445000 ;
      RECT 1.415000 1.445000 3.560000 1.450000 ;
      RECT 1.420000 1.450000 3.560000 1.615000 ;
      RECT 1.440000 1.785000 3.030000 1.955000 ;
      RECT 1.440000 1.955000 1.715000 1.995000 ;
      RECT 1.985000 0.305000 2.155000 0.735000 ;
      RECT 2.860000 1.955000 3.030000 2.215000 ;
      RECT 2.860000 2.215000 3.345000 2.385000 ;
      RECT 2.885000 0.305000 3.055000 0.735000 ;
      RECT 3.225000 1.615000 3.560000 1.815000 ;
  END
END sky130_fd_sc_hd__or4b_2
END LIBRARY

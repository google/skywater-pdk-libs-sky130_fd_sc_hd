* File: sky130_fd_sc_hd__xor3_1.pex.spice
* Created: Thu Aug 27 14:50:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_112_21# 1 2 7 9 12 14 15 16 18 19 21 23 25
+ 26 28 33 35 36
r102 38 40 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.635 $Y=1.16
+ $X2=0.655 $Y2=1.16
r103 35 36 10.5404 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=2.575 $Y=0.355
+ $X2=2.39 $Y2=0.355
r104 33 40 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.835 $Y=1.16
+ $X2=0.655 $Y2=1.16
r105 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.835
+ $Y=1.16 $X2=0.835 $Y2=1.16
r106 30 32 25.0595 $w=1.85e-07 $l=3.8e-07 $layer=LI1_cond $X=0.85 $Y=0.78
+ $X2=0.85 $Y2=1.16
r107 26 28 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.47 $Y=2.32
+ $X2=2.58 $Y2=2.32
r108 25 36 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.35 $Y=0.34
+ $X2=2.39 $Y2=0.34
r109 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.385 $Y=2.235
+ $X2=1.47 $Y2=2.32
r110 22 23 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=2.045
+ $X2=1.385 $Y2=2.235
r111 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.265 $Y=0.425
+ $X2=1.35 $Y2=0.34
r112 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.265 $Y=0.425
+ $X2=1.265 $Y2=0.695
r113 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.3 $Y=1.96
+ $X2=1.385 $Y2=2.045
r114 18 19 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.3 $Y=1.96
+ $X2=0.95 $Y2=1.96
r115 17 30 1.22693 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.95 $Y=0.78 $X2=0.85
+ $Y2=0.78
r116 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=0.78
+ $X2=1.265 $Y2=0.695
r117 16 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.18 $Y=0.78
+ $X2=0.95 $Y2=0.78
r118 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.865 $Y=1.875
+ $X2=0.95 $Y2=1.96
r119 14 32 10.9829 $w=1.85e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.865 $Y=1.325
+ $X2=0.85 $Y2=1.16
r120 14 15 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.865 $Y=1.325
+ $X2=0.865 $Y2=1.875
r121 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.325
+ $X2=0.655 $Y2=1.16
r122 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.655 $Y=1.325
+ $X2=0.655 $Y2=1.985
r123 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=1.16
r124 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=0.56
r125 2 28 600 $w=1.7e-07 $l=7.79824e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.625 $X2=2.58 $Y2=2.32
r126 1 35 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.245 $X2=2.575 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%C 1 3 4 6 7 11 13 15 16 17 20 21
c68 4 0 8.31677e-20 $X=1.255 $Y=1.325
r69 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.31
+ $Y=1.16 $X2=2.31 $Y2=1.16
r70 17 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.07 $Y=1.16 $X2=2.31
+ $Y2=1.16
r71 13 20 37.0704 $w=1.5e-07 $l=1.19896e-07 $layer=POLY_cond $X=2.365 $Y=0.985
+ $X2=2.25 $Y2=0.995
r72 13 15 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.365 $Y=0.985
+ $X2=2.365 $Y2=0.565
r73 9 20 37.0704 $w=1.5e-07 $l=3.95727e-07 $layer=POLY_cond $X=2.325 $Y=1.355
+ $X2=2.25 $Y2=0.995
r74 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.325 $Y=1.355
+ $X2=2.325 $Y2=2.045
r75 8 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.255 $Y2=1.16
r76 7 20 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.25 $Y2=0.995
r77 7 8 160.872 $w=3.3e-07 $l=9.2e-07 $layer=POLY_cond $X=2.25 $Y=1.16 $X2=1.33
+ $Y2=1.16
r78 4 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.255 $Y=1.325
+ $X2=1.255 $Y2=1.16
r79 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.255 $Y=1.325
+ $X2=1.255 $Y2=1.805
r80 1 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.255 $Y=0.995
+ $X2=1.255 $Y2=1.16
r81 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.255 $Y=0.995
+ $X2=1.255 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_266_93# 1 2 9 13 14 19 21 24 25 29 30 33
r78 30 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.16
+ $X2=2.855 $Y2=0.995
r79 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.855
+ $Y=1.16 $X2=2.855 $Y2=1.16
r80 26 29 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.75 $Y=1.16
+ $X2=2.855 $Y2=1.16
r81 23 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=1.325
+ $X2=2.75 $Y2=1.16
r82 23 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.75 $Y=1.325
+ $X2=2.75 $Y2=1.535
r83 22 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=1.62
+ $X2=1.605 $Y2=1.62
r84 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.665 $Y=1.62
+ $X2=2.75 $Y2=1.535
r85 21 22 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=2.665 $Y=1.62
+ $X2=1.69 $Y2=1.62
r86 17 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.535
+ $X2=1.605 $Y2=1.62
r87 17 19 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.605 $Y=1.535
+ $X2=1.605 $Y2=0.76
r88 14 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.62
+ $X2=1.605 $Y2=1.62
r89 14 16 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=1.52 $Y=1.62
+ $X2=1.465 $Y2=1.62
r90 13 33 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.915 $Y=0.565
+ $X2=2.915 $Y2=0.995
r91 7 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.325
+ $X2=2.855 $Y2=1.16
r92 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.855 $Y=1.325
+ $X2=2.855 $Y2=2.045
r93 2 16 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.33
+ $Y=1.485 $X2=1.465 $Y2=1.62
r94 1 19 182 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_NDIFF $count=1 $X=1.33
+ $Y=0.465 $X2=1.605 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_827_297# 1 2 9 13 15 17 19 21 22 23 27 35
+ 37 38 39 40 47 49 50 58
c169 49 0 1.83334e-19 $X=7.13 $Y=0.85
c170 15 0 1.24749e-19 $X=7.305 $Y=1.28
r171 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.11 $X2=7.25 $Y2=1.11
r172 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.18 $Y=0.85
+ $X2=7.18 $Y2=1.11
r173 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.85
+ $X2=7.13 $Y2=0.85
r174 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0.85
+ $X2=5.75 $Y2=0.85
r175 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0.85
+ $X2=4.37 $Y2=0.85
r176 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.895 $Y=0.85
+ $X2=5.75 $Y2=0.85
r177 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=7.13 $Y2=0.85
r178 39 40 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=5.895 $Y2=0.85
r179 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=0.85
+ $X2=4.37 $Y2=0.85
r180 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.605 $Y=0.85
+ $X2=5.75 $Y2=0.85
r181 37 38 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=5.605 $Y=0.85
+ $X2=4.515 $Y2=0.85
r182 35 47 7.77229 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=5.727 $Y=0.995
+ $X2=5.727 $Y2=0.85
r183 31 35 6.36987 $w=2.73e-07 $l=1.52e-07 $layer=LI1_cond $X=5.575 $Y=1.132
+ $X2=5.727 $Y2=1.132
r184 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.575
+ $Y=1.16 $X2=5.575 $Y2=1.16
r185 28 58 34.8134 $w=2.38e-07 $l=7.25e-07 $layer=LI1_cond $X=4.4 $Y=1.445
+ $X2=4.4 $Y2=0.72
r186 27 28 1.42499 $w=2.4e-07 $l=1.35e-07 $layer=LI1_cond $X=4.4 $Y=1.58 $X2=4.4
+ $Y2=1.445
r187 25 27 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.27 $Y=1.58 $X2=4.4
+ $Y2=1.58
r188 22 32 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=5.84 $Y=1.16
+ $X2=5.575 $Y2=1.16
r189 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.84 $Y=1.16
+ $X2=5.915 $Y2=1.16
r190 19 55 38.945 $w=2.68e-07 $l=1.92678e-07 $layer=POLY_cond $X=7.31 $Y=0.945
+ $X2=7.25 $Y2=1.11
r191 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.31 $Y=0.945
+ $X2=7.31 $Y2=0.535
r192 15 55 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=7.305 $Y=1.28
+ $X2=7.25 $Y2=1.11
r193 15 17 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=7.305 $Y=1.28
+ $X2=7.305 $Y2=2.065
r194 11 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.325
+ $X2=5.915 $Y2=1.16
r195 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.915 $Y=1.325
+ $X2=5.915 $Y2=1.805
r196 7 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=0.995
+ $X2=5.915 $Y2=1.16
r197 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.915 $Y=0.995
+ $X2=5.915 $Y2=0.455
r198 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.27 $Y2=1.63
r199 1 58 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.235 $X2=4.435 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%B 3 7 9 10 13 18 19 20 23 27 31 34 35 37 38
+ 41
r122 37 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=1.53
+ $X2=7.13 $Y2=1.53
r123 35 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.16
+ $X2=6.77 $Y2=1.325
r124 35 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.16
+ $X2=6.77 $Y2=0.995
r125 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.16 $X2=6.77 $Y2=1.16
r126 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.77 $Y=1.445
+ $X2=6.855 $Y2=1.53
r127 32 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.77 $Y=1.445
+ $X2=6.77 $Y2=1.16
r128 28 30 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.16
+ $X2=4.225 $Y2=1.16
r129 27 42 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.79 $Y=1.965
+ $X2=6.79 $Y2=1.325
r130 25 27 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.79 $Y=2.465
+ $X2=6.79 $Y2=1.965
r131 23 41 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.71 $Y=0.565
+ $X2=6.71 $Y2=0.995
r132 19 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.715 $Y=2.54
+ $X2=6.79 $Y2=2.465
r133 19 20 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=6.715 $Y=2.54
+ $X2=5.23 $Y2=2.54
r134 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.155 $Y=2.465
+ $X2=5.23 $Y2=2.54
r135 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.155 $Y=2.465
+ $X2=5.155 $Y2=1.905
r136 15 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.155 $Y=1.235
+ $X2=5.155 $Y2=1.16
r137 15 18 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.155 $Y=1.235
+ $X2=5.155 $Y2=1.905
r138 11 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.155 $Y=1.085
+ $X2=5.155 $Y2=1.16
r139 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.155 $Y=1.085
+ $X2=5.155 $Y2=0.565
r140 10 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.3 $Y=1.16
+ $X2=4.225 $Y2=1.16
r141 9 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.08 $Y=1.16
+ $X2=5.155 $Y2=1.16
r142 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.08 $Y=1.16 $X2=4.3
+ $Y2=1.16
r143 5 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.225 $Y=1.085
+ $X2=4.225 $Y2=1.16
r144 5 7 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.225 $Y=1.085
+ $X2=4.225 $Y2=0.56
r145 1 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.06 $Y=1.235
+ $X2=4.06 $Y2=1.16
r146 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.06 $Y=1.235
+ $X2=4.06 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A 3 6 8 11 12 13
c44 13 0 1.83334e-19 $X=7.74 $Y=0.995
r45 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.74 $Y=1.16
+ $X2=7.74 $Y2=1.325
r46 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.74 $Y=1.16
+ $X2=7.74 $Y2=0.995
r47 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.73
+ $Y=1.16 $X2=7.73 $Y2=1.16
r48 8 12 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=7.59 $Y=1.2 $X2=7.73
+ $Y2=1.2
r49 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.81 $Y=1.985
+ $X2=7.81 $Y2=1.325
r50 3 13 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.81 $Y=0.555
+ $X2=7.81 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_931_365# 1 2 3 4 13 15 18 22 24 28 29 30 31
+ 36 37 38 41 44 45
c135 36 0 1.4656e-19 $X=8.23 $Y=1.16
c136 31 0 1.06604e-19 $X=8.17 $Y=1.495
c137 30 0 1.40536e-19 $X=8.17 $Y=1.325
r138 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0.51
+ $X2=7.59 $Y2=0.51
r139 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0.51
+ $X2=4.83 $Y2=0.51
r140 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=0.51
+ $X2=4.83 $Y2=0.51
r141 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=0.51
+ $X2=7.59 $Y2=0.51
r142 37 38 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=7.445 $Y=0.51
+ $X2=4.975 $Y2=0.51
r143 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=1.16 $X2=8.23 $Y2=1.16
r144 33 35 20.4335 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=8.2 $Y=0.82 $X2=8.2
+ $Y2=1.16
r145 32 45 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=7.62 $Y=0.735
+ $X2=7.62 $Y2=0.51
r146 30 35 10.2745 $w=2.03e-07 $l=1.79374e-07 $layer=LI1_cond $X=8.17 $Y=1.325
+ $X2=8.2 $Y2=1.16
r147 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.17 $Y=1.325
+ $X2=8.17 $Y2=1.495
r148 29 32 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.765 $Y=0.82
+ $X2=7.62 $Y2=0.735
r149 28 33 1.77774 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.085 $Y=0.82
+ $X2=8.2 $Y2=0.82
r150 28 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.085 $Y=0.82
+ $X2=7.765 $Y2=0.82
r151 24 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.085 $Y=1.6
+ $X2=8.17 $Y2=1.495
r152 24 26 25.6147 $w=2.08e-07 $l=4.85e-07 $layer=LI1_cond $X=8.085 $Y=1.6
+ $X2=7.6 $Y2=1.6
r153 20 41 3.61456 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=0.595
+ $X2=4.78 $Y2=0.43
r154 20 22 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.78 $Y=0.595
+ $X2=4.78 $Y2=1.94
r155 16 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.16
r156 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.985
r157 13 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=1.16
r158 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=0.555
r159 4 26 600 $w=1.7e-07 $l=2.32164e-07 $layer=licon1_PDIFF $count=1 $X=7.38
+ $Y=1.645 $X2=7.6 $Y2=1.62
r160 3 22 600 $w=1.7e-07 $l=1.73205e-07 $layer=licon1_PDIFF $count=1 $X=4.655
+ $Y=1.825 $X2=4.78 $Y2=1.94
r161 2 45 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=7.385
+ $Y=0.235 $X2=7.6 $Y2=0.625
r162 1 41 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.245 $X2=4.945 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%X 1 2 10 15 16 17
c24 15 0 8.31677e-20 $X=0.445 $Y=1.62
r25 17 22 9.79645 $w=5.23e-07 $l=4.3e-07 $layer=LI1_cond $X=0.347 $Y=1.87
+ $X2=0.347 $Y2=2.3
r26 15 16 5.99972 $w=5.23e-07 $l=1.8e-07 $layer=LI1_cond $X=0.347 $Y=1.62
+ $X2=0.347 $Y2=1.44
r27 13 17 3.82745 $w=5.23e-07 $l=1.68e-07 $layer=LI1_cond $X=0.347 $Y=1.702
+ $X2=0.347 $Y2=1.87
r28 13 15 1.86816 $w=5.23e-07 $l=8.2e-08 $layer=LI1_cond $X=0.347 $Y=1.702
+ $X2=0.347 $Y2=1.62
r29 12 16 18.8415 $w=3.13e-07 $l=5.15e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.44
r30 10 12 10.3285 $w=5.03e-07 $l=3.65e-07 $layer=LI1_cond $X=0.337 $Y=0.56
+ $X2=0.337 $Y2=0.925
r31 2 22 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.445 $Y2=2.3
r32 2 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.445 $Y2=1.62
r33 1 10 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%VPWR 1 2 3 12 16 20 23 24 25 31 38 48 49 52
+ 55
c95 3 0 1.06604e-19 $X=7.885 $Y=1.485
r96 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r97 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 49 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r99 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r100 46 55 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.19 $Y=2.72
+ $X2=8.022 $Y2=2.72
r101 46 48 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.19 $Y=2.72
+ $X2=8.51 $Y2=2.72
r102 45 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r103 44 45 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r104 42 45 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=7.59 $Y2=2.72
r105 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 41 44 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=7.59 $Y2=2.72
r107 41 42 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 39 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.85 $Y2=2.72
r109 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.37 $Y2=2.72
r110 38 55 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.855 $Y=2.72
+ $X2=8.022 $Y2=2.72
r111 38 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.855 $Y=2.72
+ $X2=7.59 $Y2=2.72
r112 37 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r114 34 37 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r115 33 36 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r116 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 31 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.85 $Y2=2.72
r118 31 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 29 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 25 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 23 28 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.78 $Y=2.72 $X2=0.69
+ $Y2=2.72
r123 23 24 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.78 $Y=2.72
+ $X2=0.947 $Y2=2.72
r124 22 33 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 22 24 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.947 $Y2=2.72
r126 18 55 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.022 $Y=2.635
+ $X2=8.022 $Y2=2.72
r127 18 20 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=8.022 $Y=2.635
+ $X2=8.022 $Y2=2.36
r128 14 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.72
r129 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.32
r130 10 24 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.947 $Y=2.635
+ $X2=0.947 $Y2=2.72
r131 10 12 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.947 $Y=2.635
+ $X2=0.947 $Y2=2.3
r132 3 20 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.36
r133 2 16 600 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=3.725
+ $Y=1.485 $X2=3.85 $Y2=2.32
r134 1 12 600 $w=1.7e-07 $l=9.18436e-07 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.485 $X2=0.95 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_386_325# 1 2 3 4 13 18 21 23 25 27 30 32 34
+ 35 37 38 44 48
c141 34 0 1.24749e-19 $X=6.93 $Y=0.38
r142 47 48 11.956 $w=2.5e-07 $l=2.45e-07 $layer=LI1_cond $X=3.09 $Y=1.535
+ $X2=3.335 $Y2=1.535
r143 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.53
+ $X2=5.75 $Y2=1.53
r144 41 48 5.612 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=3.45 $Y=1.535
+ $X2=3.335 $Y2=1.535
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=1.53
+ $X2=3.45 $Y2=1.53
r146 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.595 $Y=1.53
+ $X2=3.45 $Y2=1.53
r147 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.605 $Y=1.53
+ $X2=5.75 $Y2=1.53
r148 37 38 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=5.605 $Y=1.53
+ $X2=3.595 $Y2=1.53
r149 34 35 13.3743 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=6.93 $Y=0.36
+ $X2=6.685 $Y2=0.36
r150 32 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.175 $Y=0.34
+ $X2=6.685 $Y2=0.34
r151 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.09 $Y=0.425
+ $X2=6.175 $Y2=0.34
r152 29 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.09 $Y=0.425
+ $X2=6.09 $Y2=1.445
r153 28 45 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=5.81 $Y=1.53
+ $X2=5.602 $Y2=1.53
r154 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.005 $Y=1.53
+ $X2=6.09 $Y2=1.445
r155 27 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.005 $Y=1.53
+ $X2=5.81 $Y2=1.53
r156 23 45 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.602 $Y=1.615
+ $X2=5.602 $Y2=1.53
r157 23 25 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=5.602 $Y=1.615
+ $X2=5.602 $Y2=1.62
r158 19 48 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.335 $Y=1.375
+ $X2=3.335 $Y2=1.535
r159 19 21 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.335 $Y=1.375
+ $X2=3.335 $Y2=0.76
r160 17 47 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.09 $Y=1.695
+ $X2=3.09 $Y2=1.535
r161 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.09 $Y=1.695
+ $X2=3.09 $Y2=1.895
r162 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.005 $Y=1.98
+ $X2=3.09 $Y2=1.895
r163 13 15 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.005 $Y=1.98
+ $X2=2.115 $Y2=1.98
r164 4 25 300 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=2 $X=5.23
+ $Y=1.485 $X2=5.57 $Y2=1.62
r165 3 15 600 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.625 $X2=2.115 $Y2=1.98
r166 2 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.245 $X2=6.93 $Y2=0.38
r167 1 21 182 $w=1.7e-07 $l=6.65507e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.245 $X2=3.335 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_404_49# 1 2 3 4 13 18 19 20 22 23 24 26 28
+ 29 32 33 34 36 39 43 48 52 54 55 57
r181 55 56 15.25 $w=1.96e-07 $l=2.45e-07 $layer=LI1_cond $X=5.12 $Y=0.772
+ $X2=5.365 $Y2=0.772
r182 50 52 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.675 $Y=1.12
+ $X2=3.79 $Y2=1.12
r183 46 48 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.315 $Y=2.32
+ $X2=3.43 $Y2=2.32
r184 41 56 1.57051 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=5.365 $Y=0.655
+ $X2=5.365 $Y2=0.772
r185 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.365 $Y=0.655
+ $X2=5.365 $Y2=0.545
r186 37 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=2.36
+ $X2=5.12 $Y2=2.36
r187 37 39 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=5.205 $Y=2.36
+ $X2=7.085 $Y2=2.36
r188 36 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.275
+ $X2=5.12 $Y2=2.36
r189 35 55 1.57051 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=5.12 $Y=0.89
+ $X2=5.12 $Y2=0.772
r190 35 36 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.12 $Y=0.89
+ $X2=5.12 $Y2=2.275
r191 33 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=2.36
+ $X2=5.12 $Y2=2.36
r192 33 34 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.035 $Y=2.36
+ $X2=4.52 $Y2=2.36
r193 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=2.275
+ $X2=4.52 $Y2=2.36
r194 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.435 $Y=2.065
+ $X2=4.435 $Y2=2.275
r195 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=1.98
+ $X2=3.79 $Y2=1.98
r196 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=1.98
+ $X2=4.435 $Y2=2.065
r197 29 30 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.35 $Y=1.98
+ $X2=3.875 $Y2=1.98
r198 28 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=1.895
+ $X2=3.79 $Y2=1.98
r199 27 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=1.205
+ $X2=3.79 $Y2=1.12
r200 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.79 $Y=1.205
+ $X2=3.79 $Y2=1.895
r201 26 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.035
+ $X2=3.675 $Y2=1.12
r202 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.675 $Y=0.425
+ $X2=3.675 $Y2=1.035
r203 23 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=1.98
+ $X2=3.79 $Y2=1.98
r204 23 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.705 $Y=1.98
+ $X2=3.515 $Y2=1.98
r205 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=2.235
+ $X2=3.43 $Y2=2.32
r206 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=2.065
+ $X2=3.515 $Y2=1.98
r207 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.43 $Y=2.065
+ $X2=3.43 $Y2=2.235
r208 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=0.34
+ $X2=3.675 $Y2=0.425
r209 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.59 $Y=0.34
+ $X2=3.08 $Y2=0.34
r210 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=0.425
+ $X2=3.08 $Y2=0.34
r211 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.995 $Y=0.425
+ $X2=2.995 $Y2=0.655
r212 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.91 $Y=0.74
+ $X2=2.995 $Y2=0.655
r213 13 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.91 $Y=0.74
+ $X2=2.155 $Y2=0.74
r214 4 39 600 $w=1.7e-07 $l=8.17634e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=1.645 $X2=7.085 $Y2=2.36
r215 3 46 600 $w=1.7e-07 $l=8.66372e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.625 $X2=3.315 $Y2=2.32
r216 2 43 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=5.23
+ $Y=0.245 $X2=5.365 $Y2=0.545
r217 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.245 $X2=2.155 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%A_1198_49# 1 2 3 4 15 18 23 26 29 31 36
c67 29 0 1.17772e-19 $X=8.17 $Y=1.99
r68 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.44 $Y=0.42
+ $X2=8.57 $Y2=0.42
r69 28 29 14.5869 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.445 $Y=1.99
+ $X2=8.17 $Y2=1.99
r70 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.57 $Y=1.875
+ $X2=8.57 $Y2=1.99
r71 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=0.585
+ $X2=8.57 $Y2=0.42
r72 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=8.57 $Y=0.585
+ $X2=8.57 $Y2=1.875
r73 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=8.507 $Y=1.99
+ $X2=8.57 $Y2=1.99
r74 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=8.507 $Y=1.99
+ $X2=8.445 $Y2=1.99
r75 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=8.507 $Y=2.105
+ $X2=8.507 $Y2=2.3
r76 20 29 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=6.58 $Y=2.02
+ $X2=8.17 $Y2=2.02
r77 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.515 $Y=2.02
+ $X2=6.58 $Y2=2.02
r78 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.43 $Y=1.935
+ $X2=6.515 $Y2=2.02
r79 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.43 $Y=1.935
+ $X2=6.43 $Y2=0.76
r80 4 28 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.445 $Y2=1.96
r81 4 23 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.445 $Y2=2.3
r82 3 20 600 $w=1.7e-07 $l=8.14709e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.485 $X2=6.58 $Y2=2.02
r83 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.42
r84 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.245 $X2=6.43 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_1%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 50
+ 51
c103 20 0 2.87884e-20 $X=8.02 $Y=0.4
c104 3 0 1.40536e-19 $X=7.885 $Y=0.235
r105 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r106 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r107 47 48 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r108 45 48 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=7.59 $Y2=0
r109 44 47 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=7.59
+ $Y2=0
r110 44 45 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r111 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r112 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r113 39 42 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=3.91 $Y2=0
r114 38 41 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.91
+ $Y2=0
r115 38 39 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r116 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r117 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r118 31 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 29 47 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.59
+ $Y2=0
r120 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=0 $X2=8.02
+ $Y2=0
r121 28 50 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=8.51 $Y2=0
r122 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.02
+ $Y2=0
r123 26 41 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.91
+ $Y2=0
r124 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=0 $X2=4.015
+ $Y2=0
r125 25 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.1 $Y=0 $X2=4.37
+ $Y2=0
r126 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=0 $X2=4.015
+ $Y2=0
r127 23 34 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.69
+ $Y2=0
r128 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.885
+ $Y2=0
r129 22 38 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.15
+ $Y2=0
r130 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.885
+ $Y2=0
r131 18 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0
r132 18 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0.4
r133 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0
r134 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.36
r135 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0.085
+ $X2=0.885 $Y2=0
r136 10 12 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.885 $Y=0.085
+ $X2=0.885 $Y2=0.36
r137 3 20 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.4
r138 2 16 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=3.85
+ $Y=0.235 $X2=4.015 $Y2=0.36
r139 1 12 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.71
+ $Y=0.235 $X2=0.925 $Y2=0.36
.ends


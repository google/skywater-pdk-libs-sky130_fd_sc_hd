* File: sky130_fd_sc_hd__mux2_8.spice
* Created: Thu Aug 27 14:27:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2_8.spice.pex"
.subckt sky130_fd_sc_hd__mux2_8  VNB VPB S A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_79_21#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75008.8 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_79_21#_M1013_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75008.4 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1013_d N_A_79_21#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75008 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_A_79_21#_M1017_g N_X_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75007.6 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1017_d N_A_79_21#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75007.1 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1026_d N_A_79_21#_M1026_g N_X_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75006.7 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1026_d N_A_79_21#_M1027_g N_X_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_A_79_21#_M1031_g N_X_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.106066 AS=0.08775 PD=0.982558 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1005 N_A_792_47#_M1005_d N_S_M1005_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0944 AS=0.104434 PD=0.935 PS=0.967442 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75003.6 SB=75005.5 A=0.096 P=1.58 MULT=1
MM1022 N_A_79_21#_M1022_d N_A1_M1022_g N_A_792_47#_M1005_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.0944 PD=0.91 PS=0.935 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75005 A=0.096 P=1.58 MULT=1
MM1032 N_A_79_21#_M1022_d N_A1_M1032_g N_A_792_47#_M1032_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.336 PD=0.91 PS=1.69 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.5
+ SB=75004.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_792_47#_M1032_s N_S_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.64
+ AD=0.336 AS=0.1072 PD=1.69 PS=0.975 NRD=145.308 NRS=11.244 M=1 R=4.26667
+ SA=75005.7 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_1302_47#_M1006_d N_A_1259_199#_M1006_g N_VGND_M1011_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1552 AS=0.1072 PD=1.125 PS=0.975 NRD=16.872 NRS=0 M=1
+ R=4.26667 SA=75006.1 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1015 N_A_1302_47#_M1006_d N_A0_M1015_g N_A_79_21#_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1552 AS=0.0864 PD=1.125 PS=0.91 NRD=21.552 NRS=0 M=1 R=4.26667
+ SA=75006.8 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1018 N_A_1302_47#_M1018_d N_A0_M1018_g N_A_79_21#_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.336 AS=0.0864 PD=1.69 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75007.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1028 N_A_1302_47#_M1018_d N_A_1259_199#_M1028_g N_VGND_M1028_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.336 AS=0.112372 PD=1.69 PS=0.992248 NRD=145.308 NRS=14.052
+ M=1 R=4.26667 SA=75008.4 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1023 N_A_1259_199#_M1023_d N_S_M1023_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.114128 PD=1.82 PS=1.00775 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_X_M1000_d N_A_79_21#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75008.9 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1000_d N_A_79_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75008.5 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_79_21#_M1003_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75008.1 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1003_d N_A_79_21#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75007.6 A=0.15 P=2.3 MULT=1
MM1019 N_X_M1019_d N_A_79_21#_M1019_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75007.2 A=0.15 P=2.3 MULT=1
MM1024 N_X_M1019_d N_A_79_21#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75006.8 A=0.15 P=2.3 MULT=1
MM1029 N_X_M1029_d N_A_79_21#_M1029_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75006.4 A=0.15 P=2.3 MULT=1
MM1030 N_X_M1029_d N_A_79_21#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1625 PD=1.27 PS=1.325 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75006 A=0.15 P=2.3 MULT=1
MM1010 N_A_792_297#_M1010_d N_S_M1010_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.5375 AS=0.1625 PD=2.075 PS=1.325 NRD=3.9203 NRS=9.8303 M=1 R=6.66667
+ SA=75003.6 SB=75005.5 A=0.15 P=2.3 MULT=1
MM1001 N_A_792_297#_M1010_d N_A0_M1001_g N_A_79_21#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.5375 AS=0.135 PD=2.075 PS=1.27 NRD=152.655 NRS=0 M=1 R=6.66667
+ SA=75004.8 SB=75004.3 A=0.15 P=2.3 MULT=1
MM1020 N_A_792_297#_M1020_d N_A0_M1020_g N_A_79_21#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2
+ SB=75003.8 A=0.15 P=2.3 MULT=1
MM1033 N_A_792_297#_M1020_d N_S_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1675 PD=1.27 PS=1.335 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.7
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1007 N_A_1302_297#_M1007_d N_A_1259_199#_M1007_g N_VPWR_M1033_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.6325 AS=0.1675 PD=2.265 PS=1.335 NRD=0 NRS=11.8003 M=1
+ R=6.66667 SA=75006.1 SB=75002.9 A=0.15 P=2.3 MULT=1
MM1016 N_A_1302_297#_M1007_d N_A1_M1016_g N_A_79_21#_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.6325 AS=0.135 PD=2.265 PS=1.27 NRD=195.01 NRS=0 M=1 R=6.66667
+ SA=75007.6 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1025 N_A_1302_297#_M1025_d N_A1_M1025_g N_A_79_21#_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 N_A_1302_297#_M1025_d N_A_1259_199#_M1008_g N_VPWR_M1008_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=14.7553 M=1 R=6.66667
+ SA=75008.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_1259_199#_M1012_d N_S_M1012_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.175 PD=2.52 PS=1.35 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX34_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_67 VNB 0 2.41285e-19 $X=0.15 $Y=-0.085
c_129 VPB 0 1.83894e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__mux2_8.spice.SKY130_FD_SC_HD__MUX2_8.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__nor4bb_2.pxi.spice
* Created: Tue Sep  1 19:19:39 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4BB_2%D_N N_D_N_M1015_g N_D_N_c_103_n N_D_N_M1003_g D_N
+ D_N N_D_N_c_104_n N_D_N_c_105_n PM_SKY130_FD_SC_HD__NOR4BB_2%D_N
x_PM_SKY130_FD_SC_HD__NOR4BB_2%C_N N_C_N_M1016_g N_C_N_M1018_g C_N N_C_N_c_137_n
+ N_C_N_c_138_n C_N PM_SKY130_FD_SC_HD__NOR4BB_2%C_N
x_PM_SKY130_FD_SC_HD__NOR4BB_2%A_201_93# N_A_201_93#_M1016_d N_A_201_93#_M1018_d
+ N_A_201_93#_c_173_n N_A_201_93#_M1002_g N_A_201_93#_M1001_g
+ N_A_201_93#_c_174_n N_A_201_93#_M1005_g N_A_201_93#_M1019_g
+ N_A_201_93#_c_183_n N_A_201_93#_c_175_n N_A_201_93#_c_176_n
+ N_A_201_93#_c_177_n N_A_201_93#_c_178_n N_A_201_93#_c_179_n
+ N_A_201_93#_c_180_n PM_SKY130_FD_SC_HD__NOR4BB_2%A_201_93#
x_PM_SKY130_FD_SC_HD__NOR4BB_2%A_27_410# N_A_27_410#_M1003_s N_A_27_410#_M1015_s
+ N_A_27_410#_c_258_n N_A_27_410#_M1006_g N_A_27_410#_M1008_g
+ N_A_27_410#_c_259_n N_A_27_410#_M1007_g N_A_27_410#_M1011_g
+ N_A_27_410#_c_260_n N_A_27_410#_c_269_n N_A_27_410#_c_270_n
+ N_A_27_410#_c_293_n N_A_27_410#_c_271_n N_A_27_410#_c_272_n
+ N_A_27_410#_c_261_n N_A_27_410#_c_262_n N_A_27_410#_c_263_n
+ N_A_27_410#_c_264_n N_A_27_410#_c_274_n N_A_27_410#_c_265_n
+ PM_SKY130_FD_SC_HD__NOR4BB_2%A_27_410#
x_PM_SKY130_FD_SC_HD__NOR4BB_2%B N_B_c_364_n N_B_M1000_g N_B_M1009_g N_B_c_365_n
+ N_B_M1017_g N_B_M1013_g B N_B_c_366_n N_B_c_367_n
+ PM_SKY130_FD_SC_HD__NOR4BB_2%B
x_PM_SKY130_FD_SC_HD__NOR4BB_2%A N_A_c_411_n N_A_M1010_g N_A_M1004_g N_A_c_412_n
+ N_A_M1014_g N_A_M1012_g A N_A_c_414_n PM_SKY130_FD_SC_HD__NOR4BB_2%A
x_PM_SKY130_FD_SC_HD__NOR4BB_2%VPWR N_VPWR_M1015_d N_VPWR_M1004_d N_VPWR_c_450_n
+ N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n VPWR N_VPWR_c_454_n
+ N_VPWR_c_455_n N_VPWR_c_449_n N_VPWR_c_457_n PM_SKY130_FD_SC_HD__NOR4BB_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR4BB_2%A_336_297# N_A_336_297#_M1001_s
+ N_A_336_297#_M1019_s N_A_336_297#_M1011_d N_A_336_297#_c_511_n
+ N_A_336_297#_c_509_n N_A_336_297#_c_510_n N_A_336_297#_c_515_n
+ PM_SKY130_FD_SC_HD__NOR4BB_2%A_336_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_2%A_418_297# N_A_418_297#_M1001_d
+ N_A_418_297#_M1009_s N_A_418_297#_c_540_n N_A_418_297#_c_551_n
+ N_A_418_297#_c_541_n N_A_418_297#_c_548_n
+ PM_SKY130_FD_SC_HD__NOR4BB_2%A_418_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_2%Y N_Y_M1002_s N_Y_M1006_s N_Y_M1000_s N_Y_M1010_s
+ N_Y_M1008_s N_Y_c_586_n N_Y_c_575_n N_Y_c_576_n N_Y_c_596_n N_Y_c_577_n
+ N_Y_c_578_n N_Y_c_624_n N_Y_c_579_n N_Y_c_628_n N_Y_c_580_n N_Y_c_581_n
+ N_Y_c_582_n Y Y N_Y_c_585_n PM_SKY130_FD_SC_HD__NOR4BB_2%Y
x_PM_SKY130_FD_SC_HD__NOR4BB_2%A_776_297# N_A_776_297#_M1009_d
+ N_A_776_297#_M1013_d N_A_776_297#_M1012_s N_A_776_297#_c_689_n
+ N_A_776_297#_c_690_n N_A_776_297#_c_708_n N_A_776_297#_c_691_n
+ N_A_776_297#_c_692_n PM_SKY130_FD_SC_HD__NOR4BB_2%A_776_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_2%VGND N_VGND_M1003_d N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_M1007_d N_VGND_M1000_d N_VGND_M1017_d N_VGND_M1014_d N_VGND_c_723_n
+ N_VGND_c_724_n N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n
+ N_VGND_c_729_n N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n VGND
+ N_VGND_c_733_n N_VGND_c_734_n N_VGND_c_735_n N_VGND_c_736_n N_VGND_c_737_n
+ N_VGND_c_738_n N_VGND_c_739_n PM_SKY130_FD_SC_HD__NOR4BB_2%VGND
cc_1 VNB N_D_N_c_103_n 0.0206607f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_2 VNB N_D_N_c_104_n 0.0224517f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_D_N_c_105_n 0.00532549f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_4 VNB N_C_N_c_137_n 0.0292119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_C_N_c_138_n 0.0189345f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_6 VNB C_N 0.00255344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_201_93#_c_173_n 0.0195354f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.675
cc_8 VNB N_A_201_93#_c_174_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_9 VNB N_A_201_93#_c_175_n 0.00651919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_201_93#_c_176_n 0.00128587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_201_93#_c_177_n 0.00556811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_201_93#_c_178_n 0.0147975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_201_93#_c_179_n 0.00209682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_201_93#_c_180_n 0.0473019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_410#_c_258_n 0.0160118f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.675
cc_16 VNB N_A_27_410#_c_259_n 0.0193055f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_17 VNB N_A_27_410#_c_260_n 0.0223059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_410#_c_261_n 5.25319e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_410#_c_262_n 0.00297898f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_410#_c_263_n 0.00326724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_410#_c_264_n 0.0192081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_410#_c_265_n 0.036201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B_c_364_n 0.0192306f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_24 VNB N_B_c_365_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_25 VNB N_B_c_366_n 0.00701525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B_c_367_n 0.0334867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_c_411_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_28 VNB N_A_c_412_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_29 VNB A 0.0171554f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.325
cc_30 VNB N_A_c_414_n 0.0384775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_449_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_575_n 0.00270239f $X=-0.19 $Y=-0.24 $X2=0.602 $Y2=1.53
cc_33 VNB N_Y_c_576_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_577_n 0.00268301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_578_n 0.00567378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_579_n 0.00494428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_580_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_581_n 0.00424437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_582_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB Y 0.0127995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_723_n 0.015023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_724_n 0.0213884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_725_n 0.0115094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_726_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_727_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_728_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_729_n 0.0101986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_730_n 0.0330496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_731_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_732_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_733_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_734_n 0.0231858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_735_n 0.00631201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_736_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_737_n 0.0259444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_738_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_739_n 0.313097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VPB N_D_N_M1015_g 0.0560989f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.26
cc_59 VPB N_D_N_c_104_n 0.00472275f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_60 VPB N_D_N_c_105_n 0.00236867f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_61 VPB N_C_N_M1018_g 0.0219484f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_62 VPB N_C_N_c_137_n 0.0065137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB C_N 4.8227e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_201_93#_M1001_g 0.0224069f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_65 VPB N_A_201_93#_M1019_g 0.0180556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_201_93#_c_183_n 0.009855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_201_93#_c_176_n 0.00555828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_201_93#_c_180_n 0.00904094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_410#_M1008_g 0.0185874f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_70 VPB N_A_27_410#_M1011_g 0.0221343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_410#_c_260_n 0.0272058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_410#_c_269_n 0.0155282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_410#_c_270_n 0.0203127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_410#_c_271_n 0.00362779f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_410#_c_272_n 0.00172096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_410#_c_261_n 0.00197688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_410#_c_274_n 0.011274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_410#_c_265_n 0.00537609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_B_M1009_g 0.022023f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_80 VPB N_B_M1013_g 0.0186831f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_81 VPB N_B_c_367_n 0.00423903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_M1004_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_83 VPB N_A_M1012_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_84 VPB N_A_c_414_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_450_n 0.0127939f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_86 VPB N_VPWR_c_451_n 0.00489695f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_87 VPB N_VPWR_c_452_n 0.102776f $X=-0.19 $Y=1.305 $X2=0.602 $Y2=1.16
cc_88 VPB N_VPWR_c_453_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_454_n 0.0144832f $X=-0.19 $Y=1.305 $X2=0.602 $Y2=1.53
cc_90 VPB N_VPWR_c_455_n 0.0183432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_449_n 0.0599656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_457_n 0.00518909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_336_297#_c_509_n 0.00297507f $X=-0.19 $Y=1.305 $X2=0.602 $Y2=1.16
cc_94 VPB N_A_336_297#_c_510_n 0.0104647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_418_297#_c_540_n 0.00749495f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_96 VPB N_A_418_297#_c_541_n 0.00246174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB Y 0.0108304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_585_n 0.00491927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_776_297#_c_689_n 0.00246327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_776_297#_c_690_n 0.0023993f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_101 VPB N_A_776_297#_c_691_n 0.0124129f $X=-0.19 $Y=1.305 $X2=0.602 $Y2=1.16
cc_102 VPB N_A_776_297#_c_692_n 0.0321878f $X=-0.19 $Y=1.305 $X2=0.602 $Y2=1.53
cc_103 N_D_N_M1015_g N_C_N_M1018_g 0.0242958f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_104 N_D_N_c_105_n N_C_N_M1018_g 0.00412572f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_105 N_D_N_c_104_n N_C_N_c_137_n 0.0204437f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_106 N_D_N_c_105_n N_C_N_c_137_n 0.00229322f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_107 N_D_N_c_103_n N_C_N_c_138_n 0.0116141f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_108 N_D_N_c_104_n C_N 2.74648e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_109 N_D_N_c_105_n C_N 0.0259606f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_110 N_D_N_M1015_g N_A_201_93#_c_183_n 2.24045e-19 $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_111 N_D_N_c_105_n N_A_201_93#_c_183_n 0.0115316f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_112 N_D_N_c_105_n N_A_201_93#_c_176_n 0.00632295f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_113 N_D_N_M1015_g N_A_27_410#_c_260_n 0.014005f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_114 N_D_N_c_103_n N_A_27_410#_c_260_n 0.00523955f $X=0.51 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_D_N_c_104_n N_A_27_410#_c_260_n 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_116 N_D_N_c_105_n N_A_27_410#_c_260_n 0.0528642f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_117 N_D_N_M1015_g N_A_27_410#_c_270_n 0.0145821f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_118 N_D_N_c_104_n N_A_27_410#_c_270_n 8.23566e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_119 N_D_N_c_105_n N_A_27_410#_c_270_n 0.0261108f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_120 N_D_N_c_103_n N_A_27_410#_c_264_n 0.00496254f $X=0.51 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_D_N_c_104_n N_A_27_410#_c_264_n 0.0012161f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_122 N_D_N_c_105_n N_A_27_410#_c_264_n 0.00276502f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_123 N_D_N_c_105_n N_VPWR_M1015_d 0.00454642f $X=0.51 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_124 N_D_N_M1015_g N_VPWR_c_450_n 0.00964097f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_125 N_D_N_M1015_g N_VPWR_c_454_n 0.00332796f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_126 N_D_N_M1015_g N_VPWR_c_449_n 0.00485312f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_127 N_D_N_c_103_n N_VGND_c_723_n 0.00286444f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_128 N_D_N_c_105_n N_VGND_c_723_n 0.0128638f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_129 N_D_N_c_103_n N_VGND_c_734_n 0.00483235f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_130 N_D_N_c_103_n N_VGND_c_739_n 0.00512902f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_131 N_C_N_M1018_g N_A_201_93#_c_183_n 0.00340004f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_132 N_C_N_c_137_n N_A_201_93#_c_183_n 0.0036075f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_133 C_N N_A_201_93#_c_183_n 0.013928f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_134 N_C_N_c_137_n N_A_201_93#_c_175_n 2.76201e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_C_N_c_138_n N_A_201_93#_c_175_n 0.00413818f $X=1.027 $Y=0.995 $X2=0
+ $Y2=0
cc_136 C_N N_A_201_93#_c_175_n 0.00618183f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_137 N_C_N_M1018_g N_A_201_93#_c_176_n 0.00309661f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_138 N_C_N_c_137_n N_A_201_93#_c_176_n 2.76201e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_139 C_N N_A_201_93#_c_176_n 0.00618183f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_140 N_C_N_c_137_n N_A_201_93#_c_178_n 0.0032984f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_141 N_C_N_c_138_n N_A_201_93#_c_178_n 3.46718e-19 $X=1.027 $Y=0.995 $X2=0
+ $Y2=0
cc_142 C_N N_A_201_93#_c_178_n 0.0140382f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_143 N_C_N_c_137_n N_A_201_93#_c_179_n 7.34273e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_144 C_N N_A_201_93#_c_179_n 0.0149497f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_145 N_C_N_c_137_n N_A_201_93#_c_180_n 0.00540018f $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_146 C_N N_A_201_93#_c_180_n 5.37965e-19 $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_147 N_C_N_M1018_g N_A_27_410#_c_270_n 0.0145954f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_148 C_N N_A_27_410#_c_270_n 0.00120587f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_149 N_C_N_M1018_g N_VPWR_c_452_n 5.4793e-19 $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_150 N_C_N_c_138_n N_VGND_c_723_n 0.00286381f $X=1.027 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C_N_c_138_n N_VGND_c_724_n 0.00510437f $X=1.027 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C_N_c_138_n N_VGND_c_725_n 0.0029214f $X=1.027 $Y=0.995 $X2=0 $Y2=0
cc_153 N_C_N_c_138_n N_VGND_c_739_n 0.00512902f $X=1.027 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_201_93#_c_174_n N_A_27_410#_c_258_n 0.0258694f $X=2.435 $Y=0.995
+ $X2=0 $Y2=0
cc_155 N_A_201_93#_M1019_g N_A_27_410#_M1008_g 0.0423624f $X=2.435 $Y=1.985
+ $X2=0 $Y2=0
cc_156 N_A_201_93#_M1018_d N_A_27_410#_c_270_n 0.00213259f $X=1.03 $Y=1.485
+ $X2=0 $Y2=0
cc_157 N_A_201_93#_c_183_n N_A_27_410#_c_270_n 0.040187f $X=1.405 $Y=1.62 $X2=0
+ $Y2=0
cc_158 N_A_201_93#_c_177_n N_A_27_410#_c_270_n 0.00495382f $X=2.225 $Y=1.16
+ $X2=0 $Y2=0
cc_159 N_A_201_93#_c_183_n N_A_27_410#_c_293_n 0.0106276f $X=1.405 $Y=1.62 $X2=0
+ $Y2=0
cc_160 N_A_201_93#_M1001_g N_A_27_410#_c_271_n 0.0155522f $X=2.015 $Y=1.985
+ $X2=0 $Y2=0
cc_161 N_A_201_93#_M1019_g N_A_27_410#_c_271_n 0.011895f $X=2.435 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_201_93#_c_177_n N_A_27_410#_c_271_n 0.0332646f $X=2.225 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_201_93#_c_180_n N_A_27_410#_c_271_n 0.00283185f $X=2.435 $Y=1.16
+ $X2=0 $Y2=0
cc_164 N_A_201_93#_c_183_n N_A_27_410#_c_272_n 0.00545025f $X=1.405 $Y=1.62
+ $X2=0 $Y2=0
cc_165 N_A_201_93#_c_176_n N_A_27_410#_c_272_n 0.00918169f $X=1.49 $Y=1.525
+ $X2=0 $Y2=0
cc_166 N_A_201_93#_c_177_n N_A_27_410#_c_272_n 0.0136617f $X=2.225 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_201_93#_c_180_n N_A_27_410#_c_272_n 0.00422084f $X=2.435 $Y=1.16
+ $X2=0 $Y2=0
cc_168 N_A_201_93#_c_180_n N_A_27_410#_c_261_n 0.00337404f $X=2.435 $Y=1.16
+ $X2=0 $Y2=0
cc_169 N_A_201_93#_c_177_n N_A_27_410#_c_262_n 0.0149758f $X=2.225 $Y=1.16 $X2=0
+ $Y2=0
cc_170 N_A_201_93#_c_180_n N_A_27_410#_c_262_n 0.00265637f $X=2.435 $Y=1.16
+ $X2=0 $Y2=0
cc_171 N_A_201_93#_c_180_n N_A_27_410#_c_265_n 0.0182371f $X=2.435 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_201_93#_M1001_g N_VPWR_c_452_n 0.00357877f $X=2.015 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_201_93#_M1019_g N_VPWR_c_452_n 0.00357877f $X=2.435 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_201_93#_M1001_g N_VPWR_c_449_n 0.00655123f $X=2.015 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_201_93#_M1019_g N_VPWR_c_449_n 0.00525237f $X=2.435 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_201_93#_M1001_g N_A_336_297#_c_511_n 2.50677e-19 $X=2.015 $Y=1.985
+ $X2=0 $Y2=0
cc_177 N_A_201_93#_M1019_g N_A_336_297#_c_511_n 0.00251788f $X=2.435 $Y=1.985
+ $X2=0 $Y2=0
cc_178 N_A_201_93#_M1001_g N_A_336_297#_c_510_n 0.00274596f $X=2.015 $Y=1.985
+ $X2=0 $Y2=0
cc_179 N_A_201_93#_M1019_g N_A_336_297#_c_510_n 2.02748e-19 $X=2.435 $Y=1.985
+ $X2=0 $Y2=0
cc_180 N_A_201_93#_M1001_g N_A_336_297#_c_515_n 0.0101149f $X=2.015 $Y=1.985
+ $X2=0 $Y2=0
cc_181 N_A_201_93#_M1019_g N_A_336_297#_c_515_n 0.00685285f $X=2.435 $Y=1.985
+ $X2=0 $Y2=0
cc_182 N_A_201_93#_M1019_g N_A_418_297#_c_540_n 0.00936118f $X=2.435 $Y=1.985
+ $X2=0 $Y2=0
cc_183 N_A_201_93#_c_173_n N_Y_c_586_n 0.0116673f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_201_93#_c_174_n N_Y_c_586_n 0.00630972f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_201_93#_c_178_n N_Y_c_586_n 0.00261667f $X=1.14 $Y=0.66 $X2=0 $Y2=0
cc_186 N_A_201_93#_c_174_n N_Y_c_575_n 0.0100105f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_201_93#_c_173_n N_Y_c_576_n 0.00403778f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_201_93#_c_174_n N_Y_c_576_n 0.00113286f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_201_93#_c_175_n N_Y_c_576_n 0.00287104f $X=1.49 $Y=1.075 $X2=0 $Y2=0
cc_190 N_A_201_93#_c_177_n N_Y_c_576_n 0.026256f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_201_93#_c_178_n N_Y_c_576_n 0.00395529f $X=1.14 $Y=0.66 $X2=0 $Y2=0
cc_192 N_A_201_93#_c_180_n N_Y_c_576_n 0.00230339f $X=2.435 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_201_93#_c_174_n N_Y_c_596_n 5.22228e-19 $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_201_93#_M1019_g N_Y_c_585_n 6.8816e-19 $X=2.435 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_201_93#_c_178_n N_VGND_c_723_n 8.15804e-19 $X=1.14 $Y=0.66 $X2=0
+ $Y2=0
cc_196 N_A_201_93#_c_178_n N_VGND_c_724_n 0.0116706f $X=1.14 $Y=0.66 $X2=0 $Y2=0
cc_197 N_A_201_93#_c_173_n N_VGND_c_725_n 0.00795516f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_201_93#_c_177_n N_VGND_c_725_n 0.0097255f $X=2.225 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_201_93#_c_178_n N_VGND_c_725_n 0.00276945f $X=1.14 $Y=0.66 $X2=0
+ $Y2=0
cc_200 N_A_201_93#_c_180_n N_VGND_c_725_n 0.0025888f $X=2.435 $Y=1.16 $X2=0
+ $Y2=0
cc_201 N_A_201_93#_c_174_n N_VGND_c_726_n 0.00146448f $X=2.435 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_201_93#_c_173_n N_VGND_c_731_n 0.00541359f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_201_93#_c_174_n N_VGND_c_731_n 0.00423334f $X=2.435 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_201_93#_c_173_n N_VGND_c_739_n 0.0109543f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_201_93#_c_174_n N_VGND_c_739_n 0.0057435f $X=2.435 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_201_93#_c_178_n N_VGND_c_739_n 0.015582f $X=1.14 $Y=0.66 $X2=0 $Y2=0
cc_207 N_A_27_410#_c_270_n N_VPWR_M1015_d 0.0055834f $X=1.745 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_208 N_A_27_410#_c_270_n N_VPWR_c_450_n 0.0192998f $X=1.745 $Y=1.97 $X2=0
+ $Y2=0
cc_209 N_A_27_410#_M1008_g N_VPWR_c_452_n 0.00357877f $X=2.855 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_27_410#_M1011_g N_VPWR_c_452_n 0.00357877f $X=3.275 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_27_410#_c_270_n N_VPWR_c_452_n 0.0136387f $X=1.745 $Y=1.97 $X2=0
+ $Y2=0
cc_212 N_A_27_410#_c_269_n N_VPWR_c_454_n 0.0168497f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_213 N_A_27_410#_c_270_n N_VPWR_c_454_n 0.00227656f $X=1.745 $Y=1.97 $X2=0
+ $Y2=0
cc_214 N_A_27_410#_M1008_g N_VPWR_c_449_n 0.00525237f $X=2.855 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_27_410#_M1011_g N_VPWR_c_449_n 0.00655123f $X=3.275 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_27_410#_c_269_n N_VPWR_c_449_n 0.00987287f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_217 N_A_27_410#_c_270_n N_VPWR_c_449_n 0.0277909f $X=1.745 $Y=1.97 $X2=0
+ $Y2=0
cc_218 N_A_27_410#_c_270_n N_A_336_297#_M1001_s 0.00528853f $X=1.745 $Y=1.97
+ $X2=-0.19 $Y2=-0.24
cc_219 N_A_27_410#_c_293_n N_A_336_297#_M1001_s 0.00886748f $X=1.83 $Y=1.885
+ $X2=-0.19 $Y2=-0.24
cc_220 N_A_27_410#_c_272_n N_A_336_297#_M1001_s 0.00119074f $X=1.915 $Y=1.5
+ $X2=-0.19 $Y2=-0.24
cc_221 N_A_27_410#_c_271_n N_A_336_297#_M1019_s 0.00236076f $X=2.56 $Y=1.5 $X2=0
+ $Y2=0
cc_222 N_A_27_410#_M1008_g N_A_336_297#_c_509_n 0.00970685f $X=2.855 $Y=1.985
+ $X2=0 $Y2=0
cc_223 N_A_27_410#_M1011_g N_A_336_297#_c_509_n 0.00970685f $X=3.275 $Y=1.985
+ $X2=0 $Y2=0
cc_224 N_A_27_410#_c_270_n N_A_336_297#_c_510_n 0.0184288f $X=1.745 $Y=1.97
+ $X2=0 $Y2=0
cc_225 N_A_27_410#_c_271_n N_A_336_297#_c_510_n 6.81309e-19 $X=2.56 $Y=1.5 $X2=0
+ $Y2=0
cc_226 N_A_27_410#_c_271_n N_A_418_297#_M1001_d 0.00181725f $X=2.56 $Y=1.5
+ $X2=-0.19 $Y2=-0.24
cc_227 N_A_27_410#_M1008_g N_A_418_297#_c_540_n 0.011938f $X=2.855 $Y=1.985
+ $X2=0 $Y2=0
cc_228 N_A_27_410#_M1011_g N_A_418_297#_c_540_n 0.0124526f $X=3.275 $Y=1.985
+ $X2=0 $Y2=0
cc_229 N_A_27_410#_c_271_n N_A_418_297#_c_540_n 0.0149682f $X=2.56 $Y=1.5 $X2=0
+ $Y2=0
cc_230 N_A_27_410#_c_263_n N_A_418_297#_c_540_n 0.00363217f $X=3.24 $Y=1.16
+ $X2=0 $Y2=0
cc_231 N_A_27_410#_c_271_n N_A_418_297#_c_548_n 0.0102367f $X=2.56 $Y=1.5 $X2=0
+ $Y2=0
cc_232 N_A_27_410#_c_258_n N_Y_c_586_n 5.22228e-19 $X=2.855 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_27_410#_c_258_n N_Y_c_575_n 0.00865686f $X=2.855 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_27_410#_c_271_n N_Y_c_575_n 0.00506789f $X=2.56 $Y=1.5 $X2=0 $Y2=0
cc_235 N_A_27_410#_c_262_n N_Y_c_575_n 0.0140787f $X=2.73 $Y=1.175 $X2=0 $Y2=0
cc_236 N_A_27_410#_c_263_n N_Y_c_575_n 0.0119703f $X=3.24 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_27_410#_c_265_n N_Y_c_575_n 3.70222e-19 $X=3.275 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_27_410#_c_258_n N_Y_c_596_n 0.00630972f $X=2.855 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_27_410#_c_259_n N_Y_c_596_n 0.0109565f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_27_410#_c_259_n N_Y_c_577_n 0.0109318f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_27_410#_c_263_n N_Y_c_577_n 0.0123531f $X=3.24 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_27_410#_c_265_n N_Y_c_577_n 6.17037e-19 $X=3.275 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_27_410#_c_258_n N_Y_c_580_n 0.00113286f $X=2.855 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_27_410#_c_259_n N_Y_c_580_n 0.00113286f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_27_410#_c_263_n N_Y_c_580_n 0.0265405f $X=3.24 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_27_410#_c_265_n N_Y_c_580_n 0.00230339f $X=3.275 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_27_410#_c_259_n Y 0.00320826f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_27_410#_M1011_g Y 0.00428969f $X=3.275 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_27_410#_c_263_n Y 0.0178198f $X=3.24 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_27_410#_c_265_n Y 0.00706473f $X=3.275 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_27_410#_M1008_g N_Y_c_585_n 0.00508901f $X=2.855 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_27_410#_M1011_g N_Y_c_585_n 0.0143034f $X=3.275 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_27_410#_c_271_n N_Y_c_585_n 0.00766226f $X=2.56 $Y=1.5 $X2=0 $Y2=0
cc_254 N_A_27_410#_c_263_n N_Y_c_585_n 0.037224f $X=3.24 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_27_410#_c_265_n N_Y_c_585_n 0.00276353f $X=3.275 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_27_410#_c_264_n N_VGND_c_723_n 0.0148719f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_257 N_A_27_410#_c_258_n N_VGND_c_726_n 0.00146339f $X=2.855 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_27_410#_c_264_n N_VGND_c_734_n 0.0114766f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_259 N_A_27_410#_c_258_n N_VGND_c_736_n 0.00423334f $X=2.855 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_27_410#_c_259_n N_VGND_c_736_n 0.00423334f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_27_410#_c_259_n N_VGND_c_737_n 0.00336341f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_27_410#_c_258_n N_VGND_c_739_n 0.0057435f $X=2.855 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A_27_410#_c_259_n N_VGND_c_739_n 0.0070399f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_27_410#_c_264_n N_VGND_c_739_n 0.0127086f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_265 N_B_c_365_n N_A_c_411_n 0.0194576f $X=4.655 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_266 N_B_M1013_g N_A_M1004_g 0.0194576f $X=4.655 $Y=1.985 $X2=0 $Y2=0
cc_267 N_B_c_366_n A 0.0175712f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B_c_366_n N_A_c_414_n 0.00192044f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B_c_367_n N_A_c_414_n 0.0194576f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B_M1009_g N_VPWR_c_452_n 0.00357877f $X=4.235 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B_M1013_g N_VPWR_c_452_n 0.00357877f $X=4.655 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B_M1009_g N_VPWR_c_449_n 0.00655123f $X=4.235 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B_M1013_g N_VPWR_c_449_n 0.00525237f $X=4.655 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B_M1009_g N_A_418_297#_c_540_n 0.0125772f $X=4.235 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B_c_366_n N_A_418_297#_c_540_n 0.00361768f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B_M1013_g N_A_418_297#_c_551_n 0.00218056f $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_277 N_B_M1009_g N_A_418_297#_c_541_n 3.11936e-19 $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_B_M1013_g N_A_418_297#_c_541_n 0.00505833f $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_279 N_B_c_366_n N_A_418_297#_c_541_n 0.0220991f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B_c_367_n N_A_418_297#_c_541_n 0.00220262f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_281 N_B_c_364_n N_Y_c_578_n 0.0110858f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_c_366_n N_Y_c_578_n 0.00789367f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_283 N_B_c_364_n N_Y_c_624_n 0.0109565f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B_c_365_n N_Y_c_624_n 0.00630972f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B_c_365_n N_Y_c_579_n 0.00865686f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B_c_366_n N_Y_c_579_n 0.0258498f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_287 N_B_c_365_n N_Y_c_628_n 5.22228e-19 $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B_c_364_n N_Y_c_582_n 0.00113286f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B_c_365_n N_Y_c_582_n 0.00113286f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B_c_366_n N_Y_c_582_n 0.0265405f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_291 N_B_c_367_n N_Y_c_582_n 0.00230339f $X=4.655 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B_c_364_n Y 0.0189704f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B_M1009_g Y 0.00604746f $X=4.235 $Y=1.985 $X2=0 $Y2=0
cc_294 N_B_c_366_n Y 0.0169224f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_295 N_B_M1009_g N_A_776_297#_c_689_n 0.00964167f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_B_M1013_g N_A_776_297#_c_689_n 0.0135526f $X=4.655 $Y=1.985 $X2=0 $Y2=0
cc_297 N_B_M1013_g N_A_776_297#_c_690_n 2.36936e-19 $X=4.655 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_B_c_366_n N_A_776_297#_c_690_n 0.0147624f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_299 N_B_c_364_n N_VGND_c_727_n 0.00423334f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B_c_365_n N_VGND_c_727_n 0.00423334f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B_c_365_n N_VGND_c_728_n 0.00146339f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B_c_364_n N_VGND_c_737_n 0.00336341f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B_c_364_n N_VGND_c_739_n 0.0070399f $X=4.235 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B_c_365_n N_VGND_c_739_n 0.0057435f $X=4.655 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_M1004_g N_VPWR_c_451_n 0.00296718f $X=5.075 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A_M1012_g N_VPWR_c_451_n 0.00274642f $X=5.495 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A_M1004_g N_VPWR_c_452_n 0.00585385f $X=5.075 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_M1012_g N_VPWR_c_455_n 0.00541359f $X=5.495 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_M1004_g N_VPWR_c_449_n 0.010464f $X=5.075 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_M1012_g N_VPWR_c_449_n 0.0104699f $X=5.495 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A_c_411_n N_Y_c_624_n 5.22228e-19 $X=5.075 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_c_411_n N_Y_c_579_n 0.0113987f $X=5.075 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_c_412_n N_Y_c_579_n 0.0026268f $X=5.495 $Y=0.995 $X2=0 $Y2=0
cc_314 A N_Y_c_579_n 0.0258288f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_315 N_A_c_414_n N_Y_c_579_n 0.00230167f $X=5.495 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_c_411_n N_Y_c_628_n 0.00630972f $X=5.075 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_c_412_n N_Y_c_628_n 0.00539651f $X=5.495 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A_M1004_g N_A_776_297#_c_691_n 0.0148206f $X=5.075 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A_M1012_g N_A_776_297#_c_691_n 0.0122159f $X=5.495 $Y=1.985 $X2=0 $Y2=0
cc_320 A N_A_776_297#_c_691_n 0.0548813f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_321 N_A_c_414_n N_A_776_297#_c_691_n 0.00212548f $X=5.495 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_M1004_g N_A_776_297#_c_692_n 6.39954e-19 $X=5.075 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_M1012_g N_A_776_297#_c_692_n 0.0102794f $X=5.495 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A_c_411_n N_VGND_c_728_n 0.00146448f $X=5.075 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_c_412_n N_VGND_c_730_n 0.00366968f $X=5.495 $Y=0.995 $X2=0 $Y2=0
cc_326 A N_VGND_c_730_n 0.0234299f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_327 N_A_c_411_n N_VGND_c_733_n 0.00423334f $X=5.075 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_c_412_n N_VGND_c_733_n 0.00541359f $X=5.495 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_c_411_n N_VGND_c_739_n 0.0057435f $X=5.075 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_c_412_n N_VGND_c_739_n 0.0104699f $X=5.495 $Y=0.995 $X2=0 $Y2=0
cc_331 N_VPWR_c_449_n N_A_336_297#_M1001_s 0.00209344f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_332 N_VPWR_c_449_n N_A_336_297#_M1019_s 0.00215227f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_449_n N_A_336_297#_M1011_d 0.00209344f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_452_n N_A_336_297#_c_510_n 0.115227f $X=5.16 $Y=2.72 $X2=0 $Y2=0
cc_335 N_VPWR_c_449_n N_A_336_297#_c_510_n 0.0722978f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_449_n N_A_418_297#_M1001_d 0.0021603f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_337 N_VPWR_c_449_n N_A_418_297#_M1009_s 0.00216833f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_452_n N_A_418_297#_c_540_n 0.00353234f $X=5.16 $Y=2.72 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_449_n N_A_418_297#_c_540_n 0.00893405f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_449_n N_Y_M1008_s 0.00216833f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_341 N_VPWR_c_449_n N_A_776_297#_M1009_d 0.00225742f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_342 N_VPWR_c_449_n N_A_776_297#_M1013_d 0.0024645f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_449_n N_A_776_297#_M1012_s 0.00221616f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_452_n N_A_776_297#_c_689_n 0.0526575f $X=5.16 $Y=2.72 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_449_n N_A_776_297#_c_689_n 0.0330421f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_452_n N_A_776_297#_c_708_n 0.012886f $X=5.16 $Y=2.72 $X2=0 $Y2=0
cc_347 N_VPWR_c_449_n N_A_776_297#_c_708_n 0.00808224f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_M1004_d N_A_776_297#_c_691_n 0.00165831f $X=5.15 $Y=1.485 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_451_n N_A_776_297#_c_691_n 0.0126919f $X=5.285 $Y=1.96 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_455_n N_A_776_297#_c_692_n 0.0210175f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_449_n N_A_776_297#_c_692_n 0.0124268f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_352 N_A_336_297#_c_515_n N_A_418_297#_M1001_d 0.00312348f $X=2.48 $Y=2.34
+ $X2=-0.19 $Y2=1.305
cc_353 N_A_336_297#_M1019_s N_A_418_297#_c_540_n 0.00372891f $X=2.51 $Y=1.485
+ $X2=0 $Y2=0
cc_354 N_A_336_297#_M1011_d N_A_418_297#_c_540_n 0.00500159f $X=3.35 $Y=1.485
+ $X2=0 $Y2=0
cc_355 N_A_336_297#_c_511_n N_A_418_297#_c_540_n 0.0617287f $X=2.605 $Y=2.34
+ $X2=0 $Y2=0
cc_356 N_A_336_297#_c_515_n N_A_418_297#_c_540_n 0.00535822f $X=2.48 $Y=2.34
+ $X2=0 $Y2=0
cc_357 N_A_336_297#_c_515_n N_A_418_297#_c_548_n 0.0112564f $X=2.48 $Y=2.34
+ $X2=0 $Y2=0
cc_358 N_A_336_297#_c_509_n N_Y_M1008_s 0.00316492f $X=3.485 $Y=2.3 $X2=0 $Y2=0
cc_359 N_A_336_297#_M1011_d Y 8.14469e-19 $X=3.35 $Y=1.485 $X2=0 $Y2=0
cc_360 N_A_336_297#_M1011_d N_Y_c_585_n 0.00233638f $X=3.35 $Y=1.485 $X2=0 $Y2=0
cc_361 N_A_336_297#_c_509_n N_A_776_297#_c_689_n 0.0200043f $X=3.485 $Y=2.3
+ $X2=0 $Y2=0
cc_362 N_A_418_297#_c_540_n N_Y_M1008_s 0.00317879f $X=4.32 $Y=1.96 $X2=0 $Y2=0
cc_363 N_A_418_297#_c_540_n Y 0.0350081f $X=4.32 $Y=1.96 $X2=0 $Y2=0
cc_364 N_A_418_297#_c_541_n Y 0.00776062f $X=4.445 $Y=1.62 $X2=0 $Y2=0
cc_365 N_A_418_297#_c_540_n N_Y_c_585_n 0.0368071f $X=4.32 $Y=1.96 $X2=0 $Y2=0
cc_366 N_A_418_297#_c_540_n N_A_776_297#_M1009_d 0.008575f $X=4.32 $Y=1.96
+ $X2=-0.19 $Y2=1.305
cc_367 N_A_418_297#_M1009_s N_A_776_297#_c_689_n 0.00316082f $X=4.31 $Y=1.485
+ $X2=0 $Y2=0
cc_368 N_A_418_297#_c_540_n N_A_776_297#_c_689_n 0.0273995f $X=4.32 $Y=1.96
+ $X2=0 $Y2=0
cc_369 N_A_418_297#_c_551_n N_A_776_297#_c_689_n 0.0144551f $X=4.465 $Y=1.875
+ $X2=0 $Y2=0
cc_370 N_A_418_297#_c_541_n N_A_776_297#_c_690_n 0.00763548f $X=4.445 $Y=1.62
+ $X2=0 $Y2=0
cc_371 Y N_A_776_297#_M1009_d 0.00517093f $X=3.825 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_372 N_Y_c_579_n N_A_776_297#_c_690_n 0.00112383f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_373 N_Y_c_579_n N_A_776_297#_c_691_n 0.0037385f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_374 N_Y_c_575_n N_VGND_M1005_d 0.00162089f $X=2.9 $Y=0.815 $X2=0 $Y2=0
cc_375 N_Y_c_577_n N_VGND_M1007_d 0.00212652f $X=3.575 $Y=0.815 $X2=0 $Y2=0
cc_376 N_Y_c_581_n N_VGND_M1007_d 6.88755e-19 $X=3.785 $Y=0.815 $X2=0 $Y2=0
cc_377 N_Y_c_578_n N_VGND_M1000_d 0.00111439f $X=4.28 $Y=0.815 $X2=0 $Y2=0
cc_378 N_Y_c_581_n N_VGND_M1000_d 0.00213021f $X=3.785 $Y=0.815 $X2=0 $Y2=0
cc_379 N_Y_c_579_n N_VGND_M1017_d 0.00162089f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_380 N_Y_c_575_n N_VGND_c_726_n 0.0122559f $X=2.9 $Y=0.815 $X2=0 $Y2=0
cc_381 N_Y_c_578_n N_VGND_c_727_n 0.00198695f $X=4.28 $Y=0.815 $X2=0 $Y2=0
cc_382 N_Y_c_624_n N_VGND_c_727_n 0.0188551f $X=4.445 $Y=0.39 $X2=0 $Y2=0
cc_383 N_Y_c_579_n N_VGND_c_727_n 0.00198695f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_384 N_Y_c_579_n N_VGND_c_728_n 0.0122559f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_385 N_Y_c_579_n N_VGND_c_730_n 0.00835456f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_386 N_Y_c_586_n N_VGND_c_731_n 0.0188551f $X=2.225 $Y=0.39 $X2=0 $Y2=0
cc_387 N_Y_c_575_n N_VGND_c_731_n 0.00198695f $X=2.9 $Y=0.815 $X2=0 $Y2=0
cc_388 N_Y_c_579_n N_VGND_c_733_n 0.00198695f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_389 N_Y_c_628_n N_VGND_c_733_n 0.0188551f $X=5.285 $Y=0.39 $X2=0 $Y2=0
cc_390 N_Y_c_575_n N_VGND_c_736_n 0.00198695f $X=2.9 $Y=0.815 $X2=0 $Y2=0
cc_391 N_Y_c_596_n N_VGND_c_736_n 0.0188551f $X=3.065 $Y=0.39 $X2=0 $Y2=0
cc_392 N_Y_c_577_n N_VGND_c_736_n 0.00198695f $X=3.575 $Y=0.815 $X2=0 $Y2=0
cc_393 N_Y_c_577_n N_VGND_c_737_n 0.0130966f $X=3.575 $Y=0.815 $X2=0 $Y2=0
cc_394 N_Y_c_578_n N_VGND_c_737_n 0.00840711f $X=4.28 $Y=0.815 $X2=0 $Y2=0
cc_395 N_Y_c_581_n N_VGND_c_737_n 0.0370461f $X=3.785 $Y=0.815 $X2=0 $Y2=0
cc_396 N_Y_M1002_s N_VGND_c_739_n 0.00215201f $X=2.09 $Y=0.235 $X2=0 $Y2=0
cc_397 N_Y_M1006_s N_VGND_c_739_n 0.00215201f $X=2.93 $Y=0.235 $X2=0 $Y2=0
cc_398 N_Y_M1000_s N_VGND_c_739_n 0.00215201f $X=4.31 $Y=0.235 $X2=0 $Y2=0
cc_399 N_Y_M1010_s N_VGND_c_739_n 0.00215201f $X=5.15 $Y=0.235 $X2=0 $Y2=0
cc_400 N_Y_c_586_n N_VGND_c_739_n 0.0122069f $X=2.225 $Y=0.39 $X2=0 $Y2=0
cc_401 N_Y_c_575_n N_VGND_c_739_n 0.00835832f $X=2.9 $Y=0.815 $X2=0 $Y2=0
cc_402 N_Y_c_596_n N_VGND_c_739_n 0.0122069f $X=3.065 $Y=0.39 $X2=0 $Y2=0
cc_403 N_Y_c_577_n N_VGND_c_739_n 0.00450968f $X=3.575 $Y=0.815 $X2=0 $Y2=0
cc_404 N_Y_c_578_n N_VGND_c_739_n 0.00427976f $X=4.28 $Y=0.815 $X2=0 $Y2=0
cc_405 N_Y_c_624_n N_VGND_c_739_n 0.0122069f $X=4.445 $Y=0.39 $X2=0 $Y2=0
cc_406 N_Y_c_579_n N_VGND_c_739_n 0.00835832f $X=5.12 $Y=0.815 $X2=0 $Y2=0
cc_407 N_Y_c_628_n N_VGND_c_739_n 0.0122069f $X=5.285 $Y=0.39 $X2=0 $Y2=0
cc_408 N_Y_c_581_n N_VGND_c_739_n 0.00181962f $X=3.785 $Y=0.815 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__inv_12.spice
* Created: Tue Sep  1 19:09:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__inv_12.pex.spice"
.subckt sky130_fd_sc_hd__inv_12  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1001_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75004.2 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1008_d N_A_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1010_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1013_d N_A_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1020_d N_A_M1020_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1022 N_Y_M1020_d N_A_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.33475 PD=0.92 PS=2.33 NRD=0 NRS=46.152 M=1 R=4.33333
+ SA=75004.8 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75005.1 A=0.15
+ P=2.3 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75004.6
+ A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75004.2 A=0.15
+ P=2.3 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75003.8
+ A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75003.4
+ A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1012_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75003 A=0.15
+ P=2.3 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75002.5
+ A=0.15 P=2.3 MULT=1
MM1017 N_Y_M1016_d N_A_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75002.1
+ A=0.15 P=2.3 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5 SB=75001.7
+ A=0.15 P=2.3 MULT=1
MM1019 N_Y_M1018_d N_A_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004 SB=75001.3 A=0.15
+ P=2.3 MULT=1
MM1021 N_Y_M1021_d N_A_M1021_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4 SB=75000.9
+ A=0.15 P=2.3 MULT=1
MM1023 N_Y_M1021_d N_A_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.515 PD=1.27 PS=3.03 NRD=0 NRS=49.2303 M=1 R=6.66667 SA=75004.8 SB=75000.4
+ A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__inv_12.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.890000 1.495000 7.300000 1.575000 ;
        RECT 6.890000 1.575000 7.220000 2.420000 ;
        RECT 6.900000 0.305000 7.230000 0.740000 ;
        RECT 6.900000 0.740000 7.300000 0.825000 ;
        RECT 7.055000 0.825000 7.300000 0.865000 ;
        RECT 7.065000 1.445000 7.300000 1.495000 ;
        RECT 7.110000 0.865000 7.300000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.810000 1.495000 9.145000 2.465000 ;
        RECT 8.890000 0.265000 9.145000 0.885000 ;
        RECT 8.930000 0.885000 9.145000 1.495000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.020000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.380000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.040000  1.905000 6.380000 2.465000 ;
      RECT 6.060000  0.300000 6.390000 0.825000 ;
      RECT 6.190000  0.825000 6.390000 0.995000 ;
      RECT 6.190000  0.995000 6.940000 1.325000 ;
      RECT 6.190000  1.325000 6.380000 1.530000 ;
      RECT 6.550000  1.625000 6.720000 2.635000 ;
      RECT 6.560000  0.085000 6.730000 0.695000 ;
      RECT 7.390000  1.720000 7.565000 2.635000 ;
      RECT 7.400000  0.085000 7.570000 0.600000 ;
      RECT 7.905000  0.345000 8.165000 0.615000 ;
      RECT 7.905000  1.715000 8.235000 2.445000 ;
      RECT 7.965000  0.615000 8.165000 0.995000 ;
      RECT 7.965000  0.995000 8.760000 1.325000 ;
      RECT 7.965000  1.325000 8.235000 1.715000 ;
      RECT 8.390000  0.085000 8.720000 0.825000 ;
      RECT 8.425000  1.495000 8.640000 2.635000 ;
      RECT 9.315000  0.085000 9.565000 0.905000 ;
      RECT 9.315000  1.495000 9.565000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxbp_2
END LIBRARY

* File: sky130_fd_sc_hd__a41oi_1.pex.spice
* Created: Tue Sep  1 18:56:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A41OI_1%B1 3 6 8 9 13 15
c29 15 0 1.90117e-19 $X=0.577 $Y=0.995
c30 8 0 9.80834e-20 $X=0.695 $Y=1.19
r31 13 16 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.16
+ $X2=0.577 $Y2=1.325
r32 13 15 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.16
+ $X2=0.577 $Y2=0.995
r33 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.66 $Y=1.16 $X2=0.66
+ $Y2=1.53
r34 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.16 $X2=0.625 $Y2=1.16
r35 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r36 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%A4 3 5 7 8 9 13
c38 8 0 1.69815e-19 $X=1.155 $Y=1.19
c39 5 0 9.80834e-20 $X=1.105 $Y=0.995
c40 3 0 1.95659e-19 $X=1.045 $Y=1.985
r41 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.16
+ $X2=1.105 $Y2=1.325
r42 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.105 $Y=1.16
+ $X2=1.105 $Y2=1.53
r43 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.16 $X2=1.105 $Y2=1.16
r44 5 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=1.16
r45 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=0.56
r46 3 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.045 $Y=1.985
+ $X2=1.045 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%A3 3 6 8 9 10 15 17
c41 17 0 9.9429e-20 $X=1.615 $Y=0.995
r42 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.16
+ $X2=1.615 $Y2=1.325
r43 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.16
+ $X2=1.615 $Y2=0.995
r44 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.59 $Y=1.16 $X2=1.59
+ $Y2=1.53
r45 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.615
+ $Y=1.16 $X2=1.615 $Y2=1.16
r46 8 9 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=1.59 $Y=0.85 $X2=1.59
+ $Y2=1.16
r47 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.605 $Y=1.985
+ $X2=1.605 $Y2=1.325
r48 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.605 $Y=0.56
+ $X2=1.605 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%A2 3 6 8 9 10 15 17
r42 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.125 $Y=1.16
+ $X2=2.125 $Y2=1.325
r43 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.125 $Y=1.16
+ $X2=2.125 $Y2=0.995
r44 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.05 $Y=1.16 $X2=2.05
+ $Y2=1.53
r45 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.16 $X2=2.125 $Y2=1.16
r46 8 9 11.1643 $w=3.18e-07 $l=3.1e-07 $layer=LI1_cond $X=2.05 $Y=0.85 $X2=2.05
+ $Y2=1.16
r47 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.065 $Y=1.985
+ $X2=2.065 $Y2=1.325
r48 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.065 $Y=0.56
+ $X2=2.065 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%A1 1 3 6 8 9 15 16
r27 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.16 $X2=2.865 $Y2=1.16
r28 12 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.64 $Y=1.16
+ $X2=2.865 $Y2=1.16
r29 8 9 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=2.932 $Y=1.19
+ $X2=2.932 $Y2=1.53
r30 8 16 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=2.932 $Y=1.19 $X2=2.932
+ $Y2=1.16
r31 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.325
+ $X2=2.64 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.64 $Y=1.325 $X2=2.64
+ $Y2=1.985
r33 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=0.995
+ $X2=2.64 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.64 $Y=0.995 $X2=2.64
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%Y 1 2 3 10 13 14 15 20 22 23 24 25 36 43
c60 43 0 1.11467e-19 $X=0.235 $Y=1.87
c61 25 0 8.4192e-20 $X=0.235 $Y=2.21
c62 15 0 1.19731e-19 $X=1.29 $Y=0.38
r63 43 44 1.32747 $w=3.33e-07 $l=2.5e-08 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=1.845
r64 38 47 0.412815 $w=3.33e-07 $l=1.2e-08 $layer=LI1_cond $X=0.257 $Y=2.012
+ $X2=0.257 $Y2=2
r65 25 38 6.81145 $w=3.33e-07 $l=1.98e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.012
r66 24 47 3.44013 $w=3.33e-07 $l=1e-07 $layer=LI1_cond $X=0.257 $Y=1.9 $X2=0.257
+ $Y2=2
r67 24 43 1.03204 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=0.257 $Y=1.9 $X2=0.257
+ $Y2=1.87
r68 24 44 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.225 $Y=1.815
+ $X2=0.225 $Y2=1.845
r69 24 36 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.225 $Y=1.815
+ $X2=0.225 $Y2=1.66
r70 19 36 37.3477 $w=2.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.225 $Y=0.785
+ $X2=0.225 $Y2=1.66
r71 19 20 3.55013 $w=2.62e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=0.785
+ $X2=0.225 $Y2=0.7
r72 18 23 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.217 $Y=0.615
+ $X2=0.217 $Y2=0.45
r73 18 20 3.55013 $w=2.62e-07 $l=8.89101e-08 $layer=LI1_cond $X=0.217 $Y=0.615
+ $X2=0.225 $Y2=0.7
r74 14 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=0.38
+ $X2=2.85 $Y2=0.38
r75 14 15 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.685 $Y=0.38
+ $X2=1.29 $Y2=0.38
r76 12 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.205 $Y=0.465
+ $X2=1.29 $Y2=0.38
r77 12 13 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.205 $Y=0.465
+ $X2=1.205 $Y2=0.615
r78 11 20 2.9446 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.36 $Y=0.7 $X2=0.225
+ $Y2=0.7
r79 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.7
+ $X2=1.205 $Y2=0.615
r80 10 11 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.12 $Y=0.7 $X2=0.36
+ $Y2=0.7
r81 3 47 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r82 3 36 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r83 2 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.715
+ $Y=0.235 $X2=2.85 $Y2=0.38
r84 1 23 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%A_109_297# 1 2 3 10 12 14 18 20 22 24 29
r41 22 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=2.015
+ $X2=2.89 $Y2=1.93
r42 22 24 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=2.89 $Y=2.015
+ $X2=2.89 $Y2=2.3
r43 21 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=1.93
+ $X2=1.845 $Y2=1.93
r44 20 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=1.93
+ $X2=2.89 $Y2=1.93
r45 20 21 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.765 $Y=1.93
+ $X2=1.93 $Y2=1.93
r46 16 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=2.015
+ $X2=1.845 $Y2=1.93
r47 16 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.845 $Y=2.015
+ $X2=1.845 $Y2=2.3
r48 15 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=1.93
+ $X2=0.72 $Y2=1.93
r49 14 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=1.93
+ $X2=1.845 $Y2=1.93
r50 14 15 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.76 $Y=1.93
+ $X2=0.845 $Y2=1.93
r51 10 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.015
+ $X2=0.72 $Y2=1.93
r52 10 12 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=2.015
+ $X2=0.72 $Y2=2.3
r53 3 31 600 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.485 $X2=2.85 $Y2=1.93
r54 3 24 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.485 $X2=2.85 $Y2=2.3
r55 2 29 600 $w=1.7e-07 $l=5.21009e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.485 $X2=1.845 $Y2=1.93
r56 2 18 600 $w=1.7e-07 $l=8.937e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.485 $X2=1.845 $Y2=2.3
r57 1 27 600 $w=1.7e-07 $l=5.41941e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.76 $Y2=1.93
r58 1 12 600 $w=1.7e-07 $l=9.16215e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.76 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%VPWR 1 2 9 13 16 17 18 20 30 31 34
r51 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 28 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.285 $Y2=2.72
r57 25 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=2.72
+ $X2=1.285 $Y2=2.72
r59 20 22 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.12 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 18 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 18 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 16 27 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.38 $Y2=2.72
r64 15 30 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.99 $Y2=2.72
r65 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.38 $Y2=2.72
r66 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2.72
r67 11 13 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2.28
r68 7 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.72
r69 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.28
r70 2 13 600 $w=1.7e-07 $l=9.07097e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.485 $X2=2.38 $Y2=2.28
r71 1 9 600 $w=1.7e-07 $l=8.73613e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.285 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_1%VGND 1 8 10 17 18 21 24
r36 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r37 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r38 15 18 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r39 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r40 14 17 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r41 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r42 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r43 12 14 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.15
+ $Y2=0
r44 10 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r45 10 24 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r46 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r47 6 8 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.32
r48 1 8 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.785 $Y2=0.32
.ends


* File: sky130_fd_sc_hd__a2111o_2.spice
* Created: Thu Aug 27 13:58:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111o_2.spice.pex"
.subckt sky130_fd_sc_hd__a2111o_2  VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_A_86_235#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.18525 PD=0.93 PS=1.87 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75000.2
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1004_d N_A_86_235#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.290875 PD=0.93 PS=1.545 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1008 N_A_86_235#_M1008_d N_D1_M1008_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.290875 PD=0.93 PS=1.545 NRD=0 NRS=56.76 M=1 R=4.33333 SA=75001.7
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_C1_M1011_g N_A_86_235#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.091 PD=1.025 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1001 N_A_86_235#_M1001_d N_B1_M1001_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.121875 PD=0.985 PS=1.025 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.6 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1013 A_715_47# N_A1_M1013_g N_A_86_235#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.108875 PD=1.04 PS=0.985 NRD=25.836 NRS=10.152 M=1 R=4.33333
+ SA=75003.1 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g A_715_47# VNB NSHORT L=0.15 W=0.65 AD=0.221
+ AS=0.12675 PD=1.98 PS=1.04 NRD=13.836 NRS=25.836 M=1 R=4.33333 SA=75003.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_86_235#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A_86_235#_M1012_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 A_427_297# N_D1_M1002_g N_A_86_235#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.41 PD=1.21 PS=2.82 NRD=9.8303 NRS=28.565 M=1 R=6.66667
+ SA=75000.3 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1006 A_499_297# N_C1_M1006_g A_427_297# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.105 PD=1.39 PS=1.21 NRD=27.5603 NRS=9.8303 M=1 R=6.66667 SA=75000.7
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1010 N_A_607_297#_M1010_d N_B1_M1010_g A_499_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=11.8003 NRS=27.5603 M=1 R=6.66667
+ SA=75001.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_607_297#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=7.8603 NRS=9.8303 M=1 R=6.66667
+ SA=75001.8 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_A_607_297#_M1007_d N_A2_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.195 PD=2.53 PS=1.39 NRD=0 NRS=13.7703 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_73 VPB 0 1.96852e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a2111o_2.spice.SKY130_FD_SC_HD__A2111O_2.pxi"
*
.ends
*
*

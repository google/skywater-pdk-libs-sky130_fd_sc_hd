* File: sky130_fd_sc_hd__a41oi_1.spice.SKY130_FD_SC_HD__A41OI_1.pxi
* Created: Thu Aug 27 14:06:22 2020
* 
x_PM_SKY130_FD_SC_HD__A41OI_1%B1 N_B1_M1008_g N_B1_M1006_g B1 B1 N_B1_c_51_n
+ N_B1_c_52_n PM_SKY130_FD_SC_HD__A41OI_1%B1
x_PM_SKY130_FD_SC_HD__A41OI_1%A4 N_A4_M1000_g N_A4_c_79_n N_A4_M1009_g A4 A4
+ N_A4_c_81_n PM_SKY130_FD_SC_HD__A41OI_1%A4
x_PM_SKY130_FD_SC_HD__A41OI_1%A3 N_A3_M1007_g N_A3_M1005_g A3 A3 A3 N_A3_c_118_n
+ N_A3_c_119_n PM_SKY130_FD_SC_HD__A41OI_1%A3
x_PM_SKY130_FD_SC_HD__A41OI_1%A2 N_A2_M1001_g N_A2_M1002_g A2 A2 A2 N_A2_c_159_n
+ N_A2_c_160_n PM_SKY130_FD_SC_HD__A41OI_1%A2
x_PM_SKY130_FD_SC_HD__A41OI_1%A1 N_A1_c_200_n N_A1_M1004_g N_A1_M1003_g A1 A1
+ N_A1_c_201_n N_A1_c_202_n PM_SKY130_FD_SC_HD__A41OI_1%A1
x_PM_SKY130_FD_SC_HD__A41OI_1%Y N_Y_M1008_s N_Y_M1004_d N_Y_M1006_s N_Y_c_233_n
+ N_Y_c_236_n N_Y_c_249_n N_Y_c_245_n N_Y_c_227_n N_Y_c_255_n Y Y Y N_Y_c_229_n
+ Y PM_SKY130_FD_SC_HD__A41OI_1%Y
x_PM_SKY130_FD_SC_HD__A41OI_1%A_109_297# N_A_109_297#_M1006_d
+ N_A_109_297#_M1005_d N_A_109_297#_M1003_d N_A_109_297#_c_288_n
+ N_A_109_297#_c_290_n N_A_109_297#_c_291_n N_A_109_297#_c_310_p
+ N_A_109_297#_c_298_n N_A_109_297#_c_304_n N_A_109_297#_c_319_p
+ N_A_109_297#_c_301_n PM_SKY130_FD_SC_HD__A41OI_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A41OI_1%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_c_329_n
+ N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n VPWR N_VPWR_c_333_n
+ N_VPWR_c_334_n N_VPWR_c_328_n N_VPWR_c_336_n PM_SKY130_FD_SC_HD__A41OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A41OI_1%VGND N_VGND_M1008_d N_VGND_c_379_n VGND
+ N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n VGND
+ PM_SKY130_FD_SC_HD__A41OI_1%VGND
cc_1 VNB B1 0.00435769f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_2 VNB N_B1_c_51_n 0.0285048f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_3 VNB N_B1_c_52_n 0.0209454f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=0.995
cc_4 VNB N_A4_c_79_n 0.0185554f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_5 VNB A4 0.00578139f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_6 VNB N_A4_c_81_n 0.0190644f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_7 VNB A3 0.00389447f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_A3_c_118_n 0.0214994f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=0.995
cc_9 VNB N_A3_c_119_n 0.0162759f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_10 VNB A2 0.00391785f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_11 VNB N_A2_c_159_n 0.0223731f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=0.995
cc_12 VNB N_A2_c_160_n 0.0168429f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_13 VNB N_A1_c_200_n 0.0234935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A1_c_201_n 0.0374287f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=0.995
cc_15 VNB N_A1_c_202_n 0.0165274f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.325
cc_16 VNB N_Y_c_227_n 0.00720662f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.53
cc_17 VNB Y 0.0127532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_229_n 0.0255445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_328_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_379_n 0.00517457f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_21 VNB N_VGND_c_380_n 0.0571348f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_22 VNB N_VGND_c_381_n 0.18244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_382_n 0.0246618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_B1_M1006_g 0.0228129f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_25 VPB B1 0.00111708f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_26 VPB N_B1_c_51_n 0.00758906f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_27 VPB N_A4_M1000_g 0.0202357f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_28 VPB A4 0.00249512f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_29 VPB N_A4_c_81_n 0.00443649f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_30 VPB N_A3_M1005_g 0.0191547f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_31 VPB A3 0.00232601f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_32 VPB N_A3_c_118_n 0.00468956f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=0.995
cc_33 VPB N_A2_M1002_g 0.019282f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_34 VPB A2 0.0028135f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_35 VPB N_A2_c_159_n 0.00476865f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=0.995
cc_36 VPB N_A1_M1003_g 0.023744f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A1_c_201_n 0.0102155f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=0.995
cc_38 VPB N_A1_c_202_n 0.00809613f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=1.325
cc_39 VPB Y 0.0163973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_Y_c_229_n 0.0230268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB Y 0.0065071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_329_n 0.00562862f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_43 VPB N_VPWR_c_330_n 0.00562936f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_44 VPB N_VPWR_c_331_n 0.0203824f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=1.325
cc_45 VPB N_VPWR_c_332_n 0.00631792f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_46 VPB N_VPWR_c_333_n 0.031482f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.53
cc_47 VPB N_VPWR_c_334_n 0.0204309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_328_n 0.0455315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_336_n 0.00631792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 N_B1_M1006_g N_A4_M1000_g 0.0308234f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_51 N_B1_c_52_n N_A4_c_79_n 0.0190742f $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_52 N_B1_M1006_g A4 4.80108e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_53 B1 A4 0.0467526f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_54 N_B1_c_51_n A4 0.00102893f $X=0.625 $Y=1.16 $X2=0 $Y2=0
cc_55 B1 N_A4_c_81_n 0.00227893f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_56 N_B1_c_51_n N_A4_c_81_n 0.0214015f $X=0.625 $Y=1.16 $X2=0 $Y2=0
cc_57 B1 N_Y_c_233_n 0.0170065f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_58 N_B1_c_51_n N_Y_c_233_n 0.00125782f $X=0.625 $Y=1.16 $X2=0 $Y2=0
cc_59 N_B1_c_52_n N_Y_c_233_n 0.0178575f $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_60 N_B1_c_52_n N_Y_c_236_n 6.99813e-19 $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_61 N_B1_M1006_g Y 0.00466652f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_62 B1 N_Y_c_229_n 0.0439433f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_63 N_B1_c_52_n N_Y_c_229_n 0.0186511f $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_64 N_B1_M1006_g Y 0.00319579f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_65 B1 N_A_109_297#_M1006_d 0.00405343f $X=0.61 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_66 B1 N_A_109_297#_c_288_n 0.0152156f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_67 N_B1_c_51_n N_A_109_297#_c_288_n 6.20416e-19 $X=0.625 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B1_M1006_g N_VPWR_c_333_n 0.00542953f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 N_B1_M1006_g N_VPWR_c_328_n 0.0110323f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_70 N_B1_c_52_n N_VGND_c_379_n 0.00619328f $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_71 N_B1_c_52_n N_VGND_c_381_n 0.00724497f $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B1_c_52_n N_VGND_c_382_n 0.00422112f $X=0.577 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A4_M1000_g N_A3_M1005_g 0.0307726f $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_74 A4 N_A3_M1005_g 0.00117514f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A4_M1000_g A3 9.79093e-19 $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A4_c_79_n A3 0.00373303f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_77 A4 A3 0.0464786f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A4_c_81_n A3 0.00110247f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_79 A4 N_A3_c_118_n 0.00114173f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A4_c_81_n N_A3_c_118_n 0.0181138f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A4_c_79_n N_A3_c_119_n 0.0293515f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A4_c_79_n N_Y_c_233_n 0.0107279f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_83 A4 N_Y_c_233_n 0.0184065f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A4_c_81_n N_Y_c_233_n 5.24803e-19 $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A4_c_79_n N_Y_c_236_n 0.00451172f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A4_c_79_n N_Y_c_245_n 0.00543517f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A4_M1000_g N_A_109_297#_c_290_n 0.0070123f $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A4_M1000_g N_A_109_297#_c_291_n 0.0132426f $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_89 A4 N_A_109_297#_c_291_n 0.016564f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A4_c_81_n N_A_109_297#_c_291_n 3.37823e-19 $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_91 A4 N_VPWR_M1000_d 0.00258719f $X=1.07 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_92 N_A4_M1000_g N_VPWR_c_329_n 0.00345703f $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A4_M1000_g N_VPWR_c_333_n 0.00434333f $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A4_M1000_g N_VPWR_c_328_n 0.00652115f $X=1.045 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A4_c_79_n N_VGND_c_379_n 0.0060603f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A4_c_79_n N_VGND_c_380_n 0.00399631f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A4_c_79_n N_VGND_c_381_n 0.00626591f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A3_M1005_g N_A2_M1002_g 0.0224765f $X=1.605 $Y=1.985 $X2=0 $Y2=0
cc_99 A3 N_A2_M1002_g 5.6481e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A3_M1005_g A2 0.0011506f $X=1.605 $Y=1.985 $X2=0 $Y2=0
cc_101 A3 A2 0.0572068f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_102 N_A3_c_118_n A2 0.00210141f $X=1.615 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A3_c_119_n A2 8.1192e-19 $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_104 A3 N_A2_c_159_n 3.28462e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A3_c_118_n N_A2_c_159_n 0.0170396f $X=1.615 $Y=1.16 $X2=0 $Y2=0
cc_106 A3 N_A2_c_160_n 3.91932e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_107 N_A3_c_119_n N_A2_c_160_n 0.0377808f $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_108 A3 N_Y_c_233_n 0.00239414f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_109 N_A3_c_119_n N_Y_c_233_n 0.00375247f $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A3_c_119_n N_Y_c_236_n 0.00291437f $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_111 A3 N_Y_c_249_n 0.0066556f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_112 N_A3_c_118_n N_Y_c_249_n 7.23908e-19 $X=1.615 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A3_c_119_n N_Y_c_249_n 0.0111389f $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A3_M1005_g N_A_109_297#_c_291_n 0.0107643f $X=1.605 $Y=1.985 $X2=0
+ $Y2=0
cc_115 A3 N_A_109_297#_c_291_n 0.0108789f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_116 N_A3_c_118_n N_A_109_297#_c_291_n 7.31249e-19 $X=1.615 $Y=1.16 $X2=0
+ $Y2=0
cc_117 A3 N_VPWR_M1000_d 0.0018094f $X=1.53 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_118 N_A3_M1005_g N_VPWR_c_329_n 0.00631231f $X=1.605 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A3_M1005_g N_VPWR_c_331_n 0.00435108f $X=1.605 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A3_M1005_g N_VPWR_c_328_n 0.00642518f $X=1.605 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A3_c_119_n N_VGND_c_380_n 0.00366111f $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A3_c_119_n N_VGND_c_381_n 0.00562591f $X=1.615 $Y=0.995 $X2=0 $Y2=0
cc_123 A3 A_236_47# 0.00159995f $X=1.53 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_124 A2 N_A1_c_200_n 0.00417243f $X=1.99 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_125 N_A2_c_160_n N_A1_c_200_n 0.0246512f $X=2.125 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_126 N_A2_M1002_g N_A1_M1003_g 0.0286719f $X=2.065 $Y=1.985 $X2=0 $Y2=0
cc_127 A2 N_A1_M1003_g 0.00349754f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_128 A2 N_A1_c_201_n 0.00138802f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_129 N_A2_c_159_n N_A1_c_201_n 0.0136914f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_130 A2 N_A1_c_202_n 0.0188964f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_131 N_A2_c_159_n N_A1_c_202_n 9.30906e-19 $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_132 A2 N_Y_c_249_n 0.00923588f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_133 N_A2_c_159_n N_Y_c_249_n 0.00148654f $X=2.125 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A2_c_160_n N_Y_c_249_n 0.0114751f $X=2.125 $Y=0.995 $X2=0 $Y2=0
cc_135 A2 N_Y_c_255_n 0.00174707f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_136 N_A2_c_160_n N_Y_c_255_n 0.00137739f $X=2.125 $Y=0.995 $X2=0 $Y2=0
cc_137 A2 N_A_109_297#_M1005_d 0.00203449f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_138 N_A2_M1002_g N_A_109_297#_c_298_n 0.0108264f $X=2.065 $Y=1.985 $X2=0
+ $Y2=0
cc_139 A2 N_A_109_297#_c_298_n 0.0119433f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_140 N_A2_c_159_n N_A_109_297#_c_298_n 0.00149472f $X=2.125 $Y=1.16 $X2=0
+ $Y2=0
cc_141 A2 N_A_109_297#_c_301_n 0.00334593f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_142 A2 N_VPWR_M1002_d 0.00287622f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_143 N_A2_M1002_g N_VPWR_c_330_n 0.00634039f $X=2.065 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A2_M1002_g N_VPWR_c_331_n 0.00435108f $X=2.065 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A2_M1002_g N_VPWR_c_328_n 0.00644211f $X=2.065 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A2_c_160_n N_VGND_c_380_n 0.00366111f $X=2.125 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A2_c_160_n N_VGND_c_381_n 0.00578162f $X=2.125 $Y=0.995 $X2=0 $Y2=0
cc_148 A2 A_336_47# 0.00172874f $X=1.99 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_149 A2 A_428_47# 0.00204636f $X=1.99 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_150 N_A1_c_200_n N_Y_c_249_n 0.0110597f $X=2.64 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_200_n N_Y_c_255_n 0.00904309f $X=2.64 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_201_n N_Y_c_255_n 0.00316009f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A1_c_202_n N_Y_c_255_n 0.0182076f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A1_c_202_n N_A_109_297#_M1003_d 0.0149832f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A1_M1003_g N_A_109_297#_c_298_n 0.0153222f $X=2.64 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A1_c_201_n N_A_109_297#_c_304_n 0.00130134f $X=2.865 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A1_c_202_n N_A_109_297#_c_304_n 0.0166084f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A1_M1003_g N_VPWR_c_330_n 0.00334605f $X=2.64 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A1_M1003_g N_VPWR_c_334_n 0.00435108f $X=2.64 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A1_M1003_g N_VPWR_c_328_n 0.00722573f $X=2.64 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A1_c_200_n N_VGND_c_380_n 0.00366071f $X=2.64 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A1_c_200_n N_VGND_c_381_n 0.00665943f $X=2.64 $Y=0.995 $X2=0 $Y2=0
cc_163 Y N_VPWR_c_333_n 0.0170261f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_164 N_Y_M1006_s N_VPWR_c_328_n 0.00211564f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_165 Y N_VPWR_c_328_n 0.0123418f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_166 N_Y_c_233_n N_VGND_M1008_d 0.0138191f $X=1.12 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_167 N_Y_c_233_n N_VGND_c_379_n 0.0248651f $X=1.12 $Y=0.7 $X2=0 $Y2=0
cc_168 N_Y_c_245_n N_VGND_c_379_n 0.0123605f $X=1.29 $Y=0.38 $X2=0 $Y2=0
cc_169 N_Y_c_233_n N_VGND_c_380_n 0.00253538f $X=1.12 $Y=0.7 $X2=0 $Y2=0
cc_170 N_Y_c_249_n N_VGND_c_380_n 0.063522f $X=2.685 $Y=0.38 $X2=0 $Y2=0
cc_171 N_Y_c_245_n N_VGND_c_380_n 0.00769612f $X=1.29 $Y=0.38 $X2=0 $Y2=0
cc_172 N_Y_c_255_n N_VGND_c_380_n 0.0165116f $X=2.85 $Y=0.38 $X2=0 $Y2=0
cc_173 N_Y_M1008_s N_VGND_c_381_n 0.00227275f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_174 N_Y_M1004_d N_VGND_c_381_n 0.00545098f $X=2.715 $Y=0.235 $X2=0 $Y2=0
cc_175 N_Y_c_233_n N_VGND_c_381_n 0.0127494f $X=1.12 $Y=0.7 $X2=0 $Y2=0
cc_176 N_Y_c_249_n N_VGND_c_381_n 0.0487326f $X=2.685 $Y=0.38 $X2=0 $Y2=0
cc_177 N_Y_c_245_n N_VGND_c_381_n 0.00607559f $X=1.29 $Y=0.38 $X2=0 $Y2=0
cc_178 N_Y_c_227_n N_VGND_c_381_n 4.57985e-19 $X=0.225 $Y=0.7 $X2=0 $Y2=0
cc_179 N_Y_c_255_n N_VGND_c_381_n 0.012143f $X=2.85 $Y=0.38 $X2=0 $Y2=0
cc_180 Y N_VGND_c_381_n 0.00960102f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_181 N_Y_c_233_n N_VGND_c_382_n 0.00383395f $X=1.12 $Y=0.7 $X2=0 $Y2=0
cc_182 Y N_VGND_c_382_n 0.0147961f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_183 N_Y_c_233_n A_236_47# 0.00417428f $X=1.12 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_184 N_Y_c_236_n A_236_47# 0.00180838f $X=1.205 $Y=0.615 $X2=-0.19 $Y2=-0.24
cc_185 N_Y_c_249_n A_236_47# 0.00872992f $X=2.685 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_186 N_Y_c_245_n A_236_47# 5.59311e-19 $X=1.29 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_187 N_Y_c_249_n A_336_47# 0.00816103f $X=2.685 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_188 N_Y_c_249_n A_428_47# 0.0141986f $X=2.685 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_189 N_A_109_297#_c_291_n N_VPWR_M1000_d 0.0129209f $X=1.76 $Y=1.93 $X2=0.47
+ $Y2=0.995
cc_190 N_A_109_297#_c_298_n N_VPWR_M1002_d 0.0144132f $X=2.765 $Y=1.93 $X2=0.47
+ $Y2=0.56
cc_191 N_A_109_297#_c_290_n N_VPWR_c_329_n 0.0153186f $X=0.76 $Y=2.3 $X2=0.61
+ $Y2=1.445
cc_192 N_A_109_297#_c_291_n N_VPWR_c_329_n 0.0201519f $X=1.76 $Y=1.93 $X2=0.61
+ $Y2=1.445
cc_193 N_A_109_297#_c_310_p N_VPWR_c_329_n 0.0132577f $X=1.845 $Y=2.3 $X2=0.61
+ $Y2=1.445
cc_194 N_A_109_297#_c_310_p N_VPWR_c_330_n 0.014102f $X=1.845 $Y=2.3 $X2=0.625
+ $Y2=1.16
cc_195 N_A_109_297#_c_298_n N_VPWR_c_330_n 0.0216336f $X=2.765 $Y=1.93 $X2=0.625
+ $Y2=1.16
cc_196 N_A_109_297#_c_291_n N_VPWR_c_331_n 0.00368641f $X=1.76 $Y=1.93 $X2=0.577
+ $Y2=1.325
cc_197 N_A_109_297#_c_310_p N_VPWR_c_331_n 0.0117342f $X=1.845 $Y=2.3 $X2=0.577
+ $Y2=1.325
cc_198 N_A_109_297#_c_298_n N_VPWR_c_331_n 0.00330939f $X=2.765 $Y=1.93
+ $X2=0.577 $Y2=1.325
cc_199 N_A_109_297#_c_290_n N_VPWR_c_333_n 0.0171158f $X=0.76 $Y=2.3 $X2=0.66
+ $Y2=1.53
cc_200 N_A_109_297#_c_291_n N_VPWR_c_333_n 0.00357266f $X=1.76 $Y=1.93 $X2=0.66
+ $Y2=1.53
cc_201 N_A_109_297#_c_298_n N_VPWR_c_334_n 0.00265435f $X=2.765 $Y=1.93 $X2=0
+ $Y2=0
cc_202 N_A_109_297#_c_319_p N_VPWR_c_334_n 0.0171158f $X=2.85 $Y=2.3 $X2=0 $Y2=0
cc_203 N_A_109_297#_M1006_d N_VPWR_c_328_n 0.00577035f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_A_109_297#_M1005_d N_VPWR_c_328_n 0.00310215f $X=1.68 $Y=1.485 $X2=0
+ $Y2=0
cc_205 N_A_109_297#_M1003_d N_VPWR_c_328_n 0.00568078f $X=2.715 $Y=1.485 $X2=0
+ $Y2=0
cc_206 N_A_109_297#_c_290_n N_VPWR_c_328_n 0.00952784f $X=0.76 $Y=2.3 $X2=0
+ $Y2=0
cc_207 N_A_109_297#_c_291_n N_VPWR_c_328_n 0.0155097f $X=1.76 $Y=1.93 $X2=0
+ $Y2=0
cc_208 N_A_109_297#_c_310_p N_VPWR_c_328_n 0.00645434f $X=1.845 $Y=2.3 $X2=0
+ $Y2=0
cc_209 N_A_109_297#_c_298_n N_VPWR_c_328_n 0.0132928f $X=2.765 $Y=1.93 $X2=0
+ $Y2=0
cc_210 N_A_109_297#_c_319_p N_VPWR_c_328_n 0.00952784f $X=2.85 $Y=2.3 $X2=0
+ $Y2=0
cc_211 N_VGND_c_381_n A_236_47# 0.00284162f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_212 N_VGND_c_381_n A_336_47# 0.00251719f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_213 N_VGND_c_381_n A_428_47# 0.00346192f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__or2_4.pex.spice
* Created: Tue Sep  1 19:27:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR2_4%B 1 3 6 8 9 17
r30 16 17 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.53
+ $Y2=1.16
r31 13 16 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r32 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r33 8 9 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=1.16
r34 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.325
+ $X2=0.53 $Y2=1.16
r35 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.53 $Y=1.325 $X2=0.53
+ $Y2=1.985
r36 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_4%A 3 6 8 11 13
c34 11 0 2.05872e-19 $X=0.95 $Y=1.16
r35 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=1.325
r36 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r38 8 12 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=0.95 $Y2=1.16
r39 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.56 $X2=0.89
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_4%A_35_297# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 41 44 45 47 48 51 55 56 66
c126 48 0 1.69595e-19 $X=1.512 $Y=1.495
c127 47 0 1.40228e-19 $X=1.512 $Y=1.245
c128 44 0 1.02064e-19 $X=0.605 $Y=1.495
r129 63 64 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=2.235 $Y2=1.16
r130 59 63 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.575 $Y=1.16
+ $X2=1.815 $Y2=1.16
r131 59 60 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.575 $Y=1.16
+ $X2=1.395 $Y2=1.16
r132 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.16 $X2=1.575 $Y2=1.16
r133 52 66 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.655 $Y2=1.16
r134 52 64 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.235 $Y2=1.16
r135 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=1.16 $X2=2.255 $Y2=1.16
r136 49 58 3.77704 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.512 $Y2=1.16
r137 49 51 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=2.255 $Y2=1.16
r138 47 58 3.11697 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.512 $Y=1.245
+ $X2=1.512 $Y2=1.16
r139 47 48 13.5255 $w=2.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.512 $Y=1.245
+ $X2=1.512 $Y2=1.495
r140 46 55 3.05049 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=0.695 $Y=1.58
+ $X2=0.425 $Y2=1.58
r141 45 48 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=1.41 $Y=1.58
+ $X2=1.512 $Y2=1.495
r142 45 46 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.41 $Y=1.58
+ $X2=0.695 $Y2=1.58
r143 44 55 3.46198 $w=2.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.425 $Y2=1.58
r144 44 56 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.605 $Y2=0.825
r145 39 56 8.12648 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.66
+ $X2=0.68 $Y2=0.825
r146 39 41 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.68 $Y=0.66
+ $X2=0.68 $Y2=0.4
r147 35 55 3.46198 $w=2.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.335 $Y=1.665
+ $X2=0.425 $Y2=1.58
r148 35 37 20.3278 $w=3.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.335 $Y=1.665
+ $X2=0.335 $Y2=2.3
r149 31 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.325
+ $X2=2.655 $Y2=1.16
r150 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.655 $Y=1.325
+ $X2=2.655 $Y2=1.985
r151 28 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=0.995
+ $X2=2.655 $Y2=1.16
r152 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.655 $Y=0.995
+ $X2=2.655 $Y2=0.56
r153 24 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.325
+ $X2=2.235 $Y2=1.16
r154 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.235 $Y=1.325
+ $X2=2.235 $Y2=1.985
r155 21 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=0.995
+ $X2=2.235 $Y2=1.16
r156 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.235 $Y=0.995
+ $X2=2.235 $Y2=0.56
r157 17 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.16
r158 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.985
r159 14 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r160 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=0.56
r161 10 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.16
r162 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.985
r163 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=1.16
r164 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=0.56
r165 2 55 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.485 $X2=0.32 $Y2=1.62
r166 2 37 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.485 $X2=0.32 $Y2=2.3
r167 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_4%VPWR 1 2 3 12 16 20 23 24 26 27 28 37 43 44
c49 3 0 1.57649e-19 $X=2.73 $Y=1.485
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 41 43 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 40 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 37 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.865 $Y2=2.72
r55 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.78 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 36 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r58 32 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 28 32 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 26 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=2.025 $Y2=2.72
r63 25 39 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=2.72
+ $X2=2.025 $Y2=2.72
r65 23 31 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=2.72 $X2=0.69
+ $Y2=2.72
r66 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=2.72
+ $X2=1.145 $Y2=2.72
r67 22 35 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.72
+ $X2=1.145 $Y2=2.72
r69 18 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.635
+ $X2=2.865 $Y2=2.72
r70 18 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.865 $Y=2.635
+ $X2=2.865 $Y2=2
r71 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.635
+ $X2=2.025 $Y2=2.72
r72 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.025 $Y=2.635
+ $X2=2.025 $Y2=2.34
r73 10 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.72
r74 10 12 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.01
r75 3 20 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=1.485 $X2=2.865 $Y2=2
r76 2 16 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.025 $Y2=2.34
r77 1 12 300 $w=1.7e-07 $l=6.08379e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.145 $Y2=2.01
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_4%X 1 2 3 4 15 19 20 21 25 27 28 31 33 35 38 39
+ 42 44 47
c90 44 0 1.57649e-19 $X=2.995 $Y=1.53
c91 3 0 1.03951e-19 $X=1.47 $Y=1.485
r92 44 47 2.61083 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.962 $Y=1.58
+ $X2=2.962 $Y2=1.495
r93 44 47 0.835104 $w=3.43e-07 $l=2.5e-08 $layer=LI1_cond $X=2.962 $Y=1.47
+ $X2=2.962 $Y2=1.495
r94 43 44 18.8733 $w=3.43e-07 $l=5.65e-07 $layer=LI1_cond $X=2.962 $Y=0.905
+ $X2=2.962 $Y2=1.47
r95 36 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.58
+ $X2=2.445 $Y2=1.58
r96 35 44 5.28309 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.79 $Y=1.58
+ $X2=2.962 $Y2=1.58
r97 35 36 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.79 $Y=1.58
+ $X2=2.61 $Y2=1.58
r98 34 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=0.82
+ $X2=2.445 $Y2=0.82
r99 33 43 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=2.79 $Y=0.82
+ $X2=2.962 $Y2=0.905
r100 33 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.79 $Y=0.82
+ $X2=2.61 $Y2=0.82
r101 29 42 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=2.005
+ $X2=2.445 $Y2=1.92
r102 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.445 $Y=2.005
+ $X2=2.445 $Y2=2.34
r103 28 42 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.835
+ $X2=2.445 $Y2=1.92
r104 27 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.665
+ $X2=2.445 $Y2=1.58
r105 27 28 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.445 $Y=1.665
+ $X2=2.445 $Y2=1.835
r106 23 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0.735
+ $X2=2.445 $Y2=0.82
r107 23 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.445 $Y=0.735
+ $X2=2.445 $Y2=0.4
r108 22 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=1.92
+ $X2=1.605 $Y2=1.92
r109 21 42 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=1.92
+ $X2=2.445 $Y2=1.92
r110 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.28 $Y=1.92
+ $X2=1.77 $Y2=1.92
r111 19 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=0.82
+ $X2=2.445 $Y2=0.82
r112 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.28 $Y=0.82
+ $X2=1.77 $Y2=0.82
r113 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.605 $Y=0.735
+ $X2=1.77 $Y2=0.82
r114 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.605 $Y=0.735
+ $X2=1.605 $Y2=0.4
r115 4 41 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.485 $X2=2.445 $Y2=1.66
r116 4 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.485 $X2=2.445 $Y2=2.34
r117 3 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=1.485 $X2=1.605 $Y2=2
r118 2 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.31
+ $Y=0.235 $X2=2.445 $Y2=0.4
r119 1 15 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.47
+ $Y=0.235 $X2=1.605 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__OR2_4%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34 35 44
+ 53 54
r59 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r60 51 53 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.99
+ $Y2=0
r61 47 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r62 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r63 44 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.865
+ $Y2=0
r64 44 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.53
+ $Y2=0
r65 43 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r66 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r67 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r68 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 37 49 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r70 37 39 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r71 35 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r72 35 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 33 42 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.61
+ $Y2=0
r74 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.025
+ $Y2=0
r75 32 46 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.53
+ $Y2=0
r76 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.025
+ $Y2=0
r77 30 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.69
+ $Y2=0
r78 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0 $X2=1.145
+ $Y2=0
r79 29 42 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.61
+ $Y2=0
r80 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.145
+ $Y2=0
r81 25 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0
r82 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0.4
r83 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r84 21 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.4
r85 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r86 17 19 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.575
r87 13 49 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r88 13 15 15.606 $w=2.38e-07 $l=3.25e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.41
r89 4 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.235 $X2=2.865 $Y2=0.4
r90 3 23 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.235 $X2=2.025 $Y2=0.4
r91 2 19 182 $w=1.7e-07 $l=4.20476e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.145 $Y2=0.575
r92 1 15 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.41
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__nor2_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__nor2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 3.530000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.800000 1.075000 6.540000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 7.275000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.895000 0.255000 4.225000 0.725000 ;
        RECT 3.935000 1.445000 7.275000 1.615000 ;
        RECT 3.935000 1.615000 4.185000 2.125000 ;
        RECT 4.735000 0.255000 5.065000 0.725000 ;
        RECT 4.775000 1.615000 5.025000 2.125000 ;
        RECT 5.575000 0.255000 5.905000 0.725000 ;
        RECT 5.615000 1.615000 5.865000 2.125000 ;
        RECT 6.415000 0.255000 6.745000 0.725000 ;
        RECT 6.455000 1.615000 6.705000 2.125000 ;
        RECT 6.710000 0.905000 7.275000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 3.765000 1.665000 ;
      RECT 0.090000  1.665000 0.405000 2.465000 ;
      RECT 0.575000  1.835000 0.825000 2.635000 ;
      RECT 0.995000  1.665000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.835000 1.665000 2.635000 ;
      RECT 1.835000  1.665000 2.085000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.835000 2.505000 2.635000 ;
      RECT 2.675000  1.665000 2.925000 2.465000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.835000 3.345000 2.635000 ;
      RECT 3.515000  1.665000 3.765000 2.295000 ;
      RECT 3.515000  2.295000 7.125000 2.465000 ;
      RECT 3.555000  0.085000 3.725000 0.555000 ;
      RECT 4.355000  1.785000 4.605000 2.295000 ;
      RECT 4.395000  0.085000 4.565000 0.555000 ;
      RECT 5.195000  1.785000 5.445000 2.295000 ;
      RECT 5.235000  0.085000 5.405000 0.555000 ;
      RECT 6.035000  1.785000 6.285000 2.295000 ;
      RECT 6.075000  0.085000 6.245000 0.555000 ;
      RECT 6.875000  1.785000 7.125000 2.295000 ;
      RECT 6.915000  0.085000 7.205000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_8

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o22ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.075000 4.165000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.075000 3.225000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 0.985000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.075000 1.925000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 2.340000 0.905000 ;
        RECT 1.375000 0.645000 1.705000 0.725000 ;
        RECT 1.415000 1.445000 3.065000 1.625000 ;
        RECT 1.415000 1.625000 1.665000 2.125000 ;
        RECT 2.095000 0.905000 2.340000 1.445000 ;
        RECT 2.815000 1.625000 3.065000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 2.855000  0.085000 3.025000 0.555000 ;
        RECT 3.695000  0.085000 3.865000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.575000 1.795000 0.825000 2.635000 ;
        RECT 3.655000 1.795000 3.905000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.305000 2.680000 0.475000 ;
      RECT 0.090000 0.475000 0.365000 0.905000 ;
      RECT 0.150000 1.455000 1.245000 1.625000 ;
      RECT 0.150000 1.625000 0.405000 2.465000 ;
      RECT 0.995000 1.625000 1.245000 2.295000 ;
      RECT 0.995000 2.295000 2.085000 2.465000 ;
      RECT 1.835000 1.795000 2.085000 2.295000 ;
      RECT 2.395000 1.795000 2.645000 2.295000 ;
      RECT 2.395000 2.295000 3.485000 2.465000 ;
      RECT 2.510000 0.475000 2.680000 0.725000 ;
      RECT 2.510000 0.725000 4.365000 0.905000 ;
      RECT 3.195000 0.255000 3.525000 0.725000 ;
      RECT 3.235000 1.455000 4.330000 1.625000 ;
      RECT 3.235000 1.625000 3.485000 2.295000 ;
      RECT 4.035000 0.255000 4.365000 0.725000 ;
      RECT 4.075000 1.625000 4.330000 2.465000 ;
  END
END sky130_fd_sc_hd__o22ai_2
END LIBRARY

* File: sky130_fd_sc_hd__sdfxtp_1.pex.spice
* Created: Tue Sep  1 19:31:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%CLK 1 2 3 5 6 8 11 13
c42 1 0 2.71124e-20 $X=0.31 $Y=1.325
r43 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.475 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=1.74
+ $X2=0.475 $Y2=2.135
r47 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r50 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_27_47# 1 2 9 13 17 19 20 25 29 31 35 39
+ 43 44 45 49 50 52 55 56 57 58 59 60 67 69 75 78 80 82 86
c247 86 0 1.77381e-19 $X=6.665 $Y=1.41
c248 57 0 1.65095e-19 $X=5.145 $Y=1.87
c249 52 0 8.70797e-20 $X=0.76 $Y=1.235
c250 50 0 1.81794e-19 $X=0.73 $Y=1.795
c251 45 0 3.29888e-20 $X=0.615 $Y=1.88
c252 29 0 4.21632e-20 $X=6.67 $Y=2.275
c253 19 0 1.57835e-19 $X=4.98 $Y=1.32
r254 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.665 $Y=1.41
+ $X2=6.665 $Y2=1.575
r255 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.665
+ $Y=1.41 $X2=6.665 $Y2=1.41
r256 82 85 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.665 $Y=1.32
+ $X2=6.665 $Y2=1.41
r257 78 81 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.74
+ $X2=5.115 $Y2=1.905
r258 78 80 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.74
+ $X2=5.115 $Y2=1.575
r259 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.74 $X2=5.115 $Y2=1.74
r260 74 75 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=0.89 $Y=1.235
+ $X2=0.895 $Y2=1.235
r261 70 86 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.675 $Y=1.87
+ $X2=6.675 $Y2=1.41
r262 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.675 $Y=1.87
+ $X2=6.675 $Y2=1.87
r263 67 79 5.68106 $w=3.53e-07 $l=1.75e-07 $layer=LI1_cond $X=5.29 $Y=1.832
+ $X2=5.115 $Y2=1.832
r264 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r265 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=1.87
+ $X2=0.725 $Y2=1.87
r266 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r267 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.53 $Y=1.87
+ $X2=6.675 $Y2=1.87
r268 59 60 1.3552 $w=1.4e-07 $l=1.095e-06 $layer=MET1_cond $X=6.53 $Y=1.87
+ $X2=5.435 $Y2=1.87
r269 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.87 $Y=1.87
+ $X2=0.725 $Y2=1.87
r270 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r271 57 58 5.29083 $w=1.4e-07 $l=4.275e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=0.87 $Y2=1.87
r272 53 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r273 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r274 50 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r275 50 52 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r276 49 56 6.0623 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=0.97
r277 49 52 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=1.235
r278 47 56 9.38461 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=0.805
+ $X2=0.712 $Y2=0.97
r279 46 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r280 45 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r281 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.35 $Y2=1.88
r282 43 47 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.712 $Y2=0.805
r283 43 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r284 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r285 37 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r286 33 35 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.315 $Y=1.245
+ $X2=7.315 $Y2=0.415
r287 32 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.8 $Y=1.32
+ $X2=6.665 $Y2=1.32
r288 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.24 $Y=1.32
+ $X2=7.315 $Y2=1.245
r289 31 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.24 $Y=1.32
+ $X2=6.8 $Y2=1.32
r290 29 87 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.67 $Y=2.275
+ $X2=6.67 $Y2=1.575
r291 25 81 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.055 $Y=2.275
+ $X2=5.055 $Y2=1.905
r292 21 80 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.055 $Y=1.395
+ $X2=5.055 $Y2=1.575
r293 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.98 $Y=1.32
+ $X2=5.055 $Y2=1.395
r294 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=4.98 $Y=1.32
+ $X2=4.67 $Y2=1.32
r295 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.595 $Y=1.245
+ $X2=4.67 $Y2=1.32
r296 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.595 $Y=1.245
+ $X2=4.595 $Y2=0.415
r297 11 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=1.235
r298 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.895 $Y=1.37
+ $X2=0.895 $Y2=2.135
r299 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r300 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r301 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r302 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%SCE 5 9 10 14 18 19 20 23 24 26 27 28 32 33
+ 37 38 41 45
c124 33 0 1.39399e-19 $X=3.15 $Y=0.93
c125 28 0 1.93564e-19 $X=3.065 $Y=0.7
c126 27 0 8.19616e-20 $X=1.99 $Y=0.7
r127 42 43 29.3768 $w=3.1e-07 $l=7.5e-08 $layer=POLY_cond $X=1.855 $Y=1.58
+ $X2=1.855 $Y2=1.655
r128 36 38 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.51
r129 36 37 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.562 $Y=0.615
+ $X2=2.562 $Y2=0.7
r130 33 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=0.93
+ $X2=3.15 $Y2=0.765
r131 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=0.93 $X2=3.15 $Y2=0.93
r132 30 32 8.69287 $w=1.83e-07 $l=1.45e-07 $layer=LI1_cond $X=3.157 $Y=0.785
+ $X2=3.157 $Y2=0.93
r133 29 37 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.65 $Y=0.7
+ $X2=2.562 $Y2=0.7
r134 28 30 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.065 $Y=0.7
+ $X2=3.157 $Y2=0.785
r135 28 29 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.065 $Y=0.7
+ $X2=2.65 $Y2=0.7
r136 27 35 8.90217 $w=2.1e-07 $l=1.57003e-07 $layer=LI1_cond $X=1.99 $Y=0.7
+ $X2=1.845 $Y2=0.725
r137 26 37 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=2.562 $Y2=0.7
r138 26 27 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.475 $Y=0.7
+ $X2=1.99 $Y2=0.7
r139 24 42 11.1686 $w=3.1e-07 $l=6e-08 $layer=POLY_cond $X=1.855 $Y=1.52
+ $X2=1.855 $Y2=1.58
r140 24 41 40.5454 $w=3.1e-07 $l=1.35e-07 $layer=POLY_cond $X=1.855 $Y=1.52
+ $X2=1.855 $Y2=1.385
r141 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.52 $X2=1.845 $Y2=1.52
r142 21 35 1.9771 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.845 $Y=0.835
+ $X2=1.845 $Y2=0.725
r143 21 23 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.845 $Y=0.835
+ $X2=1.845 $Y2=1.52
r144 20 41 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.83 $Y=0.815
+ $X2=1.83 $Y2=1.385
r145 19 20 35.9386 $w=1.7e-07 $l=8.5e-08 $layer=POLY_cond $X=1.84 $Y=0.73
+ $X2=1.84 $Y2=0.815
r146 18 45 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.21 $Y=0.445
+ $X2=3.21 $Y2=0.765
r147 12 14 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.26 $Y=1.655
+ $X2=2.26 $Y2=2.165
r148 11 42 19.7411 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.01 $Y=1.58
+ $X2=1.855 $Y2=1.58
r149 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.185 $Y=1.58
+ $X2=2.26 $Y2=1.655
r150 10 11 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.185 $Y=1.58
+ $X2=2.01 $Y2=1.58
r151 9 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.85 $Y=0.445
+ $X2=1.85 $Y2=0.73
r152 5 43 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.835 $Y=2.165
+ $X2=1.835 $Y2=1.655
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_299_47# 1 2 9 13 16 19 21 24 25 28 32 34
+ 37 38 40 42 43
c139 43 0 1.99235e-20 $X=3.185 $Y=1.47
c140 40 0 1.27981e-19 $X=2.202 $Y=1.967
c141 28 0 5.65856e-20 $X=3.135 $Y=1.86
c142 24 0 1.62582e-19 $X=2.202 $Y=1.86
c143 13 0 2.43768e-20 $X=3.125 $Y=2.165
r144 43 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.185 $Y=1.47
+ $X2=3.185 $Y2=1.635
r145 42 45 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=1.47
+ $X2=3.16 $Y2=1.635
r146 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.47 $X2=3.185 $Y2=1.47
r147 38 47 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.28 $Y=1.045
+ $X2=2.28 $Y2=0.91
r148 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.045 $X2=2.28 $Y2=1.045
r149 29 32 6.49224 $w=2.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.505 $Y=0.362
+ $X2=1.625 $Y2=0.362
r150 28 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.135 $Y=1.86
+ $X2=3.135 $Y2=1.635
r151 26 40 4.33859 $w=2.15e-07 $l=8.8e-08 $layer=LI1_cond $X=2.29 $Y=1.967
+ $X2=2.202 $Y2=1.967
r152 25 28 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.05 $Y=1.967
+ $X2=3.135 $Y2=1.86
r153 25 26 40.7375 $w=2.13e-07 $l=7.6e-07 $layer=LI1_cond $X=3.05 $Y=1.967
+ $X2=2.29 $Y2=1.967
r154 24 40 2.09329 $w=1.75e-07 $l=1.07e-07 $layer=LI1_cond $X=2.202 $Y=1.86
+ $X2=2.202 $Y2=1.967
r155 23 37 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.202 $Y=1.13
+ $X2=2.202 $Y2=1.045
r156 23 24 46.2649 $w=1.73e-07 $l=7.3e-07 $layer=LI1_cond $X=2.202 $Y=1.13
+ $X2=2.202 $Y2=1.86
r157 22 34 1.58651 $w=2.15e-07 $l=1.45e-07 $layer=LI1_cond $X=1.71 $Y=1.967
+ $X2=1.565 $Y2=1.967
r158 21 40 4.33859 $w=2.15e-07 $l=8.7e-08 $layer=LI1_cond $X=2.115 $Y=1.967
+ $X2=2.202 $Y2=1.967
r159 21 22 21.7088 $w=2.13e-07 $l=4.05e-07 $layer=LI1_cond $X=2.115 $Y=1.967
+ $X2=1.71 $Y2=1.967
r160 17 34 4.8823 $w=2.3e-07 $l=1.08e-07 $layer=LI1_cond $X=1.565 $Y=2.075
+ $X2=1.565 $Y2=1.967
r161 17 19 3.97394 $w=2.88e-07 $l=1e-07 $layer=LI1_cond $X=1.565 $Y=2.075
+ $X2=1.565 $Y2=2.175
r162 16 34 4.8823 $w=2.3e-07 $l=1.33675e-07 $layer=LI1_cond $X=1.505 $Y=1.86
+ $X2=1.565 $Y2=1.967
r163 15 29 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.505 $Y=0.465
+ $X2=1.505 $Y2=0.362
r164 15 16 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=1.505 $Y=0.465
+ $X2=1.505 $Y2=1.86
r165 13 51 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.125 $Y=2.165
+ $X2=3.125 $Y2=1.635
r166 9 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.34 $Y=0.445
+ $X2=2.34 $Y2=0.91
r167 2 19 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.845 $X2=1.625 $Y2=2.175
r168 1 32 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.625 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%D 3 7 9 12 13
r51 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.52
+ $X2=2.705 $Y2=1.355
r52 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.52 $X2=2.705 $Y2=1.52
r53 9 13 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.59 $Y=1.52
+ $X2=2.705 $Y2=1.52
r54 7 14 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.73 $Y=0.445
+ $X2=2.73 $Y2=1.355
r55 1 12 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.685
+ $X2=2.705 $Y2=1.52
r56 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.705 $Y=1.685
+ $X2=2.705 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%SCD 3 7 12 13 14 16 17 20
c56 17 0 1.63776e-19 $X=3.83 $Y=1.19
c57 14 0 5.65856e-20 $X=3.6 $Y=1.77
c58 12 0 3.56153e-19 $X=3.657 $Y=1.19
c59 3 0 1.73641e-19 $X=3.59 $Y=0.445
r60 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.665
+ $Y=1.355 $X2=3.665 $Y2=1.355
r61 17 21 4.29028 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=1.19
+ $X2=3.76 $Y2=1.355
r62 15 20 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=3.665 $Y=1.385
+ $X2=3.665 $Y2=1.355
r63 15 16 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=3.665 $Y=1.385
+ $X2=3.665 $Y2=1.52
r64 13 14 25.4904 $w=1.6e-07 $l=5.5e-08 $layer=POLY_cond $X=3.6 $Y=1.715 $X2=3.6
+ $Y2=1.77
r65 13 16 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.605 $Y=1.715
+ $X2=3.605 $Y2=1.52
r66 12 20 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.19
+ $X2=3.665 $Y2=1.355
r67 11 12 31.7529 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=3.657 $Y=1.1 $X2=3.657
+ $Y2=1.19
r68 7 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.595 $Y=2.165
+ $X2=3.595 $Y2=1.77
r69 3 11 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.59 $Y=0.445
+ $X2=3.59 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_193_47# 1 2 9 13 14 16 19 23 24 27 30 33
+ 34 38 39 41 42 43 44 47 53 60 61 62 67
c216 67 0 1.77381e-19 $X=6.895 $Y=0.87
c217 43 0 1.57835e-19 $X=6.57 $Y=0.85
r218 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.895
+ $Y=0.87 $X2=6.895 $Y2=0.87
r219 64 67 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.8 $Y=0.87
+ $X2=6.895 $Y2=0.87
r220 60 62 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.015 $Y=0.87
+ $X2=5.015 $Y2=0.705
r221 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.015
+ $Y=0.87 $X2=5.015 $Y2=0.87
r222 54 68 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=6.715 $Y=0.87
+ $X2=6.895 $Y2=0.87
r223 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.715 $Y=0.85
+ $X2=6.715 $Y2=0.85
r224 51 61 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.83 $Y=0.87
+ $X2=5.015 $Y2=0.87
r225 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0.85
+ $X2=4.83 $Y2=0.85
r226 47 76 58.6234 $w=2.08e-07 $l=1.11e-06 $layer=LI1_cond $X=1.125 $Y=0.85
+ $X2=1.125 $Y2=1.96
r227 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.125 $Y=0.85
+ $X2=1.125 $Y2=0.85
r228 44 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=0.85
+ $X2=4.83 $Y2=0.85
r229 43 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.57 $Y=0.85
+ $X2=6.715 $Y2=0.85
r230 43 44 1.97401 $w=1.4e-07 $l=1.595e-06 $layer=MET1_cond $X=6.57 $Y=0.85
+ $X2=4.975 $Y2=0.85
r231 42 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.27 $Y=0.85
+ $X2=1.125 $Y2=0.85
r232 41 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=4.83 $Y2=0.85
r233 41 42 4.22648 $w=1.4e-07 $l=3.415e-06 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=1.27 $Y2=0.85
r234 39 70 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=7.175 $Y=1.74
+ $X2=7.09 $Y2=1.74
r235 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.175
+ $Y=1.74 $X2=7.175 $Y2=1.74
r236 35 38 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.035 $Y=1.74
+ $X2=7.175 $Y2=1.74
r237 34 68 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.94 $Y=0.87
+ $X2=6.895 $Y2=0.87
r238 33 51 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=4.76 $Y=0.87 $X2=4.83
+ $Y2=0.87
r239 32 47 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.125 $Y=0.715
+ $X2=1.125 $Y2=0.85
r240 30 32 10.9884 $w=2.13e-07 $l=2.05e-07 $layer=LI1_cond $X=1.122 $Y=0.51
+ $X2=1.122 $Y2=0.715
r241 27 35 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.035 $Y=1.575
+ $X2=7.035 $Y2=1.74
r242 26 34 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.035 $Y=1.035
+ $X2=6.94 $Y2=0.87
r243 26 27 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.035 $Y=1.035
+ $X2=7.035 $Y2=1.575
r244 24 58 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.605 $Y=1.74
+ $X2=4.605 $Y2=1.875
r245 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.605
+ $Y=1.74 $X2=4.605 $Y2=1.74
r246 21 33 5.71525 $w=3.51e-07 $l=2.16852e-07 $layer=LI1_cond $X=4.64 $Y=1.035
+ $X2=4.76 $Y2=0.87
r247 21 23 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.64 $Y=1.035
+ $X2=4.64 $Y2=1.74
r248 17 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.09 $Y=1.875
+ $X2=7.09 $Y2=1.74
r249 17 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.09 $Y=1.875
+ $X2=7.09 $Y2=2.275
r250 14 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=0.705
+ $X2=6.8 $Y2=0.87
r251 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.8 $Y=0.705
+ $X2=6.8 $Y2=0.415
r252 13 62 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.075 $Y=0.415
+ $X2=5.075 $Y2=0.705
r253 9 58 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.59 $Y=2.275 $X2=4.59
+ $Y2=1.875
r254 2 76 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.815 $X2=1.105 $Y2=1.96
r255 1 30 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_1092_183# 1 2 9 13 15 18 21 23 29 30 32
+ 33 36
r95 35 36 5.54023 $w=2.61e-07 $l=3e-08 $layer=POLY_cond $X=5.535 $Y=0.93
+ $X2=5.565 $Y2=0.93
r96 32 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.365 $Y=2.3
+ $X2=6.365 $Y2=2.135
r97 27 36 24.0077 $w=2.61e-07 $l=1.3e-07 $layer=POLY_cond $X=5.695 $Y=0.93
+ $X2=5.565 $Y2=0.93
r98 26 29 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=0.93
+ $X2=5.78 $Y2=0.93
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.695
+ $Y=0.93 $X2=5.695 $Y2=0.93
r100 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=0.45
+ $X2=6.535 $Y2=0.45
r101 19 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.325 $Y=1.065
+ $X2=6.325 $Y2=0.915
r102 19 33 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.325 $Y=1.065
+ $X2=6.325 $Y2=2.135
r103 18 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.325 $Y=0.765
+ $X2=6.325 $Y2=0.915
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.325 $Y=0.535
+ $X2=6.41 $Y2=0.45
r105 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.325 $Y=0.535
+ $X2=6.325 $Y2=0.765
r106 15 30 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=0.915
+ $X2=6.325 $Y2=0.915
r107 15 29 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.24 $Y=0.915
+ $X2=5.78 $Y2=0.915
r108 11 36 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.565 $Y=0.795
+ $X2=5.565 $Y2=0.93
r109 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.565 $Y=0.795
+ $X2=5.565 $Y2=0.445
r110 7 35 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.535 $Y=1.065
+ $X2=5.535 $Y2=0.93
r111 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.535 $Y=1.065
+ $X2=5.535 $Y2=2.275
r112 2 32 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.735 $X2=6.405 $Y2=2.3
r113 1 23 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.37
+ $Y=0.235 $X2=6.535 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_933_413# 1 2 8 11 13 15 18 20 21 22 26 31
+ 33 35
c110 31 0 1.42307e-19 $X=5.355 $Y=1.315
r111 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=1.41 $X2=5.985 $Y2=1.41
r112 35 37 17.1405 $w=2.42e-07 $l=3.4e-07 $layer=LI1_cond $X=5.645 $Y=1.41
+ $X2=5.985 $Y2=1.41
r113 32 35 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=1.575
+ $X2=5.645 $Y2=1.41
r114 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.645 $Y=1.575
+ $X2=5.645 $Y2=2.19
r115 31 35 14.6198 $w=2.42e-07 $l=2.9e-07 $layer=LI1_cond $X=5.355 $Y=1.41
+ $X2=5.645 $Y2=1.41
r116 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.355 $Y=0.535
+ $X2=5.355 $Y2=1.315
r117 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.27 $Y=0.45
+ $X2=5.355 $Y2=0.535
r118 26 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.27 $Y=0.45
+ $X2=4.865 $Y2=0.45
r119 22 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.56 $Y=2.275
+ $X2=5.645 $Y2=2.19
r120 22 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.56 $Y=2.275
+ $X2=4.825 $Y2=2.275
r121 20 38 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.12 $Y=1.41
+ $X2=5.985 $Y2=1.41
r122 20 21 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.12 $Y=1.41
+ $X2=6.195 $Y2=1.41
r123 16 18 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.195 $Y=1.025
+ $X2=6.295 $Y2=1.025
r124 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.295 $Y=0.95
+ $X2=6.295 $Y2=1.025
r125 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.295 $Y=0.95
+ $X2=6.295 $Y2=0.555
r126 9 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.195 $Y=1.545
+ $X2=6.195 $Y2=1.41
r127 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.195 $Y=1.545
+ $X2=6.195 $Y2=2.11
r128 8 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.195 $Y=1.275
+ $X2=6.195 $Y2=1.41
r129 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.195 $Y=1.1
+ $X2=6.195 $Y2=1.025
r130 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.195 $Y=1.1
+ $X2=6.195 $Y2=1.275
r131 2 24 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=2.065 $X2=4.825 $Y2=2.275
r132 1 28 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.235 $X2=4.865 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_1520_315# 1 2 9 13 17 20 22 25 29 32 34
+ 37 38 41 45 46 53
c86 38 0 1.12296e-19 $X=9.15 $Y=1.16
r87 47 49 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.675 $Y=1.74
+ $X2=7.79 $Y2=1.74
r88 41 43 17.5434 $w=3.48e-07 $l=4.4e-07 $layer=LI1_cond $X=8.53 $Y=0.385
+ $X2=8.53 $Y2=0.825
r89 38 54 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=1.16
+ $X2=9.175 $Y2=1.325
r90 38 53 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=1.16
+ $X2=9.175 $Y2=0.995
r91 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.15
+ $Y=1.16 $X2=9.15 $Y2=1.16
r92 35 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.705 $Y=1.16
+ $X2=8.62 $Y2=1.16
r93 35 37 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.705 $Y=1.16
+ $X2=9.15 $Y2=1.16
r94 34 45 7.13466 $w=2.2e-07 $l=1.88348e-07 $layer=LI1_cond $X=8.62 $Y=1.575
+ $X2=8.57 $Y2=1.74
r95 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=1.325
+ $X2=8.62 $Y2=1.16
r96 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.62 $Y=1.325
+ $X2=8.62 $Y2=1.575
r97 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=0.995
+ $X2=8.62 $Y2=1.16
r98 32 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.62 $Y=0.995
+ $X2=8.62 $Y2=0.825
r99 27 45 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=1.905
+ $X2=8.57 $Y2=1.74
r100 27 29 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.57 $Y=1.905
+ $X2=8.57 $Y2=2.29
r101 25 49 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.855 $Y=1.74
+ $X2=7.79 $Y2=1.74
r102 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.855
+ $Y=1.74 $X2=7.855 $Y2=1.74
r103 22 45 0.067832 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=8.435 $Y=1.74
+ $X2=8.57 $Y2=1.74
r104 22 24 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=8.435 $Y=1.74
+ $X2=7.855 $Y2=1.74
r105 20 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.185 $Y=1.985
+ $X2=9.185 $Y2=1.325
r106 17 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.185 $Y=0.56
+ $X2=9.185 $Y2=0.995
r107 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.575
+ $X2=7.79 $Y2=1.74
r108 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.79 $Y=1.575
+ $X2=7.79 $Y2=0.445
r109 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.675 $Y=1.905
+ $X2=7.675 $Y2=1.74
r110 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.675 $Y=1.905
+ $X2=7.675 $Y2=2.275
r111 2 45 600 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=8.395
+ $Y=1.485 $X2=8.52 $Y2=1.68
r112 2 29 600 $w=1.7e-07 $l=8.65246e-07 $layer=licon1_PDIFF $count=1 $X=8.395
+ $Y=1.485 $X2=8.52 $Y2=2.29
r113 1 41 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=8.395
+ $Y=0.235 $X2=8.52 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_1349_413# 1 2 7 9 12 14 15 16 20 27 30 33
+ 34
c88 30 0 1.12296e-19 $X=8.28 $Y=1.16
c89 27 0 4.21632e-20 $X=7.515 $Y=2.165
r90 33 35 11.5578 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=7.45 $Y=1.16
+ $X2=7.45 $Y2=1.405
r91 33 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=1.16
+ $X2=7.45 $Y2=0.995
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.28
+ $Y=1.16 $X2=8.28 $Y2=1.16
r93 28 33 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.6 $Y=1.16 $X2=7.45
+ $Y2=1.16
r94 28 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.6 $Y=1.16 $X2=8.28
+ $Y2=1.16
r95 27 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.515 $Y=2.165
+ $X2=7.515 $Y2=1.405
r96 24 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.385 $Y=0.535
+ $X2=7.385 $Y2=0.995
r97 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=0.45
+ $X2=7.385 $Y2=0.535
r98 20 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.3 $Y=0.45
+ $X2=7.095 $Y2=0.45
r99 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.43 $Y=2.25
+ $X2=7.515 $Y2=2.165
r100 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.43 $Y=2.25
+ $X2=6.88 $Y2=2.25
r101 14 31 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=8.655 $Y=1.16
+ $X2=8.28 $Y2=1.16
r102 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.655 $Y=1.16
+ $X2=8.73 $Y2=1.16
r103 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=1.325
+ $X2=8.73 $Y2=1.16
r104 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.73 $Y=1.325
+ $X2=8.73 $Y2=1.985
r105 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=0.995
+ $X2=8.73 $Y2=1.16
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.73 $Y=0.995
+ $X2=8.73 $Y2=0.56
r107 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=2.065 $X2=6.88 $Y2=2.25
r108 1 22 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=6.875
+ $Y=0.235 $X2=7.095 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 52 54 59 64 86 87 90 93 96
c156 87 0 1.81794e-19 $X=9.43 $Y=2.72
c157 2 0 2.90563e-19 $X=1.91 $Y=1.845
c158 1 0 3.29888e-20 $X=0.55 $Y=1.815
r159 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r160 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r161 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r162 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r163 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r164 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r165 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r166 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r167 78 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r168 77 80 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r169 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r170 75 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r171 75 97 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r172 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r173 72 96 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=3.827 $Y2=2.72
r174 72 74 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r175 71 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r176 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r177 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r178 68 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r179 67 70 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r180 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r181 65 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.045 $Y2=2.72
r182 65 67 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.53 $Y2=2.72
r183 64 96 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.827 $Y2=2.72
r184 64 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r185 63 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r186 63 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r187 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r188 60 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=0.685 $Y2=2.72
r189 60 62 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r190 59 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=2.045 $Y2=2.72
r191 59 62 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.88 $Y=2.72
+ $X2=1.61 $Y2=2.72
r192 54 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.685 $Y2=2.72
r193 54 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r194 52 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r195 52 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r196 50 83 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.875 $Y=2.72
+ $X2=8.51 $Y2=2.72
r197 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.875 $Y=2.72
+ $X2=8.96 $Y2=2.72
r198 49 86 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.045 $Y=2.72
+ $X2=9.43 $Y2=2.72
r199 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.045 $Y=2.72
+ $X2=8.96 $Y2=2.72
r200 47 80 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.79 $Y=2.72 $X2=7.59
+ $Y2=2.72
r201 47 48 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.79 $Y=2.72
+ $X2=7.942 $Y2=2.72
r202 46 83 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.095 $Y=2.72
+ $X2=8.51 $Y2=2.72
r203 46 48 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.095 $Y=2.72
+ $X2=7.942 $Y2=2.72
r204 44 74 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.9 $Y=2.72 $X2=5.75
+ $Y2=2.72
r205 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.72
+ $X2=5.985 $Y2=2.72
r206 43 77 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.07 $Y=2.72
+ $X2=6.21 $Y2=2.72
r207 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=2.72
+ $X2=5.985 $Y2=2.72
r208 39 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=2.635
+ $X2=8.96 $Y2=2.72
r209 39 41 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.96 $Y=2.635
+ $X2=8.96 $Y2=1.79
r210 35 48 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.942 $Y=2.635
+ $X2=7.942 $Y2=2.72
r211 35 37 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=7.942 $Y=2.635
+ $X2=7.942 $Y2=2.3
r212 31 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=2.635
+ $X2=5.985 $Y2=2.72
r213 31 33 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.985 $Y=2.635
+ $X2=5.985 $Y2=2
r214 27 96 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.827 $Y=2.635
+ $X2=3.827 $Y2=2.72
r215 27 29 17.3473 $w=1.93e-07 $l=3.05e-07 $layer=LI1_cond $X=3.827 $Y=2.635
+ $X2=3.827 $Y2=2.33
r216 23 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.72
r217 23 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.045 $Y=2.635
+ $X2=2.045 $Y2=2.33
r218 19 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.72
r219 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.22
r220 6 41 300 $w=1.7e-07 $l=3.74566e-07 $layer=licon1_PDIFF $count=2 $X=8.805
+ $Y=1.485 $X2=8.96 $Y2=1.79
r221 5 37 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=2.065 $X2=7.995 $Y2=2.3
r222 4 33 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=5.61
+ $Y=2.065 $X2=5.985 $Y2=2
r223 3 29 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.845 $X2=3.815 $Y2=2.33
r224 2 25 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.845 $X2=2.045 $Y2=2.33
r225 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.815 $X2=0.685 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%A_556_369# 1 2 3 4 13 17 22 24 25 26 27 28
+ 29 30 34
c106 26 0 1.91058e-19 $X=3.56 $Y=1.91
r107 34 36 21.0047 $w=2.12e-07 $l=3.65e-07 $layer=LI1_cond $X=4.3 $Y=1.91
+ $X2=4.3 $Y2=2.275
r108 32 33 18.5652 $w=2.3e-07 $l=3.5e-07 $layer=LI1_cond $X=4.32 $Y=0.45
+ $X2=4.32 $Y2=0.8
r109 30 34 5.40561 $w=2.12e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.265 $Y=1.825
+ $X2=4.3 $Y2=1.91
r110 29 33 5.36376 $w=2.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.265 $Y=0.885
+ $X2=4.32 $Y2=0.8
r111 29 30 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.265 $Y=0.885
+ $X2=4.265 $Y2=1.825
r112 27 33 2.50919 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.18 $Y=0.8 $X2=4.32
+ $Y2=0.8
r113 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.18 $Y=0.8 $X2=3.59
+ $Y2=0.8
r114 25 34 2.03271 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.18 $Y=1.91 $X2=4.3
+ $Y2=1.91
r115 25 26 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.18 $Y=1.91
+ $X2=3.56 $Y2=1.91
r116 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=0.715
+ $X2=3.59 $Y2=0.8
r117 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.505 $Y=0.445
+ $X2=3.505 $Y2=0.715
r118 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.475 $Y=1.995
+ $X2=3.56 $Y2=1.91
r119 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.475 $Y=1.995
+ $X2=3.475 $Y2=2.245
r120 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=0.36
+ $X2=3.505 $Y2=0.445
r121 17 19 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.42 $Y=0.36
+ $X2=2.995 $Y2=0.36
r122 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.39 $Y=2.33
+ $X2=3.475 $Y2=2.245
r123 13 15 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.39 $Y=2.33
+ $X2=2.915 $Y2=2.33
r124 4 36 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.21
+ $Y=2.065 $X2=4.335 $Y2=2.275
r125 3 15 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.845 $X2=2.915 $Y2=2.33
r126 2 32 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.245
+ $Y=0.235 $X2=4.37 $Y2=0.45
r127 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.235 $X2=2.995 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%Q 1 2 11 12 13 14 15 27
r27 15 24 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=9.402 $Y=2.21
+ $X2=9.402 $Y2=2.31
r28 14 15 11.3574 $w=3.43e-07 $l=3.4e-07 $layer=LI1_cond $X=9.402 $Y=1.87
+ $X2=9.402 $Y2=2.21
r29 13 31 13.323 $w=3.43e-07 $l=3.1e-07 $layer=LI1_cond $X=9.402 $Y=0.51
+ $X2=9.402 $Y2=0.82
r30 13 27 3.84148 $w=3.43e-07 $l=1.15e-07 $layer=LI1_cond $X=9.402 $Y=0.51
+ $X2=9.402 $Y2=0.395
r31 12 31 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=9.49 $Y=1.505
+ $X2=9.49 $Y2=0.82
r32 11 12 7.14324 $w=3.43e-07 $l=1.25e-07 $layer=LI1_cond $X=9.402 $Y=1.63
+ $X2=9.402 $Y2=1.505
r33 9 14 6.447 $w=3.43e-07 $l=1.93e-07 $layer=LI1_cond $X=9.402 $Y=1.677
+ $X2=9.402 $Y2=1.87
r34 9 11 1.56999 $w=3.43e-07 $l=4.7e-08 $layer=LI1_cond $X=9.402 $Y=1.677
+ $X2=9.402 $Y2=1.63
r35 2 24 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=1.485 $X2=9.395 $Y2=2.31
r36 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=1.485 $X2=9.395 $Y2=1.63
r37 1 27 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=9.26
+ $Y=0.235 $X2=9.395 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXTP_1%VGND 1 2 3 4 5 6 21 25 29 31 35 39 43 46 47
+ 49 50 51 53 58 63 82 83 86 89 92 95
c157 83 0 2.71124e-20 $X=9.43 $Y=0
c158 2 0 8.19616e-20 $X=1.925 $Y=0.235
r159 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r160 93 96 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r161 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r162 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r163 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r164 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r165 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r166 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r167 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r168 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r169 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r170 74 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r171 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=7.59
+ $Y2=0
r172 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r173 71 95 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=5.875
+ $Y2=0
r174 71 73 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=6.21
+ $Y2=0
r175 70 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r176 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r177 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r178 67 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r179 66 69 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r180 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r181 64 89 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.132 $Y2=0
r182 64 66 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.53 $Y2=0
r183 63 92 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.86
+ $Y2=0
r184 63 69 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.45
+ $Y2=0
r185 62 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r186 62 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r187 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r188 59 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r189 59 61 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r190 58 89 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=2.132
+ $Y2=0
r191 58 61 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=1.61
+ $Y2=0
r192 53 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r193 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r194 51 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r195 51 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r196 49 79 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.875 $Y=0
+ $X2=8.51 $Y2=0
r197 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.875 $Y=0 $X2=8.96
+ $Y2=0
r198 48 82 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=9.43 $Y2=0
r199 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.045 $Y=0 $X2=8.96
+ $Y2=0
r200 46 76 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.59 $Y2=0
r201 46 47 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.715 $Y=0 $X2=7.9
+ $Y2=0
r202 45 79 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.085 $Y=0
+ $X2=8.51 $Y2=0
r203 45 47 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.085 $Y=0 $X2=7.9
+ $Y2=0
r204 41 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0
r205 41 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0.53
r206 37 47 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.085 $X2=7.9
+ $Y2=0
r207 37 39 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.9 $Y=0.085
+ $X2=7.9 $Y2=0.45
r208 33 95 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=0.085
+ $X2=5.875 $Y2=0
r209 33 35 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.875 $Y=0.085
+ $X2=5.875 $Y2=0.42
r210 32 92 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.86
+ $Y2=0
r211 31 95 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.875
+ $Y2=0
r212 31 32 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=5.69 $Y=0 $X2=3.96
+ $Y2=0
r213 27 92 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0
r214 27 29 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0.38
r215 23 89 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.132 $Y=0.085
+ $X2=2.132 $Y2=0
r216 23 25 9.18614 $w=3.43e-07 $l=2.75e-07 $layer=LI1_cond $X=2.132 $Y=0.085
+ $X2=2.132 $Y2=0.36
r217 19 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r218 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r219 6 43 182 $w=1.7e-07 $l=3.64349e-07 $layer=licon1_NDIFF $count=1 $X=8.805
+ $Y=0.235 $X2=8.96 $Y2=0.53
r220 5 39 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=7.865
+ $Y=0.235 $X2=8 $Y2=0.45
r221 4 35 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.945 $Y2=0.42
r222 3 29 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.235 $X2=3.85 $Y2=0.38
r223 2 25 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.125 $Y2=0.36
r224 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


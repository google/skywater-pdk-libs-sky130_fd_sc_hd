* File: sky130_fd_sc_hd__a41o_4.spice.SKY130_FD_SC_HD__A41O_4.pxi
* Created: Thu Aug 27 14:06:15 2020
* 
x_PM_SKY130_FD_SC_HD__A41O_4%A_79_21# N_A_79_21#_M1013_s N_A_79_21#_M1001_s
+ N_A_79_21#_M1010_s N_A_79_21#_c_103_n N_A_79_21#_M1012_g N_A_79_21#_M1000_g
+ N_A_79_21#_c_104_n N_A_79_21#_M1015_g N_A_79_21#_M1004_g N_A_79_21#_c_105_n
+ N_A_79_21#_M1017_g N_A_79_21#_M1018_g N_A_79_21#_c_106_n N_A_79_21#_M1025_g
+ N_A_79_21#_M1023_g N_A_79_21#_c_169_p N_A_79_21#_c_107_n N_A_79_21#_c_108_n
+ N_A_79_21#_c_121_p N_A_79_21#_c_194_p N_A_79_21#_c_117_n N_A_79_21#_c_147_p
+ N_A_79_21#_c_210_p N_A_79_21#_c_109_n N_A_79_21#_c_110_n N_A_79_21#_c_133_p
+ N_A_79_21#_c_125_p N_A_79_21#_c_111_n PM_SKY130_FD_SC_HD__A41O_4%A_79_21#
x_PM_SKY130_FD_SC_HD__A41O_4%B1 N_B1_c_228_n N_B1_M1013_g N_B1_c_229_n
+ N_B1_M1016_g N_B1_M1010_g N_B1_M1014_g B1 B1 N_B1_c_230_n
+ PM_SKY130_FD_SC_HD__A41O_4%B1
x_PM_SKY130_FD_SC_HD__A41O_4%A1 N_A1_c_280_n N_A1_M1001_g N_A1_M1005_g
+ N_A1_c_281_n N_A1_M1026_g N_A1_M1009_g A1 A1 N_A1_c_283_n
+ PM_SKY130_FD_SC_HD__A41O_4%A1
x_PM_SKY130_FD_SC_HD__A41O_4%A2 N_A2_M1006_g N_A2_M1002_g N_A2_M1008_g
+ N_A2_M1024_g A2 A2 N_A2_c_327_n PM_SKY130_FD_SC_HD__A41O_4%A2
x_PM_SKY130_FD_SC_HD__A41O_4%A3 N_A3_M1003_g N_A3_M1020_g N_A3_M1027_g
+ N_A3_M1007_g N_A3_c_369_n A3 A3 N_A3_c_370_n N_A3_c_371_n N_A3_c_372_n
+ PM_SKY130_FD_SC_HD__A41O_4%A3
x_PM_SKY130_FD_SC_HD__A41O_4%A4 N_A4_M1021_g N_A4_M1011_g N_A4_M1022_g
+ N_A4_M1019_g A4 A4 N_A4_c_418_n N_A4_c_419_n N_A4_c_420_n
+ PM_SKY130_FD_SC_HD__A41O_4%A4
x_PM_SKY130_FD_SC_HD__A41O_4%VPWR N_VPWR_M1000_s N_VPWR_M1004_s N_VPWR_M1023_s
+ N_VPWR_M1005_s N_VPWR_M1002_d N_VPWR_M1003_d N_VPWR_M1011_s N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n
+ N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_463_n
+ N_VPWR_c_464_n N_VPWR_c_465_n VPWR N_VPWR_c_466_n N_VPWR_c_467_n
+ N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_452_n N_VPWR_c_471_n N_VPWR_c_472_n
+ N_VPWR_c_473_n N_VPWR_c_474_n PM_SKY130_FD_SC_HD__A41O_4%VPWR
x_PM_SKY130_FD_SC_HD__A41O_4%X N_X_M1012_s N_X_M1017_s N_X_M1000_d N_X_M1018_d
+ N_X_c_614_p N_X_c_594_n N_X_c_574_n N_X_c_578_n N_X_c_613_p N_X_c_598_n
+ N_X_c_582_n N_X_c_584_n N_X_c_586_n N_X_c_588_n X X X N_X_c_606_p N_X_c_602_n
+ X X PM_SKY130_FD_SC_HD__A41O_4%X
x_PM_SKY130_FD_SC_HD__A41O_4%A_467_297# N_A_467_297#_M1010_d
+ N_A_467_297#_M1014_d N_A_467_297#_M1009_d N_A_467_297#_M1024_s
+ N_A_467_297#_M1007_s N_A_467_297#_M1019_d N_A_467_297#_c_626_n
+ N_A_467_297#_c_628_n N_A_467_297#_c_666_n N_A_467_297#_c_631_n
+ N_A_467_297#_c_636_n N_A_467_297#_c_635_n N_A_467_297#_c_671_n
+ N_A_467_297#_c_641_n N_A_467_297#_c_645_n N_A_467_297#_c_648_n
+ N_A_467_297#_c_680_n N_A_467_297#_c_624_n N_A_467_297#_c_684_n
+ N_A_467_297#_c_646_n PM_SKY130_FD_SC_HD__A41O_4%A_467_297#
x_PM_SKY130_FD_SC_HD__A41O_4%VGND N_VGND_M1012_d N_VGND_M1015_d N_VGND_M1025_d
+ N_VGND_M1016_d N_VGND_M1021_s N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n N_VGND_c_695_n VGND N_VGND_c_696_n N_VGND_c_697_n
+ N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n
+ PM_SKY130_FD_SC_HD__A41O_4%VGND
x_PM_SKY130_FD_SC_HD__A41O_4%A_639_47# N_A_639_47#_M1001_d N_A_639_47#_M1026_d
+ N_A_639_47#_M1008_d N_A_639_47#_c_805_n N_A_639_47#_c_806_n
+ PM_SKY130_FD_SC_HD__A41O_4%A_639_47#
x_PM_SKY130_FD_SC_HD__A41O_4%A_889_47# N_A_889_47#_M1006_s N_A_889_47#_M1020_d
+ N_A_889_47#_c_831_n PM_SKY130_FD_SC_HD__A41O_4%A_889_47#
x_PM_SKY130_FD_SC_HD__A41O_4%A_1079_47# N_A_1079_47#_M1020_s
+ N_A_1079_47#_M1027_s N_A_1079_47#_M1022_d N_A_1079_47#_c_850_n
+ N_A_1079_47#_c_869_n PM_SKY130_FD_SC_HD__A41O_4%A_1079_47#
cc_1 VNB N_A_79_21#_c_103_n 0.0182854f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_104_n 0.0157741f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_105_n 0.0157701f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_106_n 0.0155194f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_107_n 0.00179069f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.075
cc_6 VNB N_A_79_21#_c_108_n 4.49304e-19 $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.455
cc_7 VNB N_A_79_21#_c_109_n 0.00757042f $X=-0.19 $Y=-0.24 $X2=3.74 $Y2=0.73
cc_8 VNB N_A_79_21#_c_110_n 0.00106277f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.16
cc_9 VNB N_A_79_21#_c_111_n 0.0675919f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_10 VNB N_B1_c_228_n 0.0161338f $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=0.235
cc_11 VNB N_B1_c_229_n 0.0210848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_230_n 0.0618675f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_13 VNB N_A1_c_280_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=0.235
cc_14 VNB N_A1_c_281_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB A1 0.00313855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_283_n 0.0370014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A2_M1006_g 0.017802f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=1.485
cc_18 VNB N_A2_M1002_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_M1008_g 0.0243831f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_A2_M1024_g 4.72682e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_21 VNB A2 0.00333599f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_22 VNB N_A2_c_327_n 0.0348155f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_23 VNB N_A3_M1003_g 7.42991e-19 $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=1.485
cc_24 VNB N_A3_M1020_g 0.0243831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A3_M1027_g 0.017802f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_26 VNB N_A3_M1007_g 7.36106e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_27 VNB N_A3_c_369_n 0.0124857f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_28 VNB N_A3_c_370_n 0.0254321f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_29 VNB N_A3_c_371_n 0.00143932f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_30 VNB N_A3_c_372_n 0.0325605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A4_M1021_g 0.0175748f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=1.485
cc_32 VNB N_A4_M1011_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A4_M1022_g 0.0241559f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_34 VNB N_A4_M1019_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_35 VNB N_A4_c_418_n 0.024556f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_36 VNB N_A4_c_419_n 0.0522022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A4_c_420_n 0.0106086f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_38 VNB N_VPWR_c_452_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB X 0.0198276f $X=-0.19 $Y=-0.24 $X2=2.295 $Y2=0.73
cc_40 VNB N_VGND_c_686_n 0.010303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_687_n 0.0130541f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_42 VNB N_VGND_c_688_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_43 VNB N_VGND_c_689_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_44 VNB N_VGND_c_690_n 0.00543973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_691_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_46 VNB N_VGND_c_692_n 0.0117278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_693_n 0.00462744f $X=-0.19 $Y=-0.24 $X2=1.775 $Y2=1.16
cc_48 VNB N_VGND_c_694_n 0.0109937f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_49 VNB N_VGND_c_695_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_50 VNB N_VGND_c_696_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=1.16
cc_51 VNB N_VGND_c_697_n 0.0871172f $X=-0.19 $Y=-0.24 $X2=2.38 $Y2=0.42
cc_52 VNB N_VGND_c_698_n 0.0266114f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=1.625
cc_53 VNB N_VGND_c_699_n 0.392193f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=1.955
cc_54 VNB N_VGND_c_700_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=2.04
cc_55 VNB N_VGND_c_701_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_56 VNB N_A_639_47#_c_805_n 0.00217698f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_57 VNB N_A_639_47#_c_806_n 0.00295274f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_58 VNB N_A_889_47#_c_831_n 0.00667811f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_59 VNB N_A_1079_47#_c_850_n 0.00213317f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_60 VPB N_A_79_21#_M1000_g 0.0210031f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_A_79_21#_M1004_g 0.0182735f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_A_79_21#_M1018_g 0.0182675f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_63 VPB N_A_79_21#_M1023_g 0.0220963f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_64 VPB N_A_79_21#_c_108_n 0.00207061f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.455
cc_65 VPB N_A_79_21#_c_117_n 0.01709f $X=-0.19 $Y=1.305 $X2=2.795 $Y2=1.54
cc_66 VPB N_A_79_21#_c_111_n 0.0106359f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_67 VPB N_B1_M1010_g 0.0231641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_B1_M1014_g 0.0190537f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_69 VPB N_B1_c_230_n 0.0178517f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_70 VPB N_A1_M1005_g 0.0188339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A1_M1009_g 0.0186099f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_72 VPB N_A1_c_283_n 0.0042353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A2_M1002_g 0.0196968f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A2_M1024_g 0.0199383f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_75 VPB N_A3_M1003_g 0.028274f $X=-0.19 $Y=1.305 $X2=2.745 $Y2=1.485
cc_76 VPB N_A3_M1007_g 0.0280325f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_77 VPB N_A4_M1011_g 0.0196968f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A4_M1019_g 0.0274383f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_79 VPB N_VPWR_c_453_n 0.0103102f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_80 VPB N_VPWR_c_454_n 0.0262563f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_81 VPB N_VPWR_c_455_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_82 VPB N_VPWR_c_456_n 0.00941534f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_83 VPB N_VPWR_c_457_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_84 VPB N_VPWR_c_458_n 3.1722e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_85 VPB N_VPWR_c_459_n 0.00635696f $X=-0.19 $Y=1.305 $X2=1.675 $Y2=1.16
cc_86 VPB N_VPWR_c_460_n 0.0157658f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=0.815
cc_87 VPB N_VPWR_c_461_n 4.07719e-19 $X=-0.19 $Y=1.305 $X2=2.295 $Y2=0.73
cc_88 VPB N_VPWR_c_462_n 0.0350797f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=1.54
cc_89 VPB N_VPWR_c_463_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.38 $Y2=0.645
cc_90 VPB N_VPWR_c_464_n 0.0124915f $X=-0.19 $Y=1.305 $X2=2.38 $Y2=0.42
cc_91 VPB N_VPWR_c_465_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_466_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.74 $Y2=0.73
cc_93 VPB N_VPWR_c_467_n 0.0124915f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=1.7
cc_94 VPB N_VPWR_c_468_n 0.0164023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_469_n 0.0273603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_452_n 0.0691293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_471_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_472_n 0.00546352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_473_n 0.0132461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_474_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB X 0.00857396f $X=-0.19 $Y=1.305 $X2=2.295 $Y2=0.73
cc_102 VPB N_A_467_297#_c_624_n 0.00906696f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.075
cc_103 N_A_79_21#_c_106_n N_B1_c_228_n 0.011972f $X=1.73 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_79_21#_c_107_n N_B1_c_228_n 0.00559518f $X=1.86 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_79_21#_c_121_p N_B1_c_228_n 0.0124284f $X=2.295 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_106 N_A_79_21#_c_109_n N_B1_c_229_n 0.0141261f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_108_n N_B1_M1010_g 0.0026904f $X=1.86 $Y=1.455 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_117_n N_B1_M1010_g 0.0129283f $X=2.795 $Y=1.54 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_125_p N_B1_M1010_g 0.00275882f $X=2.88 $Y=2.04 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_117_n N_B1_M1014_g 0.00100609f $X=2.795 $Y=1.54 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_125_p N_B1_M1014_g 0.00304537f $X=2.88 $Y=2.04 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_108_n B1 0.00246196f $X=1.86 $Y=1.455 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_121_p B1 0.00662939f $X=2.295 $Y=0.73 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_117_n B1 0.0597946f $X=2.795 $Y=1.54 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_109_n B1 0.0320578f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_110_n B1 0.0138466f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_133_p B1 0.00920238f $X=2.38 $Y=0.73 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_125_p B1 0.00117101f $X=2.88 $Y=2.04 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_111_n B1 2.00657e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_108_n N_B1_c_230_n 0.00128032f $X=1.86 $Y=1.455 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_117_n N_B1_c_230_n 0.0158714f $X=2.795 $Y=1.54 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_109_n N_B1_c_230_n 0.0132852f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_110_n N_B1_c_230_n 0.00139404f $X=1.86 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_133_p N_B1_c_230_n 0.00217728f $X=2.38 $Y=0.73 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_111_n N_B1_c_230_n 0.0272253f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_109_n N_A1_c_280_n 0.0110418f $X=3.74 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_79_21#_c_109_n N_A1_c_281_n 0.00265854f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_109_n A1 0.0213252f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_109_n N_A1_c_283_n 0.00320521f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_117_n N_VPWR_M1023_s 0.00223165f $X=2.795 $Y=1.54 $X2=0
+ $Y2=0
cc_131 N_A_79_21#_c_147_p N_VPWR_M1023_s 0.00117638f $X=1.945 $Y=1.54 $X2=0
+ $Y2=0
cc_132 N_A_79_21#_M1000_g N_VPWR_c_454_n 0.0112954f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_79_21#_M1004_g N_VPWR_c_454_n 6.0901e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_79_21#_M1000_g N_VPWR_c_455_n 6.0901e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_79_21#_M1004_g N_VPWR_c_455_n 0.0101939f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_79_21#_M1018_g N_VPWR_c_455_n 0.0101939f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_79_21#_M1023_g N_VPWR_c_455_n 6.0901e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_79_21#_M1018_g N_VPWR_c_456_n 6.10071e-19 $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_79_21#_M1023_g N_VPWR_c_456_n 0.0114703f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_117_n N_VPWR_c_456_n 0.00998872f $X=2.795 $Y=1.54 $X2=0
+ $Y2=0
cc_141 N_A_79_21#_c_147_p N_VPWR_c_456_n 0.0066017f $X=1.945 $Y=1.54 $X2=0 $Y2=0
cc_142 N_A_79_21#_M1000_g N_VPWR_c_466_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_79_21#_M1004_g N_VPWR_c_466_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_79_21#_M1018_g N_VPWR_c_467_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_79_21#_M1023_g N_VPWR_c_467_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_79_21#_M1010_s N_VPWR_c_452_n 0.00216833f $X=2.745 $Y=1.485 $X2=0
+ $Y2=0
cc_147 N_A_79_21#_M1000_g N_VPWR_c_452_n 0.00789179f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_79_21#_M1004_g N_VPWR_c_452_n 0.00789179f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_79_21#_M1018_g N_VPWR_c_452_n 0.00789179f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_79_21#_M1023_g N_VPWR_c_452_n 0.00789179f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_79_21#_c_104_n N_X_c_574_n 0.0119428f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_105_n N_X_c_574_n 0.0115547f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_169_p N_X_c_574_n 0.0355556f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_111_n N_X_c_574_n 0.00423243f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_79_21#_M1004_g N_X_c_578_n 0.0148668f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_79_21#_M1018_g N_X_c_578_n 0.0144787f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_169_p N_X_c_578_n 0.0304888f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_111_n N_X_c_578_n 0.00408007f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_103_n N_X_c_582_n 0.0158497f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_79_21#_c_169_p N_X_c_582_n 0.00374684f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_169_p N_X_c_584_n 0.00881067f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_111_n N_X_c_584_n 0.00216182f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_79_21#_M1000_g N_X_c_586_n 0.0185751f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_79_21#_c_169_p N_X_c_586_n 0.0031876f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_169_p N_X_c_588_n 0.00768518f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_111_n N_X_c_588_n 0.00210139f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_103_n X 0.0290345f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_169_p X 0.0134244f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_117_n N_A_467_297#_M1010_d 0.00390196f $X=2.795 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_170 N_A_79_21#_M1023_g N_A_467_297#_c_626_n 0.00148337f $X=1.73 $Y=1.985
+ $X2=0 $Y2=0
cc_171 N_A_79_21#_c_117_n N_A_467_297#_c_626_n 0.0131641f $X=2.795 $Y=1.54 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_M1010_s N_A_467_297#_c_628_n 0.00312348f $X=2.745 $Y=1.485
+ $X2=0 $Y2=0
cc_173 N_A_79_21#_c_117_n N_A_467_297#_c_628_n 0.00259534f $X=2.795 $Y=1.54
+ $X2=0 $Y2=0
cc_174 N_A_79_21#_c_125_p N_A_467_297#_c_628_n 0.0155384f $X=2.88 $Y=2.04 $X2=0
+ $Y2=0
cc_175 N_A_79_21#_c_125_p N_A_467_297#_c_631_n 0.011519f $X=2.88 $Y=2.04 $X2=0
+ $Y2=0
cc_176 N_A_79_21#_c_107_n N_VGND_M1025_d 7.90193e-19 $X=1.86 $Y=1.075 $X2=0
+ $Y2=0
cc_177 N_A_79_21#_c_121_p N_VGND_M1025_d 0.00275654f $X=2.295 $Y=0.73 $X2=0
+ $Y2=0
cc_178 N_A_79_21#_c_194_p N_VGND_M1025_d 9.05974e-19 $X=1.945 $Y=0.73 $X2=0
+ $Y2=0
cc_179 N_A_79_21#_c_109_n N_VGND_M1016_d 0.00489262f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_180 N_A_79_21#_c_103_n N_VGND_c_687_n 0.00774571f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_79_21#_c_104_n N_VGND_c_687_n 5.08801e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_79_21#_c_103_n N_VGND_c_688_n 5.08801e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_79_21#_c_104_n N_VGND_c_688_n 0.00664421f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_79_21#_c_105_n N_VGND_c_688_n 0.00664421f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_79_21#_c_106_n N_VGND_c_688_n 5.08801e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_79_21#_c_105_n N_VGND_c_689_n 5.10011e-19 $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_79_21#_c_106_n N_VGND_c_689_n 0.00671223f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_79_21#_c_121_p N_VGND_c_689_n 0.00866404f $X=2.295 $Y=0.73 $X2=0
+ $Y2=0
cc_189 N_A_79_21#_c_194_p N_VGND_c_689_n 0.00880282f $X=1.945 $Y=0.73 $X2=0
+ $Y2=0
cc_190 N_A_79_21#_c_109_n N_VGND_c_690_n 0.0196494f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_105_n N_VGND_c_692_n 0.00339367f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_79_21#_c_106_n N_VGND_c_692_n 0.0046653f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_121_p N_VGND_c_694_n 0.00238578f $X=2.295 $Y=0.73 $X2=0
+ $Y2=0
cc_194 N_A_79_21#_c_210_p N_VGND_c_694_n 0.0112415f $X=2.38 $Y=0.42 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_109_n N_VGND_c_694_n 0.00238578f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_103_n N_VGND_c_696_n 0.00339367f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_79_21#_c_104_n N_VGND_c_696_n 0.00339367f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_79_21#_c_109_n N_VGND_c_697_n 0.00339034f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_199 N_A_79_21#_M1013_s N_VGND_c_699_n 0.00250764f $X=2.245 $Y=0.235 $X2=0
+ $Y2=0
cc_200 N_A_79_21#_M1001_s N_VGND_c_699_n 0.00219239f $X=3.605 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_A_79_21#_c_103_n N_VGND_c_699_n 0.00394406f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_79_21#_c_104_n N_VGND_c_699_n 0.00394406f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_79_21#_c_105_n N_VGND_c_699_n 0.00394406f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_79_21#_c_106_n N_VGND_c_699_n 0.00789179f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_79_21#_c_121_p N_VGND_c_699_n 0.00495288f $X=2.295 $Y=0.73 $X2=0
+ $Y2=0
cc_206 N_A_79_21#_c_194_p N_VGND_c_699_n 8.47467e-19 $X=1.945 $Y=0.73 $X2=0
+ $Y2=0
cc_207 N_A_79_21#_c_210_p N_VGND_c_699_n 0.00643744f $X=2.38 $Y=0.42 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_109_n N_VGND_c_699_n 0.0124405f $X=3.74 $Y=0.73 $X2=0 $Y2=0
cc_209 N_A_79_21#_c_109_n N_A_639_47#_M1001_d 0.010508f $X=3.74 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_210 N_A_79_21#_M1001_s N_A_639_47#_c_805_n 0.003196f $X=3.605 $Y=0.235 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_c_109_n N_A_639_47#_c_805_n 0.0372327f $X=3.74 $Y=0.73 $X2=0
+ $Y2=0
cc_212 N_B1_M1014_g N_A1_M1005_g 0.0132702f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_213 B1 A1 0.0125741f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_214 N_B1_c_230_n A1 9.74533e-19 $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_215 B1 N_A1_c_283_n 2.4642e-19 $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_216 N_B1_c_230_n N_A1_c_283_n 0.0321413f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B1_M1010_g N_VPWR_c_456_n 0.00244463f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_M1014_g N_VPWR_c_457_n 0.00107061f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B1_M1010_g N_VPWR_c_462_n 0.00357877f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B1_M1014_g N_VPWR_c_462_n 0.00357877f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B1_M1010_g N_VPWR_c_452_n 0.00655123f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_222 N_B1_M1014_g N_VPWR_c_452_n 0.00530095f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B1_M1010_g N_A_467_297#_c_628_n 0.00940156f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_B1_M1014_g N_A_467_297#_c_628_n 0.0112437f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B1_M1014_g N_A_467_297#_c_631_n 0.00504295f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_B1_M1014_g N_A_467_297#_c_635_n 0.00168107f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_B1_c_228_n N_VGND_c_689_n 0.00671343f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_229_n N_VGND_c_689_n 5.10011e-19 $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_228_n N_VGND_c_690_n 5.08801e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_229_n N_VGND_c_690_n 0.00775781f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_228_n N_VGND_c_694_n 0.00340533f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B1_c_229_n N_VGND_c_694_n 0.00340533f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_228_n N_VGND_c_699_n 0.00396343f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B1_c_229_n N_VGND_c_699_n 0.00396343f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A1_c_281_n N_A2_M1006_g 0.0262473f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A1_c_283_n N_A2_M1002_g 0.0297623f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_237 A1 A2 0.0148574f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_238 N_A1_c_283_n A2 2.58364e-19 $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_239 A1 N_A2_c_327_n 3.34282e-19 $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_240 N_A1_c_283_n N_A2_c_327_n 0.0185615f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_M1005_g N_VPWR_c_457_n 0.0114515f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A1_M1009_g N_VPWR_c_457_n 0.0102418f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A1_M1009_g N_VPWR_c_458_n 6.0901e-19 $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A1_M1005_g N_VPWR_c_462_n 0.0046653f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A1_M1009_g N_VPWR_c_464_n 0.0046653f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A1_M1005_g N_VPWR_c_452_n 0.00796757f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A1_M1009_g N_VPWR_c_452_n 0.007919f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A1_M1005_g N_A_467_297#_c_636_n 0.0141246f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A1_M1009_g N_A_467_297#_c_636_n 0.0144336f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_250 A1 N_A_467_297#_c_636_n 0.0297787f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_251 N_A1_c_283_n N_A_467_297#_c_636_n 0.00199384f $X=3.95 $Y=1.16 $X2=0 $Y2=0
cc_252 A1 N_A_467_297#_c_635_n 3.72838e-19 $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A1_c_280_n N_VGND_c_690_n 0.00294182f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_280_n N_VGND_c_697_n 0.00366111f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_281_n N_VGND_c_697_n 0.00366111f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A1_c_280_n N_VGND_c_699_n 0.00656615f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A1_c_281_n N_VGND_c_699_n 0.00530732f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_c_280_n N_A_639_47#_c_805_n 0.00790826f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_281_n N_A_639_47#_c_805_n 0.0109652f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_260 A1 N_A_639_47#_c_805_n 0.00335763f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_261 N_A2_M1024_g N_A3_M1003_g 0.0273833f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_262 A2 N_A3_c_369_n 7.93071e-19 $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_263 N_A2_c_327_n N_A3_c_369_n 0.0185903f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_264 A2 N_A3_c_371_n 0.0177963f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_265 N_A2_c_327_n N_A3_c_371_n 3.16775e-19 $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A2_M1002_g N_VPWR_c_457_n 6.0901e-19 $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A2_M1002_g N_VPWR_c_458_n 0.0102418f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A2_M1024_g N_VPWR_c_458_n 0.0107237f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A2_M1002_g N_VPWR_c_464_n 0.0046653f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A2_M1024_g N_VPWR_c_468_n 0.0046653f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A2_M1002_g N_VPWR_c_452_n 0.007919f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A2_M1024_g N_VPWR_c_452_n 0.00796757f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A2_M1002_g N_A_467_297#_c_641_n 0.0145338f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A2_M1024_g N_A_467_297#_c_641_n 0.0146524f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_275 A2 N_A_467_297#_c_641_n 0.0290418f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_276 N_A2_c_327_n N_A_467_297#_c_641_n 0.00314532f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A2_M1024_g N_A_467_297#_c_645_n 0.00593237f $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_278 A2 N_A_467_297#_c_646_n 0.00250121f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_279 N_A2_c_327_n N_A_467_297#_c_646_n 2.17302e-19 $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A2_M1006_g N_VGND_c_697_n 0.00414474f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A2_M1008_g N_VGND_c_697_n 0.00366111f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A2_M1006_g N_VGND_c_699_n 0.00576602f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A2_M1008_g N_VGND_c_699_n 0.00661716f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A2_M1006_g N_A_639_47#_c_806_n 0.0100379f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A2_M1008_g N_A_639_47#_c_806_n 0.00889468f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_286 A2 N_A_639_47#_c_806_n 0.0303153f $X=4.79 $Y=1.105 $X2=0 $Y2=0
cc_287 N_A2_c_327_n N_A_639_47#_c_806_n 0.00348379f $X=4.79 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A2_M1006_g N_A_889_47#_c_831_n 0.00246655f $X=4.37 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A2_M1008_g N_A_889_47#_c_831_n 0.0100554f $X=4.79 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A3_M1027_g N_A4_M1021_g 0.0238565f $X=6.15 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A3_M1007_g N_A4_M1011_g 0.0238565f $X=6.15 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A3_c_371_n N_A4_c_418_n 2.58387e-19 $X=6.02 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A3_c_372_n N_A4_c_418_n 0.0238565f $X=6.15 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A3_c_371_n N_A4_c_420_n 0.0113623f $X=6.02 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A3_c_372_n N_A4_c_420_n 9.89829e-19 $X=6.15 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A3_M1003_g N_VPWR_c_458_n 6.42981e-19 $X=5.23 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A3_M1003_g N_VPWR_c_459_n 0.0144145f $X=5.23 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A3_M1007_g N_VPWR_c_459_n 0.0143861f $X=6.15 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A3_M1007_g N_VPWR_c_460_n 0.00585385f $X=6.15 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A3_M1007_g N_VPWR_c_461_n 6.37932e-19 $X=6.15 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A3_M1003_g N_VPWR_c_468_n 0.00585385f $X=5.23 $Y=1.985 $X2=0 $Y2=0
cc_302 N_A3_M1003_g N_VPWR_c_452_n 0.0120405f $X=5.23 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A3_M1007_g N_VPWR_c_452_n 0.0119919f $X=6.15 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A3_M1003_g N_A_467_297#_c_648_n 0.0175396f $X=5.23 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A3_M1007_g N_A_467_297#_c_648_n 0.0185325f $X=6.15 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A3_c_370_n N_A_467_297#_c_648_n 0.0131832f $X=5.655 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A3_c_371_n N_A_467_297#_c_648_n 0.0526793f $X=6.02 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A3_M1027_g N_VGND_c_691_n 0.0018398f $X=6.15 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A3_M1020_g N_VGND_c_697_n 0.00366111f $X=5.73 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A3_M1027_g N_VGND_c_697_n 0.00414474f $X=6.15 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A3_M1020_g N_VGND_c_699_n 0.00661716f $X=5.73 $Y=0.56 $X2=0 $Y2=0
cc_312 N_A3_M1027_g N_VGND_c_699_n 0.00576602f $X=6.15 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A3_c_369_n N_A_639_47#_c_806_n 2.61353e-19 $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A3_c_371_n N_A_639_47#_c_806_n 5.30975e-19 $X=6.02 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A3_M1020_g N_A_889_47#_c_831_n 0.0100554f $X=5.73 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A3_M1027_g N_A_889_47#_c_831_n 0.0036428f $X=6.15 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A3_c_369_n N_A_889_47#_c_831_n 0.00397513f $X=5.305 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A3_c_371_n N_A_889_47#_c_831_n 0.00525016f $X=6.02 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A3_M1020_g N_A_1079_47#_c_850_n 0.00893883f $X=5.73 $Y=0.56 $X2=0 $Y2=0
cc_320 N_A3_M1027_g N_A_1079_47#_c_850_n 0.0110926f $X=6.15 $Y=0.56 $X2=0 $Y2=0
cc_321 N_A3_c_370_n N_A_1079_47#_c_850_n 0.00644521f $X=5.655 $Y=1.16 $X2=0
+ $Y2=0
cc_322 N_A3_c_371_n N_A_1079_47#_c_850_n 0.0377211f $X=6.02 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A3_c_372_n N_A_1079_47#_c_850_n 0.00193451f $X=6.15 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A4_M1011_g N_VPWR_c_460_n 0.0046653f $X=6.57 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A4_M1011_g N_VPWR_c_461_n 0.0104049f $X=6.57 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A4_M1019_g N_VPWR_c_461_n 0.0121374f $X=6.99 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A4_M1019_g N_VPWR_c_469_n 0.0046653f $X=6.99 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A4_M1011_g N_VPWR_c_452_n 0.007919f $X=6.57 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A4_M1019_g N_VPWR_c_452_n 0.00921786f $X=6.99 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A4_M1011_g N_A_467_297#_c_624_n 0.0144777f $X=6.57 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A4_M1019_g N_A_467_297#_c_624_n 0.0159719f $X=6.99 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A4_c_418_n N_A_467_297#_c_624_n 0.0018492f $X=7.065 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A4_c_419_n N_A_467_297#_c_624_n 0.00539341f $X=7.34 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A4_c_420_n N_A_467_297#_c_624_n 0.0436638f $X=7.34 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A4_M1021_g N_VGND_c_691_n 0.0093539f $X=6.57 $Y=0.56 $X2=0 $Y2=0
cc_336 N_A4_M1022_g N_VGND_c_691_n 0.00835959f $X=6.99 $Y=0.56 $X2=0 $Y2=0
cc_337 N_A4_M1021_g N_VGND_c_697_n 0.00340533f $X=6.57 $Y=0.56 $X2=0 $Y2=0
cc_338 N_A4_M1022_g N_VGND_c_698_n 0.00340533f $X=6.99 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A4_M1021_g N_VGND_c_699_n 0.00403482f $X=6.57 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A4_M1022_g N_VGND_c_699_n 0.0052895f $X=6.99 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A4_M1021_g N_A_889_47#_c_831_n 4.913e-19 $X=6.57 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A4_M1021_g N_A_1079_47#_c_850_n 0.00997866f $X=6.57 $Y=0.56 $X2=0 $Y2=0
cc_343 N_A4_M1022_g N_A_1079_47#_c_850_n 0.0132313f $X=6.99 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A4_c_418_n N_A_1079_47#_c_850_n 0.00193451f $X=7.065 $Y=1.16 $X2=0
+ $Y2=0
cc_345 N_A4_c_419_n N_A_1079_47#_c_850_n 0.00378971f $X=7.34 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A4_c_420_n N_A_1079_47#_c_850_n 0.0363753f $X=7.34 $Y=1.16 $X2=0 $Y2=0
cc_347 N_VPWR_c_452_n N_X_M1000_d 0.00562358f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_348 N_VPWR_c_452_n N_X_M1018_d 0.00562358f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_349 N_VPWR_c_466_n N_X_c_594_n 0.0113958f $X=0.935 $Y=2.72 $X2=0 $Y2=0
cc_350 N_VPWR_c_452_n N_X_c_594_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_351 N_VPWR_M1004_s N_X_c_578_n 0.00363759f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_352 N_VPWR_c_455_n N_X_c_578_n 0.0170259f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_353 N_VPWR_c_467_n N_X_c_598_n 0.0113958f $X=1.775 $Y=2.72 $X2=0 $Y2=0
cc_354 N_VPWR_c_452_n N_X_c_598_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_355 N_VPWR_M1000_s N_X_c_586_n 8.29358e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_356 N_VPWR_c_454_n N_X_c_586_n 0.00359494f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_357 N_VPWR_M1000_s N_X_c_602_n 0.0101395f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_358 N_VPWR_c_454_n N_X_c_602_n 0.0152373f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_359 N_VPWR_M1000_s X 0.00469457f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_360 N_VPWR_c_452_n N_A_467_297#_M1010_d 0.00348186f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_361 N_VPWR_c_452_n N_A_467_297#_M1014_d 0.00401374f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_452_n N_A_467_297#_M1009_d 0.00562358f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_452_n N_A_467_297#_M1024_s 0.00647849f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_364 N_VPWR_c_452_n N_A_467_297#_M1007_s 0.00562358f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_452_n N_A_467_297#_M1019_d 0.00525232f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_456_n N_A_467_297#_c_626_n 0.0225594f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_367 N_VPWR_c_462_n N_A_467_297#_c_628_n 0.0485926f $X=3.575 $Y=2.72 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_452_n N_A_467_297#_c_628_n 0.0307343f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_456_n N_A_467_297#_c_666_n 0.0112071f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_370 N_VPWR_c_462_n N_A_467_297#_c_666_n 0.0116982f $X=3.575 $Y=2.72 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_452_n N_A_467_297#_c_666_n 0.00654447f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_372 N_VPWR_M1005_s N_A_467_297#_c_636_n 0.00351266f $X=3.605 $Y=1.485 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_457_n N_A_467_297#_c_636_n 0.0145016f $X=3.74 $Y=2 $X2=0 $Y2=0
cc_374 N_VPWR_c_464_n N_A_467_297#_c_671_n 0.0113958f $X=4.415 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_452_n N_A_467_297#_c_671_n 0.00646998f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_376 N_VPWR_M1002_d N_A_467_297#_c_641_n 0.00355451f $X=4.445 $Y=1.485 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_458_n N_A_467_297#_c_641_n 0.0145016f $X=4.58 $Y=2 $X2=0 $Y2=0
cc_378 N_VPWR_c_458_n N_A_467_297#_c_645_n 0.0372674f $X=4.58 $Y=2 $X2=0 $Y2=0
cc_379 N_VPWR_c_468_n N_A_467_297#_c_645_n 0.0116048f $X=5.345 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_452_n N_A_467_297#_c_645_n 0.00646998f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_M1003_d N_A_467_297#_c_648_n 0.0180859f $X=5.305 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_459_n N_A_467_297#_c_648_n 0.045605f $X=5.87 $Y=2 $X2=0 $Y2=0
cc_383 N_VPWR_c_460_n N_A_467_297#_c_680_n 0.0113958f $X=6.615 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_452_n N_A_467_297#_c_680_n 0.00646998f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_M1011_s N_A_467_297#_c_624_n 0.0035232f $X=6.645 $Y=1.485 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_461_n N_A_467_297#_c_624_n 0.0145016f $X=6.78 $Y=2 $X2=0 $Y2=0
cc_387 N_VPWR_c_469_n N_A_467_297#_c_684_n 0.0116048f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_452_n N_A_467_297#_c_684_n 0.00646998f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_X_c_582_n N_VGND_M1012_d 8.22501e-19 $X=0.595 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_390 N_X_c_606_p N_VGND_M1012_d 0.0100901f $X=0.235 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_391 X N_VGND_M1012_d 0.00416709f $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_392 N_X_c_574_n N_VGND_M1015_d 0.00337587f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_393 N_X_c_582_n N_VGND_c_687_n 0.00337064f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_394 N_X_c_606_p N_VGND_c_687_n 0.0143265f $X=0.235 $Y=0.805 $X2=0 $Y2=0
cc_395 N_X_c_574_n N_VGND_c_688_n 0.0159625f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_396 N_X_c_574_n N_VGND_c_692_n 0.00244309f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_397 N_X_c_613_p N_VGND_c_692_n 0.0112274f $X=1.52 $Y=0.42 $X2=0 $Y2=0
cc_398 N_X_c_614_p N_VGND_c_696_n 0.0112274f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_399 N_X_c_574_n N_VGND_c_696_n 0.00244309f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_400 N_X_c_582_n N_VGND_c_696_n 0.00244309f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_401 N_X_M1012_s N_VGND_c_699_n 0.00249348f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_402 N_X_M1017_s N_VGND_c_699_n 0.00405853f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_403 N_X_c_614_p N_VGND_c_699_n 0.00643448f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_404 N_X_c_574_n N_VGND_c_699_n 0.00984256f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_405 N_X_c_613_p N_VGND_c_699_n 0.00643448f $X=1.52 $Y=0.42 $X2=0 $Y2=0
cc_406 N_X_c_582_n N_VGND_c_699_n 0.00465289f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_407 N_X_c_606_p N_VGND_c_699_n 8.57032e-19 $X=0.235 $Y=0.805 $X2=0 $Y2=0
cc_408 N_VGND_c_699_n N_A_639_47#_M1001_d 0.00211652f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_409 N_VGND_c_699_n N_A_639_47#_M1026_d 0.00237695f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_699_n N_A_639_47#_M1008_d 0.00212464f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_690_n N_A_639_47#_c_805_n 0.0137364f $X=2.8 $Y=0.38 $X2=0 $Y2=0
cc_412 N_VGND_c_697_n N_A_639_47#_c_805_n 0.0501343f $X=6.615 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_699_n N_A_639_47#_c_805_n 0.0383323f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_697_n N_A_639_47#_c_806_n 0.00238885f $X=6.615 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_699_n N_A_639_47#_c_806_n 0.00560614f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_699_n N_A_889_47#_M1006_s 0.00217615f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_417 N_VGND_c_699_n N_A_889_47#_M1020_d 0.00217615f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_691_n N_A_889_47#_c_831_n 0.00545039f $X=6.78 $Y=0.38 $X2=0
+ $Y2=0
cc_419 N_VGND_c_697_n N_A_889_47#_c_831_n 0.0775216f $X=6.615 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_699_n N_A_889_47#_c_831_n 0.0594678f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_699_n N_A_1079_47#_M1020_s 0.00212464f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_422 N_VGND_c_699_n N_A_1079_47#_M1027_s 0.00319211f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_699_n N_A_1079_47#_M1022_d 0.00369435f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_M1021_s N_A_1079_47#_c_850_n 0.00339267f $X=6.645 $Y=0.235 $X2=0
+ $Y2=0
cc_425 N_VGND_c_691_n N_A_1079_47#_c_850_n 0.0152077f $X=6.78 $Y=0.38 $X2=0
+ $Y2=0
cc_426 N_VGND_c_697_n N_A_1079_47#_c_850_n 0.00757283f $X=6.615 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_698_n N_A_1079_47#_c_850_n 0.00238578f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_699_n N_A_1079_47#_c_850_n 0.020203f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_698_n N_A_1079_47#_c_869_n 0.0114446f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_699_n N_A_1079_47#_c_869_n 0.00643744f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_431 N_A_639_47#_c_806_n N_A_889_47#_M1006_s 0.00339635f $X=5 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_432 N_A_639_47#_M1008_d N_A_889_47#_c_831_n 0.00501197f $X=4.865 $Y=0.235
+ $X2=0 $Y2=0
cc_433 N_A_639_47#_c_806_n N_A_889_47#_c_831_n 0.0372291f $X=5 $Y=0.73 $X2=0
+ $Y2=0
cc_434 N_A_639_47#_c_806_n N_A_1079_47#_c_850_n 0.0145425f $X=5 $Y=0.73 $X2=0
+ $Y2=0
cc_435 N_A_889_47#_c_831_n N_A_1079_47#_M1020_s 0.00482233f $X=5.94 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_436 N_A_889_47#_M1020_d N_A_1079_47#_c_850_n 0.00339635f $X=5.805 $Y=0.235
+ $X2=0 $Y2=0
cc_437 N_A_889_47#_c_831_n N_A_1079_47#_c_850_n 0.0372291f $X=5.94 $Y=0.38 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__dfxtp_4.pxi.spice
* Created: Thu Aug 27 14:16:04 2020
* 
x_PM_SKY130_FD_SC_HD__DFXTP_4%CLK N_CLK_c_179_n N_CLK_c_183_n N_CLK_c_180_n
+ N_CLK_M1024_g N_CLK_c_184_n N_CLK_M1011_g N_CLK_c_185_n CLK CLK
+ PM_SKY130_FD_SC_HD__DFXTP_4%CLK
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_27_47# N_A_27_47#_M1024_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1014_g N_A_27_47#_M1000_g N_A_27_47#_M1022_g N_A_27_47#_c_221_n
+ N_A_27_47#_c_222_n N_A_27_47#_M1006_g N_A_27_47#_M1019_g N_A_27_47#_c_223_n
+ N_A_27_47#_M1027_g N_A_27_47#_c_422_p N_A_27_47#_c_225_n N_A_27_47#_c_226_n
+ N_A_27_47#_c_237_n N_A_27_47#_c_334_p N_A_27_47#_c_227_n N_A_27_47#_c_239_n
+ N_A_27_47#_c_240_n N_A_27_47#_c_241_n N_A_27_47#_c_242_n N_A_27_47#_c_243_n
+ N_A_27_47#_c_244_n N_A_27_47#_c_245_n N_A_27_47#_c_228_n N_A_27_47#_c_247_n
+ N_A_27_47#_c_248_n N_A_27_47#_c_229_n N_A_27_47#_c_230_n
+ PM_SKY130_FD_SC_HD__DFXTP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__DFXTP_4%D N_D_M1001_g N_D_M1018_g D D N_D_c_438_n
+ PM_SKY130_FD_SC_HD__DFXTP_4%D
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_193_47# N_A_193_47#_M1014_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1012_g N_A_193_47#_M1026_g N_A_193_47#_c_473_n
+ N_A_193_47#_M1003_g N_A_193_47#_M1013_g N_A_193_47#_c_474_n
+ N_A_193_47#_c_489_n N_A_193_47#_c_475_n N_A_193_47#_c_476_n
+ N_A_193_47#_c_491_n N_A_193_47#_c_492_n N_A_193_47#_c_477_n
+ N_A_193_47#_c_478_n N_A_193_47#_c_479_n N_A_193_47#_c_591_p
+ N_A_193_47#_c_480_n N_A_193_47#_c_481_n N_A_193_47#_c_482_n
+ N_A_193_47#_c_483_n N_A_193_47#_c_484_n N_A_193_47#_c_485_n
+ PM_SKY130_FD_SC_HD__DFXTP_4%A_193_47#
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_634_183# N_A_634_183#_M1016_d
+ N_A_634_183#_M1002_d N_A_634_183#_M1028_g N_A_634_183#_M1009_g
+ N_A_634_183#_c_660_n N_A_634_183#_c_686_n N_A_634_183#_c_706_p
+ N_A_634_183#_c_687_n N_A_634_183#_c_661_n N_A_634_183#_c_662_n
+ N_A_634_183#_c_674_n N_A_634_183#_c_663_n N_A_634_183#_c_664_n
+ PM_SKY130_FD_SC_HD__DFXTP_4%A_634_183#
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_475_413# N_A_475_413#_M1022_d
+ N_A_475_413#_M1012_d N_A_475_413#_c_753_n N_A_475_413#_M1002_g
+ N_A_475_413#_c_754_n N_A_475_413#_M1016_g N_A_475_413#_c_755_n
+ N_A_475_413#_c_756_n N_A_475_413#_c_757_n N_A_475_413#_c_771_n
+ N_A_475_413#_c_797_n N_A_475_413#_c_758_n N_A_475_413#_c_763_n
+ N_A_475_413#_c_759_n PM_SKY130_FD_SC_HD__DFXTP_4%A_475_413#
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_1062_300# N_A_1062_300#_M1017_s
+ N_A_1062_300#_M1023_s N_A_1062_300#_M1020_g N_A_1062_300#_M1008_g
+ N_A_1062_300#_c_863_n N_A_1062_300#_M1004_g N_A_1062_300#_M1007_g
+ N_A_1062_300#_c_864_n N_A_1062_300#_M1005_g N_A_1062_300#_M1015_g
+ N_A_1062_300#_c_865_n N_A_1062_300#_M1010_g N_A_1062_300#_M1021_g
+ N_A_1062_300#_c_866_n N_A_1062_300#_M1029_g N_A_1062_300#_M1025_g
+ N_A_1062_300#_c_878_n N_A_1062_300#_c_879_n N_A_1062_300#_c_914_p
+ N_A_1062_300#_c_867_n N_A_1062_300#_c_868_n N_A_1062_300#_c_869_n
+ N_A_1062_300#_c_870_n N_A_1062_300#_c_890_p N_A_1062_300#_c_897_p
+ N_A_1062_300#_c_871_n PM_SKY130_FD_SC_HD__DFXTP_4%A_1062_300#
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_891_413# N_A_891_413#_M1003_d
+ N_A_891_413#_M1019_d N_A_891_413#_c_999_n N_A_891_413#_M1017_g
+ N_A_891_413#_M1023_g N_A_891_413#_c_1000_n N_A_891_413#_c_1001_n
+ N_A_891_413#_c_1010_n N_A_891_413#_c_1013_n N_A_891_413#_c_1002_n
+ N_A_891_413#_c_1003_n N_A_891_413#_c_1004_n N_A_891_413#_c_1005_n
+ PM_SKY130_FD_SC_HD__DFXTP_4%A_891_413#
x_PM_SKY130_FD_SC_HD__DFXTP_4%VPWR N_VPWR_M1011_d N_VPWR_M1018_s N_VPWR_M1028_d
+ N_VPWR_M1020_d N_VPWR_M1023_d N_VPWR_M1015_d N_VPWR_M1025_d N_VPWR_c_1081_n
+ N_VPWR_c_1082_n N_VPWR_c_1083_n N_VPWR_c_1084_n N_VPWR_c_1085_n
+ N_VPWR_c_1086_n N_VPWR_c_1087_n N_VPWR_c_1088_n N_VPWR_c_1089_n
+ N_VPWR_c_1090_n N_VPWR_c_1091_n N_VPWR_c_1092_n N_VPWR_c_1093_n
+ N_VPWR_c_1094_n VPWR N_VPWR_c_1095_n N_VPWR_c_1096_n N_VPWR_c_1097_n
+ N_VPWR_c_1098_n N_VPWR_c_1099_n N_VPWR_c_1100_n N_VPWR_c_1101_n
+ N_VPWR_c_1080_n PM_SKY130_FD_SC_HD__DFXTP_4%VPWR
x_PM_SKY130_FD_SC_HD__DFXTP_4%A_381_47# N_A_381_47#_M1001_d N_A_381_47#_M1018_d
+ N_A_381_47#_c_1221_n N_A_381_47#_c_1215_n N_A_381_47#_c_1214_n
+ PM_SKY130_FD_SC_HD__DFXTP_4%A_381_47#
x_PM_SKY130_FD_SC_HD__DFXTP_4%Q N_Q_M1004_s N_Q_M1010_s N_Q_M1007_s N_Q_M1021_s
+ N_Q_c_1249_n N_Q_c_1250_n N_Q_c_1254_n N_Q_c_1272_n N_Q_c_1275_n N_Q_c_1255_n
+ N_Q_c_1251_n N_Q_c_1252_n N_Q_c_1257_n N_Q_c_1253_n N_Q_c_1258_n Q Q Q
+ N_Q_c_1300_n PM_SKY130_FD_SC_HD__DFXTP_4%Q
x_PM_SKY130_FD_SC_HD__DFXTP_4%VGND N_VGND_M1024_d N_VGND_M1001_s N_VGND_M1009_d
+ N_VGND_M1008_d N_VGND_M1017_d N_VGND_M1005_d N_VGND_M1029_d N_VGND_c_1336_n
+ N_VGND_c_1337_n N_VGND_c_1338_n N_VGND_c_1339_n N_VGND_c_1340_n
+ N_VGND_c_1341_n N_VGND_c_1342_n N_VGND_c_1343_n N_VGND_c_1344_n
+ N_VGND_c_1345_n N_VGND_c_1346_n VGND N_VGND_c_1347_n N_VGND_c_1348_n
+ N_VGND_c_1349_n N_VGND_c_1350_n N_VGND_c_1351_n N_VGND_c_1352_n
+ N_VGND_c_1353_n N_VGND_c_1354_n N_VGND_c_1355_n N_VGND_c_1356_n
+ N_VGND_c_1357_n PM_SKY130_FD_SC_HD__DFXTP_4%VGND
cc_1 VNB N_CLK_c_179_n 0.0577303f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.325
cc_2 VNB N_CLK_c_180_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0187424f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1014_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_5 VNB N_A_27_47#_M1022_g 0.0447392f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_6 VNB N_A_27_47#_c_221_n 0.0136466f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_7 VNB N_A_27_47#_c_222_n 0.00223524f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_8 VNB N_A_27_47#_c_223_n 0.0162028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1027_g 0.0472613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_225_n 0.00174761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_226_n 0.00642437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_227_n 0.00246672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_228_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_229_n 0.00980165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_230_n 0.00148891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1001_g 0.0512268f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_17 VNB D 0.00726464f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_18 VNB N_A_193_47#_c_473_n 0.0180517f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_19 VNB N_A_193_47#_c_474_n 0.00330484f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_20 VNB N_A_193_47#_c_475_n 0.00393307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_193_47#_c_476_n 0.00674234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_193_47#_c_477_n 0.0192896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_193_47#_c_478_n 0.00615268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_193_47#_c_479_n 0.0101801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_c_480_n 0.00510919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_481_n 9.18319e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_482_n 0.0266741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_483_n 0.0176138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_c_484_n 0.0285203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_485_n 0.0178295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_634_183#_M1028_g 0.0146965f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_32 VNB N_A_634_183#_M1009_g 0.0210316f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_33 VNB N_A_634_183#_c_660_n 0.00354578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_634_183#_c_661_n 0.00364457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_634_183#_c_662_n 0.00130441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_634_183#_c_663_n 0.00302393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_634_183#_c_664_n 0.0338642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_475_413#_c_753_n 0.0118275f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_39 VNB N_A_475_413#_c_754_n 0.0158415f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_40 VNB N_A_475_413#_c_755_n 0.0152351f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_41 VNB N_A_475_413#_c_756_n 0.00913873f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_42 VNB N_A_475_413#_c_757_n 8.51874e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_475_413#_c_758_n 0.0118177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_475_413#_c_759_n 0.00180949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_1062_300#_M1008_g 0.0534651f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_46 VNB N_A_1062_300#_c_863_n 0.0166449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1062_300#_c_864_n 0.0159904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1062_300#_c_865_n 0.0159887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1062_300#_c_866_n 0.019173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1062_300#_c_867_n 0.010614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1062_300#_c_868_n 0.00175203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1062_300#_c_869_n 6.15295e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1062_300#_c_870_n 0.0122441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1062_300#_c_871_n 0.0669861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_891_413#_c_999_n 0.0216567f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_56 VNB N_A_891_413#_c_1000_n 0.0361219f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_57 VNB N_A_891_413#_c_1001_n 0.00956995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_891_413#_c_1002_n 0.00923386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_891_413#_c_1003_n 0.00118662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_891_413#_c_1004_n 0.0171922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_891_413#_c_1005_n 0.00187583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_1080_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_381_47#_c_1214_n 0.00364179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_Q_c_1249_n 0.00228841f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_65 VNB N_Q_c_1250_n 0.00224394f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_66 VNB N_Q_c_1251_n 0.0102934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_Q_c_1252_n 0.020942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_Q_c_1253_n 0.00224394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1336_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1337_n 0.00817148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1338_n 0.0058544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1339_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1340_n 0.022706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1341_n 0.00472373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1342_n 0.00470426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1343_n 0.0121044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1344_n 0.00469613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1345_n 0.0187183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1346_n 0.0032431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1347_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1348_n 0.0165418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1349_n 0.0450336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1350_n 0.0495175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1351_n 0.0174478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1352_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1353_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1354_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1355_n 0.00324452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1356_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1357_n 0.423948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VPB N_CLK_c_179_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.325
cc_92 VPB N_CLK_c_183_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_93 VPB N_CLK_c_184_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_94 VPB N_CLK_c_185_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_95 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_96 VPB N_A_27_47#_M1000_g 0.037921f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_97 VPB N_A_27_47#_c_221_n 0.0143056f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_98 VPB N_A_27_47#_c_222_n 0.00486539f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_99 VPB N_A_27_47#_M1006_g 0.0191311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_M1019_g 0.033754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_47#_c_223_n 0.023202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_c_237_n 0.00121034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_47#_c_227_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_47#_c_239_n 0.00356676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_c_240_n 0.0259282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_47#_c_241_n 0.00241912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_47#_c_242_n 8.44137e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_c_243_n 0.00143033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_c_244_n 0.00853784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_c_245_n 0.00536377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_228_n 0.0117132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_c_247_n 0.0266783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_27_47#_c_248_n 0.0106236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_27_47#_c_229_n 0.020895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_230_n 0.00437972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_D_M1001_g 0.00151446f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_117 VPB N_D_M1018_g 0.03733f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_118 VPB D 0.00598733f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_119 VPB N_D_c_438_n 0.0438829f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_120 VPB N_A_193_47#_M1012_g 0.0211778f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_121 VPB N_A_193_47#_M1013_g 0.0221869f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_122 VPB N_A_193_47#_c_474_n 0.00406692f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_123 VPB N_A_193_47#_c_489_n 0.0301652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_193_47#_c_475_n 0.00308137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_193_47#_c_491_n 0.00568216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_193_47#_c_492_n 0.0266712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_193_47#_c_485_n 0.0195113f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_634_183#_M1028_g 0.049805f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_129 VPB N_A_634_183#_c_663_n 0.00255179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_475_413#_M1002_g 0.0226707f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_131 VPB N_A_475_413#_c_756_n 0.0189969f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_132 VPB N_A_475_413#_c_757_n 0.00681499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_475_413#_c_763_n 0.00161138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_475_413#_c_759_n 0.00885027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_1062_300#_M1020_g 0.0340711f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_136 VPB N_A_1062_300#_M1008_g 0.0158134f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_137 VPB N_A_1062_300#_M1007_g 0.0193028f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_138 VPB N_A_1062_300#_M1015_g 0.0184805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_1062_300#_M1021_g 0.0184779f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_1062_300#_M1025_g 0.021922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_1062_300#_c_878_n 0.0216566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_1062_300#_c_879_n 0.0418129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_1062_300#_c_869_n 0.00183059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_1062_300#_c_871_n 0.0107424f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_891_413#_M1023_g 0.025978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_891_413#_c_1000_n 0.0125514f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_147 VPB N_A_891_413#_c_1001_n 6.19358e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_891_413#_c_1003_n 0.0155887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_1081_n 0.00105771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_1082_n 0.0082753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_1083_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_1084_n 0.00498288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_1085_n 0.00479834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_1086_n 0.0041827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1087_n 0.0127816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_1088_n 0.0041827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_1089_n 0.0502868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1090_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1091_n 0.0449679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1092_n 0.00410926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1093_n 0.0193207f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1094_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1095_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1096_n 0.0159233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1097_n 0.0276627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1098_n 0.0185662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1099_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1100_n 0.00506925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1101_n 0.00343636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1080_n 0.0718731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_381_47#_c_1215_n 7.45986e-19 $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_172 VPB N_A_381_47#_c_1214_n 0.00511751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_Q_c_1254_n 0.00248773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_Q_c_1255_n 0.0125754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_Q_c_1252_n 0.00834441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_Q_c_1257_n 0.00244705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_Q_c_1258_n 0.00244705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 N_CLK_c_179_n N_A_27_47#_M1014_g 0.00510767f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_179 N_CLK_c_180_n N_A_27_47#_M1014_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_180 CLK N_A_27_47#_M1014_g 3.09846e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_181 N_CLK_c_183_n N_A_27_47#_M1000_g 0.00531917f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_182 N_CLK_c_185_n N_A_27_47#_M1000_g 0.0276478f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_183 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_184 N_CLK_c_179_n N_A_27_47#_c_225_n 0.00787672f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_185 N_CLK_c_180_n N_A_27_47#_c_225_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_186 CLK N_A_27_47#_c_225_n 0.00736322f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_187 N_CLK_c_179_n N_A_27_47#_c_226_n 0.00639426f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_188 CLK N_A_27_47#_c_226_n 0.0144136f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_189 N_CLK_c_184_n N_A_27_47#_c_237_n 0.0128144f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_190 N_CLK_c_185_n N_A_27_47#_c_237_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_191 CLK N_A_27_47#_c_237_n 0.00728212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_192 N_CLK_c_179_n N_A_27_47#_c_227_n 0.00466159f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_193 N_CLK_c_183_n N_A_27_47#_c_227_n 7.09762e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_194 N_CLK_c_185_n N_A_27_47#_c_227_n 0.00440146f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_195 CLK N_A_27_47#_c_227_n 0.0517133f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_196 N_CLK_c_179_n N_A_27_47#_c_239_n 2.26313e-19 $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_197 N_CLK_c_184_n N_A_27_47#_c_239_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_198 N_CLK_c_185_n N_A_27_47#_c_239_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_199 CLK N_A_27_47#_c_239_n 0.0153364f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_200 N_CLK_c_184_n N_A_27_47#_c_241_n 0.00103212f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_201 N_CLK_c_179_n N_A_27_47#_c_228_n 0.0169285f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_202 CLK N_A_27_47#_c_228_n 0.00161876f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_203 N_CLK_c_184_n N_VPWR_c_1081_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_204 N_CLK_c_184_n N_VPWR_c_1095_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_205 N_CLK_c_184_n N_VPWR_c_1080_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_206 N_CLK_c_180_n N_VGND_c_1336_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_207 N_CLK_c_179_n N_VGND_c_1347_n 4.74473e-19 $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_208 N_CLK_c_180_n N_VGND_c_1347_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_209 N_CLK_c_180_n N_VGND_c_1357_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1022_g N_D_M1001_g 0.0168666f $X=2.305 $Y=0.415 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_240_n N_D_M1018_g 0.0103159f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_240_n D 0.00929587f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_222_n N_D_c_438_n 0.0168666f $X=2.38 $Y=1.32 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_240_n N_D_c_438_n 8.87075e-19 $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_228_n N_D_c_438_n 0.00497342f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_240_n N_A_193_47#_M1000_d 6.81311e-19 $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_240_n N_A_193_47#_M1012_g 0.00313687f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_244_n N_A_193_47#_M1012_g 9.6099e-19 $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_247_n N_A_193_47#_M1012_g 0.0144171f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1027_g N_A_193_47#_c_473_n 0.0146445f $X=5.025 $Y=0.415 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_M1019_g N_A_193_47#_M1013_g 0.0175056f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_245_n N_A_193_47#_M1013_g 0.00136781f $X=4.395 $Y=1.87 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_230_n N_A_193_47#_M1013_g 5.16255e-19 $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_M1022_g N_A_193_47#_c_474_n 0.00764677f $X=2.305 $Y=0.415
+ $X2=0 $Y2=0
cc_225 N_A_27_47#_c_221_n N_A_193_47#_c_474_n 0.00687115f $X=2.69 $Y=1.32 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_222_n N_A_193_47#_c_474_n 0.00412863f $X=2.38 $Y=1.32 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_240_n N_A_193_47#_c_474_n 0.0139233f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_244_n N_A_193_47#_c_474_n 0.016922f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_247_n N_A_193_47#_c_474_n 7.29366e-19 $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_248_n N_A_193_47#_c_474_n 0.00604391f $X=2.825 $Y=1.575
+ $X2=0 $Y2=0
cc_231 N_A_27_47#_c_222_n N_A_193_47#_c_489_n 0.0162569f $X=2.38 $Y=1.32 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_240_n N_A_193_47#_c_489_n 0.00465146f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_244_n N_A_193_47#_c_489_n 0.00118389f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_247_n N_A_193_47#_c_489_n 0.0174998f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_223_n N_A_193_47#_c_475_n 0.0118376f $X=4.95 $Y=1.32 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_M1027_g N_A_193_47#_c_475_n 0.00465209f $X=5.025 $Y=0.415
+ $X2=0 $Y2=0
cc_237 N_A_27_47#_c_229_n N_A_193_47#_c_475_n 0.00402309f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_230_n N_A_193_47#_c_475_n 0.0234373f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1027_g N_A_193_47#_c_476_n 0.00274371f $X=5.025 $Y=0.415
+ $X2=0 $Y2=0
cc_240 N_A_27_47#_c_229_n N_A_193_47#_c_476_n 0.00222109f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_230_n N_A_193_47#_c_476_n 0.0119224f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1019_g N_A_193_47#_c_491_n 0.00117691f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_223_n N_A_193_47#_c_491_n 0.00338756f $X=4.95 $Y=1.32 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_245_n N_A_193_47#_c_491_n 0.00513984f $X=4.395 $Y=1.87 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_230_n N_A_193_47#_c_491_n 0.0245563f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_M1019_g N_A_193_47#_c_492_n 0.0130792f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_223_n N_A_193_47#_c_492_n 0.0218248f $X=4.95 $Y=1.32 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_230_n N_A_193_47#_c_492_n 6.54911e-19 $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1022_g N_A_193_47#_c_477_n 9.97044e-19 $X=2.305 $Y=0.415
+ $X2=0 $Y2=0
cc_250 N_A_27_47#_M1014_g N_A_193_47#_c_478_n 0.00654297f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_225_n N_A_193_47#_c_478_n 0.00215348f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_227_n N_A_193_47#_c_478_n 0.00507209f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_229_n N_A_193_47#_c_479_n 2.10748e-19 $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1022_g N_A_193_47#_c_480_n 0.011756f $X=2.305 $Y=0.415 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_221_n N_A_193_47#_c_480_n 0.00587088f $X=2.69 $Y=1.32 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_244_n N_A_193_47#_c_480_n 0.00398178f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_229_n N_A_193_47#_c_481_n 9.82747e-19 $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_230_n N_A_193_47#_c_481_n 0.00125233f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1022_g N_A_193_47#_c_482_n 0.0213105f $X=2.305 $Y=0.415 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_221_n N_A_193_47#_c_482_n 0.0174066f $X=2.69 $Y=1.32 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_244_n N_A_193_47#_c_482_n 4.76262e-19 $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_247_n N_A_193_47#_c_482_n 5.43883e-19 $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1022_g N_A_193_47#_c_483_n 0.0102605f $X=2.305 $Y=0.415 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1027_g N_A_193_47#_c_484_n 0.0193601f $X=5.025 $Y=0.415 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_229_n N_A_193_47#_c_484_n 0.020308f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1014_g N_A_193_47#_c_485_n 0.0232514f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_225_n N_A_193_47#_c_485_n 0.011891f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_334_p N_A_193_47#_c_485_n 0.00826851f $X=0.725 $Y=1.795
+ $X2=0 $Y2=0
cc_269 N_A_27_47#_c_227_n N_A_193_47#_c_485_n 0.0701354f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_240_n N_A_193_47#_c_485_n 0.0267497f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_241_n N_A_193_47#_c_485_n 0.00185693f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_242_n N_A_634_183#_M1002_d 0.00523078f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_221_n N_A_634_183#_M1028_g 0.0113457f $X=2.69 $Y=1.32 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1006_g N_A_634_183#_M1028_g 0.0276008f $X=2.765 $Y=2.275
+ $X2=0 $Y2=0
cc_275 N_A_27_47#_c_242_n N_A_634_183#_M1028_g 0.00281129f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_243_n N_A_634_183#_M1028_g 0.00153318f $X=3.16 $Y=1.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_244_n N_A_634_183#_M1028_g 0.0022f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_247_n N_A_634_183#_M1028_g 0.0206011f $X=2.825 $Y=1.74 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_242_n N_A_634_183#_c_674_n 0.00261642f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1019_g N_A_634_183#_c_663_n 0.00455971f $X=4.38 $Y=2.275
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_242_n N_A_634_183#_c_663_n 0.0193938f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_245_n N_A_634_183#_c_663_n 0.00311096f $X=4.395 $Y=1.87
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_229_n N_A_634_183#_c_663_n 0.00225153f $X=4.375 $Y=1.32
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_c_230_n N_A_634_183#_c_663_n 0.0517157f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_229_n N_A_475_413#_c_753_n 0.0158005f $X=4.375 $Y=1.32 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_230_n N_A_475_413#_c_753_n 3.03019e-19 $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_M1019_g N_A_475_413#_M1002_g 0.0247799f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_242_n N_A_475_413#_M1002_g 0.00700233f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_230_n N_A_475_413#_M1002_g 8.29633e-19 $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_242_n N_A_475_413#_c_756_n 0.00109659f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_M1006_g N_A_475_413#_c_771_n 0.00859956f $X=2.765 $Y=2.275
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_240_n N_A_475_413#_c_771_n 0.00714382f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_242_n N_A_475_413#_c_771_n 0.00257439f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_243_n N_A_475_413#_c_771_n 0.00275128f $X=3.16 $Y=1.87 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_244_n N_A_475_413#_c_771_n 0.0252894f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_247_n N_A_475_413#_c_771_n 5.38487e-19 $X=2.825 $Y=1.74
+ $X2=0 $Y2=0
cc_297 N_A_27_47#_M1022_g N_A_475_413#_c_758_n 9.86268e-19 $X=2.305 $Y=0.415
+ $X2=0 $Y2=0
cc_298 N_A_27_47#_c_221_n N_A_475_413#_c_758_n 8.14452e-19 $X=2.69 $Y=1.32 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1006_g N_A_475_413#_c_763_n 9.97608e-19 $X=2.765 $Y=2.275
+ $X2=0 $Y2=0
cc_300 N_A_27_47#_c_242_n N_A_475_413#_c_763_n 0.0183205f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_243_n N_A_475_413#_c_763_n 0.00270727f $X=3.16 $Y=1.87 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_244_n N_A_475_413#_c_763_n 0.0249708f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_247_n N_A_475_413#_c_763_n 7.00613e-19 $X=2.825 $Y=1.74
+ $X2=0 $Y2=0
cc_304 N_A_27_47#_c_221_n N_A_475_413#_c_759_n 0.00225879f $X=2.69 $Y=1.32 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_242_n N_A_475_413#_c_759_n 0.0156267f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_243_n N_A_475_413#_c_759_n 0.00371621f $X=3.16 $Y=1.87 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_244_n N_A_475_413#_c_759_n 0.00980238f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_248_n N_A_475_413#_c_759_n 4.44848e-19 $X=2.825 $Y=1.575
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_M1027_g N_A_1062_300#_M1008_g 0.0419344f $X=5.025 $Y=0.415
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_M1019_g N_A_891_413#_c_1010_n 0.00281529f $X=4.38 $Y=2.275
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_245_n N_A_891_413#_c_1010_n 0.00241029f $X=4.395 $Y=1.87
+ $X2=0 $Y2=0
cc_312 N_A_27_47#_c_230_n N_A_891_413#_c_1010_n 0.0022468f $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_M1027_g N_A_891_413#_c_1013_n 0.0125837f $X=5.025 $Y=0.415
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_M1027_g N_A_891_413#_c_1002_n 0.00659966f $X=5.025 $Y=0.415
+ $X2=0 $Y2=0
cc_315 N_A_27_47#_c_223_n N_A_891_413#_c_1003_n 0.00176978f $X=4.95 $Y=1.32
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_245_n N_A_891_413#_c_1003_n 0.00230468f $X=4.395 $Y=1.87
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_c_230_n N_A_891_413#_c_1003_n 9.59883e-19 $X=4.375 $Y=1.41
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_M1027_g N_A_891_413#_c_1005_n 0.00196411f $X=5.025 $Y=0.415
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_334_p N_VPWR_M1011_d 6.91013e-19 $X=0.725 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_320 N_A_27_47#_c_241_n N_VPWR_M1011_d 0.00195102f $X=0.84 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_321 N_A_27_47#_c_242_n N_VPWR_M1028_d 0.00678497f $X=4.25 $Y=1.87 $X2=0 $Y2=0
cc_322 N_A_27_47#_M1000_g N_VPWR_c_1081_n 0.0082523f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_237_n N_VPWR_c_1081_n 0.00355272f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_334_p N_VPWR_c_1081_n 0.0133497f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_239_n N_VPWR_c_1081_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_241_n N_VPWR_c_1081_n 0.00347913f $X=0.84 $Y=1.87 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_M1000_g N_VPWR_c_1082_n 0.00180698f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_240_n N_VPWR_c_1082_n 0.00413138f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_242_n N_VPWR_c_1083_n 0.00950843f $X=4.25 $Y=1.87 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_M1006_g N_VPWR_c_1089_n 0.0037886f $X=2.765 $Y=2.275 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_M1019_g N_VPWR_c_1091_n 0.00430107f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_230_n N_VPWR_c_1091_n 0.00157744f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_237_n N_VPWR_c_1095_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_239_n N_VPWR_c_1095_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_335 N_A_27_47#_M1000_g N_VPWR_c_1096_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_M1000_g N_VPWR_c_1080_n 0.00536257f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_M1006_g N_VPWR_c_1080_n 0.00557714f $X=2.765 $Y=2.275 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_M1019_g N_VPWR_c_1080_n 0.0057371f $X=4.38 $Y=2.275 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_237_n N_VPWR_c_1080_n 0.00396423f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_239_n N_VPWR_c_1080_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_240_n N_VPWR_c_1080_n 0.0988846f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_342 N_A_27_47#_c_241_n N_VPWR_c_1080_n 0.0144757f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_242_n N_VPWR_c_1080_n 0.0515095f $X=4.25 $Y=1.87 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_243_n N_VPWR_c_1080_n 0.0149246f $X=3.16 $Y=1.87 $X2=0 $Y2=0
cc_345 N_A_27_47#_c_245_n N_VPWR_c_1080_n 0.0159163f $X=4.395 $Y=1.87 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_230_n N_VPWR_c_1080_n 0.00100625f $X=4.375 $Y=1.41 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_240_n N_A_381_47#_c_1215_n 0.00234842f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_M1022_g N_A_381_47#_c_1214_n 0.00680074f $X=2.305 $Y=0.415
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_240_n N_A_381_47#_c_1214_n 0.0214082f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_244_n N_A_381_47#_c_1214_n 0.00292246f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_225_n N_VGND_M1024_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_352 N_A_27_47#_M1014_g N_VGND_c_1336_n 0.0078844f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_225_n N_VGND_c_1336_n 0.0170164f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_228_n N_VGND_c_1336_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_M1014_g N_VGND_c_1337_n 0.00304372f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_422_p N_VGND_c_1347_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_225_n N_VGND_c_1347_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1014_g N_VGND_c_1348_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1022_g N_VGND_c_1349_n 0.00435108f $X=2.305 $Y=0.415 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_M1027_g N_VGND_c_1350_n 0.0037981f $X=5.025 $Y=0.415 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_M1024_s N_VGND_c_1357_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_M1014_g N_VGND_c_1357_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_M1022_g N_VGND_c_1357_n 0.006034f $X=2.305 $Y=0.415 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_M1027_g N_VGND_c_1357_n 0.00575801f $X=5.025 $Y=0.415 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_422_p N_VGND_c_1357_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_225_n N_VGND_c_1357_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_367 N_D_M1018_g N_A_193_47#_M1012_g 0.013616f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_368 N_D_M1001_g N_A_193_47#_c_474_n 3.61314e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_369 N_D_c_438_n N_A_193_47#_c_474_n 0.00134637f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_370 N_D_c_438_n N_A_193_47#_c_489_n 0.0140728f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_371 N_D_M1001_g N_A_193_47#_c_477_n 0.0103159f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_372 D N_A_193_47#_c_477_n 0.00986021f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_373 N_D_c_438_n N_A_193_47#_c_477_n 7.52422e-19 $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_374 N_D_M1001_g N_A_193_47#_c_478_n 0.00181416f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_375 N_D_M1001_g N_A_193_47#_c_480_n 3.97833e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_376 N_D_M1001_g N_A_193_47#_c_485_n 0.0075997f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_377 N_D_M1018_g N_A_193_47#_c_485_n 0.00729808f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_378 D N_A_193_47#_c_485_n 0.0427669f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_379 N_D_c_438_n N_A_193_47#_c_485_n 0.00114684f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_380 N_D_M1018_g N_VPWR_c_1082_n 0.00451231f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_381 D N_VPWR_c_1082_n 0.00430704f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_382 N_D_c_438_n N_VPWR_c_1082_n 0.00130415f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_383 N_D_M1018_g N_VPWR_c_1089_n 0.00564615f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_384 N_D_M1018_g N_VPWR_c_1080_n 0.00763133f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_385 N_D_M1001_g N_A_381_47#_c_1221_n 0.00197415f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_386 N_D_M1018_g N_A_381_47#_c_1215_n 0.00535586f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_387 N_D_M1001_g N_A_381_47#_c_1214_n 0.0187795f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_388 N_D_M1018_g N_A_381_47#_c_1214_n 0.0104656f $X=1.83 $Y=2.275 $X2=0 $Y2=0
cc_389 D N_A_381_47#_c_1214_n 0.0433322f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_390 N_D_c_438_n N_A_381_47#_c_1214_n 0.00952781f $X=1.83 $Y=1.5 $X2=0 $Y2=0
cc_391 N_D_M1001_g N_VGND_c_1337_n 0.0044954f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_392 D N_VGND_c_1337_n 0.00430459f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_393 N_D_M1001_g N_VGND_c_1349_n 0.00564827f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_394 N_D_M1001_g N_VGND_c_1357_n 0.00763092f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_395 N_A_193_47#_c_476_n N_A_634_183#_M1016_d 0.00133652f $X=4.65 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_396 N_A_193_47#_c_479_n N_A_634_183#_M1016_d 9.65449e-19 $X=4.25 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_397 N_A_193_47#_c_481_n N_A_634_183#_M1016_d 6.4695e-19 $X=4.395 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_398 N_A_193_47#_c_479_n N_A_634_183#_M1009_g 0.00208483f $X=4.25 $Y=0.85
+ $X2=0 $Y2=0
cc_399 N_A_193_47#_c_483_n N_A_634_183#_M1009_g 0.013781f $X=2.725 $Y=0.705
+ $X2=0 $Y2=0
cc_400 N_A_193_47#_c_479_n N_A_634_183#_c_660_n 0.0221014f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_401 N_A_193_47#_c_481_n N_A_634_183#_c_686_n 8.93965e-19 $X=4.395 $Y=0.85
+ $X2=0 $Y2=0
cc_402 N_A_193_47#_c_476_n N_A_634_183#_c_687_n 0.00716698f $X=4.65 $Y=0.87
+ $X2=0 $Y2=0
cc_403 N_A_193_47#_c_479_n N_A_634_183#_c_687_n 0.00363224f $X=4.25 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_193_47#_c_481_n N_A_634_183#_c_687_n 0.00168986f $X=4.395 $Y=0.85
+ $X2=0 $Y2=0
cc_405 N_A_193_47#_c_479_n N_A_634_183#_c_661_n 0.00899288f $X=4.25 $Y=0.85
+ $X2=0 $Y2=0
cc_406 N_A_193_47#_c_475_n N_A_634_183#_c_662_n 0.00114045f $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_407 N_A_193_47#_c_476_n N_A_634_183#_c_662_n 0.018732f $X=4.65 $Y=0.87 $X2=0
+ $Y2=0
cc_408 N_A_193_47#_c_479_n N_A_634_183#_c_662_n 0.0176435f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_409 N_A_193_47#_c_481_n N_A_634_183#_c_662_n 0.00185392f $X=4.395 $Y=0.85
+ $X2=0 $Y2=0
cc_410 N_A_193_47#_c_484_n N_A_634_183#_c_662_n 5.82389e-19 $X=4.605 $Y=0.87
+ $X2=0 $Y2=0
cc_411 N_A_193_47#_c_475_n N_A_634_183#_c_663_n 0.00620052f $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_412 N_A_193_47#_c_479_n N_A_634_183#_c_664_n 0.00299829f $X=4.25 $Y=0.85
+ $X2=0 $Y2=0
cc_413 N_A_193_47#_c_482_n N_A_634_183#_c_664_n 0.0179412f $X=2.725 $Y=0.87
+ $X2=0 $Y2=0
cc_414 N_A_193_47#_c_475_n N_A_475_413#_c_753_n 6.31337e-19 $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_415 N_A_193_47#_c_473_n N_A_475_413#_c_754_n 0.00957285f $X=4.51 $Y=0.705
+ $X2=0 $Y2=0
cc_416 N_A_193_47#_c_476_n N_A_475_413#_c_754_n 0.00100831f $X=4.65 $Y=0.87
+ $X2=0 $Y2=0
cc_417 N_A_193_47#_c_475_n N_A_475_413#_c_755_n 3.37852e-19 $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_418 N_A_193_47#_c_484_n N_A_475_413#_c_755_n 0.00957285f $X=4.605 $Y=0.87
+ $X2=0 $Y2=0
cc_419 N_A_193_47#_M1012_g N_A_475_413#_c_771_n 0.0017787f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_420 N_A_193_47#_c_474_n N_A_475_413#_c_771_n 0.00286257f $X=2.315 $Y=1.74
+ $X2=0 $Y2=0
cc_421 N_A_193_47#_c_489_n N_A_475_413#_c_771_n 6.94615e-19 $X=2.315 $Y=1.74
+ $X2=0 $Y2=0
cc_422 N_A_193_47#_c_479_n N_A_475_413#_c_797_n 0.00489874f $X=4.25 $Y=0.85
+ $X2=0 $Y2=0
cc_423 N_A_193_47#_c_591_p N_A_475_413#_c_797_n 0.00119052f $X=2.7 $Y=0.85 $X2=0
+ $Y2=0
cc_424 N_A_193_47#_c_480_n N_A_475_413#_c_797_n 0.0241387f $X=2.555 $Y=0.85
+ $X2=0 $Y2=0
cc_425 N_A_193_47#_c_482_n N_A_475_413#_c_797_n 0.00256542f $X=2.725 $Y=0.87
+ $X2=0 $Y2=0
cc_426 N_A_193_47#_c_483_n N_A_475_413#_c_797_n 0.00840911f $X=2.725 $Y=0.705
+ $X2=0 $Y2=0
cc_427 N_A_193_47#_c_474_n N_A_475_413#_c_758_n 0.00981359f $X=2.315 $Y=1.74
+ $X2=0 $Y2=0
cc_428 N_A_193_47#_c_479_n N_A_475_413#_c_758_n 0.0188221f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_429 N_A_193_47#_c_591_p N_A_475_413#_c_758_n 5.13248e-19 $X=2.7 $Y=0.85 $X2=0
+ $Y2=0
cc_430 N_A_193_47#_c_480_n N_A_475_413#_c_758_n 0.0239322f $X=2.555 $Y=0.85
+ $X2=0 $Y2=0
cc_431 N_A_193_47#_c_483_n N_A_475_413#_c_758_n 0.00604394f $X=2.725 $Y=0.705
+ $X2=0 $Y2=0
cc_432 N_A_193_47#_c_474_n N_A_475_413#_c_759_n 0.00649323f $X=2.315 $Y=1.74
+ $X2=0 $Y2=0
cc_433 N_A_193_47#_c_479_n N_A_475_413#_c_759_n 0.00803733f $X=4.25 $Y=0.85
+ $X2=0 $Y2=0
cc_434 N_A_193_47#_M1013_g N_A_1062_300#_M1020_g 0.0179923f $X=4.8 $Y=2.275
+ $X2=0 $Y2=0
cc_435 N_A_193_47#_c_492_n N_A_1062_300#_c_879_n 0.0118218f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_436 N_A_193_47#_M1013_g N_A_891_413#_c_1010_n 0.00974744f $X=4.8 $Y=2.275
+ $X2=0 $Y2=0
cc_437 N_A_193_47#_c_491_n N_A_891_413#_c_1010_n 0.012999f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_438 N_A_193_47#_c_492_n N_A_891_413#_c_1010_n 0.00300896f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_439 N_A_193_47#_c_476_n N_A_891_413#_c_1013_n 0.0153172f $X=4.65 $Y=0.87
+ $X2=0 $Y2=0
cc_440 N_A_193_47#_c_484_n N_A_891_413#_c_1013_n 8.54271e-19 $X=4.605 $Y=0.87
+ $X2=0 $Y2=0
cc_441 N_A_193_47#_c_475_n N_A_891_413#_c_1002_n 0.00199251f $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_442 N_A_193_47#_c_476_n N_A_891_413#_c_1002_n 0.017354f $X=4.65 $Y=0.87 $X2=0
+ $Y2=0
cc_443 N_A_193_47#_c_481_n N_A_891_413#_c_1002_n 9.56356e-19 $X=4.395 $Y=0.85
+ $X2=0 $Y2=0
cc_444 N_A_193_47#_M1013_g N_A_891_413#_c_1003_n 0.0046302f $X=4.8 $Y=2.275
+ $X2=0 $Y2=0
cc_445 N_A_193_47#_c_475_n N_A_891_413#_c_1003_n 0.0162763f $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_446 N_A_193_47#_c_491_n N_A_891_413#_c_1003_n 0.024681f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_447 N_A_193_47#_c_492_n N_A_891_413#_c_1003_n 0.00187857f $X=4.885 $Y=1.74
+ $X2=0 $Y2=0
cc_448 N_A_193_47#_c_475_n N_A_891_413#_c_1005_n 0.00971483f $X=4.745 $Y=1.575
+ $X2=0 $Y2=0
cc_449 N_A_193_47#_c_485_n N_VPWR_c_1081_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_450 N_A_193_47#_c_485_n N_VPWR_c_1082_n 0.0205851f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_451 N_A_193_47#_M1012_g N_VPWR_c_1089_n 0.005785f $X=2.3 $Y=2.275 $X2=0 $Y2=0
cc_452 N_A_193_47#_M1013_g N_VPWR_c_1091_n 0.00383564f $X=4.8 $Y=2.275 $X2=0
+ $Y2=0
cc_453 N_A_193_47#_c_485_n N_VPWR_c_1096_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_454 N_A_193_47#_M1012_g N_VPWR_c_1080_n 0.00612376f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_455 N_A_193_47#_M1013_g N_VPWR_c_1080_n 0.00579176f $X=4.8 $Y=2.275 $X2=0
+ $Y2=0
cc_456 N_A_193_47#_c_474_n N_VPWR_c_1080_n 0.00189161f $X=2.315 $Y=1.74 $X2=0
+ $Y2=0
cc_457 N_A_193_47#_c_489_n N_VPWR_c_1080_n 4.15345e-19 $X=2.315 $Y=1.74 $X2=0
+ $Y2=0
cc_458 N_A_193_47#_c_485_n N_VPWR_c_1080_n 0.00409094f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_459 N_A_193_47#_c_477_n N_A_381_47#_c_1221_n 0.0047557f $X=2.41 $Y=0.85 $X2=0
+ $Y2=0
cc_460 N_A_193_47#_M1012_g N_A_381_47#_c_1215_n 0.0048729f $X=2.3 $Y=2.275 $X2=0
+ $Y2=0
cc_461 N_A_193_47#_M1012_g N_A_381_47#_c_1214_n 0.00231702f $X=2.3 $Y=2.275
+ $X2=0 $Y2=0
cc_462 N_A_193_47#_c_474_n N_A_381_47#_c_1214_n 0.0640433f $X=2.315 $Y=1.74
+ $X2=0 $Y2=0
cc_463 N_A_193_47#_c_489_n N_A_381_47#_c_1214_n 0.00171737f $X=2.315 $Y=1.74
+ $X2=0 $Y2=0
cc_464 N_A_193_47#_c_477_n N_A_381_47#_c_1214_n 0.0193509f $X=2.41 $Y=0.85 $X2=0
+ $Y2=0
cc_465 N_A_193_47#_c_478_n N_A_381_47#_c_1214_n 0.00189056f $X=1.3 $Y=0.85 $X2=0
+ $Y2=0
cc_466 N_A_193_47#_c_591_p N_A_381_47#_c_1214_n 4.43882e-19 $X=2.7 $Y=0.85 $X2=0
+ $Y2=0
cc_467 N_A_193_47#_c_480_n N_A_381_47#_c_1214_n 0.0240253f $X=2.555 $Y=0.85
+ $X2=0 $Y2=0
cc_468 N_A_193_47#_c_485_n N_A_381_47#_c_1214_n 0.022122f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_469 N_A_193_47#_c_477_n N_VGND_c_1337_n 0.0039309f $X=2.41 $Y=0.85 $X2=0
+ $Y2=0
cc_470 N_A_193_47#_c_485_n N_VGND_c_1337_n 0.0134396f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_471 N_A_193_47#_c_479_n N_VGND_c_1338_n 0.00197288f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_472 N_A_193_47#_c_485_n N_VGND_c_1348_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_473 N_A_193_47#_c_480_n N_VGND_c_1349_n 0.00252373f $X=2.555 $Y=0.85 $X2=0
+ $Y2=0
cc_474 N_A_193_47#_c_483_n N_VGND_c_1349_n 0.0037981f $X=2.725 $Y=0.705 $X2=0
+ $Y2=0
cc_475 N_A_193_47#_c_473_n N_VGND_c_1350_n 0.00435108f $X=4.51 $Y=0.705 $X2=0
+ $Y2=0
cc_476 N_A_193_47#_c_476_n N_VGND_c_1350_n 0.00341023f $X=4.65 $Y=0.87 $X2=0
+ $Y2=0
cc_477 N_A_193_47#_c_484_n N_VGND_c_1350_n 8.04624e-19 $X=4.605 $Y=0.87 $X2=0
+ $Y2=0
cc_478 N_A_193_47#_M1014_d N_VGND_c_1357_n 0.0033946f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_479 N_A_193_47#_c_473_n N_VGND_c_1357_n 0.00623562f $X=4.51 $Y=0.705 $X2=0
+ $Y2=0
cc_480 N_A_193_47#_c_476_n N_VGND_c_1357_n 0.00402561f $X=4.65 $Y=0.87 $X2=0
+ $Y2=0
cc_481 N_A_193_47#_c_477_n N_VGND_c_1357_n 0.0536241f $X=2.41 $Y=0.85 $X2=0
+ $Y2=0
cc_482 N_A_193_47#_c_478_n N_VGND_c_1357_n 0.0151433f $X=1.3 $Y=0.85 $X2=0 $Y2=0
cc_483 N_A_193_47#_c_479_n N_VGND_c_1357_n 0.0711725f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_484 N_A_193_47#_c_591_p N_VGND_c_1357_n 0.0146104f $X=2.7 $Y=0.85 $X2=0 $Y2=0
cc_485 N_A_193_47#_c_480_n N_VGND_c_1357_n 0.00247006f $X=2.555 $Y=0.85 $X2=0
+ $Y2=0
cc_486 N_A_193_47#_c_481_n N_VGND_c_1357_n 0.0147739f $X=4.395 $Y=0.85 $X2=0
+ $Y2=0
cc_487 N_A_193_47#_c_483_n N_VGND_c_1357_n 0.00563926f $X=2.725 $Y=0.705 $X2=0
+ $Y2=0
cc_488 N_A_193_47#_c_484_n N_VGND_c_1357_n 0.00134095f $X=4.605 $Y=0.87 $X2=0
+ $Y2=0
cc_489 N_A_193_47#_c_485_n N_VGND_c_1357_n 0.00372614f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_490 N_A_634_183#_c_663_n N_A_475_413#_c_753_n 0.00595764f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_491 N_A_634_183#_M1028_g N_A_475_413#_M1002_g 0.0139082f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_492 N_A_634_183#_c_674_n N_A_475_413#_M1002_g 0.00378805f $X=4.115 $Y=2.3
+ $X2=0 $Y2=0
cc_493 N_A_634_183#_c_663_n N_A_475_413#_M1002_g 0.0122998f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_494 N_A_634_183#_M1009_g N_A_475_413#_c_754_n 0.0109128f $X=3.275 $Y=0.445
+ $X2=0 $Y2=0
cc_495 N_A_634_183#_c_660_n N_A_475_413#_c_754_n 0.00351053f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_496 N_A_634_183#_c_686_n N_A_475_413#_c_754_n 0.00675936f $X=4.035 $Y=0.765
+ $X2=0 $Y2=0
cc_497 N_A_634_183#_c_706_p N_A_475_413#_c_754_n 0.004701f $X=4.12 $Y=0.45 $X2=0
+ $Y2=0
cc_498 N_A_634_183#_c_662_n N_A_475_413#_c_754_n 0.00333126f $X=4.035 $Y=0.915
+ $X2=0 $Y2=0
cc_499 N_A_634_183#_c_664_n N_A_475_413#_c_754_n 0.00500517f $X=3.275 $Y=0.93
+ $X2=0 $Y2=0
cc_500 N_A_634_183#_M1028_g N_A_475_413#_c_755_n 0.00398999f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_501 N_A_634_183#_c_660_n N_A_475_413#_c_755_n 0.00996228f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_502 N_A_634_183#_c_661_n N_A_475_413#_c_755_n 2.46578e-19 $X=3.49 $Y=0.93
+ $X2=0 $Y2=0
cc_503 N_A_634_183#_c_662_n N_A_475_413#_c_755_n 0.00234347f $X=4.035 $Y=0.915
+ $X2=0 $Y2=0
cc_504 N_A_634_183#_c_663_n N_A_475_413#_c_755_n 0.00394884f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_505 N_A_634_183#_c_664_n N_A_475_413#_c_755_n 0.00573363f $X=3.275 $Y=0.93
+ $X2=0 $Y2=0
cc_506 N_A_634_183#_M1028_g N_A_475_413#_c_756_n 0.0173592f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_507 N_A_634_183#_c_660_n N_A_475_413#_c_756_n 0.00400764f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_508 N_A_634_183#_c_664_n N_A_475_413#_c_756_n 0.00238133f $X=3.275 $Y=0.93
+ $X2=0 $Y2=0
cc_509 N_A_634_183#_c_663_n N_A_475_413#_c_757_n 0.00611615f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_510 N_A_634_183#_M1028_g N_A_475_413#_c_771_n 0.0101048f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_511 N_A_634_183#_M1009_g N_A_475_413#_c_758_n 0.00441151f $X=3.275 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_634_183#_c_661_n N_A_475_413#_c_758_n 0.0242417f $X=3.49 $Y=0.93
+ $X2=0 $Y2=0
cc_513 N_A_634_183#_c_664_n N_A_475_413#_c_758_n 0.0095167f $X=3.275 $Y=0.93
+ $X2=0 $Y2=0
cc_514 N_A_634_183#_M1028_g N_A_475_413#_c_763_n 0.0153748f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_515 N_A_634_183#_c_663_n N_A_475_413#_c_763_n 0.00754007f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_516 N_A_634_183#_M1028_g N_A_475_413#_c_759_n 0.0138593f $X=3.245 $Y=2.275
+ $X2=0 $Y2=0
cc_517 N_A_634_183#_c_660_n N_A_475_413#_c_759_n 0.0186614f $X=3.95 $Y=0.915
+ $X2=0 $Y2=0
cc_518 N_A_634_183#_c_661_n N_A_475_413#_c_759_n 0.0112018f $X=3.49 $Y=0.93
+ $X2=0 $Y2=0
cc_519 N_A_634_183#_c_663_n N_A_475_413#_c_759_n 0.0245884f $X=4.075 $Y=2.135
+ $X2=0 $Y2=0
cc_520 N_A_634_183#_c_664_n N_A_475_413#_c_759_n 0.00213749f $X=3.275 $Y=0.93
+ $X2=0 $Y2=0
cc_521 N_A_634_183#_c_674_n N_A_891_413#_c_1010_n 0.0109209f $X=4.115 $Y=2.3
+ $X2=0 $Y2=0
cc_522 N_A_634_183#_M1028_g N_VPWR_c_1083_n 0.0057281f $X=3.245 $Y=2.275 $X2=0
+ $Y2=0
cc_523 N_A_634_183#_c_663_n N_VPWR_c_1083_n 0.0237f $X=4.075 $Y=2.135 $X2=0
+ $Y2=0
cc_524 N_A_634_183#_M1028_g N_VPWR_c_1089_n 0.00378797f $X=3.245 $Y=2.275 $X2=0
+ $Y2=0
cc_525 N_A_634_183#_c_674_n N_VPWR_c_1091_n 0.015079f $X=4.115 $Y=2.3 $X2=0
+ $Y2=0
cc_526 N_A_634_183#_M1002_d N_VPWR_c_1080_n 0.00285796f $X=3.98 $Y=1.735 $X2=0
+ $Y2=0
cc_527 N_A_634_183#_M1028_g N_VPWR_c_1080_n 0.00596544f $X=3.245 $Y=2.275 $X2=0
+ $Y2=0
cc_528 N_A_634_183#_c_674_n N_VPWR_c_1080_n 0.00439826f $X=4.115 $Y=2.3 $X2=0
+ $Y2=0
cc_529 N_A_634_183#_c_660_n N_VGND_M1009_d 0.00306998f $X=3.95 $Y=0.915 $X2=0
+ $Y2=0
cc_530 N_A_634_183#_M1009_g N_VGND_c_1338_n 0.00603751f $X=3.275 $Y=0.445 $X2=0
+ $Y2=0
cc_531 N_A_634_183#_c_686_n N_VGND_c_1338_n 0.00354103f $X=4.035 $Y=0.765 $X2=0
+ $Y2=0
cc_532 N_A_634_183#_c_706_p N_VGND_c_1338_n 0.013122f $X=4.12 $Y=0.45 $X2=0
+ $Y2=0
cc_533 N_A_634_183#_c_661_n N_VGND_c_1338_n 0.0258565f $X=3.49 $Y=0.93 $X2=0
+ $Y2=0
cc_534 N_A_634_183#_c_664_n N_VGND_c_1338_n 0.00122075f $X=3.275 $Y=0.93 $X2=0
+ $Y2=0
cc_535 N_A_634_183#_M1009_g N_VGND_c_1349_n 0.00585385f $X=3.275 $Y=0.445 $X2=0
+ $Y2=0
cc_536 N_A_634_183#_c_706_p N_VGND_c_1350_n 0.00594819f $X=4.12 $Y=0.45 $X2=0
+ $Y2=0
cc_537 N_A_634_183#_c_687_n N_VGND_c_1350_n 0.0100275f $X=4.245 $Y=0.45 $X2=0
+ $Y2=0
cc_538 N_A_634_183#_M1016_d N_VGND_c_1357_n 0.00246577f $X=4.08 $Y=0.235 $X2=0
+ $Y2=0
cc_539 N_A_634_183#_M1009_g N_VGND_c_1357_n 0.0070154f $X=3.275 $Y=0.445 $X2=0
+ $Y2=0
cc_540 N_A_634_183#_c_660_n N_VGND_c_1357_n 0.0042145f $X=3.95 $Y=0.915 $X2=0
+ $Y2=0
cc_541 N_A_634_183#_c_706_p N_VGND_c_1357_n 0.00261981f $X=4.12 $Y=0.45 $X2=0
+ $Y2=0
cc_542 N_A_634_183#_c_687_n N_VGND_c_1357_n 0.00441842f $X=4.245 $Y=0.45 $X2=0
+ $Y2=0
cc_543 N_A_634_183#_c_661_n N_VGND_c_1357_n 0.00269026f $X=3.49 $Y=0.93 $X2=0
+ $Y2=0
cc_544 N_A_475_413#_c_771_n N_VPWR_M1028_d 0.00236303f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_545 N_A_475_413#_c_763_n N_VPWR_M1028_d 0.00412006f $X=3.355 $Y=2.19 $X2=0
+ $Y2=0
cc_546 N_A_475_413#_M1002_g N_VPWR_c_1083_n 0.00314007f $X=3.905 $Y=2.11 $X2=0
+ $Y2=0
cc_547 N_A_475_413#_c_756_n N_VPWR_c_1083_n 9.53331e-19 $X=3.83 $Y=1.41 $X2=0
+ $Y2=0
cc_548 N_A_475_413#_c_771_n N_VPWR_c_1083_n 0.0138309f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_549 N_A_475_413#_c_763_n N_VPWR_c_1083_n 0.0252179f $X=3.355 $Y=2.19 $X2=0
+ $Y2=0
cc_550 N_A_475_413#_c_759_n N_VPWR_c_1083_n 0.00741701f $X=3.355 $Y=1.41 $X2=0
+ $Y2=0
cc_551 N_A_475_413#_c_771_n N_VPWR_c_1089_n 0.0359536f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_552 N_A_475_413#_M1002_g N_VPWR_c_1091_n 0.00541359f $X=3.905 $Y=2.11 $X2=0
+ $Y2=0
cc_553 N_A_475_413#_M1012_d N_VPWR_c_1080_n 0.00217001f $X=2.375 $Y=2.065 $X2=0
+ $Y2=0
cc_554 N_A_475_413#_M1002_g N_VPWR_c_1080_n 0.00665748f $X=3.905 $Y=2.11 $X2=0
+ $Y2=0
cc_555 N_A_475_413#_c_771_n N_VPWR_c_1080_n 0.0161651f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_556 N_A_475_413#_c_771_n N_A_381_47#_c_1215_n 0.0101821f $X=3.27 $Y=2.275
+ $X2=0 $Y2=0
cc_557 N_A_475_413#_c_771_n A_568_413# 0.0045944f $X=3.27 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_558 N_A_475_413#_c_754_n N_VGND_c_1338_n 0.00816054f $X=4.005 $Y=0.95 $X2=0
+ $Y2=0
cc_559 N_A_475_413#_c_797_n N_VGND_c_1349_n 0.0258035f $X=2.98 $Y=0.45 $X2=0
+ $Y2=0
cc_560 N_A_475_413#_c_754_n N_VGND_c_1350_n 0.00407056f $X=4.005 $Y=0.95 $X2=0
+ $Y2=0
cc_561 N_A_475_413#_M1022_d N_VGND_c_1357_n 0.00225806f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_562 N_A_475_413#_c_754_n N_VGND_c_1357_n 0.00620172f $X=4.005 $Y=0.95 $X2=0
+ $Y2=0
cc_563 N_A_475_413#_c_797_n N_VGND_c_1357_n 0.0114499f $X=2.98 $Y=0.45 $X2=0
+ $Y2=0
cc_564 N_A_475_413#_c_797_n A_572_47# 0.00455507f $X=2.98 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_565 N_A_475_413#_c_758_n A_572_47# 0.00200718f $X=3.065 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_566 N_A_1062_300#_c_863_n N_A_891_413#_c_999_n 0.018057f $X=6.94 $Y=0.995
+ $X2=0 $Y2=0
cc_567 N_A_1062_300#_c_867_n N_A_891_413#_c_999_n 0.0142803f $X=6.505 $Y=0.905
+ $X2=0 $Y2=0
cc_568 N_A_1062_300#_c_868_n N_A_891_413#_c_999_n 0.00471713f $X=6.505 $Y=1.075
+ $X2=0 $Y2=0
cc_569 N_A_1062_300#_M1007_g N_A_891_413#_M1023_g 0.018057f $X=6.94 $Y=1.985
+ $X2=0 $Y2=0
cc_570 N_A_1062_300#_c_869_n N_A_891_413#_M1023_g 0.00927345f $X=6.505 $Y=1.5
+ $X2=0 $Y2=0
cc_571 N_A_1062_300#_c_890_p N_A_891_413#_M1023_g 0.0115645f $X=6.255 $Y=1.61
+ $X2=0 $Y2=0
cc_572 N_A_1062_300#_M1008_g N_A_891_413#_c_1000_n 0.0121715f $X=5.5 $Y=0.445
+ $X2=0 $Y2=0
cc_573 N_A_1062_300#_c_878_n N_A_891_413#_c_1000_n 0.00570311f $X=6.17 $Y=1.665
+ $X2=0 $Y2=0
cc_574 N_A_1062_300#_c_867_n N_A_891_413#_c_1000_n 0.0087082f $X=6.505 $Y=0.905
+ $X2=0 $Y2=0
cc_575 N_A_1062_300#_c_890_p N_A_891_413#_c_1000_n 0.00559631f $X=6.255 $Y=1.61
+ $X2=0 $Y2=0
cc_576 N_A_1062_300#_c_868_n N_A_891_413#_c_1001_n 0.00461715f $X=6.505 $Y=1.075
+ $X2=0 $Y2=0
cc_577 N_A_1062_300#_c_869_n N_A_891_413#_c_1001_n 0.00461715f $X=6.505 $Y=1.5
+ $X2=0 $Y2=0
cc_578 N_A_1062_300#_c_897_p N_A_891_413#_c_1001_n 0.00678299f $X=6.505 $Y=1.16
+ $X2=0 $Y2=0
cc_579 N_A_1062_300#_c_871_n N_A_891_413#_c_1001_n 0.018057f $X=8.215 $Y=1.16
+ $X2=0 $Y2=0
cc_580 N_A_1062_300#_M1020_g N_A_891_413#_c_1010_n 0.00194535f $X=5.385 $Y=2.275
+ $X2=0 $Y2=0
cc_581 N_A_1062_300#_M1008_g N_A_891_413#_c_1013_n 0.00171633f $X=5.5 $Y=0.445
+ $X2=0 $Y2=0
cc_582 N_A_1062_300#_M1008_g N_A_891_413#_c_1002_n 0.011078f $X=5.5 $Y=0.445
+ $X2=0 $Y2=0
cc_583 N_A_1062_300#_M1008_g N_A_891_413#_c_1003_n 0.00717747f $X=5.5 $Y=0.445
+ $X2=0 $Y2=0
cc_584 N_A_1062_300#_c_878_n N_A_891_413#_c_1003_n 0.0262086f $X=6.17 $Y=1.665
+ $X2=0 $Y2=0
cc_585 N_A_1062_300#_c_879_n N_A_891_413#_c_1003_n 0.012028f $X=5.565 $Y=1.665
+ $X2=0 $Y2=0
cc_586 N_A_1062_300#_M1008_g N_A_891_413#_c_1004_n 0.0172589f $X=5.5 $Y=0.445
+ $X2=0 $Y2=0
cc_587 N_A_1062_300#_c_878_n N_A_891_413#_c_1004_n 0.0388789f $X=6.17 $Y=1.665
+ $X2=0 $Y2=0
cc_588 N_A_1062_300#_c_879_n N_A_891_413#_c_1004_n 0.00698627f $X=5.565 $Y=1.665
+ $X2=0 $Y2=0
cc_589 N_A_1062_300#_c_867_n N_A_891_413#_c_1004_n 0.0111887f $X=6.505 $Y=0.905
+ $X2=0 $Y2=0
cc_590 N_A_1062_300#_c_890_p N_A_891_413#_c_1004_n 0.00346944f $X=6.255 $Y=1.61
+ $X2=0 $Y2=0
cc_591 N_A_1062_300#_c_897_p N_A_891_413#_c_1004_n 0.0129954f $X=6.505 $Y=1.16
+ $X2=0 $Y2=0
cc_592 N_A_1062_300#_M1020_g N_VPWR_c_1084_n 0.00461184f $X=5.385 $Y=2.275 $X2=0
+ $Y2=0
cc_593 N_A_1062_300#_c_878_n N_VPWR_c_1084_n 0.0104755f $X=6.17 $Y=1.665 $X2=0
+ $Y2=0
cc_594 N_A_1062_300#_c_879_n N_VPWR_c_1084_n 0.00467318f $X=5.565 $Y=1.665 $X2=0
+ $Y2=0
cc_595 N_A_1062_300#_c_914_p N_VPWR_c_1084_n 0.0112508f $X=6.255 $Y=1.95 $X2=0
+ $Y2=0
cc_596 N_A_1062_300#_M1007_g N_VPWR_c_1085_n 0.00604944f $X=6.94 $Y=1.985 $X2=0
+ $Y2=0
cc_597 N_A_1062_300#_c_870_n N_VPWR_c_1085_n 0.00582033f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_598 N_A_1062_300#_M1015_g N_VPWR_c_1086_n 0.00602529f $X=7.36 $Y=1.985 $X2=0
+ $Y2=0
cc_599 N_A_1062_300#_M1021_g N_VPWR_c_1086_n 0.00148704f $X=7.795 $Y=1.985 $X2=0
+ $Y2=0
cc_600 N_A_1062_300#_M1025_g N_VPWR_c_1088_n 0.00316354f $X=8.215 $Y=1.985 $X2=0
+ $Y2=0
cc_601 N_A_1062_300#_M1020_g N_VPWR_c_1091_n 0.00585385f $X=5.385 $Y=2.275 $X2=0
+ $Y2=0
cc_602 N_A_1062_300#_M1007_g N_VPWR_c_1093_n 0.0054411f $X=6.94 $Y=1.985 $X2=0
+ $Y2=0
cc_603 N_A_1062_300#_M1015_g N_VPWR_c_1093_n 0.00536993f $X=7.36 $Y=1.985 $X2=0
+ $Y2=0
cc_604 N_A_1062_300#_c_914_p N_VPWR_c_1097_n 0.0109058f $X=6.255 $Y=1.95 $X2=0
+ $Y2=0
cc_605 N_A_1062_300#_M1021_g N_VPWR_c_1098_n 0.0054411f $X=7.795 $Y=1.985 $X2=0
+ $Y2=0
cc_606 N_A_1062_300#_M1025_g N_VPWR_c_1098_n 0.0054411f $X=8.215 $Y=1.985 $X2=0
+ $Y2=0
cc_607 N_A_1062_300#_M1023_s N_VPWR_c_1080_n 0.00611269f $X=6.11 $Y=1.485 $X2=0
+ $Y2=0
cc_608 N_A_1062_300#_M1020_g N_VPWR_c_1080_n 0.0122833f $X=5.385 $Y=2.275 $X2=0
+ $Y2=0
cc_609 N_A_1062_300#_M1007_g N_VPWR_c_1080_n 0.00969004f $X=6.94 $Y=1.985 $X2=0
+ $Y2=0
cc_610 N_A_1062_300#_M1015_g N_VPWR_c_1080_n 0.00940158f $X=7.36 $Y=1.985 $X2=0
+ $Y2=0
cc_611 N_A_1062_300#_M1021_g N_VPWR_c_1080_n 0.00954766f $X=7.795 $Y=1.985 $X2=0
+ $Y2=0
cc_612 N_A_1062_300#_M1025_g N_VPWR_c_1080_n 0.0105113f $X=8.215 $Y=1.985 $X2=0
+ $Y2=0
cc_613 N_A_1062_300#_c_914_p N_VPWR_c_1080_n 0.00643939f $X=6.255 $Y=1.95 $X2=0
+ $Y2=0
cc_614 N_A_1062_300#_c_864_n N_Q_c_1249_n 0.00832844f $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_615 N_A_1062_300#_c_865_n N_Q_c_1249_n 0.00860437f $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_616 N_A_1062_300#_c_870_n N_Q_c_1249_n 0.0354432f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_617 N_A_1062_300#_c_871_n N_Q_c_1249_n 0.00257975f $X=8.215 $Y=1.16 $X2=0
+ $Y2=0
cc_618 N_A_1062_300#_c_863_n N_Q_c_1250_n 0.00324219f $X=6.94 $Y=0.995 $X2=0
+ $Y2=0
cc_619 N_A_1062_300#_c_864_n N_Q_c_1250_n 0.00120512f $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_620 N_A_1062_300#_c_867_n N_Q_c_1250_n 0.00402715f $X=6.505 $Y=0.905 $X2=0
+ $Y2=0
cc_621 N_A_1062_300#_c_870_n N_Q_c_1250_n 0.0258576f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_622 N_A_1062_300#_c_871_n N_Q_c_1250_n 0.00229134f $X=8.215 $Y=1.16 $X2=0
+ $Y2=0
cc_623 N_A_1062_300#_M1015_g N_Q_c_1254_n 0.0106705f $X=7.36 $Y=1.985 $X2=0
+ $Y2=0
cc_624 N_A_1062_300#_M1021_g N_Q_c_1254_n 0.0110491f $X=7.795 $Y=1.985 $X2=0
+ $Y2=0
cc_625 N_A_1062_300#_c_870_n N_Q_c_1254_n 0.029722f $X=8.075 $Y=1.16 $X2=0 $Y2=0
cc_626 N_A_1062_300#_c_871_n N_Q_c_1254_n 0.00250357f $X=8.215 $Y=1.16 $X2=0
+ $Y2=0
cc_627 N_A_1062_300#_c_864_n N_Q_c_1272_n 5.11724e-19 $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_628 N_A_1062_300#_c_865_n N_Q_c_1272_n 0.00597981f $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_629 N_A_1062_300#_c_866_n N_Q_c_1272_n 0.0107208f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_630 N_A_1062_300#_M1015_g N_Q_c_1275_n 6.04594e-19 $X=7.36 $Y=1.985 $X2=0
+ $Y2=0
cc_631 N_A_1062_300#_M1021_g N_Q_c_1275_n 0.00947724f $X=7.795 $Y=1.985 $X2=0
+ $Y2=0
cc_632 N_A_1062_300#_M1025_g N_Q_c_1275_n 0.0142067f $X=8.215 $Y=1.985 $X2=0
+ $Y2=0
cc_633 N_A_1062_300#_M1025_g N_Q_c_1255_n 0.0129914f $X=8.215 $Y=1.985 $X2=0
+ $Y2=0
cc_634 N_A_1062_300#_c_870_n N_Q_c_1255_n 0.00383323f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_635 N_A_1062_300#_c_866_n N_Q_c_1251_n 0.0104229f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_636 N_A_1062_300#_c_870_n N_Q_c_1251_n 0.00427132f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_637 N_A_1062_300#_c_866_n N_Q_c_1252_n 0.0208834f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_638 N_A_1062_300#_c_870_n N_Q_c_1252_n 0.0137873f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_639 N_A_1062_300#_M1007_g N_Q_c_1257_n 0.00336273f $X=6.94 $Y=1.985 $X2=0
+ $Y2=0
cc_640 N_A_1062_300#_M1015_g N_Q_c_1257_n 0.00134785f $X=7.36 $Y=1.985 $X2=0
+ $Y2=0
cc_641 N_A_1062_300#_c_869_n N_Q_c_1257_n 0.00114511f $X=6.505 $Y=1.5 $X2=0
+ $Y2=0
cc_642 N_A_1062_300#_c_870_n N_Q_c_1257_n 0.0220011f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_643 N_A_1062_300#_c_871_n N_Q_c_1257_n 0.00225167f $X=8.215 $Y=1.16 $X2=0
+ $Y2=0
cc_644 N_A_1062_300#_c_865_n N_Q_c_1253_n 0.00105193f $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_645 N_A_1062_300#_c_866_n N_Q_c_1253_n 0.0011466f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_646 N_A_1062_300#_c_870_n N_Q_c_1253_n 0.0258576f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_647 N_A_1062_300#_c_871_n N_Q_c_1253_n 0.00229134f $X=8.215 $Y=1.16 $X2=0
+ $Y2=0
cc_648 N_A_1062_300#_M1021_g N_Q_c_1258_n 0.0011847f $X=7.795 $Y=1.985 $X2=0
+ $Y2=0
cc_649 N_A_1062_300#_M1025_g N_Q_c_1258_n 0.0011847f $X=8.215 $Y=1.985 $X2=0
+ $Y2=0
cc_650 N_A_1062_300#_c_870_n N_Q_c_1258_n 0.0216915f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_651 N_A_1062_300#_c_871_n N_Q_c_1258_n 0.00225167f $X=8.215 $Y=1.16 $X2=0
+ $Y2=0
cc_652 N_A_1062_300#_M1007_g Q 0.0103228f $X=6.94 $Y=1.985 $X2=0 $Y2=0
cc_653 N_A_1062_300#_M1015_g Q 0.00992901f $X=7.36 $Y=1.985 $X2=0 $Y2=0
cc_654 N_A_1062_300#_M1021_g Q 6.20474e-19 $X=7.795 $Y=1.985 $X2=0 $Y2=0
cc_655 N_A_1062_300#_c_863_n N_Q_c_1300_n 0.00612348f $X=6.94 $Y=0.995 $X2=0
+ $Y2=0
cc_656 N_A_1062_300#_c_864_n N_Q_c_1300_n 0.00617761f $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_657 N_A_1062_300#_c_865_n N_Q_c_1300_n 5.17178e-19 $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_658 N_A_1062_300#_c_867_n N_Q_c_1300_n 0.00487223f $X=6.505 $Y=0.905 $X2=0
+ $Y2=0
cc_659 N_A_1062_300#_M1008_g N_VGND_c_1339_n 0.00475832f $X=5.5 $Y=0.445 $X2=0
+ $Y2=0
cc_660 N_A_1062_300#_c_867_n N_VGND_c_1339_n 0.0170073f $X=6.505 $Y=0.905 $X2=0
+ $Y2=0
cc_661 N_A_1062_300#_c_867_n N_VGND_c_1340_n 0.0200466f $X=6.505 $Y=0.905 $X2=0
+ $Y2=0
cc_662 N_A_1062_300#_c_863_n N_VGND_c_1341_n 0.00474311f $X=6.94 $Y=0.995 $X2=0
+ $Y2=0
cc_663 N_A_1062_300#_c_867_n N_VGND_c_1341_n 0.0197221f $X=6.505 $Y=0.905 $X2=0
+ $Y2=0
cc_664 N_A_1062_300#_c_870_n N_VGND_c_1341_n 0.00626932f $X=8.075 $Y=1.16 $X2=0
+ $Y2=0
cc_665 N_A_1062_300#_c_864_n N_VGND_c_1342_n 0.00469816f $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_666 N_A_1062_300#_c_865_n N_VGND_c_1342_n 0.0026837f $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_667 N_A_1062_300#_c_866_n N_VGND_c_1344_n 0.00434782f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_668 N_A_1062_300#_c_863_n N_VGND_c_1345_n 0.00543342f $X=6.94 $Y=0.995 $X2=0
+ $Y2=0
cc_669 N_A_1062_300#_c_864_n N_VGND_c_1345_n 0.00423505f $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_670 N_A_1062_300#_M1008_g N_VGND_c_1350_n 0.00585385f $X=5.5 $Y=0.445 $X2=0
+ $Y2=0
cc_671 N_A_1062_300#_c_865_n N_VGND_c_1351_n 0.00425859f $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_672 N_A_1062_300#_c_866_n N_VGND_c_1351_n 0.00423505f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_673 N_A_1062_300#_M1017_s N_VGND_c_1357_n 0.00211564f $X=6.13 $Y=0.235 $X2=0
+ $Y2=0
cc_674 N_A_1062_300#_M1008_g N_VGND_c_1357_n 0.0122284f $X=5.5 $Y=0.445 $X2=0
+ $Y2=0
cc_675 N_A_1062_300#_c_863_n N_VGND_c_1357_n 0.00971227f $X=6.94 $Y=0.995 $X2=0
+ $Y2=0
cc_676 N_A_1062_300#_c_864_n N_VGND_c_1357_n 0.005767f $X=7.36 $Y=0.995 $X2=0
+ $Y2=0
cc_677 N_A_1062_300#_c_865_n N_VGND_c_1357_n 0.00578199f $X=7.795 $Y=0.995 $X2=0
+ $Y2=0
cc_678 N_A_1062_300#_c_866_n N_VGND_c_1357_n 0.00671804f $X=8.215 $Y=0.995 $X2=0
+ $Y2=0
cc_679 N_A_1062_300#_c_867_n N_VGND_c_1357_n 0.0166104f $X=6.505 $Y=0.905 $X2=0
+ $Y2=0
cc_680 N_A_891_413#_M1023_g N_VPWR_c_1084_n 0.00248819f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_681 N_A_891_413#_M1023_g N_VPWR_c_1085_n 0.00565423f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_682 N_A_891_413#_c_1010_n N_VPWR_c_1091_n 0.0273845f $X=5.14 $Y=2.25 $X2=0
+ $Y2=0
cc_683 N_A_891_413#_M1023_g N_VPWR_c_1097_n 0.00585385f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_684 N_A_891_413#_M1019_d N_VPWR_c_1080_n 0.00217593f $X=4.455 $Y=2.065 $X2=0
+ $Y2=0
cc_685 N_A_891_413#_M1023_g N_VPWR_c_1080_n 0.0121077f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_686 N_A_891_413#_c_1010_n N_VPWR_c_1080_n 0.0274677f $X=5.14 $Y=2.25 $X2=0
+ $Y2=0
cc_687 N_A_891_413#_c_1010_n A_975_413# 0.0105858f $X=5.14 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_688 N_A_891_413#_c_1003_n A_975_413# 0.00184879f $X=5.225 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_689 N_A_891_413#_M1023_g Q 6.91159e-19 $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_690 N_A_891_413#_c_999_n N_Q_c_1300_n 5.01503e-19 $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_691 N_A_891_413#_c_999_n N_VGND_c_1339_n 0.00231174f $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_692 N_A_891_413#_c_1004_n N_VGND_c_1339_n 0.00667571f $X=6.065 $Y=1.16 $X2=0
+ $Y2=0
cc_693 N_A_891_413#_c_999_n N_VGND_c_1340_n 0.00409806f $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_694 N_A_891_413#_c_999_n N_VGND_c_1341_n 0.00439958f $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_695 N_A_891_413#_c_1013_n N_VGND_c_1350_n 0.0234603f $X=5.14 $Y=0.45 $X2=0
+ $Y2=0
cc_696 N_A_891_413#_M1003_d N_VGND_c_1357_n 0.00333348f $X=4.585 $Y=0.235 $X2=0
+ $Y2=0
cc_697 N_A_891_413#_c_999_n N_VGND_c_1357_n 0.00714808f $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_698 N_A_891_413#_c_1013_n N_VGND_c_1357_n 0.0227598f $X=5.14 $Y=0.45 $X2=0
+ $Y2=0
cc_699 N_A_891_413#_c_1013_n A_1020_47# 0.00400578f $X=5.14 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_700 N_A_891_413#_c_1002_n A_1020_47# 0.00147605f $X=5.225 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_701 N_VPWR_c_1080_n N_A_381_47#_M1018_d 0.00274646f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_1089_n N_A_381_47#_c_1215_n 0.0122088f $X=3.61 $Y=2.72 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_1080_n N_A_381_47#_c_1215_n 0.00414216f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_1080_n A_568_413# 0.00220276f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_705 N_VPWR_c_1080_n A_975_413# 0.00377587f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_706 N_VPWR_c_1080_n N_Q_M1007_s 0.00220947f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_707 N_VPWR_c_1080_n N_Q_M1021_s 0.00220947f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_708 N_VPWR_M1015_d N_Q_c_1254_n 0.00206549f $X=7.435 $Y=1.485 $X2=0 $Y2=0
cc_709 N_VPWR_c_1086_n N_Q_c_1254_n 0.0131801f $X=7.585 $Y=1.97 $X2=0 $Y2=0
cc_710 N_VPWR_c_1098_n N_Q_c_1275_n 0.013082f $X=8.34 $Y=2.72 $X2=0 $Y2=0
cc_711 N_VPWR_c_1080_n N_Q_c_1275_n 0.0117641f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_712 N_VPWR_M1025_d N_Q_c_1255_n 0.00533663f $X=8.29 $Y=1.485 $X2=0 $Y2=0
cc_713 N_VPWR_c_1088_n N_Q_c_1255_n 0.0140151f $X=8.425 $Y=1.97 $X2=0 $Y2=0
cc_714 N_VPWR_c_1085_n Q 0.0383541f $X=6.71 $Y=2.02 $X2=0 $Y2=0
cc_715 N_VPWR_c_1086_n Q 0.0417286f $X=7.585 $Y=1.97 $X2=0 $Y2=0
cc_716 N_VPWR_c_1093_n Q 0.0133145f $X=7.5 $Y=2.72 $X2=0 $Y2=0
cc_717 N_VPWR_c_1080_n Q 0.0119259f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_718 N_A_381_47#_c_1221_n N_VGND_c_1349_n 0.0106218f $X=2.055 $Y=0.45 $X2=0
+ $Y2=0
cc_719 N_A_381_47#_M1001_d N_VGND_c_1357_n 0.00232113f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_720 N_A_381_47#_c_1221_n N_VGND_c_1357_n 0.0051217f $X=2.055 $Y=0.45 $X2=0
+ $Y2=0
cc_721 N_Q_c_1249_n N_VGND_M1005_d 0.00173322f $X=7.84 $Y=0.815 $X2=0 $Y2=0
cc_722 N_Q_c_1251_n N_VGND_M1029_d 0.00388224f $X=8.41 $Y=0.815 $X2=0 $Y2=0
cc_723 N_Q_c_1300_n N_VGND_c_1341_n 0.0176379f $X=7.15 $Y=0.395 $X2=0 $Y2=0
cc_724 N_Q_c_1249_n N_VGND_c_1342_n 0.0130881f $X=7.84 $Y=0.815 $X2=0 $Y2=0
cc_725 N_Q_c_1300_n N_VGND_c_1342_n 0.0184321f $X=7.15 $Y=0.395 $X2=0 $Y2=0
cc_726 N_Q_c_1251_n N_VGND_c_1343_n 0.00230956f $X=8.41 $Y=0.815 $X2=0 $Y2=0
cc_727 N_Q_c_1251_n N_VGND_c_1344_n 0.013909f $X=8.41 $Y=0.815 $X2=0 $Y2=0
cc_728 N_Q_c_1249_n N_VGND_c_1345_n 0.00198954f $X=7.84 $Y=0.815 $X2=0 $Y2=0
cc_729 N_Q_c_1300_n N_VGND_c_1345_n 0.0144978f $X=7.15 $Y=0.395 $X2=0 $Y2=0
cc_730 N_Q_c_1249_n N_VGND_c_1351_n 0.00199746f $X=7.84 $Y=0.815 $X2=0 $Y2=0
cc_731 N_Q_c_1272_n N_VGND_c_1351_n 0.0144978f $X=8.005 $Y=0.395 $X2=0 $Y2=0
cc_732 N_Q_c_1251_n N_VGND_c_1351_n 0.00193122f $X=8.41 $Y=0.815 $X2=0 $Y2=0
cc_733 N_Q_M1004_s N_VGND_c_1357_n 0.00218509f $X=7.015 $Y=0.235 $X2=0 $Y2=0
cc_734 N_Q_M1010_s N_VGND_c_1357_n 0.00218509f $X=7.87 $Y=0.235 $X2=0 $Y2=0
cc_735 N_Q_c_1249_n N_VGND_c_1357_n 0.00862624f $X=7.84 $Y=0.815 $X2=0 $Y2=0
cc_736 N_Q_c_1272_n N_VGND_c_1357_n 0.0120158f $X=8.005 $Y=0.395 $X2=0 $Y2=0
cc_737 N_Q_c_1251_n N_VGND_c_1357_n 0.00851067f $X=8.41 $Y=0.815 $X2=0 $Y2=0
cc_738 N_Q_c_1300_n N_VGND_c_1357_n 0.0120158f $X=7.15 $Y=0.395 $X2=0 $Y2=0
cc_739 N_VGND_c_1357_n A_572_47# 0.00272292f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
cc_740 N_VGND_c_1357_n A_1020_47# 0.00669936f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24

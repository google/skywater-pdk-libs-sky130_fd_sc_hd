* File: sky130_fd_sc_hd__a41oi_1.spice
* Created: Thu Aug 27 14:06:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a41oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a41oi_1  VNB VPB B1 A4 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.163425 AS=0.169 PD=1.175 PS=1.82 NRD=19.38 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1009 A_236_47# N_A4_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65 AD=0.11375
+ AS=0.163425 PD=1 PS=1.175 NRD=22.152 NRS=20.304 M=1 R=4.33333 SA=75000.8
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1007 A_336_47# N_A3_M1007_g A_236_47# VNB NSHORT L=0.15 W=0.65 AD=0.10075
+ AS=0.11375 PD=0.96 PS=1 NRD=18.456 NRS=22.152 M=1 R=4.33333 SA=75001.3
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1001 A_428_47# N_A2_M1001_g A_336_47# VNB NSHORT L=0.15 W=0.65 AD=0.138125
+ AS=0.10075 PD=1.075 PS=0.96 NRD=29.076 NRS=18.456 M=1 R=4.33333 SA=75001.8
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A1_M1004_g A_428_47# VNB NSHORT L=0.15 W=0.65 AD=0.2405
+ AS=0.138125 PD=2.04 PS=1.075 NRD=0 NRS=29.076 M=1 R=4.33333 SA=75002.4
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1006 N_A_109_297#_M1006_d N_B1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2125 AS=0.26 PD=1.425 PS=2.52 NRD=14.7553 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A4_M1000_g N_A_109_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.205 AS=0.2125 PD=1.41 PS=1.425 NRD=4.9053 NRS=13.7703 M=1 R=6.66667
+ SA=75000.8 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1005 N_A_109_297#_M1005_d N_A3_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.205 PD=1.31 PS=1.41 NRD=4.9053 NRS=20.685 M=1 R=6.66667
+ SA=75001.3 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_109_297#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.2125 AS=0.155 PD=1.425 PS=1.31 NRD=19.7 NRS=0.9653 M=1 R=6.66667
+ SA=75001.8 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1003 N_A_109_297#_M1003_d N_A1_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.37 AS=0.2125 PD=2.74 PS=1.425 NRD=0 NRS=8.8453 M=1 R=6.66667 SA=75002.4
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a41oi_1.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__mux4_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__mux4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.540000 0.375000 6.850000 0.995000 ;
        RECT 6.540000 0.995000 6.950000 1.075000 ;
        RECT 6.640000 1.075000 6.950000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 0.715000 5.120000 1.395000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 0.765000 1.240000 1.095000 ;
        RECT 1.025000 0.395000 1.240000 0.765000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 0.715000 2.620000 1.015000 ;
        RECT 2.415000 1.015000 2.620000 1.320000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.975000 0.330000 1.745000 ;
        RECT 1.010000 1.445000 1.395000 1.615000 ;
        RECT 1.225000 1.285000 1.395000 1.445000 ;
        RECT 6.130000 1.245000 6.470000 1.645000 ;
      LAYER mcon ;
        RECT 0.150000 1.445000 0.320000 1.615000 ;
        RECT 1.070000 1.445000 1.240000 1.615000 ;
        RECT 6.130000 1.445000 6.300000 1.615000 ;
      LAYER met1 ;
        RECT 0.085000 1.415000 0.380000 1.460000 ;
        RECT 0.085000 1.460000 6.360000 1.600000 ;
        RECT 0.085000 1.600000 0.380000 1.645000 ;
        RECT 1.010000 1.415000 1.300000 1.460000 ;
        RECT 1.010000 1.600000 1.300000 1.645000 ;
        RECT 6.070000 1.415000 6.360000 1.460000 ;
        RECT 6.070000 1.600000 6.360000 1.645000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.715000 3.080000 1.320000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.360000 1.835000 7.770000 2.455000 ;
        RECT 7.440000 0.265000 7.770000 0.725000 ;
        RECT 7.460000 1.495000 7.770000 1.835000 ;
        RECT 7.600000 0.725000 7.770000 1.065000 ;
        RECT 7.600000 1.065000 8.685000 1.305000 ;
        RECT 7.600000 1.305000 7.770000 1.495000 ;
        RECT 8.360000 0.265000 8.685000 1.065000 ;
        RECT 8.360000 1.305000 8.685000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.200000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 2.455000  0.085000 2.785000 0.545000 ;
        RECT 4.800000  0.085000 5.130000 0.545000 ;
        RECT 7.020000  0.085000 7.270000 0.815000 ;
        RECT 7.940000  0.085000 8.190000 0.885000 ;
        RECT 8.855000  0.085000 9.105000 0.885000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.200000 2.805000 ;
        RECT 0.515000 2.255000 0.845000 2.635000 ;
        RECT 2.600000 2.055000 2.830000 2.635000 ;
        RECT 4.760000 2.005000 5.105000 2.635000 ;
        RECT 7.020000 1.835000 7.190000 2.635000 ;
        RECT 7.940000 1.495000 8.190000 2.635000 ;
        RECT 8.855000 1.495000 9.105000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.135000 0.345000 0.345000 0.635000 ;
      RECT 0.135000 0.635000 0.670000 0.805000 ;
      RECT 0.135000 1.915000 1.905000 1.955000 ;
      RECT 0.135000 1.955000 0.670000 2.085000 ;
      RECT 0.135000 2.085000 0.345000 2.375000 ;
      RECT 0.500000 0.805000 0.670000 1.785000 ;
      RECT 0.500000 1.785000 1.905000 1.915000 ;
      RECT 1.410000 0.705000 1.735000 1.035000 ;
      RECT 1.415000 2.125000 2.245000 2.295000 ;
      RECT 1.475000 0.365000 2.075000 0.535000 ;
      RECT 1.565000 1.035000 1.735000 1.575000 ;
      RECT 1.565000 1.575000 1.905000 1.785000 ;
      RECT 1.905000 0.535000 2.075000 1.235000 ;
      RECT 1.905000 1.235000 2.245000 1.405000 ;
      RECT 2.075000 1.405000 2.245000 2.125000 ;
      RECT 2.975000 1.785000 3.320000 1.955000 ;
      RECT 2.990000 0.295000 3.420000 0.465000 ;
      RECT 3.150000 1.490000 3.420000 1.660000 ;
      RECT 3.150000 1.660000 3.320000 1.785000 ;
      RECT 3.250000 0.465000 3.420000 1.060000 ;
      RECT 3.250000 1.060000 3.485000 1.390000 ;
      RECT 3.250000 1.390000 3.420000 1.490000 ;
      RECT 3.310000 2.125000 3.825000 2.295000 ;
      RECT 3.575000 1.810000 3.825000 2.125000 ;
      RECT 3.590000 0.345000 3.825000 0.675000 ;
      RECT 3.655000 0.675000 3.825000 1.810000 ;
      RECT 3.995000 0.345000 4.185000 2.125000 ;
      RECT 3.995000 2.125000 4.520000 2.295000 ;
      RECT 4.400000 0.255000 4.605000 0.585000 ;
      RECT 4.400000 0.585000 4.570000 1.565000 ;
      RECT 4.400000 1.565000 5.500000 1.735000 ;
      RECT 4.400000 1.735000 4.590000 1.895000 ;
      RECT 5.330000 0.295000 6.225000 0.465000 ;
      RECT 5.330000 0.465000 5.500000 1.565000 ;
      RECT 5.330000 1.735000 5.500000 2.155000 ;
      RECT 5.330000 2.155000 6.280000 2.325000 ;
      RECT 5.670000 0.705000 6.290000 1.035000 ;
      RECT 5.670000 1.035000 5.960000 1.985000 ;
      RECT 6.530000 2.125000 6.850000 2.295000 ;
      RECT 6.680000 1.495000 7.290000 1.665000 ;
      RECT 6.680000 1.665000 6.850000 2.125000 ;
      RECT 7.120000 0.995000 7.430000 1.325000 ;
      RECT 7.120000 1.325000 7.290000 1.495000 ;
    LAYER mcon ;
      RECT 1.530000 1.785000 1.700000 1.955000 ;
      RECT 1.990000 2.125000 2.160000 2.295000 ;
      RECT 3.370000 2.125000 3.540000 2.295000 ;
      RECT 4.290000 2.125000 4.460000 2.295000 ;
      RECT 5.670000 1.785000 5.840000 1.955000 ;
      RECT 6.590000 2.125000 6.760000 2.295000 ;
    LAYER met1 ;
      RECT 1.470000 1.755000 1.760000 1.800000 ;
      RECT 1.470000 1.800000 5.900000 1.940000 ;
      RECT 1.470000 1.940000 1.760000 1.985000 ;
      RECT 1.930000 2.095000 2.220000 2.140000 ;
      RECT 1.930000 2.140000 3.600000 2.280000 ;
      RECT 1.930000 2.280000 2.220000 2.325000 ;
      RECT 3.310000 2.095000 3.600000 2.140000 ;
      RECT 3.310000 2.280000 3.600000 2.325000 ;
      RECT 4.230000 2.095000 4.520000 2.140000 ;
      RECT 4.230000 2.140000 6.820000 2.280000 ;
      RECT 4.230000 2.280000 4.520000 2.325000 ;
      RECT 5.610000 1.755000 5.900000 1.800000 ;
      RECT 5.610000 1.940000 5.900000 1.985000 ;
      RECT 6.530000 2.095000 6.820000 2.140000 ;
      RECT 6.530000 2.280000 6.820000 2.325000 ;
  END
END sky130_fd_sc_hd__mux4_4

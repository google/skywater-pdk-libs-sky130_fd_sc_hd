# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__sdfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.410000 0.275000 13.740000 0.825000 ;
        RECT 13.410000 1.495000 13.740000 2.450000 ;
        RECT 13.515000 0.825000 13.740000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.460000 0.255000 11.855000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
        RECT 2.405000 1.075000 2.735000 1.590000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
        RECT 8.880000 1.435000 9.115000 1.525000 ;
        RECT 8.880000 1.525000 9.935000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.100000 1.970000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.260000 0.085000 ;
        RECT  0.085000  0.085000  0.700000 0.595000 ;
        RECT  1.840000  0.085000  2.090000 0.545000 ;
        RECT  2.700000  0.085000  3.100000 0.555000 ;
        RECT  3.640000  0.085000  3.940000 0.545000 ;
        RECT  5.665000  0.085000  6.165000 0.465000 ;
        RECT  6.720000  0.085000  7.705000 0.805000 ;
        RECT 10.035000  0.085000 10.285000 0.545000 ;
        RECT 11.120000  0.085000 11.290000 0.885000 ;
        RECT 12.025000  0.085000 12.315000 0.885000 ;
        RECT 12.885000  0.085000 13.240000 0.825000 ;
        RECT 13.910000  0.085000 14.175000 0.885000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 14.260000 2.805000 ;
        RECT  0.515000 2.275000  0.845000 2.635000 ;
        RECT  2.705000 2.140000  3.100000 2.635000 ;
        RECT  3.645000 2.275000  3.975000 2.635000 ;
        RECT  6.000000 2.275000  6.330000 2.635000 ;
        RECT  7.060000 2.125000  8.015000 2.635000 ;
        RECT  9.160000 2.235000  9.490000 2.635000 ;
        RECT 10.100000 2.235000 10.430000 2.635000 ;
        RECT 11.080000 1.485000 11.290000 2.635000 ;
        RECT 12.025000 1.485000 12.315000 2.635000 ;
        RECT 12.885000 1.635000 13.240000 2.635000 ;
        RECT 13.910000 1.485000 14.175000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
        RECT 13.945000 2.635000 14.115000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 1.845000  1.185000 2.075000 ;
      RECT  0.085000 2.075000  0.345000 2.465000 ;
      RECT  0.870000 0.255000  1.670000 0.595000 ;
      RECT  1.015000 2.075000  1.185000 2.255000 ;
      RECT  1.015000 2.255000  2.105000 2.465000 ;
      RECT  1.355000 1.845000  1.695000 2.085000 ;
      RECT  1.495000 0.595000  1.670000 0.645000 ;
      RECT  1.495000 0.645000  1.695000 0.705000 ;
      RECT  1.500000 0.705000  1.695000 0.720000 ;
      RECT  1.505000 0.720000  1.695000 1.845000 ;
      RECT  1.980000 0.715000  2.530000 0.905000 ;
      RECT  1.980000 0.905000  2.235000 1.760000 ;
      RECT  1.980000 1.760000  2.535000 2.085000 ;
      RECT  2.260000 0.255000  2.530000 0.715000 ;
      RECT  2.275000 2.085000  2.535000 2.465000 ;
      RECT  3.270000 0.255000  3.470000 0.715000 ;
      RECT  3.270000 0.715000  3.995000 0.885000 ;
      RECT  3.270000 1.830000  3.995000 2.000000 ;
      RECT  3.270000 2.000000  3.475000 2.325000 ;
      RECT  3.735000 0.885000  3.995000 1.830000 ;
      RECT  4.110000 0.255000  4.335000 0.585000 ;
      RECT  4.145000 2.135000  4.440000 2.465000 ;
      RECT  4.165000 0.585000  4.335000 1.090000 ;
      RECT  4.165000 1.090000  4.490000 1.420000 ;
      RECT  4.165000 1.420000  4.440000 2.135000 ;
      RECT  4.505000 0.255000  4.885000 0.920000 ;
      RECT  4.665000 1.590000  4.970000 1.615000 ;
      RECT  4.665000 1.615000  4.890000 2.465000 ;
      RECT  4.715000 0.920000  4.885000 1.445000 ;
      RECT  4.715000 1.445000  4.970000 1.590000 ;
      RECT  5.055000 0.255000  5.450000 1.225000 ;
      RECT  5.055000 1.225000  7.705000 1.275000 ;
      RECT  5.060000 2.135000  5.805000 2.465000 ;
      RECT  5.140000 1.275000  6.475000 1.395000 ;
      RECT  5.205000 1.575000  5.465000 1.955000 ;
      RECT  5.620000 0.635000  6.550000 0.805000 ;
      RECT  5.620000 0.805000  6.015000 1.015000 ;
      RECT  5.635000 1.395000  5.805000 2.135000 ;
      RECT  5.975000 1.575000  6.145000 1.935000 ;
      RECT  5.975000 1.935000  6.820000 2.105000 ;
      RECT  6.305000 0.975000  7.705000 1.225000 ;
      RECT  6.335000 0.255000  6.550000 0.635000 ;
      RECT  6.605000 2.105000  6.820000 2.450000 ;
      RECT  7.355000 1.275000  7.705000 1.325000 ;
      RECT  7.385000 1.705000  8.055000 1.955000 ;
      RECT  7.885000 0.695000  9.085000 0.895000 ;
      RECT  7.885000 0.895000  8.055000 1.705000 ;
      RECT  8.185000 2.125000  8.990000 2.460000 ;
      RECT  8.420000 1.075000  8.650000 1.905000 ;
      RECT  8.465000 0.275000  9.855000 0.515000 ;
      RECT  8.820000 1.895000 10.430000 2.065000 ;
      RECT  8.820000 2.065000  8.990000 2.125000 ;
      RECT  8.830000 0.895000  9.085000 1.265000 ;
      RECT  9.285000 0.855000  9.515000 1.185000 ;
      RECT  9.285000 1.185000 10.910000 1.355000 ;
      RECT  9.660000 2.065000  9.930000 2.450000 ;
      RECT  9.685000 0.515000  9.855000 0.845000 ;
      RECT  9.685000 0.845000 10.560000 1.015000 ;
      RECT 10.105000 1.525000 10.430000 1.895000 ;
      RECT 10.465000 0.255000 10.910000 0.585000 ;
      RECT 10.600000 1.355000 10.845000 2.465000 ;
      RECT 10.730000 0.585000 10.910000 1.185000 ;
      RECT 12.530000 0.255000 12.715000 0.995000 ;
      RECT 12.530000 0.995000 13.345000 1.325000 ;
      RECT 12.530000 1.325000 12.715000 2.465000 ;
    LAYER mcon ;
      RECT 1.525000 1.445000 1.695000 1.615000 ;
      RECT 3.825000 1.785000 3.995000 1.955000 ;
      RECT 4.285000 1.105000 4.455000 1.275000 ;
      RECT 4.800000 1.445000 4.970000 1.615000 ;
      RECT 5.260000 1.785000 5.430000 1.955000 ;
      RECT 7.560000 1.785000 7.730000 1.955000 ;
      RECT 8.480000 1.105000 8.650000 1.275000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 5.030000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.740000 1.415000 5.030000 1.460000 ;
      RECT 4.740000 1.600000 5.030000 1.645000 ;
      RECT 5.200000 1.755000 5.490000 1.800000 ;
      RECT 5.200000 1.940000 5.490000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfsbp_2
